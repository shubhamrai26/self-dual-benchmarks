module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n524 , n525 , n526 ;
  assign n12 = ~x1 & x4 ;
  assign n13 = ~x4 & ~x8 ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = x0 & ~n14 ;
  assign n16 = x1 & x4 ;
  assign n17 = ~x0 & n16 ;
  assign n18 = ~n15 & ~n17 ;
  assign n19 = ~x6 & ~n18 ;
  assign n20 = ~x7 & n19 ;
  assign n21 = x4 & x8 ;
  assign n22 = ~n20 & ~n21 ;
  assign n23 = ~x5 & ~n22 ;
  assign n24 = ~x4 & x7 ;
  assign n25 = x1 & ~x2 ;
  assign n26 = x5 & ~x7 ;
  assign n27 = n25 & n26 ;
  assign n28 = ~n24 & ~n27 ;
  assign n29 = x3 & ~n28 ;
  assign n30 = x4 & x7 ;
  assign n31 = ~x3 & n30 ;
  assign n32 = ~n29 & ~n31 ;
  assign n33 = ~x8 & ~n32 ;
  assign n34 = x5 & x8 ;
  assign n35 = ~x4 & n34 ;
  assign n36 = ~n33 & ~n35 ;
  assign n37 = ~n23 & n36 ;
  assign n38 = ~x9 & ~n37 ;
  assign n39 = x4 & ~x8 ;
  assign n40 = ~x3 & n39 ;
  assign n41 = ~x4 & ~x7 ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = ~x2 & ~n42 ;
  assign n44 = x1 & n43 ;
  assign n45 = ~x1 & x2 ;
  assign n46 = ~x7 & ~x8 ;
  assign n47 = n45 & n46 ;
  assign n48 = ~x9 & ~n47 ;
  assign n49 = ~n44 & n48 ;
  assign n50 = ~x6 & ~n49 ;
  assign n51 = x5 & n50 ;
  assign n52 = x6 & x9 ;
  assign n53 = ~x5 & n52 ;
  assign n54 = ~n51 & ~n53 ;
  assign n55 = ~n38 & n54 ;
  assign n56 = ~x10 & ~n55 ;
  assign n57 = ~x2 & x3 ;
  assign n58 = x2 & ~x3 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = ~x9 & ~n59 ;
  assign n61 = ~x8 & n60 ;
  assign n62 = ~x10 & ~n61 ;
  assign n63 = ~x7 & ~n62 ;
  assign n64 = x9 & x10 ;
  assign n65 = x8 & n64 ;
  assign n66 = ~n63 & ~n65 ;
  assign n67 = x6 & ~n66 ;
  assign n68 = ~x6 & x10 ;
  assign n69 = x7 & n68 ;
  assign n70 = ~n67 & ~n69 ;
  assign n71 = ~n56 & n70 ;
  assign n124 = ~n71 & x11 ;
  assign n72 = x1 & ~x4 ;
  assign n73 = ~n21 & ~n72 ;
  assign n74 = ~x0 & ~n73 ;
  assign n75 = ~x1 & ~x4 ;
  assign n76 = x0 & n75 ;
  assign n77 = ~n74 & ~n76 ;
  assign n78 = x6 & ~n77 ;
  assign n79 = x7 & n78 ;
  assign n80 = ~n13 & ~n79 ;
  assign n81 = x5 & ~n80 ;
  assign n82 = x4 & ~x7 ;
  assign n83 = ~x5 & x7 ;
  assign n84 = n45 & n83 ;
  assign n85 = ~n82 & ~n84 ;
  assign n86 = ~x3 & ~n85 ;
  assign n87 = x3 & n41 ;
  assign n88 = ~n86 & ~n87 ;
  assign n89 = x8 & ~n88 ;
  assign n90 = ~x5 & ~x8 ;
  assign n91 = x4 & n90 ;
  assign n92 = ~n89 & ~n91 ;
  assign n93 = ~n81 & n92 ;
  assign n94 = x9 & ~n93 ;
  assign n95 = ~x4 & x8 ;
  assign n96 = x3 & n95 ;
  assign n97 = ~n30 & ~n96 ;
  assign n98 = x2 & ~n97 ;
  assign n99 = ~x1 & n98 ;
  assign n100 = x7 & x8 ;
  assign n101 = n25 & n100 ;
  assign n102 = x9 & ~n101 ;
  assign n103 = ~n99 & n102 ;
  assign n104 = x6 & ~n103 ;
  assign n105 = ~x5 & n104 ;
  assign n106 = ~x6 & ~x9 ;
  assign n107 = x5 & n106 ;
  assign n108 = ~n105 & ~n107 ;
  assign n109 = ~n94 & n108 ;
  assign n110 = x10 & ~n109 ;
  assign n111 = x9 & ~n59 ;
  assign n112 = x8 & n111 ;
  assign n113 = x10 & ~n112 ;
  assign n114 = x7 & ~n113 ;
  assign n115 = ~x9 & ~x10 ;
  assign n116 = ~x8 & n115 ;
  assign n117 = ~n114 & ~n116 ;
  assign n118 = ~x6 & ~n117 ;
  assign n119 = x6 & ~x10 ;
  assign n120 = ~x7 & n119 ;
  assign n121 = ~n118 & ~n120 ;
  assign n122 = ~n110 & n121 ;
  assign n125 = n122 & ~x11 ;
  assign n126 = ~n124 & ~n125 ;
  assign n127 = ~x4 & ~x9 ;
  assign n128 = ~x2 & ~x7 ;
  assign n129 = ~n127 & ~n128 ;
  assign n130 = ~x1 & ~n129 ;
  assign n131 = x1 & x2 ;
  assign n132 = x0 & n131 ;
  assign n133 = ~x0 & ~x2 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = ~x7 & ~n134 ;
  assign n136 = x4 & n135 ;
  assign n137 = x8 & ~x9 ;
  assign n138 = ~n136 & ~n137 ;
  assign n139 = ~n130 & n138 ;
  assign n140 = ~x6 & ~n139 ;
  assign n141 = x3 & x4 ;
  assign n142 = x7 & ~n141 ;
  assign n143 = ~x9 & n142 ;
  assign n144 = ~x8 & n143 ;
  assign n145 = ~x7 & x9 ;
  assign n146 = ~n144 & ~n145 ;
  assign n147 = ~n140 & n146 ;
  assign n148 = ~x5 & ~n147 ;
  assign n149 = ~x8 & ~x9 ;
  assign n150 = x4 & n149 ;
  assign n151 = ~x6 & ~x7 ;
  assign n152 = ~x4 & n151 ;
  assign n153 = ~n150 & ~n152 ;
  assign n154 = x2 & ~n153 ;
  assign n155 = x1 & n154 ;
  assign n156 = x7 & ~x9 ;
  assign n157 = n39 & n156 ;
  assign n158 = ~n155 & ~n157 ;
  assign n159 = x3 & ~n158 ;
  assign n160 = x4 & n137 ;
  assign n161 = x7 & x9 ;
  assign n162 = ~n160 & ~n161 ;
  assign n163 = x6 & ~n162 ;
  assign n164 = ~n159 & ~n163 ;
  assign n165 = x5 & ~n164 ;
  assign n166 = ~x4 & n137 ;
  assign n167 = ~n145 & ~n166 ;
  assign n168 = ~x6 & ~n167 ;
  assign n169 = ~n165 & ~n168 ;
  assign n170 = ~n148 & n169 ;
  assign n171 = ~x10 & ~n170 ;
  assign n172 = x6 & ~x9 ;
  assign n173 = ~x4 & n172 ;
  assign n174 = x5 & ~x6 ;
  assign n175 = ~x3 & n174 ;
  assign n176 = ~n173 & ~n175 ;
  assign n177 = ~x2 & ~n176 ;
  assign n178 = ~x1 & n174 ;
  assign n179 = ~n173 & ~n178 ;
  assign n180 = ~x3 & ~n179 ;
  assign n181 = x2 & x3 ;
  assign n182 = x4 & n172 ;
  assign n183 = n181 & n182 ;
  assign n184 = ~x10 & ~n183 ;
  assign n185 = ~n180 & n184 ;
  assign n186 = ~n177 & n185 ;
  assign n187 = ~x7 & ~n186 ;
  assign n188 = ~n68 & ~n187 ;
  assign n189 = ~x8 & ~n188 ;
  assign n190 = x6 & x10 ;
  assign n191 = x7 & n190 ;
  assign n192 = n137 & n191 ;
  assign n193 = ~n189 & ~n192 ;
  assign n194 = ~n171 & n193 ;
  assign n262 = n194 & x12 ;
  assign n195 = x4 & x9 ;
  assign n196 = x2 & x7 ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = x1 & ~n197 ;
  assign n199 = ~x1 & ~x2 ;
  assign n200 = ~x0 & n199 ;
  assign n201 = x0 & x2 ;
  assign n202 = ~n200 & ~n201 ;
  assign n203 = x7 & ~n202 ;
  assign n204 = ~x4 & n203 ;
  assign n205 = ~x8 & x9 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = ~n198 & n206 ;
  assign n208 = x6 & ~n207 ;
  assign n209 = ~x3 & ~x4 ;
  assign n210 = ~x7 & ~n209 ;
  assign n211 = x9 & n210 ;
  assign n212 = x8 & n211 ;
  assign n213 = ~n156 & ~n212 ;
  assign n214 = ~n208 & n213 ;
  assign n215 = x5 & ~n214 ;
  assign n216 = x8 & x9 ;
  assign n217 = ~x4 & n216 ;
  assign n218 = x6 & x7 ;
  assign n219 = x4 & n218 ;
  assign n220 = ~n217 & ~n219 ;
  assign n221 = ~x2 & ~n220 ;
  assign n222 = ~x1 & n221 ;
  assign n223 = n95 & n145 ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = ~x3 & ~n224 ;
  assign n226 = ~x4 & n205 ;
  assign n227 = ~x7 & ~x9 ;
  assign n228 = ~n226 & ~n227 ;
  assign n229 = ~x6 & ~n228 ;
  assign n230 = ~n225 & ~n229 ;
  assign n231 = ~x5 & ~n230 ;
  assign n232 = x4 & n205 ;
  assign n233 = ~n156 & ~n232 ;
  assign n234 = x6 & ~n233 ;
  assign n235 = ~n231 & ~n234 ;
  assign n236 = ~n215 & n235 ;
  assign n237 = x10 & ~n236 ;
  assign n238 = ~x6 & x9 ;
  assign n239 = x4 & n238 ;
  assign n240 = ~x5 & x6 ;
  assign n241 = x3 & n240 ;
  assign n242 = ~n239 & ~n241 ;
  assign n243 = x2 & ~n242 ;
  assign n244 = x1 & n240 ;
  assign n245 = ~n239 & ~n244 ;
  assign n246 = x3 & ~n245 ;
  assign n247 = ~x2 & ~x3 ;
  assign n248 = ~x4 & n238 ;
  assign n249 = n247 & n248 ;
  assign n250 = x10 & ~n249 ;
  assign n251 = ~n246 & n250 ;
  assign n252 = ~n243 & n251 ;
  assign n253 = x7 & ~n252 ;
  assign n254 = ~n119 & ~n253 ;
  assign n255 = x8 & ~n254 ;
  assign n256 = ~x6 & ~x10 ;
  assign n257 = ~x7 & n256 ;
  assign n258 = n205 & n257 ;
  assign n259 = ~n255 & ~n258 ;
  assign n260 = ~n237 & n259 ;
  assign n263 = ~n260 & ~x12 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = x4 & ~x6 ;
  assign n266 = x0 & ~x3 ;
  assign n267 = n265 & n266 ;
  assign n268 = ~x4 & x5 ;
  assign n269 = x3 & n268 ;
  assign n270 = ~n267 & ~n269 ;
  assign n271 = x1 & ~n270 ;
  assign n272 = ~x4 & ~x6 ;
  assign n273 = x0 & x1 ;
  assign n274 = x4 & ~n273 ;
  assign n275 = x3 & n274 ;
  assign n276 = ~n272 & ~n275 ;
  assign n277 = ~x5 & ~n276 ;
  assign n278 = ~n271 & ~n277 ;
  assign n279 = x2 & ~n278 ;
  assign n280 = x3 & ~x6 ;
  assign n281 = ~x2 & n280 ;
  assign n282 = ~x3 & x5 ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = x4 & ~n283 ;
  assign n285 = ~n279 & ~n284 ;
  assign n286 = ~x7 & ~n285 ;
  assign n287 = x2 & n240 ;
  assign n288 = ~n178 & ~n287 ;
  assign n289 = x4 & ~n288 ;
  assign n290 = x3 & n289 ;
  assign n291 = x5 & ~n141 ;
  assign n292 = x6 & n291 ;
  assign n293 = ~n290 & ~n292 ;
  assign n294 = ~n286 & n293 ;
  assign n295 = ~x8 & ~n294 ;
  assign n296 = ~x6 & x7 ;
  assign n297 = x3 & n296 ;
  assign n298 = x6 & ~x7 ;
  assign n299 = ~x2 & n298 ;
  assign n300 = ~n297 & ~n299 ;
  assign n301 = x5 & ~n300 ;
  assign n302 = x4 & n301 ;
  assign n303 = x4 & x5 ;
  assign n304 = x7 & ~n303 ;
  assign n305 = x6 & n304 ;
  assign n306 = ~n302 & ~n305 ;
  assign n307 = ~n295 & n306 ;
  assign n308 = ~x9 & ~n307 ;
  assign n309 = x4 & x6 ;
  assign n310 = n26 & n309 ;
  assign n311 = ~n296 & ~n310 ;
  assign n312 = x8 & ~n311 ;
  assign n313 = ~n308 & ~n312 ;
  assign n314 = ~x10 & ~n313 ;
  assign n315 = x8 & x10 ;
  assign n316 = x5 & n205 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = x7 & ~n317 ;
  assign n319 = x6 & n318 ;
  assign n320 = x5 & x7 ;
  assign n321 = x8 & ~n320 ;
  assign n322 = ~x10 & ~n321 ;
  assign n323 = x9 & ~n322 ;
  assign n324 = ~n319 & ~n323 ;
  assign n325 = ~n314 & n324 ;
  assign n384 = ~n325 & x13 ;
  assign n326 = ~x4 & x6 ;
  assign n327 = ~x0 & x3 ;
  assign n328 = n326 & n327 ;
  assign n329 = x4 & ~x5 ;
  assign n330 = ~x3 & n329 ;
  assign n331 = ~n328 & ~n330 ;
  assign n332 = ~x1 & ~n331 ;
  assign n333 = ~x0 & ~x1 ;
  assign n334 = ~x4 & ~n333 ;
  assign n335 = ~x3 & n334 ;
  assign n336 = ~n309 & ~n335 ;
  assign n337 = x5 & ~n336 ;
  assign n338 = ~n332 & ~n337 ;
  assign n339 = ~x2 & ~n338 ;
  assign n340 = ~x3 & x6 ;
  assign n341 = x2 & n340 ;
  assign n342 = x3 & ~x5 ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = ~x4 & ~n343 ;
  assign n345 = ~n339 & ~n344 ;
  assign n346 = x7 & ~n345 ;
  assign n347 = ~x2 & n174 ;
  assign n348 = ~n244 & ~n347 ;
  assign n349 = ~x4 & ~n348 ;
  assign n350 = ~x3 & n349 ;
  assign n351 = ~x5 & ~n209 ;
  assign n352 = ~x6 & n351 ;
  assign n353 = ~n350 & ~n352 ;
  assign n354 = ~n346 & n353 ;
  assign n355 = x8 & ~n354 ;
  assign n356 = ~x3 & n298 ;
  assign n357 = x2 & n296 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = ~x5 & ~n358 ;
  assign n360 = ~x4 & n359 ;
  assign n361 = ~x4 & ~x5 ;
  assign n362 = ~x7 & ~n361 ;
  assign n363 = ~x6 & n362 ;
  assign n364 = ~n360 & ~n363 ;
  assign n365 = ~n355 & n364 ;
  assign n366 = x9 & ~n365 ;
  assign n367 = n83 & n272 ;
  assign n368 = ~n298 & ~n367 ;
  assign n369 = ~x8 & ~n368 ;
  assign n370 = ~n366 & ~n369 ;
  assign n371 = x10 & ~n370 ;
  assign n372 = ~x8 & ~x10 ;
  assign n373 = ~x5 & n137 ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = ~x7 & ~n374 ;
  assign n376 = ~x6 & n375 ;
  assign n377 = ~x5 & ~x7 ;
  assign n378 = ~x8 & ~n377 ;
  assign n379 = x10 & ~n378 ;
  assign n380 = ~x9 & ~n379 ;
  assign n381 = ~n376 & ~n380 ;
  assign n382 = ~n371 & n381 ;
  assign n385 = n382 & ~x13 ;
  assign n386 = ~n384 & ~n385 ;
  assign n387 = ~x2 & n218 ;
  assign n388 = x5 & n21 ;
  assign n389 = n387 & n388 ;
  assign n390 = ~x5 & n13 ;
  assign n391 = n151 & n390 ;
  assign n392 = ~n389 & ~n391 ;
  assign n393 = ~x9 & ~n392 ;
  assign n394 = ~x10 & n393 ;
  assign n395 = ~x3 & n394 ;
  assign n404 = ~n395 & x14 ;
  assign n396 = x2 & n151 ;
  assign n397 = n390 & n396 ;
  assign n398 = n218 & n388 ;
  assign n399 = ~n397 & ~n398 ;
  assign n400 = x9 & ~n399 ;
  assign n401 = x10 & n400 ;
  assign n402 = x3 & n401 ;
  assign n405 = n402 & ~x14 ;
  assign n406 = ~n404 & ~n405 ;
  assign n407 = x5 & x6 ;
  assign n408 = n82 & n407 ;
  assign n409 = ~x5 & ~x6 ;
  assign n410 = n273 & n409 ;
  assign n411 = ~n408 & ~n410 ;
  assign n412 = x3 & ~n411 ;
  assign n413 = x2 & n412 ;
  assign n414 = ~x4 & ~n298 ;
  assign n415 = ~x7 & ~n174 ;
  assign n416 = ~x3 & ~n415 ;
  assign n417 = x7 & ~n407 ;
  assign n418 = ~x6 & ~n131 ;
  assign n419 = x5 & n418 ;
  assign n420 = ~x9 & ~n419 ;
  assign n421 = ~n417 & n420 ;
  assign n422 = ~n416 & n421 ;
  assign n423 = ~n414 & n422 ;
  assign n424 = ~n413 & n423 ;
  assign n425 = ~x8 & ~n424 ;
  assign n426 = x3 & x8 ;
  assign n427 = ~n58 & ~n426 ;
  assign n428 = x6 & ~n427 ;
  assign n429 = x5 & n428 ;
  assign n430 = x7 & n429 ;
  assign n431 = ~x9 & n430 ;
  assign n432 = x4 & n431 ;
  assign n433 = x7 & n407 ;
  assign n434 = x9 & ~n433 ;
  assign n435 = ~n432 & ~n434 ;
  assign n436 = ~n425 & n435 ;
  assign n437 = ~x10 & ~n436 ;
  assign n468 = ~n437 & x15 ;
  assign n438 = n24 & n409 ;
  assign n439 = n333 & n407 ;
  assign n440 = ~n438 & ~n439 ;
  assign n441 = ~x3 & ~n440 ;
  assign n442 = ~x2 & n441 ;
  assign n443 = x4 & ~n296 ;
  assign n444 = x7 & ~n240 ;
  assign n445 = x3 & ~n444 ;
  assign n446 = ~x7 & ~n409 ;
  assign n447 = x6 & ~n199 ;
  assign n448 = ~x5 & n447 ;
  assign n449 = x9 & ~n448 ;
  assign n450 = ~n446 & n449 ;
  assign n451 = ~n445 & n450 ;
  assign n452 = ~n443 & n451 ;
  assign n453 = ~n442 & n452 ;
  assign n454 = x8 & ~n453 ;
  assign n455 = ~x3 & ~x8 ;
  assign n456 = ~n57 & ~n455 ;
  assign n457 = ~x6 & ~n456 ;
  assign n458 = ~x5 & n457 ;
  assign n459 = ~x7 & n458 ;
  assign n460 = x9 & n459 ;
  assign n461 = ~x4 & n460 ;
  assign n462 = ~x7 & n409 ;
  assign n463 = ~x9 & ~n462 ;
  assign n464 = ~n461 & ~n463 ;
  assign n465 = ~n454 & n464 ;
  assign n466 = x10 & ~n465 ;
  assign n469 = n466 & ~x15 ;
  assign n470 = ~n468 & ~n469 ;
  assign n471 = x6 & x8 ;
  assign n472 = n320 & n471 ;
  assign n473 = x1 & x3 ;
  assign n474 = x0 & n473 ;
  assign n475 = ~x8 & n377 ;
  assign n476 = n474 & n475 ;
  assign n477 = ~n472 & ~n476 ;
  assign n478 = x2 & ~n477 ;
  assign n479 = x8 & n320 ;
  assign n480 = x3 & x6 ;
  assign n481 = n479 & n480 ;
  assign n482 = ~n478 & ~n481 ;
  assign n483 = x4 & ~n482 ;
  assign n484 = n181 & n309 ;
  assign n485 = x5 & ~n484 ;
  assign n486 = ~n240 & ~n485 ;
  assign n487 = ~x7 & ~n486 ;
  assign n488 = ~x8 & n487 ;
  assign n489 = n115 & ~n488 ;
  assign n490 = ~n483 & n489 ;
  assign n510 = ~n490 & x16 ;
  assign n491 = ~x6 & ~x8 ;
  assign n492 = n377 & n491 ;
  assign n493 = ~x1 & ~x3 ;
  assign n494 = ~x0 & n493 ;
  assign n495 = n479 & n494 ;
  assign n496 = ~n492 & ~n495 ;
  assign n497 = ~x2 & ~n496 ;
  assign n498 = ~x3 & ~x6 ;
  assign n499 = n475 & n498 ;
  assign n500 = ~n497 & ~n499 ;
  assign n501 = ~x4 & ~n500 ;
  assign n502 = n247 & n272 ;
  assign n503 = ~x5 & ~n502 ;
  assign n504 = ~n174 & ~n503 ;
  assign n505 = x7 & ~n504 ;
  assign n506 = x8 & n505 ;
  assign n507 = n64 & ~n506 ;
  assign n508 = ~n501 & n507 ;
  assign n511 = n508 & ~x16 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = x2 & n141 ;
  assign n514 = n407 & n513 ;
  assign n515 = ~x9 & ~n514 ;
  assign n516 = ~x10 & n515 ;
  assign n517 = n46 & n516 ;
  assign n524 = ~n517 & x17 ;
  assign n518 = ~x2 & n209 ;
  assign n519 = n409 & n518 ;
  assign n520 = x9 & ~n519 ;
  assign n521 = x10 & n520 ;
  assign n522 = n100 & n521 ;
  assign n525 = n522 & ~x17 ;
  assign n526 = ~n524 & ~n525 ;
  assign y0 = ~n126 ;
  assign y1 = ~n264 ;
  assign y2 = ~n386 ;
  assign y3 = ~n406 ;
  assign y4 = ~n470 ;
  assign y5 = ~n512 ;
  assign y6 = ~n526 ;
endmodule
