module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2426 , n2427 , n2428 ;
  assign n257 = x0 & ~x128 ;
  assign n258 = ~x0 & x128 ;
  assign n259 = ~n257 & ~n258 ;
  assign n261 = ~n259 & x256 ;
  assign n262 = n259 & ~x256 ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = x0 & x128 ;
  assign n265 = ~x1 & ~x129 ;
  assign n266 = x1 & x129 ;
  assign n267 = ~n265 & ~n266 ;
  assign n268 = n264 & ~n267 ;
  assign n269 = ~n264 & n267 ;
  assign n270 = ~n268 & ~n269 ;
  assign n276 = ~n270 & x257 ;
  assign n271 = ~x0 & ~x128 ;
  assign n272 = ~n267 & n271 ;
  assign n273 = n267 & ~n271 ;
  assign n274 = ~n272 & ~n273 ;
  assign n277 = n274 & ~x257 ;
  assign n278 = ~n276 & ~n277 ;
  assign n279 = n264 & ~n265 ;
  assign n280 = ~n266 & ~n279 ;
  assign n281 = ~x2 & ~x130 ;
  assign n282 = x2 & x130 ;
  assign n283 = ~n281 & ~n282 ;
  assign n284 = n280 & ~n283 ;
  assign n285 = ~n280 & n283 ;
  assign n286 = ~n284 & ~n285 ;
  assign n293 = n286 & x258 ;
  assign n287 = ~n266 & n271 ;
  assign n288 = ~n265 & ~n287 ;
  assign n289 = ~n283 & n288 ;
  assign n290 = n283 & ~n288 ;
  assign n291 = ~n289 & ~n290 ;
  assign n294 = ~n291 & ~x258 ;
  assign n295 = ~n293 & ~n294 ;
  assign n296 = ~n280 & ~n281 ;
  assign n297 = ~n282 & ~n296 ;
  assign n298 = ~x3 & ~x131 ;
  assign n299 = x3 & x131 ;
  assign n300 = ~n298 & ~n299 ;
  assign n301 = n297 & ~n300 ;
  assign n302 = ~n297 & n300 ;
  assign n303 = ~n301 & ~n302 ;
  assign n310 = n303 & x259 ;
  assign n304 = ~n282 & ~n288 ;
  assign n305 = ~n281 & ~n304 ;
  assign n306 = ~n300 & n305 ;
  assign n307 = n300 & ~n305 ;
  assign n308 = ~n306 & ~n307 ;
  assign n311 = ~n308 & ~x259 ;
  assign n312 = ~n310 & ~n311 ;
  assign n313 = ~n297 & ~n298 ;
  assign n314 = ~n299 & ~n313 ;
  assign n315 = ~x4 & ~x132 ;
  assign n316 = x4 & x132 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = n314 & ~n317 ;
  assign n319 = ~n314 & n317 ;
  assign n320 = ~n318 & ~n319 ;
  assign n327 = n320 & x260 ;
  assign n321 = ~n299 & ~n305 ;
  assign n322 = ~n298 & ~n321 ;
  assign n323 = ~n317 & n322 ;
  assign n324 = n317 & ~n322 ;
  assign n325 = ~n323 & ~n324 ;
  assign n328 = ~n325 & ~x260 ;
  assign n329 = ~n327 & ~n328 ;
  assign n330 = ~n314 & ~n315 ;
  assign n331 = ~n316 & ~n330 ;
  assign n332 = ~x5 & ~x133 ;
  assign n333 = x5 & x133 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = n331 & ~n334 ;
  assign n336 = ~n331 & n334 ;
  assign n337 = ~n335 & ~n336 ;
  assign n344 = n337 & x261 ;
  assign n338 = ~n316 & ~n322 ;
  assign n339 = ~n315 & ~n338 ;
  assign n340 = ~n334 & n339 ;
  assign n341 = n334 & ~n339 ;
  assign n342 = ~n340 & ~n341 ;
  assign n345 = ~n342 & ~x261 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = ~n331 & ~n332 ;
  assign n348 = ~n333 & ~n347 ;
  assign n349 = ~x6 & ~x134 ;
  assign n350 = x6 & x134 ;
  assign n351 = ~n349 & ~n350 ;
  assign n352 = n348 & ~n351 ;
  assign n353 = ~n348 & n351 ;
  assign n354 = ~n352 & ~n353 ;
  assign n361 = n354 & x262 ;
  assign n355 = ~n333 & ~n339 ;
  assign n356 = ~n332 & ~n355 ;
  assign n357 = ~n351 & n356 ;
  assign n358 = n351 & ~n356 ;
  assign n359 = ~n357 & ~n358 ;
  assign n362 = ~n359 & ~x262 ;
  assign n363 = ~n361 & ~n362 ;
  assign n364 = ~n348 & ~n349 ;
  assign n365 = ~n350 & ~n364 ;
  assign n366 = ~x7 & ~x135 ;
  assign n367 = x7 & x135 ;
  assign n368 = ~n366 & ~n367 ;
  assign n369 = n365 & ~n368 ;
  assign n370 = ~n365 & n368 ;
  assign n371 = ~n369 & ~n370 ;
  assign n378 = n371 & x263 ;
  assign n372 = ~n350 & ~n356 ;
  assign n373 = ~n349 & ~n372 ;
  assign n374 = ~n368 & n373 ;
  assign n375 = n368 & ~n373 ;
  assign n376 = ~n374 & ~n375 ;
  assign n379 = ~n376 & ~x263 ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = ~n365 & ~n366 ;
  assign n382 = ~n367 & ~n381 ;
  assign n383 = ~x8 & ~x136 ;
  assign n384 = x8 & x136 ;
  assign n385 = ~n383 & ~n384 ;
  assign n386 = n382 & ~n385 ;
  assign n387 = ~n382 & n385 ;
  assign n388 = ~n386 & ~n387 ;
  assign n395 = n388 & x264 ;
  assign n389 = ~n367 & ~n373 ;
  assign n390 = ~n366 & ~n389 ;
  assign n391 = ~n385 & n390 ;
  assign n392 = n385 & ~n390 ;
  assign n393 = ~n391 & ~n392 ;
  assign n396 = ~n393 & ~x264 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = ~n382 & ~n383 ;
  assign n399 = ~n384 & ~n398 ;
  assign n400 = ~x9 & ~x137 ;
  assign n401 = x9 & x137 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = n399 & ~n402 ;
  assign n404 = ~n399 & n402 ;
  assign n405 = ~n403 & ~n404 ;
  assign n412 = n405 & x265 ;
  assign n406 = ~n384 & ~n390 ;
  assign n407 = ~n383 & ~n406 ;
  assign n408 = ~n402 & n407 ;
  assign n409 = n402 & ~n407 ;
  assign n410 = ~n408 & ~n409 ;
  assign n413 = ~n410 & ~x265 ;
  assign n414 = ~n412 & ~n413 ;
  assign n415 = ~n399 & ~n400 ;
  assign n416 = ~n401 & ~n415 ;
  assign n417 = ~x10 & ~x138 ;
  assign n418 = x10 & x138 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = n416 & ~n419 ;
  assign n421 = ~n416 & n419 ;
  assign n422 = ~n420 & ~n421 ;
  assign n429 = n422 & x266 ;
  assign n423 = ~n401 & ~n407 ;
  assign n424 = ~n400 & ~n423 ;
  assign n425 = ~n419 & n424 ;
  assign n426 = n419 & ~n424 ;
  assign n427 = ~n425 & ~n426 ;
  assign n430 = ~n427 & ~x266 ;
  assign n431 = ~n429 & ~n430 ;
  assign n432 = ~n416 & ~n417 ;
  assign n433 = ~n418 & ~n432 ;
  assign n434 = ~x11 & ~x139 ;
  assign n435 = x11 & x139 ;
  assign n436 = ~n434 & ~n435 ;
  assign n437 = n433 & ~n436 ;
  assign n438 = ~n433 & n436 ;
  assign n439 = ~n437 & ~n438 ;
  assign n446 = n439 & x267 ;
  assign n440 = ~n418 & ~n424 ;
  assign n441 = ~n417 & ~n440 ;
  assign n442 = ~n436 & n441 ;
  assign n443 = n436 & ~n441 ;
  assign n444 = ~n442 & ~n443 ;
  assign n447 = ~n444 & ~x267 ;
  assign n448 = ~n446 & ~n447 ;
  assign n449 = ~n433 & ~n434 ;
  assign n450 = ~n435 & ~n449 ;
  assign n451 = ~x12 & ~x140 ;
  assign n452 = x12 & x140 ;
  assign n453 = ~n451 & ~n452 ;
  assign n454 = n450 & ~n453 ;
  assign n455 = ~n450 & n453 ;
  assign n456 = ~n454 & ~n455 ;
  assign n463 = n456 & x268 ;
  assign n457 = ~n435 & ~n441 ;
  assign n458 = ~n434 & ~n457 ;
  assign n459 = ~n453 & n458 ;
  assign n460 = n453 & ~n458 ;
  assign n461 = ~n459 & ~n460 ;
  assign n464 = ~n461 & ~x268 ;
  assign n465 = ~n463 & ~n464 ;
  assign n466 = ~n450 & ~n451 ;
  assign n467 = ~n452 & ~n466 ;
  assign n468 = ~x13 & ~x141 ;
  assign n469 = x13 & x141 ;
  assign n470 = ~n468 & ~n469 ;
  assign n471 = n467 & ~n470 ;
  assign n472 = ~n467 & n470 ;
  assign n473 = ~n471 & ~n472 ;
  assign n480 = n473 & x269 ;
  assign n474 = ~n452 & ~n458 ;
  assign n475 = ~n451 & ~n474 ;
  assign n476 = ~n470 & n475 ;
  assign n477 = n470 & ~n475 ;
  assign n478 = ~n476 & ~n477 ;
  assign n481 = ~n478 & ~x269 ;
  assign n482 = ~n480 & ~n481 ;
  assign n483 = ~n467 & ~n468 ;
  assign n484 = ~n469 & ~n483 ;
  assign n485 = ~x14 & ~x142 ;
  assign n486 = x14 & x142 ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = n484 & ~n487 ;
  assign n489 = ~n484 & n487 ;
  assign n490 = ~n488 & ~n489 ;
  assign n497 = n490 & x270 ;
  assign n491 = ~n469 & ~n475 ;
  assign n492 = ~n468 & ~n491 ;
  assign n493 = ~n487 & n492 ;
  assign n494 = n487 & ~n492 ;
  assign n495 = ~n493 & ~n494 ;
  assign n498 = ~n495 & ~x270 ;
  assign n499 = ~n497 & ~n498 ;
  assign n500 = ~n484 & ~n485 ;
  assign n501 = ~n486 & ~n500 ;
  assign n502 = ~x15 & ~x143 ;
  assign n503 = x15 & x143 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = n501 & ~n504 ;
  assign n506 = ~n501 & n504 ;
  assign n507 = ~n505 & ~n506 ;
  assign n514 = n507 & x271 ;
  assign n508 = ~n486 & ~n492 ;
  assign n509 = ~n485 & ~n508 ;
  assign n510 = ~n504 & n509 ;
  assign n511 = n504 & ~n509 ;
  assign n512 = ~n510 & ~n511 ;
  assign n515 = ~n512 & ~x271 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = ~n501 & ~n502 ;
  assign n518 = ~n503 & ~n517 ;
  assign n519 = ~x16 & ~x144 ;
  assign n520 = x16 & x144 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = n518 & ~n521 ;
  assign n523 = ~n518 & n521 ;
  assign n524 = ~n522 & ~n523 ;
  assign n531 = n524 & x272 ;
  assign n525 = ~n503 & ~n509 ;
  assign n526 = ~n502 & ~n525 ;
  assign n527 = ~n521 & n526 ;
  assign n528 = n521 & ~n526 ;
  assign n529 = ~n527 & ~n528 ;
  assign n532 = ~n529 & ~x272 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~n518 & ~n519 ;
  assign n535 = ~n520 & ~n534 ;
  assign n536 = ~x17 & ~x145 ;
  assign n537 = x17 & x145 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = n535 & ~n538 ;
  assign n540 = ~n535 & n538 ;
  assign n541 = ~n539 & ~n540 ;
  assign n548 = n541 & x273 ;
  assign n542 = ~n520 & ~n526 ;
  assign n543 = ~n519 & ~n542 ;
  assign n544 = ~n538 & n543 ;
  assign n545 = n538 & ~n543 ;
  assign n546 = ~n544 & ~n545 ;
  assign n549 = ~n546 & ~x273 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = ~n535 & ~n536 ;
  assign n552 = ~n537 & ~n551 ;
  assign n553 = ~x18 & ~x146 ;
  assign n554 = x18 & x146 ;
  assign n555 = ~n553 & ~n554 ;
  assign n556 = n552 & ~n555 ;
  assign n557 = ~n552 & n555 ;
  assign n558 = ~n556 & ~n557 ;
  assign n565 = n558 & x274 ;
  assign n559 = ~n537 & ~n543 ;
  assign n560 = ~n536 & ~n559 ;
  assign n561 = ~n555 & n560 ;
  assign n562 = n555 & ~n560 ;
  assign n563 = ~n561 & ~n562 ;
  assign n566 = ~n563 & ~x274 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = ~n552 & ~n553 ;
  assign n569 = ~n554 & ~n568 ;
  assign n570 = ~x19 & ~x147 ;
  assign n571 = x19 & x147 ;
  assign n572 = ~n570 & ~n571 ;
  assign n573 = n569 & ~n572 ;
  assign n574 = ~n569 & n572 ;
  assign n575 = ~n573 & ~n574 ;
  assign n582 = n575 & x275 ;
  assign n576 = ~n554 & ~n560 ;
  assign n577 = ~n553 & ~n576 ;
  assign n578 = ~n572 & n577 ;
  assign n579 = n572 & ~n577 ;
  assign n580 = ~n578 & ~n579 ;
  assign n583 = ~n580 & ~x275 ;
  assign n584 = ~n582 & ~n583 ;
  assign n585 = ~n569 & ~n570 ;
  assign n586 = ~n571 & ~n585 ;
  assign n587 = ~x20 & ~x148 ;
  assign n588 = x20 & x148 ;
  assign n589 = ~n587 & ~n588 ;
  assign n590 = n586 & ~n589 ;
  assign n591 = ~n586 & n589 ;
  assign n592 = ~n590 & ~n591 ;
  assign n599 = n592 & x276 ;
  assign n593 = ~n571 & ~n577 ;
  assign n594 = ~n570 & ~n593 ;
  assign n595 = ~n589 & n594 ;
  assign n596 = n589 & ~n594 ;
  assign n597 = ~n595 & ~n596 ;
  assign n600 = ~n597 & ~x276 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = ~n586 & ~n587 ;
  assign n603 = ~n588 & ~n602 ;
  assign n604 = ~x21 & ~x149 ;
  assign n605 = x21 & x149 ;
  assign n606 = ~n604 & ~n605 ;
  assign n607 = n603 & ~n606 ;
  assign n608 = ~n603 & n606 ;
  assign n609 = ~n607 & ~n608 ;
  assign n616 = n609 & x277 ;
  assign n610 = ~n588 & ~n594 ;
  assign n611 = ~n587 & ~n610 ;
  assign n612 = ~n606 & n611 ;
  assign n613 = n606 & ~n611 ;
  assign n614 = ~n612 & ~n613 ;
  assign n617 = ~n614 & ~x277 ;
  assign n618 = ~n616 & ~n617 ;
  assign n619 = ~n603 & ~n604 ;
  assign n620 = ~n605 & ~n619 ;
  assign n621 = ~x22 & ~x150 ;
  assign n622 = x22 & x150 ;
  assign n623 = ~n621 & ~n622 ;
  assign n624 = n620 & ~n623 ;
  assign n625 = ~n620 & n623 ;
  assign n626 = ~n624 & ~n625 ;
  assign n633 = n626 & x278 ;
  assign n627 = ~n605 & ~n611 ;
  assign n628 = ~n604 & ~n627 ;
  assign n629 = ~n623 & n628 ;
  assign n630 = n623 & ~n628 ;
  assign n631 = ~n629 & ~n630 ;
  assign n634 = ~n631 & ~x278 ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = ~n620 & ~n621 ;
  assign n637 = ~n622 & ~n636 ;
  assign n638 = ~x23 & ~x151 ;
  assign n639 = x23 & x151 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = n637 & ~n640 ;
  assign n642 = ~n637 & n640 ;
  assign n643 = ~n641 & ~n642 ;
  assign n650 = n643 & x279 ;
  assign n644 = ~n622 & ~n628 ;
  assign n645 = ~n621 & ~n644 ;
  assign n646 = ~n640 & n645 ;
  assign n647 = n640 & ~n645 ;
  assign n648 = ~n646 & ~n647 ;
  assign n651 = ~n648 & ~x279 ;
  assign n652 = ~n650 & ~n651 ;
  assign n653 = ~n637 & ~n638 ;
  assign n654 = ~n639 & ~n653 ;
  assign n655 = ~x24 & ~x152 ;
  assign n656 = x24 & x152 ;
  assign n657 = ~n655 & ~n656 ;
  assign n658 = n654 & ~n657 ;
  assign n659 = ~n654 & n657 ;
  assign n660 = ~n658 & ~n659 ;
  assign n667 = n660 & x280 ;
  assign n661 = ~n639 & ~n645 ;
  assign n662 = ~n638 & ~n661 ;
  assign n663 = ~n657 & n662 ;
  assign n664 = n657 & ~n662 ;
  assign n665 = ~n663 & ~n664 ;
  assign n668 = ~n665 & ~x280 ;
  assign n669 = ~n667 & ~n668 ;
  assign n670 = ~n654 & ~n655 ;
  assign n671 = ~n656 & ~n670 ;
  assign n672 = ~x25 & ~x153 ;
  assign n673 = x25 & x153 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = n671 & ~n674 ;
  assign n676 = ~n671 & n674 ;
  assign n677 = ~n675 & ~n676 ;
  assign n684 = n677 & x281 ;
  assign n678 = ~n656 & ~n662 ;
  assign n679 = ~n655 & ~n678 ;
  assign n680 = ~n674 & n679 ;
  assign n681 = n674 & ~n679 ;
  assign n682 = ~n680 & ~n681 ;
  assign n685 = ~n682 & ~x281 ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = ~n671 & ~n672 ;
  assign n688 = ~n673 & ~n687 ;
  assign n689 = ~x26 & ~x154 ;
  assign n690 = x26 & x154 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = n688 & ~n691 ;
  assign n693 = ~n688 & n691 ;
  assign n694 = ~n692 & ~n693 ;
  assign n701 = n694 & x282 ;
  assign n695 = ~n673 & ~n679 ;
  assign n696 = ~n672 & ~n695 ;
  assign n697 = ~n691 & n696 ;
  assign n698 = n691 & ~n696 ;
  assign n699 = ~n697 & ~n698 ;
  assign n702 = ~n699 & ~x282 ;
  assign n703 = ~n701 & ~n702 ;
  assign n704 = ~n688 & ~n689 ;
  assign n705 = ~n690 & ~n704 ;
  assign n706 = ~x27 & ~x155 ;
  assign n707 = x27 & x155 ;
  assign n708 = ~n706 & ~n707 ;
  assign n709 = n705 & ~n708 ;
  assign n710 = ~n705 & n708 ;
  assign n711 = ~n709 & ~n710 ;
  assign n718 = n711 & x283 ;
  assign n712 = ~n690 & ~n696 ;
  assign n713 = ~n689 & ~n712 ;
  assign n714 = ~n708 & n713 ;
  assign n715 = n708 & ~n713 ;
  assign n716 = ~n714 & ~n715 ;
  assign n719 = ~n716 & ~x283 ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = ~n705 & ~n706 ;
  assign n722 = ~n707 & ~n721 ;
  assign n723 = ~x28 & ~x156 ;
  assign n724 = x28 & x156 ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = n722 & ~n725 ;
  assign n727 = ~n722 & n725 ;
  assign n728 = ~n726 & ~n727 ;
  assign n735 = n728 & x284 ;
  assign n729 = ~n707 & ~n713 ;
  assign n730 = ~n706 & ~n729 ;
  assign n731 = ~n725 & n730 ;
  assign n732 = n725 & ~n730 ;
  assign n733 = ~n731 & ~n732 ;
  assign n736 = ~n733 & ~x284 ;
  assign n737 = ~n735 & ~n736 ;
  assign n738 = ~n722 & ~n723 ;
  assign n739 = ~n724 & ~n738 ;
  assign n740 = ~x29 & ~x157 ;
  assign n741 = x29 & x157 ;
  assign n742 = ~n740 & ~n741 ;
  assign n743 = n739 & ~n742 ;
  assign n744 = ~n739 & n742 ;
  assign n745 = ~n743 & ~n744 ;
  assign n752 = n745 & x285 ;
  assign n746 = ~n724 & ~n730 ;
  assign n747 = ~n723 & ~n746 ;
  assign n748 = ~n742 & n747 ;
  assign n749 = n742 & ~n747 ;
  assign n750 = ~n748 & ~n749 ;
  assign n753 = ~n750 & ~x285 ;
  assign n754 = ~n752 & ~n753 ;
  assign n755 = ~n739 & ~n740 ;
  assign n756 = ~n741 & ~n755 ;
  assign n757 = ~x30 & ~x158 ;
  assign n758 = x30 & x158 ;
  assign n759 = ~n757 & ~n758 ;
  assign n760 = n756 & ~n759 ;
  assign n761 = ~n756 & n759 ;
  assign n762 = ~n760 & ~n761 ;
  assign n769 = n762 & x286 ;
  assign n763 = ~n741 & ~n747 ;
  assign n764 = ~n740 & ~n763 ;
  assign n765 = ~n759 & n764 ;
  assign n766 = n759 & ~n764 ;
  assign n767 = ~n765 & ~n766 ;
  assign n770 = ~n767 & ~x286 ;
  assign n771 = ~n769 & ~n770 ;
  assign n772 = ~n756 & ~n757 ;
  assign n773 = ~n758 & ~n772 ;
  assign n774 = ~x31 & ~x159 ;
  assign n775 = x31 & x159 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = n773 & ~n776 ;
  assign n778 = ~n773 & n776 ;
  assign n779 = ~n777 & ~n778 ;
  assign n786 = n779 & x287 ;
  assign n780 = ~n758 & ~n764 ;
  assign n781 = ~n757 & ~n780 ;
  assign n782 = ~n776 & n781 ;
  assign n783 = n776 & ~n781 ;
  assign n784 = ~n782 & ~n783 ;
  assign n787 = ~n784 & ~x287 ;
  assign n788 = ~n786 & ~n787 ;
  assign n789 = ~n773 & ~n774 ;
  assign n790 = ~n775 & ~n789 ;
  assign n791 = ~x32 & ~x160 ;
  assign n792 = x32 & x160 ;
  assign n793 = ~n791 & ~n792 ;
  assign n794 = n790 & ~n793 ;
  assign n795 = ~n790 & n793 ;
  assign n796 = ~n794 & ~n795 ;
  assign n803 = n796 & x288 ;
  assign n797 = ~n775 & ~n781 ;
  assign n798 = ~n774 & ~n797 ;
  assign n799 = ~n793 & n798 ;
  assign n800 = n793 & ~n798 ;
  assign n801 = ~n799 & ~n800 ;
  assign n804 = ~n801 & ~x288 ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = ~n790 & ~n791 ;
  assign n807 = ~n792 & ~n806 ;
  assign n808 = ~x33 & ~x161 ;
  assign n809 = x33 & x161 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = n807 & ~n810 ;
  assign n812 = ~n807 & n810 ;
  assign n813 = ~n811 & ~n812 ;
  assign n820 = n813 & x289 ;
  assign n814 = ~n792 & ~n798 ;
  assign n815 = ~n791 & ~n814 ;
  assign n816 = ~n810 & n815 ;
  assign n817 = n810 & ~n815 ;
  assign n818 = ~n816 & ~n817 ;
  assign n821 = ~n818 & ~x289 ;
  assign n822 = ~n820 & ~n821 ;
  assign n823 = ~n807 & ~n808 ;
  assign n824 = ~n809 & ~n823 ;
  assign n825 = ~x34 & ~x162 ;
  assign n826 = x34 & x162 ;
  assign n827 = ~n825 & ~n826 ;
  assign n828 = n824 & ~n827 ;
  assign n829 = ~n824 & n827 ;
  assign n830 = ~n828 & ~n829 ;
  assign n837 = n830 & x290 ;
  assign n831 = ~n809 & ~n815 ;
  assign n832 = ~n808 & ~n831 ;
  assign n833 = ~n827 & n832 ;
  assign n834 = n827 & ~n832 ;
  assign n835 = ~n833 & ~n834 ;
  assign n838 = ~n835 & ~x290 ;
  assign n839 = ~n837 & ~n838 ;
  assign n840 = ~n824 & ~n825 ;
  assign n841 = ~n826 & ~n840 ;
  assign n842 = ~x35 & ~x163 ;
  assign n843 = x35 & x163 ;
  assign n844 = ~n842 & ~n843 ;
  assign n845 = n841 & ~n844 ;
  assign n846 = ~n841 & n844 ;
  assign n847 = ~n845 & ~n846 ;
  assign n854 = n847 & x291 ;
  assign n848 = ~n826 & ~n832 ;
  assign n849 = ~n825 & ~n848 ;
  assign n850 = ~n844 & n849 ;
  assign n851 = n844 & ~n849 ;
  assign n852 = ~n850 & ~n851 ;
  assign n855 = ~n852 & ~x291 ;
  assign n856 = ~n854 & ~n855 ;
  assign n857 = ~n841 & ~n842 ;
  assign n858 = ~n843 & ~n857 ;
  assign n859 = ~x36 & ~x164 ;
  assign n860 = x36 & x164 ;
  assign n861 = ~n859 & ~n860 ;
  assign n862 = n858 & ~n861 ;
  assign n863 = ~n858 & n861 ;
  assign n864 = ~n862 & ~n863 ;
  assign n871 = n864 & x292 ;
  assign n865 = ~n843 & ~n849 ;
  assign n866 = ~n842 & ~n865 ;
  assign n867 = ~n861 & n866 ;
  assign n868 = n861 & ~n866 ;
  assign n869 = ~n867 & ~n868 ;
  assign n872 = ~n869 & ~x292 ;
  assign n873 = ~n871 & ~n872 ;
  assign n874 = ~n858 & ~n859 ;
  assign n875 = ~n860 & ~n874 ;
  assign n876 = ~x37 & ~x165 ;
  assign n877 = x37 & x165 ;
  assign n878 = ~n876 & ~n877 ;
  assign n879 = n875 & ~n878 ;
  assign n880 = ~n875 & n878 ;
  assign n881 = ~n879 & ~n880 ;
  assign n888 = n881 & x293 ;
  assign n882 = ~n860 & ~n866 ;
  assign n883 = ~n859 & ~n882 ;
  assign n884 = ~n878 & n883 ;
  assign n885 = n878 & ~n883 ;
  assign n886 = ~n884 & ~n885 ;
  assign n889 = ~n886 & ~x293 ;
  assign n890 = ~n888 & ~n889 ;
  assign n891 = ~n875 & ~n876 ;
  assign n892 = ~n877 & ~n891 ;
  assign n893 = ~x38 & ~x166 ;
  assign n894 = x38 & x166 ;
  assign n895 = ~n893 & ~n894 ;
  assign n896 = n892 & ~n895 ;
  assign n897 = ~n892 & n895 ;
  assign n898 = ~n896 & ~n897 ;
  assign n905 = n898 & x294 ;
  assign n899 = ~n877 & ~n883 ;
  assign n900 = ~n876 & ~n899 ;
  assign n901 = ~n895 & n900 ;
  assign n902 = n895 & ~n900 ;
  assign n903 = ~n901 & ~n902 ;
  assign n906 = ~n903 & ~x294 ;
  assign n907 = ~n905 & ~n906 ;
  assign n908 = ~n892 & ~n893 ;
  assign n909 = ~n894 & ~n908 ;
  assign n910 = ~x39 & ~x167 ;
  assign n911 = x39 & x167 ;
  assign n912 = ~n910 & ~n911 ;
  assign n913 = n909 & ~n912 ;
  assign n914 = ~n909 & n912 ;
  assign n915 = ~n913 & ~n914 ;
  assign n922 = n915 & x295 ;
  assign n916 = ~n894 & ~n900 ;
  assign n917 = ~n893 & ~n916 ;
  assign n918 = ~n912 & n917 ;
  assign n919 = n912 & ~n917 ;
  assign n920 = ~n918 & ~n919 ;
  assign n923 = ~n920 & ~x295 ;
  assign n924 = ~n922 & ~n923 ;
  assign n925 = ~n909 & ~n910 ;
  assign n926 = ~n911 & ~n925 ;
  assign n927 = ~x40 & ~x168 ;
  assign n928 = x40 & x168 ;
  assign n929 = ~n927 & ~n928 ;
  assign n930 = n926 & ~n929 ;
  assign n931 = ~n926 & n929 ;
  assign n932 = ~n930 & ~n931 ;
  assign n939 = n932 & x296 ;
  assign n933 = ~n911 & ~n917 ;
  assign n934 = ~n910 & ~n933 ;
  assign n935 = ~n929 & n934 ;
  assign n936 = n929 & ~n934 ;
  assign n937 = ~n935 & ~n936 ;
  assign n940 = ~n937 & ~x296 ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = ~n926 & ~n927 ;
  assign n943 = ~n928 & ~n942 ;
  assign n944 = ~x41 & ~x169 ;
  assign n945 = x41 & x169 ;
  assign n946 = ~n944 & ~n945 ;
  assign n947 = n943 & ~n946 ;
  assign n948 = ~n943 & n946 ;
  assign n949 = ~n947 & ~n948 ;
  assign n956 = n949 & x297 ;
  assign n950 = ~n928 & ~n934 ;
  assign n951 = ~n927 & ~n950 ;
  assign n952 = ~n946 & n951 ;
  assign n953 = n946 & ~n951 ;
  assign n954 = ~n952 & ~n953 ;
  assign n957 = ~n954 & ~x297 ;
  assign n958 = ~n956 & ~n957 ;
  assign n959 = ~n943 & ~n944 ;
  assign n960 = ~n945 & ~n959 ;
  assign n961 = ~x42 & ~x170 ;
  assign n962 = x42 & x170 ;
  assign n963 = ~n961 & ~n962 ;
  assign n964 = n960 & ~n963 ;
  assign n965 = ~n960 & n963 ;
  assign n966 = ~n964 & ~n965 ;
  assign n973 = n966 & x298 ;
  assign n967 = ~n945 & ~n951 ;
  assign n968 = ~n944 & ~n967 ;
  assign n969 = ~n963 & n968 ;
  assign n970 = n963 & ~n968 ;
  assign n971 = ~n969 & ~n970 ;
  assign n974 = ~n971 & ~x298 ;
  assign n975 = ~n973 & ~n974 ;
  assign n976 = ~n960 & ~n961 ;
  assign n977 = ~n962 & ~n976 ;
  assign n978 = ~x43 & ~x171 ;
  assign n979 = x43 & x171 ;
  assign n980 = ~n978 & ~n979 ;
  assign n981 = n977 & ~n980 ;
  assign n982 = ~n977 & n980 ;
  assign n983 = ~n981 & ~n982 ;
  assign n990 = n983 & x299 ;
  assign n984 = ~n962 & ~n968 ;
  assign n985 = ~n961 & ~n984 ;
  assign n986 = ~n980 & n985 ;
  assign n987 = n980 & ~n985 ;
  assign n988 = ~n986 & ~n987 ;
  assign n991 = ~n988 & ~x299 ;
  assign n992 = ~n990 & ~n991 ;
  assign n993 = ~n977 & ~n978 ;
  assign n994 = ~n979 & ~n993 ;
  assign n995 = ~x44 & ~x172 ;
  assign n996 = x44 & x172 ;
  assign n997 = ~n995 & ~n996 ;
  assign n998 = n994 & ~n997 ;
  assign n999 = ~n994 & n997 ;
  assign n1000 = ~n998 & ~n999 ;
  assign n1007 = n1000 & x300 ;
  assign n1001 = ~n979 & ~n985 ;
  assign n1002 = ~n978 & ~n1001 ;
  assign n1003 = ~n997 & n1002 ;
  assign n1004 = n997 & ~n1002 ;
  assign n1005 = ~n1003 & ~n1004 ;
  assign n1008 = ~n1005 & ~x300 ;
  assign n1009 = ~n1007 & ~n1008 ;
  assign n1010 = ~n994 & ~n995 ;
  assign n1011 = ~n996 & ~n1010 ;
  assign n1012 = ~x45 & ~x173 ;
  assign n1013 = x45 & x173 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = n1011 & ~n1014 ;
  assign n1016 = ~n1011 & n1014 ;
  assign n1017 = ~n1015 & ~n1016 ;
  assign n1024 = n1017 & x301 ;
  assign n1018 = ~n996 & ~n1002 ;
  assign n1019 = ~n995 & ~n1018 ;
  assign n1020 = ~n1014 & n1019 ;
  assign n1021 = n1014 & ~n1019 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1025 = ~n1022 & ~x301 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~n1011 & ~n1012 ;
  assign n1028 = ~n1013 & ~n1027 ;
  assign n1029 = ~x46 & ~x174 ;
  assign n1030 = x46 & x174 ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = n1028 & ~n1031 ;
  assign n1033 = ~n1028 & n1031 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1041 = n1034 & x302 ;
  assign n1035 = ~n1013 & ~n1019 ;
  assign n1036 = ~n1012 & ~n1035 ;
  assign n1037 = ~n1031 & n1036 ;
  assign n1038 = n1031 & ~n1036 ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1042 = ~n1039 & ~x302 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = ~n1028 & ~n1029 ;
  assign n1045 = ~n1030 & ~n1044 ;
  assign n1046 = ~x47 & ~x175 ;
  assign n1047 = x47 & x175 ;
  assign n1048 = ~n1046 & ~n1047 ;
  assign n1049 = n1045 & ~n1048 ;
  assign n1050 = ~n1045 & n1048 ;
  assign n1051 = ~n1049 & ~n1050 ;
  assign n1058 = n1051 & x303 ;
  assign n1052 = ~n1030 & ~n1036 ;
  assign n1053 = ~n1029 & ~n1052 ;
  assign n1054 = ~n1048 & n1053 ;
  assign n1055 = n1048 & ~n1053 ;
  assign n1056 = ~n1054 & ~n1055 ;
  assign n1059 = ~n1056 & ~x303 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1061 = ~n1045 & ~n1046 ;
  assign n1062 = ~n1047 & ~n1061 ;
  assign n1063 = ~x48 & ~x176 ;
  assign n1064 = x48 & x176 ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = n1062 & ~n1065 ;
  assign n1067 = ~n1062 & n1065 ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1075 = n1068 & x304 ;
  assign n1069 = ~n1047 & ~n1053 ;
  assign n1070 = ~n1046 & ~n1069 ;
  assign n1071 = ~n1065 & n1070 ;
  assign n1072 = n1065 & ~n1070 ;
  assign n1073 = ~n1071 & ~n1072 ;
  assign n1076 = ~n1073 & ~x304 ;
  assign n1077 = ~n1075 & ~n1076 ;
  assign n1078 = ~n1062 & ~n1063 ;
  assign n1079 = ~n1064 & ~n1078 ;
  assign n1080 = ~x49 & ~x177 ;
  assign n1081 = x49 & x177 ;
  assign n1082 = ~n1080 & ~n1081 ;
  assign n1083 = n1079 & ~n1082 ;
  assign n1084 = ~n1079 & n1082 ;
  assign n1085 = ~n1083 & ~n1084 ;
  assign n1092 = n1085 & x305 ;
  assign n1086 = ~n1064 & ~n1070 ;
  assign n1087 = ~n1063 & ~n1086 ;
  assign n1088 = ~n1082 & n1087 ;
  assign n1089 = n1082 & ~n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1093 = ~n1090 & ~x305 ;
  assign n1094 = ~n1092 & ~n1093 ;
  assign n1095 = ~n1079 & ~n1080 ;
  assign n1096 = ~n1081 & ~n1095 ;
  assign n1097 = ~x50 & ~x178 ;
  assign n1098 = x50 & x178 ;
  assign n1099 = ~n1097 & ~n1098 ;
  assign n1100 = n1096 & ~n1099 ;
  assign n1101 = ~n1096 & n1099 ;
  assign n1102 = ~n1100 & ~n1101 ;
  assign n1109 = n1102 & x306 ;
  assign n1103 = ~n1081 & ~n1087 ;
  assign n1104 = ~n1080 & ~n1103 ;
  assign n1105 = ~n1099 & n1104 ;
  assign n1106 = n1099 & ~n1104 ;
  assign n1107 = ~n1105 & ~n1106 ;
  assign n1110 = ~n1107 & ~x306 ;
  assign n1111 = ~n1109 & ~n1110 ;
  assign n1112 = ~n1096 & ~n1097 ;
  assign n1113 = ~n1098 & ~n1112 ;
  assign n1114 = ~x51 & ~x179 ;
  assign n1115 = x51 & x179 ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1117 = n1113 & ~n1116 ;
  assign n1118 = ~n1113 & n1116 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1126 = n1119 & x307 ;
  assign n1120 = ~n1098 & ~n1104 ;
  assign n1121 = ~n1097 & ~n1120 ;
  assign n1122 = ~n1116 & n1121 ;
  assign n1123 = n1116 & ~n1121 ;
  assign n1124 = ~n1122 & ~n1123 ;
  assign n1127 = ~n1124 & ~x307 ;
  assign n1128 = ~n1126 & ~n1127 ;
  assign n1129 = ~n1113 & ~n1114 ;
  assign n1130 = ~n1115 & ~n1129 ;
  assign n1131 = ~x52 & ~x180 ;
  assign n1132 = x52 & x180 ;
  assign n1133 = ~n1131 & ~n1132 ;
  assign n1134 = n1130 & ~n1133 ;
  assign n1135 = ~n1130 & n1133 ;
  assign n1136 = ~n1134 & ~n1135 ;
  assign n1143 = n1136 & x308 ;
  assign n1137 = ~n1115 & ~n1121 ;
  assign n1138 = ~n1114 & ~n1137 ;
  assign n1139 = ~n1133 & n1138 ;
  assign n1140 = n1133 & ~n1138 ;
  assign n1141 = ~n1139 & ~n1140 ;
  assign n1144 = ~n1141 & ~x308 ;
  assign n1145 = ~n1143 & ~n1144 ;
  assign n1146 = ~n1130 & ~n1131 ;
  assign n1147 = ~n1132 & ~n1146 ;
  assign n1148 = ~x53 & ~x181 ;
  assign n1149 = x53 & x181 ;
  assign n1150 = ~n1148 & ~n1149 ;
  assign n1151 = n1147 & ~n1150 ;
  assign n1152 = ~n1147 & n1150 ;
  assign n1153 = ~n1151 & ~n1152 ;
  assign n1160 = n1153 & x309 ;
  assign n1154 = ~n1132 & ~n1138 ;
  assign n1155 = ~n1131 & ~n1154 ;
  assign n1156 = ~n1150 & n1155 ;
  assign n1157 = n1150 & ~n1155 ;
  assign n1158 = ~n1156 & ~n1157 ;
  assign n1161 = ~n1158 & ~x309 ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = ~n1147 & ~n1148 ;
  assign n1164 = ~n1149 & ~n1163 ;
  assign n1165 = ~x54 & ~x182 ;
  assign n1166 = x54 & x182 ;
  assign n1167 = ~n1165 & ~n1166 ;
  assign n1168 = n1164 & ~n1167 ;
  assign n1169 = ~n1164 & n1167 ;
  assign n1170 = ~n1168 & ~n1169 ;
  assign n1177 = n1170 & x310 ;
  assign n1171 = ~n1149 & ~n1155 ;
  assign n1172 = ~n1148 & ~n1171 ;
  assign n1173 = ~n1167 & n1172 ;
  assign n1174 = n1167 & ~n1172 ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1178 = ~n1175 & ~x310 ;
  assign n1179 = ~n1177 & ~n1178 ;
  assign n1180 = ~n1164 & ~n1165 ;
  assign n1181 = ~n1166 & ~n1180 ;
  assign n1182 = ~x55 & ~x183 ;
  assign n1183 = x55 & x183 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = n1181 & ~n1184 ;
  assign n1186 = ~n1181 & n1184 ;
  assign n1187 = ~n1185 & ~n1186 ;
  assign n1194 = n1187 & x311 ;
  assign n1188 = ~n1166 & ~n1172 ;
  assign n1189 = ~n1165 & ~n1188 ;
  assign n1190 = ~n1184 & n1189 ;
  assign n1191 = n1184 & ~n1189 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1195 = ~n1192 & ~x311 ;
  assign n1196 = ~n1194 & ~n1195 ;
  assign n1197 = ~n1181 & ~n1182 ;
  assign n1198 = ~n1183 & ~n1197 ;
  assign n1199 = ~x56 & ~x184 ;
  assign n1200 = x56 & x184 ;
  assign n1201 = ~n1199 & ~n1200 ;
  assign n1202 = n1198 & ~n1201 ;
  assign n1203 = ~n1198 & n1201 ;
  assign n1204 = ~n1202 & ~n1203 ;
  assign n1211 = n1204 & x312 ;
  assign n1205 = ~n1183 & ~n1189 ;
  assign n1206 = ~n1182 & ~n1205 ;
  assign n1207 = ~n1201 & n1206 ;
  assign n1208 = n1201 & ~n1206 ;
  assign n1209 = ~n1207 & ~n1208 ;
  assign n1212 = ~n1209 & ~x312 ;
  assign n1213 = ~n1211 & ~n1212 ;
  assign n1214 = ~n1198 & ~n1199 ;
  assign n1215 = ~n1200 & ~n1214 ;
  assign n1216 = ~x57 & ~x185 ;
  assign n1217 = x57 & x185 ;
  assign n1218 = ~n1216 & ~n1217 ;
  assign n1219 = n1215 & ~n1218 ;
  assign n1220 = ~n1215 & n1218 ;
  assign n1221 = ~n1219 & ~n1220 ;
  assign n1228 = n1221 & x313 ;
  assign n1222 = ~n1200 & ~n1206 ;
  assign n1223 = ~n1199 & ~n1222 ;
  assign n1224 = ~n1218 & n1223 ;
  assign n1225 = n1218 & ~n1223 ;
  assign n1226 = ~n1224 & ~n1225 ;
  assign n1229 = ~n1226 & ~x313 ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = ~n1215 & ~n1216 ;
  assign n1232 = ~n1217 & ~n1231 ;
  assign n1233 = ~x58 & ~x186 ;
  assign n1234 = x58 & x186 ;
  assign n1235 = ~n1233 & ~n1234 ;
  assign n1236 = n1232 & ~n1235 ;
  assign n1237 = ~n1232 & n1235 ;
  assign n1238 = ~n1236 & ~n1237 ;
  assign n1245 = n1238 & x314 ;
  assign n1239 = ~n1217 & ~n1223 ;
  assign n1240 = ~n1216 & ~n1239 ;
  assign n1241 = ~n1235 & n1240 ;
  assign n1242 = n1235 & ~n1240 ;
  assign n1243 = ~n1241 & ~n1242 ;
  assign n1246 = ~n1243 & ~x314 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = ~n1232 & ~n1233 ;
  assign n1249 = ~n1234 & ~n1248 ;
  assign n1250 = ~x59 & ~x187 ;
  assign n1251 = x59 & x187 ;
  assign n1252 = ~n1250 & ~n1251 ;
  assign n1253 = n1249 & ~n1252 ;
  assign n1254 = ~n1249 & n1252 ;
  assign n1255 = ~n1253 & ~n1254 ;
  assign n1262 = n1255 & x315 ;
  assign n1256 = ~n1234 & ~n1240 ;
  assign n1257 = ~n1233 & ~n1256 ;
  assign n1258 = ~n1252 & n1257 ;
  assign n1259 = n1252 & ~n1257 ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1263 = ~n1260 & ~x315 ;
  assign n1264 = ~n1262 & ~n1263 ;
  assign n1265 = ~n1249 & ~n1250 ;
  assign n1266 = ~n1251 & ~n1265 ;
  assign n1267 = ~x60 & ~x188 ;
  assign n1268 = x60 & x188 ;
  assign n1269 = ~n1267 & ~n1268 ;
  assign n1270 = n1266 & ~n1269 ;
  assign n1271 = ~n1266 & n1269 ;
  assign n1272 = ~n1270 & ~n1271 ;
  assign n1279 = n1272 & x316 ;
  assign n1273 = ~n1251 & ~n1257 ;
  assign n1274 = ~n1250 & ~n1273 ;
  assign n1275 = ~n1269 & n1274 ;
  assign n1276 = n1269 & ~n1274 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1280 = ~n1277 & ~x316 ;
  assign n1281 = ~n1279 & ~n1280 ;
  assign n1282 = ~n1266 & ~n1267 ;
  assign n1283 = ~n1268 & ~n1282 ;
  assign n1284 = ~x61 & ~x189 ;
  assign n1285 = x61 & x189 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = n1283 & ~n1286 ;
  assign n1288 = ~n1283 & n1286 ;
  assign n1289 = ~n1287 & ~n1288 ;
  assign n1296 = n1289 & x317 ;
  assign n1290 = ~n1268 & ~n1274 ;
  assign n1291 = ~n1267 & ~n1290 ;
  assign n1292 = ~n1286 & n1291 ;
  assign n1293 = n1286 & ~n1291 ;
  assign n1294 = ~n1292 & ~n1293 ;
  assign n1297 = ~n1294 & ~x317 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = ~n1283 & ~n1284 ;
  assign n1300 = ~n1285 & ~n1299 ;
  assign n1301 = ~x62 & ~x190 ;
  assign n1302 = x62 & x190 ;
  assign n1303 = ~n1301 & ~n1302 ;
  assign n1304 = n1300 & ~n1303 ;
  assign n1305 = ~n1300 & n1303 ;
  assign n1306 = ~n1304 & ~n1305 ;
  assign n1313 = n1306 & x318 ;
  assign n1307 = ~n1285 & ~n1291 ;
  assign n1308 = ~n1284 & ~n1307 ;
  assign n1309 = ~n1303 & n1308 ;
  assign n1310 = n1303 & ~n1308 ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1314 = ~n1311 & ~x318 ;
  assign n1315 = ~n1313 & ~n1314 ;
  assign n1316 = ~n1300 & ~n1301 ;
  assign n1317 = ~n1302 & ~n1316 ;
  assign n1318 = ~x63 & ~x191 ;
  assign n1319 = x63 & x191 ;
  assign n1320 = ~n1318 & ~n1319 ;
  assign n1321 = n1317 & ~n1320 ;
  assign n1322 = ~n1317 & n1320 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1330 = n1323 & x319 ;
  assign n1324 = ~n1302 & ~n1308 ;
  assign n1325 = ~n1301 & ~n1324 ;
  assign n1326 = ~n1320 & n1325 ;
  assign n1327 = n1320 & ~n1325 ;
  assign n1328 = ~n1326 & ~n1327 ;
  assign n1331 = ~n1328 & ~x319 ;
  assign n1332 = ~n1330 & ~n1331 ;
  assign n1333 = ~n1317 & ~n1318 ;
  assign n1334 = ~n1319 & ~n1333 ;
  assign n1335 = ~x64 & ~x192 ;
  assign n1336 = x64 & x192 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = n1334 & ~n1337 ;
  assign n1339 = ~n1334 & n1337 ;
  assign n1340 = ~n1338 & ~n1339 ;
  assign n1347 = n1340 & x320 ;
  assign n1341 = ~n1319 & ~n1325 ;
  assign n1342 = ~n1318 & ~n1341 ;
  assign n1343 = ~n1337 & n1342 ;
  assign n1344 = n1337 & ~n1342 ;
  assign n1345 = ~n1343 & ~n1344 ;
  assign n1348 = ~n1345 & ~x320 ;
  assign n1349 = ~n1347 & ~n1348 ;
  assign n1350 = ~n1334 & ~n1335 ;
  assign n1351 = ~n1336 & ~n1350 ;
  assign n1352 = ~x65 & ~x193 ;
  assign n1353 = x65 & x193 ;
  assign n1354 = ~n1352 & ~n1353 ;
  assign n1355 = n1351 & ~n1354 ;
  assign n1356 = ~n1351 & n1354 ;
  assign n1357 = ~n1355 & ~n1356 ;
  assign n1364 = n1357 & x321 ;
  assign n1358 = ~n1336 & ~n1342 ;
  assign n1359 = ~n1335 & ~n1358 ;
  assign n1360 = ~n1354 & n1359 ;
  assign n1361 = n1354 & ~n1359 ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1365 = ~n1362 & ~x321 ;
  assign n1366 = ~n1364 & ~n1365 ;
  assign n1367 = ~n1351 & ~n1352 ;
  assign n1368 = ~n1353 & ~n1367 ;
  assign n1369 = ~x66 & ~x194 ;
  assign n1370 = x66 & x194 ;
  assign n1371 = ~n1369 & ~n1370 ;
  assign n1372 = n1368 & ~n1371 ;
  assign n1373 = ~n1368 & n1371 ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1381 = n1374 & x322 ;
  assign n1375 = ~n1353 & ~n1359 ;
  assign n1376 = ~n1352 & ~n1375 ;
  assign n1377 = ~n1371 & n1376 ;
  assign n1378 = n1371 & ~n1376 ;
  assign n1379 = ~n1377 & ~n1378 ;
  assign n1382 = ~n1379 & ~x322 ;
  assign n1383 = ~n1381 & ~n1382 ;
  assign n1384 = ~n1368 & ~n1369 ;
  assign n1385 = ~n1370 & ~n1384 ;
  assign n1386 = ~x67 & ~x195 ;
  assign n1387 = x67 & x195 ;
  assign n1388 = ~n1386 & ~n1387 ;
  assign n1389 = n1385 & ~n1388 ;
  assign n1390 = ~n1385 & n1388 ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1398 = n1391 & x323 ;
  assign n1392 = ~n1370 & ~n1376 ;
  assign n1393 = ~n1369 & ~n1392 ;
  assign n1394 = ~n1388 & n1393 ;
  assign n1395 = n1388 & ~n1393 ;
  assign n1396 = ~n1394 & ~n1395 ;
  assign n1399 = ~n1396 & ~x323 ;
  assign n1400 = ~n1398 & ~n1399 ;
  assign n1401 = ~n1385 & ~n1386 ;
  assign n1402 = ~n1387 & ~n1401 ;
  assign n1403 = ~x68 & ~x196 ;
  assign n1404 = x68 & x196 ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = n1402 & ~n1405 ;
  assign n1407 = ~n1402 & n1405 ;
  assign n1408 = ~n1406 & ~n1407 ;
  assign n1415 = n1408 & x324 ;
  assign n1409 = ~n1387 & ~n1393 ;
  assign n1410 = ~n1386 & ~n1409 ;
  assign n1411 = ~n1405 & n1410 ;
  assign n1412 = n1405 & ~n1410 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1416 = ~n1413 & ~x324 ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = ~n1402 & ~n1403 ;
  assign n1419 = ~n1404 & ~n1418 ;
  assign n1420 = ~x69 & ~x197 ;
  assign n1421 = x69 & x197 ;
  assign n1422 = ~n1420 & ~n1421 ;
  assign n1423 = n1419 & ~n1422 ;
  assign n1424 = ~n1419 & n1422 ;
  assign n1425 = ~n1423 & ~n1424 ;
  assign n1432 = n1425 & x325 ;
  assign n1426 = ~n1404 & ~n1410 ;
  assign n1427 = ~n1403 & ~n1426 ;
  assign n1428 = ~n1422 & n1427 ;
  assign n1429 = n1422 & ~n1427 ;
  assign n1430 = ~n1428 & ~n1429 ;
  assign n1433 = ~n1430 & ~x325 ;
  assign n1434 = ~n1432 & ~n1433 ;
  assign n1435 = ~n1419 & ~n1420 ;
  assign n1436 = ~n1421 & ~n1435 ;
  assign n1437 = ~x70 & ~x198 ;
  assign n1438 = x70 & x198 ;
  assign n1439 = ~n1437 & ~n1438 ;
  assign n1440 = n1436 & ~n1439 ;
  assign n1441 = ~n1436 & n1439 ;
  assign n1442 = ~n1440 & ~n1441 ;
  assign n1449 = n1442 & x326 ;
  assign n1443 = ~n1421 & ~n1427 ;
  assign n1444 = ~n1420 & ~n1443 ;
  assign n1445 = ~n1439 & n1444 ;
  assign n1446 = n1439 & ~n1444 ;
  assign n1447 = ~n1445 & ~n1446 ;
  assign n1450 = ~n1447 & ~x326 ;
  assign n1451 = ~n1449 & ~n1450 ;
  assign n1452 = ~n1436 & ~n1437 ;
  assign n1453 = ~n1438 & ~n1452 ;
  assign n1454 = ~x71 & ~x199 ;
  assign n1455 = x71 & x199 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = n1453 & ~n1456 ;
  assign n1458 = ~n1453 & n1456 ;
  assign n1459 = ~n1457 & ~n1458 ;
  assign n1466 = n1459 & x327 ;
  assign n1460 = ~n1438 & ~n1444 ;
  assign n1461 = ~n1437 & ~n1460 ;
  assign n1462 = ~n1456 & n1461 ;
  assign n1463 = n1456 & ~n1461 ;
  assign n1464 = ~n1462 & ~n1463 ;
  assign n1467 = ~n1464 & ~x327 ;
  assign n1468 = ~n1466 & ~n1467 ;
  assign n1469 = ~n1453 & ~n1454 ;
  assign n1470 = ~n1455 & ~n1469 ;
  assign n1471 = ~x72 & ~x200 ;
  assign n1472 = x72 & x200 ;
  assign n1473 = ~n1471 & ~n1472 ;
  assign n1474 = n1470 & ~n1473 ;
  assign n1475 = ~n1470 & n1473 ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1483 = n1476 & x328 ;
  assign n1477 = ~n1455 & ~n1461 ;
  assign n1478 = ~n1454 & ~n1477 ;
  assign n1479 = ~n1473 & n1478 ;
  assign n1480 = n1473 & ~n1478 ;
  assign n1481 = ~n1479 & ~n1480 ;
  assign n1484 = ~n1481 & ~x328 ;
  assign n1485 = ~n1483 & ~n1484 ;
  assign n1486 = ~n1470 & ~n1471 ;
  assign n1487 = ~n1472 & ~n1486 ;
  assign n1488 = ~x73 & ~x201 ;
  assign n1489 = x73 & x201 ;
  assign n1490 = ~n1488 & ~n1489 ;
  assign n1491 = n1487 & ~n1490 ;
  assign n1492 = ~n1487 & n1490 ;
  assign n1493 = ~n1491 & ~n1492 ;
  assign n1500 = n1493 & x329 ;
  assign n1494 = ~n1472 & ~n1478 ;
  assign n1495 = ~n1471 & ~n1494 ;
  assign n1496 = ~n1490 & n1495 ;
  assign n1497 = n1490 & ~n1495 ;
  assign n1498 = ~n1496 & ~n1497 ;
  assign n1501 = ~n1498 & ~x329 ;
  assign n1502 = ~n1500 & ~n1501 ;
  assign n1503 = ~n1487 & ~n1488 ;
  assign n1504 = ~n1489 & ~n1503 ;
  assign n1505 = ~x74 & ~x202 ;
  assign n1506 = x74 & x202 ;
  assign n1507 = ~n1505 & ~n1506 ;
  assign n1508 = n1504 & ~n1507 ;
  assign n1509 = ~n1504 & n1507 ;
  assign n1510 = ~n1508 & ~n1509 ;
  assign n1517 = n1510 & x330 ;
  assign n1511 = ~n1489 & ~n1495 ;
  assign n1512 = ~n1488 & ~n1511 ;
  assign n1513 = ~n1507 & n1512 ;
  assign n1514 = n1507 & ~n1512 ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1518 = ~n1515 & ~x330 ;
  assign n1519 = ~n1517 & ~n1518 ;
  assign n1520 = ~n1504 & ~n1505 ;
  assign n1521 = ~n1506 & ~n1520 ;
  assign n1522 = ~x75 & ~x203 ;
  assign n1523 = x75 & x203 ;
  assign n1524 = ~n1522 & ~n1523 ;
  assign n1525 = n1521 & ~n1524 ;
  assign n1526 = ~n1521 & n1524 ;
  assign n1527 = ~n1525 & ~n1526 ;
  assign n1534 = n1527 & x331 ;
  assign n1528 = ~n1506 & ~n1512 ;
  assign n1529 = ~n1505 & ~n1528 ;
  assign n1530 = ~n1524 & n1529 ;
  assign n1531 = n1524 & ~n1529 ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1535 = ~n1532 & ~x331 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = ~n1521 & ~n1522 ;
  assign n1538 = ~n1523 & ~n1537 ;
  assign n1539 = ~x76 & ~x204 ;
  assign n1540 = x76 & x204 ;
  assign n1541 = ~n1539 & ~n1540 ;
  assign n1542 = n1538 & ~n1541 ;
  assign n1543 = ~n1538 & n1541 ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1551 = n1544 & x332 ;
  assign n1545 = ~n1523 & ~n1529 ;
  assign n1546 = ~n1522 & ~n1545 ;
  assign n1547 = ~n1541 & n1546 ;
  assign n1548 = n1541 & ~n1546 ;
  assign n1549 = ~n1547 & ~n1548 ;
  assign n1552 = ~n1549 & ~x332 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = ~n1538 & ~n1539 ;
  assign n1555 = ~n1540 & ~n1554 ;
  assign n1556 = ~x77 & ~x205 ;
  assign n1557 = x77 & x205 ;
  assign n1558 = ~n1556 & ~n1557 ;
  assign n1559 = n1555 & ~n1558 ;
  assign n1560 = ~n1555 & n1558 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1568 = n1561 & x333 ;
  assign n1562 = ~n1540 & ~n1546 ;
  assign n1563 = ~n1539 & ~n1562 ;
  assign n1564 = ~n1558 & n1563 ;
  assign n1565 = n1558 & ~n1563 ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1569 = ~n1566 & ~x333 ;
  assign n1570 = ~n1568 & ~n1569 ;
  assign n1571 = ~n1555 & ~n1556 ;
  assign n1572 = ~n1557 & ~n1571 ;
  assign n1573 = ~x78 & ~x206 ;
  assign n1574 = x78 & x206 ;
  assign n1575 = ~n1573 & ~n1574 ;
  assign n1576 = n1572 & ~n1575 ;
  assign n1577 = ~n1572 & n1575 ;
  assign n1578 = ~n1576 & ~n1577 ;
  assign n1585 = n1578 & x334 ;
  assign n1579 = ~n1557 & ~n1563 ;
  assign n1580 = ~n1556 & ~n1579 ;
  assign n1581 = ~n1575 & n1580 ;
  assign n1582 = n1575 & ~n1580 ;
  assign n1583 = ~n1581 & ~n1582 ;
  assign n1586 = ~n1583 & ~x334 ;
  assign n1587 = ~n1585 & ~n1586 ;
  assign n1588 = ~n1572 & ~n1573 ;
  assign n1589 = ~n1574 & ~n1588 ;
  assign n1590 = ~x79 & ~x207 ;
  assign n1591 = x79 & x207 ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = n1589 & ~n1592 ;
  assign n1594 = ~n1589 & n1592 ;
  assign n1595 = ~n1593 & ~n1594 ;
  assign n1602 = n1595 & x335 ;
  assign n1596 = ~n1574 & ~n1580 ;
  assign n1597 = ~n1573 & ~n1596 ;
  assign n1598 = ~n1592 & n1597 ;
  assign n1599 = n1592 & ~n1597 ;
  assign n1600 = ~n1598 & ~n1599 ;
  assign n1603 = ~n1600 & ~x335 ;
  assign n1604 = ~n1602 & ~n1603 ;
  assign n1605 = ~n1589 & ~n1590 ;
  assign n1606 = ~n1591 & ~n1605 ;
  assign n1607 = ~x80 & ~x208 ;
  assign n1608 = x80 & x208 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = n1606 & ~n1609 ;
  assign n1611 = ~n1606 & n1609 ;
  assign n1612 = ~n1610 & ~n1611 ;
  assign n1619 = n1612 & x336 ;
  assign n1613 = ~n1591 & ~n1597 ;
  assign n1614 = ~n1590 & ~n1613 ;
  assign n1615 = ~n1609 & n1614 ;
  assign n1616 = n1609 & ~n1614 ;
  assign n1617 = ~n1615 & ~n1616 ;
  assign n1620 = ~n1617 & ~x336 ;
  assign n1621 = ~n1619 & ~n1620 ;
  assign n1622 = ~n1606 & ~n1607 ;
  assign n1623 = ~n1608 & ~n1622 ;
  assign n1624 = ~x81 & ~x209 ;
  assign n1625 = x81 & x209 ;
  assign n1626 = ~n1624 & ~n1625 ;
  assign n1627 = n1623 & ~n1626 ;
  assign n1628 = ~n1623 & n1626 ;
  assign n1629 = ~n1627 & ~n1628 ;
  assign n1636 = n1629 & x337 ;
  assign n1630 = ~n1608 & ~n1614 ;
  assign n1631 = ~n1607 & ~n1630 ;
  assign n1632 = ~n1626 & n1631 ;
  assign n1633 = n1626 & ~n1631 ;
  assign n1634 = ~n1632 & ~n1633 ;
  assign n1637 = ~n1634 & ~x337 ;
  assign n1638 = ~n1636 & ~n1637 ;
  assign n1639 = ~n1623 & ~n1624 ;
  assign n1640 = ~n1625 & ~n1639 ;
  assign n1641 = ~x82 & ~x210 ;
  assign n1642 = x82 & x210 ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = n1640 & ~n1643 ;
  assign n1645 = ~n1640 & n1643 ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1653 = n1646 & x338 ;
  assign n1647 = ~n1625 & ~n1631 ;
  assign n1648 = ~n1624 & ~n1647 ;
  assign n1649 = ~n1643 & n1648 ;
  assign n1650 = n1643 & ~n1648 ;
  assign n1651 = ~n1649 & ~n1650 ;
  assign n1654 = ~n1651 & ~x338 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = ~n1640 & ~n1641 ;
  assign n1657 = ~n1642 & ~n1656 ;
  assign n1658 = ~x83 & ~x211 ;
  assign n1659 = x83 & x211 ;
  assign n1660 = ~n1658 & ~n1659 ;
  assign n1661 = n1657 & ~n1660 ;
  assign n1662 = ~n1657 & n1660 ;
  assign n1663 = ~n1661 & ~n1662 ;
  assign n1670 = n1663 & x339 ;
  assign n1664 = ~n1642 & ~n1648 ;
  assign n1665 = ~n1641 & ~n1664 ;
  assign n1666 = ~n1660 & n1665 ;
  assign n1667 = n1660 & ~n1665 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1671 = ~n1668 & ~x339 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = ~n1657 & ~n1658 ;
  assign n1674 = ~n1659 & ~n1673 ;
  assign n1675 = ~x84 & ~x212 ;
  assign n1676 = x84 & x212 ;
  assign n1677 = ~n1675 & ~n1676 ;
  assign n1678 = n1674 & ~n1677 ;
  assign n1679 = ~n1674 & n1677 ;
  assign n1680 = ~n1678 & ~n1679 ;
  assign n1687 = n1680 & x340 ;
  assign n1681 = ~n1659 & ~n1665 ;
  assign n1682 = ~n1658 & ~n1681 ;
  assign n1683 = ~n1677 & n1682 ;
  assign n1684 = n1677 & ~n1682 ;
  assign n1685 = ~n1683 & ~n1684 ;
  assign n1688 = ~n1685 & ~x340 ;
  assign n1689 = ~n1687 & ~n1688 ;
  assign n1690 = ~n1674 & ~n1675 ;
  assign n1691 = ~n1676 & ~n1690 ;
  assign n1692 = ~x85 & ~x213 ;
  assign n1693 = x85 & x213 ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = n1691 & ~n1694 ;
  assign n1696 = ~n1691 & n1694 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1704 = n1697 & x341 ;
  assign n1698 = ~n1676 & ~n1682 ;
  assign n1699 = ~n1675 & ~n1698 ;
  assign n1700 = ~n1694 & n1699 ;
  assign n1701 = n1694 & ~n1699 ;
  assign n1702 = ~n1700 & ~n1701 ;
  assign n1705 = ~n1702 & ~x341 ;
  assign n1706 = ~n1704 & ~n1705 ;
  assign n1707 = ~n1691 & ~n1692 ;
  assign n1708 = ~n1693 & ~n1707 ;
  assign n1709 = ~x86 & ~x214 ;
  assign n1710 = x86 & x214 ;
  assign n1711 = ~n1709 & ~n1710 ;
  assign n1712 = n1708 & ~n1711 ;
  assign n1713 = ~n1708 & n1711 ;
  assign n1714 = ~n1712 & ~n1713 ;
  assign n1721 = n1714 & x342 ;
  assign n1715 = ~n1693 & ~n1699 ;
  assign n1716 = ~n1692 & ~n1715 ;
  assign n1717 = ~n1711 & n1716 ;
  assign n1718 = n1711 & ~n1716 ;
  assign n1719 = ~n1717 & ~n1718 ;
  assign n1722 = ~n1719 & ~x342 ;
  assign n1723 = ~n1721 & ~n1722 ;
  assign n1724 = ~n1708 & ~n1709 ;
  assign n1725 = ~n1710 & ~n1724 ;
  assign n1726 = ~x87 & ~x215 ;
  assign n1727 = x87 & x215 ;
  assign n1728 = ~n1726 & ~n1727 ;
  assign n1729 = n1725 & ~n1728 ;
  assign n1730 = ~n1725 & n1728 ;
  assign n1731 = ~n1729 & ~n1730 ;
  assign n1738 = n1731 & x343 ;
  assign n1732 = ~n1710 & ~n1716 ;
  assign n1733 = ~n1709 & ~n1732 ;
  assign n1734 = ~n1728 & n1733 ;
  assign n1735 = n1728 & ~n1733 ;
  assign n1736 = ~n1734 & ~n1735 ;
  assign n1739 = ~n1736 & ~x343 ;
  assign n1740 = ~n1738 & ~n1739 ;
  assign n1741 = ~n1725 & ~n1726 ;
  assign n1742 = ~n1727 & ~n1741 ;
  assign n1743 = ~x88 & ~x216 ;
  assign n1744 = x88 & x216 ;
  assign n1745 = ~n1743 & ~n1744 ;
  assign n1746 = n1742 & ~n1745 ;
  assign n1747 = ~n1742 & n1745 ;
  assign n1748 = ~n1746 & ~n1747 ;
  assign n1755 = n1748 & x344 ;
  assign n1749 = ~n1727 & ~n1733 ;
  assign n1750 = ~n1726 & ~n1749 ;
  assign n1751 = ~n1745 & n1750 ;
  assign n1752 = n1745 & ~n1750 ;
  assign n1753 = ~n1751 & ~n1752 ;
  assign n1756 = ~n1753 & ~x344 ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = ~n1742 & ~n1743 ;
  assign n1759 = ~n1744 & ~n1758 ;
  assign n1760 = ~x89 & ~x217 ;
  assign n1761 = x89 & x217 ;
  assign n1762 = ~n1760 & ~n1761 ;
  assign n1763 = n1759 & ~n1762 ;
  assign n1764 = ~n1759 & n1762 ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1772 = n1765 & x345 ;
  assign n1766 = ~n1744 & ~n1750 ;
  assign n1767 = ~n1743 & ~n1766 ;
  assign n1768 = ~n1762 & n1767 ;
  assign n1769 = n1762 & ~n1767 ;
  assign n1770 = ~n1768 & ~n1769 ;
  assign n1773 = ~n1770 & ~x345 ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = ~n1759 & ~n1760 ;
  assign n1776 = ~n1761 & ~n1775 ;
  assign n1777 = ~x90 & ~x218 ;
  assign n1778 = x90 & x218 ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1780 = n1776 & ~n1779 ;
  assign n1781 = ~n1776 & n1779 ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1789 = n1782 & x346 ;
  assign n1783 = ~n1761 & ~n1767 ;
  assign n1784 = ~n1760 & ~n1783 ;
  assign n1785 = ~n1779 & n1784 ;
  assign n1786 = n1779 & ~n1784 ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1790 = ~n1787 & ~x346 ;
  assign n1791 = ~n1789 & ~n1790 ;
  assign n1792 = ~n1776 & ~n1777 ;
  assign n1793 = ~n1778 & ~n1792 ;
  assign n1794 = ~x91 & ~x219 ;
  assign n1795 = x91 & x219 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = n1793 & ~n1796 ;
  assign n1798 = ~n1793 & n1796 ;
  assign n1799 = ~n1797 & ~n1798 ;
  assign n1806 = n1799 & x347 ;
  assign n1800 = ~n1778 & ~n1784 ;
  assign n1801 = ~n1777 & ~n1800 ;
  assign n1802 = ~n1796 & n1801 ;
  assign n1803 = n1796 & ~n1801 ;
  assign n1804 = ~n1802 & ~n1803 ;
  assign n1807 = ~n1804 & ~x347 ;
  assign n1808 = ~n1806 & ~n1807 ;
  assign n1809 = ~n1793 & ~n1794 ;
  assign n1810 = ~n1795 & ~n1809 ;
  assign n1811 = ~x92 & ~x220 ;
  assign n1812 = x92 & x220 ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = n1810 & ~n1813 ;
  assign n1815 = ~n1810 & n1813 ;
  assign n1816 = ~n1814 & ~n1815 ;
  assign n1823 = n1816 & x348 ;
  assign n1817 = ~n1795 & ~n1801 ;
  assign n1818 = ~n1794 & ~n1817 ;
  assign n1819 = ~n1813 & n1818 ;
  assign n1820 = n1813 & ~n1818 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1824 = ~n1821 & ~x348 ;
  assign n1825 = ~n1823 & ~n1824 ;
  assign n1826 = ~n1810 & ~n1811 ;
  assign n1827 = ~n1812 & ~n1826 ;
  assign n1828 = ~x93 & ~x221 ;
  assign n1829 = x93 & x221 ;
  assign n1830 = ~n1828 & ~n1829 ;
  assign n1831 = n1827 & ~n1830 ;
  assign n1832 = ~n1827 & n1830 ;
  assign n1833 = ~n1831 & ~n1832 ;
  assign n1840 = n1833 & x349 ;
  assign n1834 = ~n1812 & ~n1818 ;
  assign n1835 = ~n1811 & ~n1834 ;
  assign n1836 = ~n1830 & n1835 ;
  assign n1837 = n1830 & ~n1835 ;
  assign n1838 = ~n1836 & ~n1837 ;
  assign n1841 = ~n1838 & ~x349 ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = ~n1827 & ~n1828 ;
  assign n1844 = ~n1829 & ~n1843 ;
  assign n1845 = ~x94 & ~x222 ;
  assign n1846 = x94 & x222 ;
  assign n1847 = ~n1845 & ~n1846 ;
  assign n1848 = n1844 & ~n1847 ;
  assign n1849 = ~n1844 & n1847 ;
  assign n1850 = ~n1848 & ~n1849 ;
  assign n1857 = n1850 & x350 ;
  assign n1851 = ~n1829 & ~n1835 ;
  assign n1852 = ~n1828 & ~n1851 ;
  assign n1853 = ~n1847 & n1852 ;
  assign n1854 = n1847 & ~n1852 ;
  assign n1855 = ~n1853 & ~n1854 ;
  assign n1858 = ~n1855 & ~x350 ;
  assign n1859 = ~n1857 & ~n1858 ;
  assign n1860 = ~n1844 & ~n1845 ;
  assign n1861 = ~n1846 & ~n1860 ;
  assign n1862 = ~x95 & ~x223 ;
  assign n1863 = x95 & x223 ;
  assign n1864 = ~n1862 & ~n1863 ;
  assign n1865 = n1861 & ~n1864 ;
  assign n1866 = ~n1861 & n1864 ;
  assign n1867 = ~n1865 & ~n1866 ;
  assign n1874 = n1867 & x351 ;
  assign n1868 = ~n1846 & ~n1852 ;
  assign n1869 = ~n1845 & ~n1868 ;
  assign n1870 = ~n1864 & n1869 ;
  assign n1871 = n1864 & ~n1869 ;
  assign n1872 = ~n1870 & ~n1871 ;
  assign n1875 = ~n1872 & ~x351 ;
  assign n1876 = ~n1874 & ~n1875 ;
  assign n1877 = ~n1861 & ~n1862 ;
  assign n1878 = ~n1863 & ~n1877 ;
  assign n1879 = ~x96 & ~x224 ;
  assign n1880 = x96 & x224 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = n1878 & ~n1881 ;
  assign n1883 = ~n1878 & n1881 ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1891 = n1884 & x352 ;
  assign n1885 = ~n1863 & ~n1869 ;
  assign n1886 = ~n1862 & ~n1885 ;
  assign n1887 = ~n1881 & n1886 ;
  assign n1888 = n1881 & ~n1886 ;
  assign n1889 = ~n1887 & ~n1888 ;
  assign n1892 = ~n1889 & ~x352 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = ~n1878 & ~n1879 ;
  assign n1895 = ~n1880 & ~n1894 ;
  assign n1896 = ~x97 & ~x225 ;
  assign n1897 = x97 & x225 ;
  assign n1898 = ~n1896 & ~n1897 ;
  assign n1899 = n1895 & ~n1898 ;
  assign n1900 = ~n1895 & n1898 ;
  assign n1901 = ~n1899 & ~n1900 ;
  assign n1908 = n1901 & x353 ;
  assign n1902 = ~n1880 & ~n1886 ;
  assign n1903 = ~n1879 & ~n1902 ;
  assign n1904 = ~n1898 & n1903 ;
  assign n1905 = n1898 & ~n1903 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1909 = ~n1906 & ~x353 ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1911 = ~n1895 & ~n1896 ;
  assign n1912 = ~n1897 & ~n1911 ;
  assign n1913 = ~x98 & ~x226 ;
  assign n1914 = x98 & x226 ;
  assign n1915 = ~n1913 & ~n1914 ;
  assign n1916 = n1912 & ~n1915 ;
  assign n1917 = ~n1912 & n1915 ;
  assign n1918 = ~n1916 & ~n1917 ;
  assign n1925 = n1918 & x354 ;
  assign n1919 = ~n1897 & ~n1903 ;
  assign n1920 = ~n1896 & ~n1919 ;
  assign n1921 = ~n1915 & n1920 ;
  assign n1922 = n1915 & ~n1920 ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1926 = ~n1923 & ~x354 ;
  assign n1927 = ~n1925 & ~n1926 ;
  assign n1928 = ~n1912 & ~n1913 ;
  assign n1929 = ~n1914 & ~n1928 ;
  assign n1930 = ~x99 & ~x227 ;
  assign n1931 = x99 & x227 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = n1929 & ~n1932 ;
  assign n1934 = ~n1929 & n1932 ;
  assign n1935 = ~n1933 & ~n1934 ;
  assign n1942 = n1935 & x355 ;
  assign n1936 = ~n1914 & ~n1920 ;
  assign n1937 = ~n1913 & ~n1936 ;
  assign n1938 = ~n1932 & n1937 ;
  assign n1939 = n1932 & ~n1937 ;
  assign n1940 = ~n1938 & ~n1939 ;
  assign n1943 = ~n1940 & ~x355 ;
  assign n1944 = ~n1942 & ~n1943 ;
  assign n1945 = ~n1929 & ~n1930 ;
  assign n1946 = ~n1931 & ~n1945 ;
  assign n1947 = ~x100 & ~x228 ;
  assign n1948 = x100 & x228 ;
  assign n1949 = ~n1947 & ~n1948 ;
  assign n1950 = n1946 & ~n1949 ;
  assign n1951 = ~n1946 & n1949 ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1959 = n1952 & x356 ;
  assign n1953 = ~n1931 & ~n1937 ;
  assign n1954 = ~n1930 & ~n1953 ;
  assign n1955 = ~n1949 & n1954 ;
  assign n1956 = n1949 & ~n1954 ;
  assign n1957 = ~n1955 & ~n1956 ;
  assign n1960 = ~n1957 & ~x356 ;
  assign n1961 = ~n1959 & ~n1960 ;
  assign n1962 = ~n1946 & ~n1947 ;
  assign n1963 = ~n1948 & ~n1962 ;
  assign n1964 = ~x101 & ~x229 ;
  assign n1965 = x101 & x229 ;
  assign n1966 = ~n1964 & ~n1965 ;
  assign n1967 = n1963 & ~n1966 ;
  assign n1968 = ~n1963 & n1966 ;
  assign n1969 = ~n1967 & ~n1968 ;
  assign n1976 = n1969 & x357 ;
  assign n1970 = ~n1948 & ~n1954 ;
  assign n1971 = ~n1947 & ~n1970 ;
  assign n1972 = ~n1966 & n1971 ;
  assign n1973 = n1966 & ~n1971 ;
  assign n1974 = ~n1972 & ~n1973 ;
  assign n1977 = ~n1974 & ~x357 ;
  assign n1978 = ~n1976 & ~n1977 ;
  assign n1979 = ~n1963 & ~n1964 ;
  assign n1980 = ~n1965 & ~n1979 ;
  assign n1981 = ~x102 & ~x230 ;
  assign n1982 = x102 & x230 ;
  assign n1983 = ~n1981 & ~n1982 ;
  assign n1984 = n1980 & ~n1983 ;
  assign n1985 = ~n1980 & n1983 ;
  assign n1986 = ~n1984 & ~n1985 ;
  assign n1993 = n1986 & x358 ;
  assign n1987 = ~n1965 & ~n1971 ;
  assign n1988 = ~n1964 & ~n1987 ;
  assign n1989 = ~n1983 & n1988 ;
  assign n1990 = n1983 & ~n1988 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1994 = ~n1991 & ~x358 ;
  assign n1995 = ~n1993 & ~n1994 ;
  assign n1996 = ~n1980 & ~n1981 ;
  assign n1997 = ~n1982 & ~n1996 ;
  assign n1998 = ~x103 & ~x231 ;
  assign n1999 = x103 & x231 ;
  assign n2000 = ~n1998 & ~n1999 ;
  assign n2001 = n1997 & ~n2000 ;
  assign n2002 = ~n1997 & n2000 ;
  assign n2003 = ~n2001 & ~n2002 ;
  assign n2010 = n2003 & x359 ;
  assign n2004 = ~n1982 & ~n1988 ;
  assign n2005 = ~n1981 & ~n2004 ;
  assign n2006 = ~n2000 & n2005 ;
  assign n2007 = n2000 & ~n2005 ;
  assign n2008 = ~n2006 & ~n2007 ;
  assign n2011 = ~n2008 & ~x359 ;
  assign n2012 = ~n2010 & ~n2011 ;
  assign n2013 = ~n1997 & ~n1998 ;
  assign n2014 = ~n1999 & ~n2013 ;
  assign n2015 = ~x104 & ~x232 ;
  assign n2016 = x104 & x232 ;
  assign n2017 = ~n2015 & ~n2016 ;
  assign n2018 = n2014 & ~n2017 ;
  assign n2019 = ~n2014 & n2017 ;
  assign n2020 = ~n2018 & ~n2019 ;
  assign n2027 = n2020 & x360 ;
  assign n2021 = ~n1999 & ~n2005 ;
  assign n2022 = ~n1998 & ~n2021 ;
  assign n2023 = ~n2017 & n2022 ;
  assign n2024 = n2017 & ~n2022 ;
  assign n2025 = ~n2023 & ~n2024 ;
  assign n2028 = ~n2025 & ~x360 ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2030 = ~n2014 & ~n2015 ;
  assign n2031 = ~n2016 & ~n2030 ;
  assign n2032 = ~x105 & ~x233 ;
  assign n2033 = x105 & x233 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = n2031 & ~n2034 ;
  assign n2036 = ~n2031 & n2034 ;
  assign n2037 = ~n2035 & ~n2036 ;
  assign n2044 = n2037 & x361 ;
  assign n2038 = ~n2016 & ~n2022 ;
  assign n2039 = ~n2015 & ~n2038 ;
  assign n2040 = ~n2034 & n2039 ;
  assign n2041 = n2034 & ~n2039 ;
  assign n2042 = ~n2040 & ~n2041 ;
  assign n2045 = ~n2042 & ~x361 ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2047 = ~n2031 & ~n2032 ;
  assign n2048 = ~n2033 & ~n2047 ;
  assign n2049 = ~x106 & ~x234 ;
  assign n2050 = x106 & x234 ;
  assign n2051 = ~n2049 & ~n2050 ;
  assign n2052 = n2048 & ~n2051 ;
  assign n2053 = ~n2048 & n2051 ;
  assign n2054 = ~n2052 & ~n2053 ;
  assign n2061 = n2054 & x362 ;
  assign n2055 = ~n2033 & ~n2039 ;
  assign n2056 = ~n2032 & ~n2055 ;
  assign n2057 = ~n2051 & n2056 ;
  assign n2058 = n2051 & ~n2056 ;
  assign n2059 = ~n2057 & ~n2058 ;
  assign n2062 = ~n2059 & ~x362 ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = ~n2048 & ~n2049 ;
  assign n2065 = ~n2050 & ~n2064 ;
  assign n2066 = ~x107 & ~x235 ;
  assign n2067 = x107 & x235 ;
  assign n2068 = ~n2066 & ~n2067 ;
  assign n2069 = n2065 & ~n2068 ;
  assign n2070 = ~n2065 & n2068 ;
  assign n2071 = ~n2069 & ~n2070 ;
  assign n2078 = n2071 & x363 ;
  assign n2072 = ~n2050 & ~n2056 ;
  assign n2073 = ~n2049 & ~n2072 ;
  assign n2074 = ~n2068 & n2073 ;
  assign n2075 = n2068 & ~n2073 ;
  assign n2076 = ~n2074 & ~n2075 ;
  assign n2079 = ~n2076 & ~x363 ;
  assign n2080 = ~n2078 & ~n2079 ;
  assign n2081 = ~n2065 & ~n2066 ;
  assign n2082 = ~n2067 & ~n2081 ;
  assign n2083 = ~x108 & ~x236 ;
  assign n2084 = x108 & x236 ;
  assign n2085 = ~n2083 & ~n2084 ;
  assign n2086 = n2082 & ~n2085 ;
  assign n2087 = ~n2082 & n2085 ;
  assign n2088 = ~n2086 & ~n2087 ;
  assign n2095 = n2088 & x364 ;
  assign n2089 = ~n2067 & ~n2073 ;
  assign n2090 = ~n2066 & ~n2089 ;
  assign n2091 = ~n2085 & n2090 ;
  assign n2092 = n2085 & ~n2090 ;
  assign n2093 = ~n2091 & ~n2092 ;
  assign n2096 = ~n2093 & ~x364 ;
  assign n2097 = ~n2095 & ~n2096 ;
  assign n2098 = ~n2082 & ~n2083 ;
  assign n2099 = ~n2084 & ~n2098 ;
  assign n2100 = ~x109 & ~x237 ;
  assign n2101 = x109 & x237 ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = n2099 & ~n2102 ;
  assign n2104 = ~n2099 & n2102 ;
  assign n2105 = ~n2103 & ~n2104 ;
  assign n2112 = n2105 & x365 ;
  assign n2106 = ~n2084 & ~n2090 ;
  assign n2107 = ~n2083 & ~n2106 ;
  assign n2108 = ~n2102 & n2107 ;
  assign n2109 = n2102 & ~n2107 ;
  assign n2110 = ~n2108 & ~n2109 ;
  assign n2113 = ~n2110 & ~x365 ;
  assign n2114 = ~n2112 & ~n2113 ;
  assign n2115 = ~n2099 & ~n2100 ;
  assign n2116 = ~n2101 & ~n2115 ;
  assign n2117 = ~x110 & ~x238 ;
  assign n2118 = x110 & x238 ;
  assign n2119 = ~n2117 & ~n2118 ;
  assign n2120 = n2116 & ~n2119 ;
  assign n2121 = ~n2116 & n2119 ;
  assign n2122 = ~n2120 & ~n2121 ;
  assign n2129 = n2122 & x366 ;
  assign n2123 = ~n2101 & ~n2107 ;
  assign n2124 = ~n2100 & ~n2123 ;
  assign n2125 = ~n2119 & n2124 ;
  assign n2126 = n2119 & ~n2124 ;
  assign n2127 = ~n2125 & ~n2126 ;
  assign n2130 = ~n2127 & ~x366 ;
  assign n2131 = ~n2129 & ~n2130 ;
  assign n2132 = ~n2116 & ~n2117 ;
  assign n2133 = ~n2118 & ~n2132 ;
  assign n2134 = ~x111 & ~x239 ;
  assign n2135 = x111 & x239 ;
  assign n2136 = ~n2134 & ~n2135 ;
  assign n2137 = n2133 & ~n2136 ;
  assign n2138 = ~n2133 & n2136 ;
  assign n2139 = ~n2137 & ~n2138 ;
  assign n2146 = n2139 & x367 ;
  assign n2140 = ~n2118 & ~n2124 ;
  assign n2141 = ~n2117 & ~n2140 ;
  assign n2142 = ~n2136 & n2141 ;
  assign n2143 = n2136 & ~n2141 ;
  assign n2144 = ~n2142 & ~n2143 ;
  assign n2147 = ~n2144 & ~x367 ;
  assign n2148 = ~n2146 & ~n2147 ;
  assign n2149 = ~n2133 & ~n2134 ;
  assign n2150 = ~n2135 & ~n2149 ;
  assign n2151 = ~x112 & ~x240 ;
  assign n2152 = x112 & x240 ;
  assign n2153 = ~n2151 & ~n2152 ;
  assign n2154 = n2150 & ~n2153 ;
  assign n2155 = ~n2150 & n2153 ;
  assign n2156 = ~n2154 & ~n2155 ;
  assign n2163 = n2156 & x368 ;
  assign n2157 = ~n2135 & ~n2141 ;
  assign n2158 = ~n2134 & ~n2157 ;
  assign n2159 = ~n2153 & n2158 ;
  assign n2160 = n2153 & ~n2158 ;
  assign n2161 = ~n2159 & ~n2160 ;
  assign n2164 = ~n2161 & ~x368 ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2166 = ~n2150 & ~n2151 ;
  assign n2167 = ~n2152 & ~n2166 ;
  assign n2168 = ~x113 & ~x241 ;
  assign n2169 = x113 & x241 ;
  assign n2170 = ~n2168 & ~n2169 ;
  assign n2171 = n2167 & ~n2170 ;
  assign n2172 = ~n2167 & n2170 ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2180 = n2173 & x369 ;
  assign n2174 = ~n2152 & ~n2158 ;
  assign n2175 = ~n2151 & ~n2174 ;
  assign n2176 = ~n2170 & n2175 ;
  assign n2177 = n2170 & ~n2175 ;
  assign n2178 = ~n2176 & ~n2177 ;
  assign n2181 = ~n2178 & ~x369 ;
  assign n2182 = ~n2180 & ~n2181 ;
  assign n2183 = ~n2167 & ~n2168 ;
  assign n2184 = ~n2169 & ~n2183 ;
  assign n2185 = ~x114 & ~x242 ;
  assign n2186 = x114 & x242 ;
  assign n2187 = ~n2185 & ~n2186 ;
  assign n2188 = n2184 & ~n2187 ;
  assign n2189 = ~n2184 & n2187 ;
  assign n2190 = ~n2188 & ~n2189 ;
  assign n2197 = n2190 & x370 ;
  assign n2191 = ~n2169 & ~n2175 ;
  assign n2192 = ~n2168 & ~n2191 ;
  assign n2193 = ~n2187 & n2192 ;
  assign n2194 = n2187 & ~n2192 ;
  assign n2195 = ~n2193 & ~n2194 ;
  assign n2198 = ~n2195 & ~x370 ;
  assign n2199 = ~n2197 & ~n2198 ;
  assign n2200 = ~n2184 & ~n2185 ;
  assign n2201 = ~n2186 & ~n2200 ;
  assign n2202 = ~x115 & ~x243 ;
  assign n2203 = x115 & x243 ;
  assign n2204 = ~n2202 & ~n2203 ;
  assign n2205 = n2201 & ~n2204 ;
  assign n2206 = ~n2201 & n2204 ;
  assign n2207 = ~n2205 & ~n2206 ;
  assign n2214 = n2207 & x371 ;
  assign n2208 = ~n2186 & ~n2192 ;
  assign n2209 = ~n2185 & ~n2208 ;
  assign n2210 = ~n2204 & n2209 ;
  assign n2211 = n2204 & ~n2209 ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2215 = ~n2212 & ~x371 ;
  assign n2216 = ~n2214 & ~n2215 ;
  assign n2217 = ~n2201 & ~n2202 ;
  assign n2218 = ~n2203 & ~n2217 ;
  assign n2219 = ~x116 & ~x244 ;
  assign n2220 = x116 & x244 ;
  assign n2221 = ~n2219 & ~n2220 ;
  assign n2222 = n2218 & ~n2221 ;
  assign n2223 = ~n2218 & n2221 ;
  assign n2224 = ~n2222 & ~n2223 ;
  assign n2231 = n2224 & x372 ;
  assign n2225 = ~n2203 & ~n2209 ;
  assign n2226 = ~n2202 & ~n2225 ;
  assign n2227 = ~n2221 & n2226 ;
  assign n2228 = n2221 & ~n2226 ;
  assign n2229 = ~n2227 & ~n2228 ;
  assign n2232 = ~n2229 & ~x372 ;
  assign n2233 = ~n2231 & ~n2232 ;
  assign n2234 = ~n2218 & ~n2219 ;
  assign n2235 = ~n2220 & ~n2234 ;
  assign n2236 = ~x117 & ~x245 ;
  assign n2237 = x117 & x245 ;
  assign n2238 = ~n2236 & ~n2237 ;
  assign n2239 = n2235 & ~n2238 ;
  assign n2240 = ~n2235 & n2238 ;
  assign n2241 = ~n2239 & ~n2240 ;
  assign n2248 = n2241 & x373 ;
  assign n2242 = ~n2220 & ~n2226 ;
  assign n2243 = ~n2219 & ~n2242 ;
  assign n2244 = ~n2238 & n2243 ;
  assign n2245 = n2238 & ~n2243 ;
  assign n2246 = ~n2244 & ~n2245 ;
  assign n2249 = ~n2246 & ~x373 ;
  assign n2250 = ~n2248 & ~n2249 ;
  assign n2251 = ~n2235 & ~n2236 ;
  assign n2252 = ~n2237 & ~n2251 ;
  assign n2253 = ~x118 & ~x246 ;
  assign n2254 = x118 & x246 ;
  assign n2255 = ~n2253 & ~n2254 ;
  assign n2256 = n2252 & ~n2255 ;
  assign n2257 = ~n2252 & n2255 ;
  assign n2258 = ~n2256 & ~n2257 ;
  assign n2265 = n2258 & x374 ;
  assign n2259 = ~n2237 & ~n2243 ;
  assign n2260 = ~n2236 & ~n2259 ;
  assign n2261 = ~n2255 & n2260 ;
  assign n2262 = n2255 & ~n2260 ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2266 = ~n2263 & ~x374 ;
  assign n2267 = ~n2265 & ~n2266 ;
  assign n2268 = ~n2252 & ~n2253 ;
  assign n2269 = ~n2254 & ~n2268 ;
  assign n2270 = ~x119 & ~x247 ;
  assign n2271 = x119 & x247 ;
  assign n2272 = ~n2270 & ~n2271 ;
  assign n2273 = n2269 & ~n2272 ;
  assign n2274 = ~n2269 & n2272 ;
  assign n2275 = ~n2273 & ~n2274 ;
  assign n2282 = n2275 & x375 ;
  assign n2276 = ~n2254 & ~n2260 ;
  assign n2277 = ~n2253 & ~n2276 ;
  assign n2278 = ~n2272 & n2277 ;
  assign n2279 = n2272 & ~n2277 ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2283 = ~n2280 & ~x375 ;
  assign n2284 = ~n2282 & ~n2283 ;
  assign n2285 = ~n2269 & ~n2270 ;
  assign n2286 = ~n2271 & ~n2285 ;
  assign n2287 = ~x120 & ~x248 ;
  assign n2288 = x120 & x248 ;
  assign n2289 = ~n2287 & ~n2288 ;
  assign n2290 = n2286 & ~n2289 ;
  assign n2291 = ~n2286 & n2289 ;
  assign n2292 = ~n2290 & ~n2291 ;
  assign n2299 = n2292 & x376 ;
  assign n2293 = ~n2271 & ~n2277 ;
  assign n2294 = ~n2270 & ~n2293 ;
  assign n2295 = ~n2289 & n2294 ;
  assign n2296 = n2289 & ~n2294 ;
  assign n2297 = ~n2295 & ~n2296 ;
  assign n2300 = ~n2297 & ~x376 ;
  assign n2301 = ~n2299 & ~n2300 ;
  assign n2302 = ~n2286 & ~n2287 ;
  assign n2303 = ~n2288 & ~n2302 ;
  assign n2304 = ~x121 & ~x249 ;
  assign n2305 = x121 & x249 ;
  assign n2306 = ~n2304 & ~n2305 ;
  assign n2307 = n2303 & ~n2306 ;
  assign n2308 = ~n2303 & n2306 ;
  assign n2309 = ~n2307 & ~n2308 ;
  assign n2316 = n2309 & x377 ;
  assign n2310 = ~n2288 & ~n2294 ;
  assign n2311 = ~n2287 & ~n2310 ;
  assign n2312 = ~n2306 & n2311 ;
  assign n2313 = n2306 & ~n2311 ;
  assign n2314 = ~n2312 & ~n2313 ;
  assign n2317 = ~n2314 & ~x377 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = ~n2303 & ~n2304 ;
  assign n2320 = ~n2305 & ~n2319 ;
  assign n2321 = ~x122 & ~x250 ;
  assign n2322 = x122 & x250 ;
  assign n2323 = ~n2321 & ~n2322 ;
  assign n2324 = n2320 & ~n2323 ;
  assign n2325 = ~n2320 & n2323 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2333 = n2326 & x378 ;
  assign n2327 = ~n2305 & ~n2311 ;
  assign n2328 = ~n2304 & ~n2327 ;
  assign n2329 = ~n2323 & n2328 ;
  assign n2330 = n2323 & ~n2328 ;
  assign n2331 = ~n2329 & ~n2330 ;
  assign n2334 = ~n2331 & ~x378 ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = ~n2320 & ~n2321 ;
  assign n2337 = ~n2322 & ~n2336 ;
  assign n2338 = ~x123 & ~x251 ;
  assign n2339 = x123 & x251 ;
  assign n2340 = ~n2338 & ~n2339 ;
  assign n2341 = n2337 & ~n2340 ;
  assign n2342 = ~n2337 & n2340 ;
  assign n2343 = ~n2341 & ~n2342 ;
  assign n2350 = n2343 & x379 ;
  assign n2344 = ~n2322 & ~n2328 ;
  assign n2345 = ~n2321 & ~n2344 ;
  assign n2346 = ~n2340 & n2345 ;
  assign n2347 = n2340 & ~n2345 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2351 = ~n2348 & ~x379 ;
  assign n2352 = ~n2350 & ~n2351 ;
  assign n2353 = ~n2337 & ~n2338 ;
  assign n2354 = ~n2339 & ~n2353 ;
  assign n2355 = ~x124 & ~x252 ;
  assign n2356 = x124 & x252 ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = n2354 & ~n2357 ;
  assign n2359 = ~n2354 & n2357 ;
  assign n2360 = ~n2358 & ~n2359 ;
  assign n2367 = n2360 & x380 ;
  assign n2361 = ~n2339 & ~n2345 ;
  assign n2362 = ~n2338 & ~n2361 ;
  assign n2363 = ~n2357 & n2362 ;
  assign n2364 = n2357 & ~n2362 ;
  assign n2365 = ~n2363 & ~n2364 ;
  assign n2368 = ~n2365 & ~x380 ;
  assign n2369 = ~n2367 & ~n2368 ;
  assign n2370 = ~n2354 & ~n2355 ;
  assign n2371 = ~n2356 & ~n2370 ;
  assign n2372 = ~x125 & ~x253 ;
  assign n2373 = x125 & x253 ;
  assign n2374 = ~n2372 & ~n2373 ;
  assign n2375 = n2371 & ~n2374 ;
  assign n2376 = ~n2371 & n2374 ;
  assign n2377 = ~n2375 & ~n2376 ;
  assign n2384 = n2377 & x381 ;
  assign n2378 = ~n2356 & ~n2362 ;
  assign n2379 = ~n2355 & ~n2378 ;
  assign n2380 = ~n2374 & n2379 ;
  assign n2381 = n2374 & ~n2379 ;
  assign n2382 = ~n2380 & ~n2381 ;
  assign n2385 = ~n2382 & ~x381 ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2387 = ~n2371 & ~n2372 ;
  assign n2388 = ~n2373 & ~n2387 ;
  assign n2389 = ~x126 & ~x254 ;
  assign n2390 = x126 & x254 ;
  assign n2391 = ~n2389 & ~n2390 ;
  assign n2392 = n2388 & ~n2391 ;
  assign n2393 = ~n2388 & n2391 ;
  assign n2394 = ~n2392 & ~n2393 ;
  assign n2401 = n2394 & x382 ;
  assign n2395 = ~n2373 & ~n2379 ;
  assign n2396 = ~n2372 & ~n2395 ;
  assign n2397 = ~n2391 & n2396 ;
  assign n2398 = n2391 & ~n2396 ;
  assign n2399 = ~n2397 & ~n2398 ;
  assign n2402 = ~n2399 & ~x382 ;
  assign n2403 = ~n2401 & ~n2402 ;
  assign n2404 = ~n2388 & ~n2389 ;
  assign n2405 = ~n2390 & ~n2404 ;
  assign n2406 = ~x127 & ~x255 ;
  assign n2407 = x127 & x255 ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = n2405 & ~n2408 ;
  assign n2410 = ~n2405 & n2408 ;
  assign n2411 = ~n2409 & ~n2410 ;
  assign n2418 = n2411 & x383 ;
  assign n2412 = ~n2390 & ~n2396 ;
  assign n2413 = ~n2389 & ~n2412 ;
  assign n2414 = ~n2408 & n2413 ;
  assign n2415 = n2408 & ~n2413 ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2419 = ~n2416 & ~x383 ;
  assign n2420 = ~n2418 & ~n2419 ;
  assign n2421 = ~n2405 & ~n2406 ;
  assign n2422 = ~n2407 & ~n2421 ;
  assign n2426 = ~n2422 & x384 ;
  assign n2423 = ~n2407 & ~n2413 ;
  assign n2424 = ~n2406 & ~n2423 ;
  assign n2427 = n2424 & ~x384 ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign y0 = ~n263 ;
  assign y1 = ~n278 ;
  assign y2 = ~n295 ;
  assign y3 = ~n312 ;
  assign y4 = ~n329 ;
  assign y5 = ~n346 ;
  assign y6 = ~n363 ;
  assign y7 = ~n380 ;
  assign y8 = ~n397 ;
  assign y9 = ~n414 ;
  assign y10 = ~n431 ;
  assign y11 = ~n448 ;
  assign y12 = ~n465 ;
  assign y13 = ~n482 ;
  assign y14 = ~n499 ;
  assign y15 = ~n516 ;
  assign y16 = ~n533 ;
  assign y17 = ~n550 ;
  assign y18 = ~n567 ;
  assign y19 = ~n584 ;
  assign y20 = ~n601 ;
  assign y21 = ~n618 ;
  assign y22 = ~n635 ;
  assign y23 = ~n652 ;
  assign y24 = ~n669 ;
  assign y25 = ~n686 ;
  assign y26 = ~n703 ;
  assign y27 = ~n720 ;
  assign y28 = ~n737 ;
  assign y29 = ~n754 ;
  assign y30 = ~n771 ;
  assign y31 = ~n788 ;
  assign y32 = ~n805 ;
  assign y33 = ~n822 ;
  assign y34 = ~n839 ;
  assign y35 = ~n856 ;
  assign y36 = ~n873 ;
  assign y37 = ~n890 ;
  assign y38 = ~n907 ;
  assign y39 = ~n924 ;
  assign y40 = ~n941 ;
  assign y41 = ~n958 ;
  assign y42 = ~n975 ;
  assign y43 = ~n992 ;
  assign y44 = ~n1009 ;
  assign y45 = ~n1026 ;
  assign y46 = ~n1043 ;
  assign y47 = ~n1060 ;
  assign y48 = ~n1077 ;
  assign y49 = ~n1094 ;
  assign y50 = ~n1111 ;
  assign y51 = ~n1128 ;
  assign y52 = ~n1145 ;
  assign y53 = ~n1162 ;
  assign y54 = ~n1179 ;
  assign y55 = ~n1196 ;
  assign y56 = ~n1213 ;
  assign y57 = ~n1230 ;
  assign y58 = ~n1247 ;
  assign y59 = ~n1264 ;
  assign y60 = ~n1281 ;
  assign y61 = ~n1298 ;
  assign y62 = ~n1315 ;
  assign y63 = ~n1332 ;
  assign y64 = ~n1349 ;
  assign y65 = ~n1366 ;
  assign y66 = ~n1383 ;
  assign y67 = ~n1400 ;
  assign y68 = ~n1417 ;
  assign y69 = ~n1434 ;
  assign y70 = ~n1451 ;
  assign y71 = ~n1468 ;
  assign y72 = ~n1485 ;
  assign y73 = ~n1502 ;
  assign y74 = ~n1519 ;
  assign y75 = ~n1536 ;
  assign y76 = ~n1553 ;
  assign y77 = ~n1570 ;
  assign y78 = ~n1587 ;
  assign y79 = ~n1604 ;
  assign y80 = ~n1621 ;
  assign y81 = ~n1638 ;
  assign y82 = ~n1655 ;
  assign y83 = ~n1672 ;
  assign y84 = ~n1689 ;
  assign y85 = ~n1706 ;
  assign y86 = ~n1723 ;
  assign y87 = ~n1740 ;
  assign y88 = ~n1757 ;
  assign y89 = ~n1774 ;
  assign y90 = ~n1791 ;
  assign y91 = ~n1808 ;
  assign y92 = ~n1825 ;
  assign y93 = ~n1842 ;
  assign y94 = ~n1859 ;
  assign y95 = ~n1876 ;
  assign y96 = ~n1893 ;
  assign y97 = ~n1910 ;
  assign y98 = ~n1927 ;
  assign y99 = ~n1944 ;
  assign y100 = ~n1961 ;
  assign y101 = ~n1978 ;
  assign y102 = ~n1995 ;
  assign y103 = ~n2012 ;
  assign y104 = ~n2029 ;
  assign y105 = ~n2046 ;
  assign y106 = ~n2063 ;
  assign y107 = ~n2080 ;
  assign y108 = ~n2097 ;
  assign y109 = ~n2114 ;
  assign y110 = ~n2131 ;
  assign y111 = ~n2148 ;
  assign y112 = ~n2165 ;
  assign y113 = ~n2182 ;
  assign y114 = ~n2199 ;
  assign y115 = ~n2216 ;
  assign y116 = ~n2233 ;
  assign y117 = ~n2250 ;
  assign y118 = ~n2267 ;
  assign y119 = ~n2284 ;
  assign y120 = ~n2301 ;
  assign y121 = ~n2318 ;
  assign y122 = ~n2335 ;
  assign y123 = ~n2352 ;
  assign y124 = ~n2369 ;
  assign y125 = ~n2386 ;
  assign y126 = ~n2403 ;
  assign y127 = ~n2420 ;
  assign y128 = ~n2428 ;
endmodule
