module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 ;
  assign n256 = ( x67 & ~x94 ) | ( x67 & x234 ) | ( ~x94 & x234 ) ;
  assign n259 = x208 ^ x187 ^ x184 ;
  assign n258 = ( x26 & ~x30 ) | ( x26 & x120 ) | ( ~x30 & x120 ) ;
  assign n257 = ( x17 & ~x77 ) | ( x17 & x191 ) | ( ~x77 & x191 ) ;
  assign n260 = n259 ^ n258 ^ n257 ;
  assign n261 = ( ~x17 & x72 ) | ( ~x17 & x194 ) | ( x72 & x194 ) ;
  assign n262 = n261 ^ n260 ^ x118 ;
  assign n263 = n262 ^ x185 ^ x175 ;
  assign n264 = x73 & ~x98 ;
  assign n265 = n264 ^ x228 ^ x44 ;
  assign n266 = x139 ^ x105 ^ 1'b0 ;
  assign n267 = x15 & x95 ;
  assign n268 = ~x252 & n267 ;
  assign n269 = ( x32 & ~x101 ) | ( x32 & n268 ) | ( ~x101 & n268 ) ;
  assign n270 = x222 & ~n269 ;
  assign n271 = ~n266 & n270 ;
  assign n273 = x236 ^ x210 ^ x68 ;
  assign n274 = n273 ^ x153 ^ x26 ;
  assign n272 = ( ~x42 & x54 ) | ( ~x42 & x158 ) | ( x54 & x158 ) ;
  assign n275 = n274 ^ n272 ^ x70 ;
  assign n276 = x205 ^ x118 ^ x1 ;
  assign n277 = x105 ^ x60 ^ x40 ;
  assign n278 = ( x41 & x83 ) | ( x41 & n277 ) | ( x83 & n277 ) ;
  assign n279 = x18 ^ x4 ^ 1'b0 ;
  assign n280 = x147 & n279 ;
  assign n281 = ( x29 & x142 ) | ( x29 & ~n280 ) | ( x142 & ~n280 ) ;
  assign n282 = n281 ^ x177 ^ x8 ;
  assign n283 = n282 ^ x234 ^ x1 ;
  assign n284 = ( x6 & x179 ) | ( x6 & n275 ) | ( x179 & n275 ) ;
  assign n285 = x204 ^ x179 ^ x175 ;
  assign n286 = ( x119 & x173 ) | ( x119 & ~n280 ) | ( x173 & ~n280 ) ;
  assign n287 = ( x1 & x19 ) | ( x1 & ~x219 ) | ( x19 & ~x219 ) ;
  assign n288 = n287 ^ x188 ^ x154 ;
  assign n289 = n288 ^ x199 ^ x196 ;
  assign n290 = ( ~x45 & n286 ) | ( ~x45 & n289 ) | ( n286 & n289 ) ;
  assign n291 = n290 ^ x85 ^ x54 ;
  assign n292 = ( x20 & ~x76 ) | ( x20 & x90 ) | ( ~x76 & x90 ) ;
  assign n293 = ( x174 & ~x186 ) | ( x174 & n269 ) | ( ~x186 & n269 ) ;
  assign n294 = ( x109 & ~n292 ) | ( x109 & n293 ) | ( ~n292 & n293 ) ;
  assign n295 = ( x88 & x221 ) | ( x88 & ~x236 ) | ( x221 & ~x236 ) ;
  assign n296 = ( x12 & ~x250 ) | ( x12 & n287 ) | ( ~x250 & n287 ) ;
  assign n297 = ( x184 & n295 ) | ( x184 & ~n296 ) | ( n295 & ~n296 ) ;
  assign n298 = x226 ^ x177 ^ x141 ;
  assign n299 = ( x84 & ~x165 ) | ( x84 & n298 ) | ( ~x165 & n298 ) ;
  assign n300 = n299 ^ x232 ^ 1'b0 ;
  assign n301 = n300 ^ x34 ^ x3 ;
  assign n303 = ( x188 & ~x212 ) | ( x188 & x248 ) | ( ~x212 & x248 ) ;
  assign n302 = x218 ^ x176 ^ x93 ;
  assign n304 = n303 ^ n302 ^ n275 ;
  assign n305 = n304 ^ x205 ^ x87 ;
  assign n306 = ( x73 & ~x109 ) | ( x73 & x149 ) | ( ~x109 & x149 ) ;
  assign n307 = x247 ^ x181 ^ 1'b0 ;
  assign n308 = n306 & n307 ;
  assign n309 = x138 ^ x97 ^ x65 ;
  assign n310 = n309 ^ x63 ^ x61 ;
  assign n311 = ( x217 & n308 ) | ( x217 & ~n310 ) | ( n308 & ~n310 ) ;
  assign n312 = ( x70 & x134 ) | ( x70 & ~x254 ) | ( x134 & ~x254 ) ;
  assign n313 = ~x118 & x138 ;
  assign n314 = ( x71 & ~n312 ) | ( x71 & n313 ) | ( ~n312 & n313 ) ;
  assign n315 = x152 ^ x78 ^ x46 ;
  assign n316 = n256 ^ x26 ^ 1'b0 ;
  assign n317 = x0 & n316 ;
  assign n318 = ( x55 & n315 ) | ( x55 & ~n317 ) | ( n315 & ~n317 ) ;
  assign n319 = n318 ^ x133 ^ 1'b0 ;
  assign n324 = ( x15 & x66 ) | ( x15 & ~x176 ) | ( x66 & ~x176 ) ;
  assign n322 = ( x15 & ~x204 ) | ( x15 & x209 ) | ( ~x204 & x209 ) ;
  assign n320 = x252 ^ x112 ^ x111 ;
  assign n321 = n320 ^ x142 ^ x61 ;
  assign n323 = n322 ^ n321 ^ x98 ;
  assign n325 = n324 ^ n323 ^ x116 ;
  assign n328 = x185 ^ x173 ^ x100 ;
  assign n327 = ( ~x7 & x147 ) | ( ~x7 & x196 ) | ( x147 & x196 ) ;
  assign n329 = n328 ^ n327 ^ x205 ;
  assign n330 = x190 ^ x106 ^ 1'b0 ;
  assign n331 = n329 & n330 ;
  assign n326 = ( x214 & ~x230 ) | ( x214 & n275 ) | ( ~x230 & n275 ) ;
  assign n332 = n331 ^ n326 ^ x115 ;
  assign n333 = n266 ^ x250 ^ x15 ;
  assign n334 = n333 ^ x238 ^ x73 ;
  assign n335 = ( n257 & n259 ) | ( n257 & n334 ) | ( n259 & n334 ) ;
  assign n336 = n335 ^ x205 ^ x50 ;
  assign n337 = ( x12 & x27 ) | ( x12 & ~x130 ) | ( x27 & ~x130 ) ;
  assign n338 = ( ~x164 & x218 ) | ( ~x164 & n337 ) | ( x218 & n337 ) ;
  assign n339 = x229 ^ x16 ^ x13 ;
  assign n340 = ( x5 & x125 ) | ( x5 & ~x233 ) | ( x125 & ~x233 ) ;
  assign n341 = n340 ^ x179 ^ x109 ;
  assign n342 = ( x136 & n339 ) | ( x136 & ~n341 ) | ( n339 & ~n341 ) ;
  assign n343 = x101 ^ x94 ^ x72 ;
  assign n345 = ( ~x16 & x160 ) | ( ~x16 & x226 ) | ( x160 & x226 ) ;
  assign n344 = x48 & x124 ;
  assign n346 = n345 ^ n344 ^ 1'b0 ;
  assign n347 = ( x174 & n343 ) | ( x174 & ~n346 ) | ( n343 & ~n346 ) ;
  assign n348 = x197 & n258 ;
  assign n349 = n348 ^ x10 ^ 1'b0 ;
  assign n352 = ( x154 & x195 ) | ( x154 & ~x242 ) | ( x195 & ~x242 ) ;
  assign n350 = x189 ^ x55 ^ x36 ;
  assign n351 = ( n260 & ~n277 ) | ( n260 & n350 ) | ( ~n277 & n350 ) ;
  assign n353 = n352 ^ n351 ^ 1'b0 ;
  assign n354 = x134 & n353 ;
  assign n357 = ( x21 & x202 ) | ( x21 & n275 ) | ( x202 & n275 ) ;
  assign n355 = ( x105 & ~x108 ) | ( x105 & x135 ) | ( ~x108 & x135 ) ;
  assign n356 = ( x36 & ~n327 ) | ( x36 & n355 ) | ( ~n327 & n355 ) ;
  assign n358 = n357 ^ n356 ^ n322 ;
  assign n363 = ( x76 & ~x147 ) | ( x76 & x235 ) | ( ~x147 & x235 ) ;
  assign n364 = ( ~x3 & x64 ) | ( ~x3 & n363 ) | ( x64 & n363 ) ;
  assign n359 = x241 ^ x186 ^ x22 ;
  assign n360 = n359 ^ n259 ^ x245 ;
  assign n361 = ( x102 & ~x153 ) | ( x102 & n359 ) | ( ~x153 & n359 ) ;
  assign n362 = ( x234 & n360 ) | ( x234 & n361 ) | ( n360 & n361 ) ;
  assign n365 = n364 ^ n362 ^ x47 ;
  assign n366 = x31 & x179 ;
  assign n367 = n366 ^ x202 ^ 1'b0 ;
  assign n368 = n367 ^ x237 ^ x98 ;
  assign n369 = n362 ^ x53 ^ x50 ;
  assign n370 = n369 ^ x120 ^ x49 ;
  assign n371 = ( x101 & ~x224 ) | ( x101 & n370 ) | ( ~x224 & n370 ) ;
  assign n372 = ( ~x69 & x209 ) | ( ~x69 & n371 ) | ( x209 & n371 ) ;
  assign n373 = x192 ^ x30 ^ 1'b0 ;
  assign n374 = ~n269 & n373 ;
  assign n375 = ( x121 & n333 ) | ( x121 & n334 ) | ( n333 & n334 ) ;
  assign n376 = x213 ^ x180 ^ x137 ;
  assign n377 = ( x88 & ~x123 ) | ( x88 & x240 ) | ( ~x123 & x240 ) ;
  assign n378 = x203 ^ x81 ^ x74 ;
  assign n379 = n378 ^ x98 ^ x27 ;
  assign n380 = ( ~x209 & n362 ) | ( ~x209 & n379 ) | ( n362 & n379 ) ;
  assign n381 = n377 & ~n380 ;
  assign n382 = n381 ^ n265 ^ 1'b0 ;
  assign n385 = x99 & x109 ;
  assign n386 = ~x156 & n385 ;
  assign n383 = x43 ^ x25 ^ x11 ;
  assign n384 = ( x232 & ~x235 ) | ( x232 & n383 ) | ( ~x235 & n383 ) ;
  assign n387 = n386 ^ n384 ^ x35 ;
  assign n396 = n287 ^ x233 ^ x77 ;
  assign n391 = ( x118 & ~x145 ) | ( x118 & n287 ) | ( ~x145 & n287 ) ;
  assign n392 = x211 ^ x52 ^ 1'b0 ;
  assign n393 = x192 & n392 ;
  assign n394 = ( x196 & n391 ) | ( x196 & ~n393 ) | ( n391 & ~n393 ) ;
  assign n388 = ( ~n303 & n308 ) | ( ~n303 & n322 ) | ( n308 & n322 ) ;
  assign n389 = ( ~x35 & x98 ) | ( ~x35 & n388 ) | ( x98 & n388 ) ;
  assign n390 = x235 & n389 ;
  assign n395 = n394 ^ n390 ^ 1'b0 ;
  assign n397 = n396 ^ n395 ^ n261 ;
  assign n398 = n322 ^ n309 ^ x131 ;
  assign n399 = ( ~x238 & n397 ) | ( ~x238 & n398 ) | ( n397 & n398 ) ;
  assign n400 = ( x202 & n311 ) | ( x202 & n399 ) | ( n311 & n399 ) ;
  assign n401 = ( x24 & ~x163 ) | ( x24 & x223 ) | ( ~x163 & x223 ) ;
  assign n402 = n401 ^ n265 ^ n259 ;
  assign n403 = ( ~x115 & x171 ) | ( ~x115 & n402 ) | ( x171 & n402 ) ;
  assign n414 = ( ~x159 & x188 ) | ( ~x159 & x229 ) | ( x188 & x229 ) ;
  assign n408 = x188 & ~n343 ;
  assign n409 = n408 ^ x209 ^ 1'b0 ;
  assign n410 = n409 ^ n277 ^ x227 ;
  assign n405 = x61 ^ x44 ^ 1'b0 ;
  assign n406 = x130 & n405 ;
  assign n407 = ( ~x78 & x198 ) | ( ~x78 & n406 ) | ( x198 & n406 ) ;
  assign n404 = n351 ^ n294 ^ x14 ;
  assign n411 = n410 ^ n407 ^ n404 ;
  assign n412 = x11 & n411 ;
  assign n413 = n412 ^ x231 ^ 1'b0 ;
  assign n415 = n414 ^ n413 ^ x1 ;
  assign n416 = x237 ^ x219 ^ x33 ;
  assign n417 = ( ~x45 & x238 ) | ( ~x45 & x245 ) | ( x238 & x245 ) ;
  assign n418 = n417 ^ x182 ^ x109 ;
  assign n419 = ( ~x23 & x240 ) | ( ~x23 & n418 ) | ( x240 & n418 ) ;
  assign n420 = ( x157 & ~x218 ) | ( x157 & n419 ) | ( ~x218 & n419 ) ;
  assign n421 = ( x3 & x248 ) | ( x3 & ~n389 ) | ( x248 & ~n389 ) ;
  assign n422 = n421 ^ x196 ^ x118 ;
  assign n423 = ( x167 & n420 ) | ( x167 & n422 ) | ( n420 & n422 ) ;
  assign n424 = x228 ^ x53 ^ x45 ;
  assign n425 = x227 & ~n424 ;
  assign n426 = ~x158 & n425 ;
  assign n427 = x254 ^ x201 ^ x63 ;
  assign n428 = n427 ^ x144 ^ x80 ;
  assign n429 = n428 ^ n298 ^ n277 ;
  assign n430 = ( x5 & x223 ) | ( x5 & n429 ) | ( x223 & n429 ) ;
  assign n431 = x217 ^ x172 ^ x75 ;
  assign n432 = n258 ^ x193 ^ 1'b0 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = ( ~x123 & x156 ) | ( ~x123 & n433 ) | ( x156 & n433 ) ;
  assign n435 = ( n426 & n430 ) | ( n426 & n434 ) | ( n430 & n434 ) ;
  assign n436 = n435 ^ n404 ^ x73 ;
  assign n437 = ( n416 & ~n423 ) | ( n416 & n436 ) | ( ~n423 & n436 ) ;
  assign n438 = ( ~x52 & x118 ) | ( ~x52 & x131 ) | ( x118 & x131 ) ;
  assign n439 = n438 ^ x27 ^ 1'b0 ;
  assign n443 = x199 & x205 ;
  assign n444 = n443 ^ x158 ^ 1'b0 ;
  assign n441 = x17 & x85 ;
  assign n442 = n441 ^ x131 ^ 1'b0 ;
  assign n445 = n444 ^ n442 ^ x0 ;
  assign n440 = n331 ^ x207 ^ x160 ;
  assign n446 = n445 ^ n440 ^ n356 ;
  assign n447 = n439 & ~n446 ;
  assign n448 = n362 & n447 ;
  assign n452 = ( x57 & ~x219 ) | ( x57 & n363 ) | ( ~x219 & n363 ) ;
  assign n449 = n308 ^ x138 ^ x6 ;
  assign n450 = n449 ^ n293 ^ x219 ;
  assign n451 = n450 ^ n406 ^ x27 ;
  assign n453 = n452 ^ n451 ^ x171 ;
  assign n454 = n453 ^ n309 ^ x68 ;
  assign n455 = n277 ^ x109 ^ 1'b0 ;
  assign n456 = x37 & ~n455 ;
  assign n457 = ( x32 & x70 ) | ( x32 & ~n456 ) | ( x70 & ~n456 ) ;
  assign n458 = x197 & x246 ;
  assign n459 = ~x176 & n458 ;
  assign n460 = n459 ^ n421 ^ x108 ;
  assign n461 = ( x179 & n305 ) | ( x179 & ~n460 ) | ( n305 & ~n460 ) ;
  assign n462 = n461 ^ n423 ^ x148 ;
  assign n463 = ( n352 & ~n457 ) | ( n352 & n462 ) | ( ~n457 & n462 ) ;
  assign n465 = ( n321 & n329 ) | ( n321 & ~n428 ) | ( n329 & ~n428 ) ;
  assign n464 = x171 & ~n299 ;
  assign n466 = n465 ^ n464 ^ x207 ;
  assign n467 = n449 ^ n442 ^ n393 ;
  assign n468 = n467 ^ x249 ^ 1'b0 ;
  assign n476 = n401 ^ x156 ^ x106 ;
  assign n477 = n476 ^ n439 ^ x64 ;
  assign n471 = ( x94 & x118 ) | ( x94 & ~n297 ) | ( x118 & ~n297 ) ;
  assign n472 = ~n450 & n471 ;
  assign n473 = n391 ^ x110 ^ x74 ;
  assign n474 = x224 & ~n473 ;
  assign n475 = ~n472 & n474 ;
  assign n469 = n266 ^ x250 ^ x10 ;
  assign n470 = n469 ^ x96 ^ x43 ;
  assign n478 = n477 ^ n475 ^ n470 ;
  assign n479 = n321 ^ x117 ^ 1'b0 ;
  assign n480 = ( x74 & x192 ) | ( x74 & ~n479 ) | ( x192 & ~n479 ) ;
  assign n482 = ( x61 & x101 ) | ( x61 & ~x239 ) | ( x101 & ~x239 ) ;
  assign n481 = ( ~x105 & n278 ) | ( ~x105 & n359 ) | ( n278 & n359 ) ;
  assign n483 = n482 ^ n481 ^ x124 ;
  assign n484 = n483 ^ n438 ^ n260 ;
  assign n485 = n484 ^ n312 ^ 1'b0 ;
  assign n486 = ( x50 & x59 ) | ( x50 & ~x118 ) | ( x59 & ~x118 ) ;
  assign n487 = ( ~x206 & x245 ) | ( ~x206 & n486 ) | ( x245 & n486 ) ;
  assign n488 = ( ~n378 & n382 ) | ( ~n378 & n487 ) | ( n382 & n487 ) ;
  assign n489 = n488 ^ n305 ^ x107 ;
  assign n490 = x222 ^ x102 ^ 1'b0 ;
  assign n491 = ( x15 & ~x148 ) | ( x15 & x219 ) | ( ~x148 & x219 ) ;
  assign n492 = n491 ^ n302 ^ 1'b0 ;
  assign n493 = n490 & ~n492 ;
  assign n494 = ( ~x167 & x209 ) | ( ~x167 & n320 ) | ( x209 & n320 ) ;
  assign n495 = ( ~n304 & n444 ) | ( ~n304 & n494 ) | ( n444 & n494 ) ;
  assign n496 = n495 ^ n371 ^ x32 ;
  assign n497 = ( x253 & n493 ) | ( x253 & n496 ) | ( n493 & n496 ) ;
  assign n498 = ( x57 & ~x96 ) | ( x57 & n262 ) | ( ~x96 & n262 ) ;
  assign n499 = n388 ^ n289 ^ x154 ;
  assign n500 = ( x233 & ~n498 ) | ( x233 & n499 ) | ( ~n498 & n499 ) ;
  assign n501 = n500 ^ n488 ^ n340 ;
  assign n502 = ( x7 & ~x147 ) | ( x7 & n431 ) | ( ~x147 & n431 ) ;
  assign n503 = x161 & n389 ;
  assign n504 = n502 & n503 ;
  assign n505 = x224 ^ x222 ^ x135 ;
  assign n506 = n505 ^ n343 ^ x103 ;
  assign n507 = n506 ^ n427 ^ 1'b0 ;
  assign n508 = ( ~x139 & n295 ) | ( ~x139 & n355 ) | ( n295 & n355 ) ;
  assign n509 = n406 ^ x212 ^ 1'b0 ;
  assign n510 = n508 & n509 ;
  assign n511 = ( x23 & n507 ) | ( x23 & ~n510 ) | ( n507 & ~n510 ) ;
  assign n512 = ( ~x81 & x188 ) | ( ~x81 & x211 ) | ( x188 & x211 ) ;
  assign n513 = ( x22 & x109 ) | ( x22 & ~n512 ) | ( x109 & ~n512 ) ;
  assign n514 = ( n504 & n511 ) | ( n504 & n513 ) | ( n511 & n513 ) ;
  assign n515 = n514 ^ n321 ^ x75 ;
  assign n518 = x208 ^ x151 ^ x46 ;
  assign n516 = x209 ^ x182 ^ x171 ;
  assign n517 = ( x70 & x75 ) | ( x70 & n516 ) | ( x75 & n516 ) ;
  assign n519 = n518 ^ n517 ^ n380 ;
  assign n520 = ( x28 & ~x99 ) | ( x28 & n510 ) | ( ~x99 & n510 ) ;
  assign n521 = ( ~x7 & x134 ) | ( ~x7 & n520 ) | ( x134 & n520 ) ;
  assign n522 = n312 ^ x200 ^ x152 ;
  assign n543 = x131 & n280 ;
  assign n544 = ~n260 & n543 ;
  assign n545 = ( x210 & ~n308 ) | ( x210 & n544 ) | ( ~n308 & n544 ) ;
  assign n546 = ( ~x39 & x173 ) | ( ~x39 & n545 ) | ( x173 & n545 ) ;
  assign n547 = ( x159 & ~x231 ) | ( x159 & n546 ) | ( ~x231 & n546 ) ;
  assign n534 = x250 ^ x186 ^ x170 ;
  assign n535 = ( x101 & n262 ) | ( x101 & ~n534 ) | ( n262 & ~n534 ) ;
  assign n536 = x19 & ~n535 ;
  assign n537 = ( x19 & ~n276 ) | ( x19 & n536 ) | ( ~n276 & n536 ) ;
  assign n539 = ( x230 & x240 ) | ( x230 & n268 ) | ( x240 & n268 ) ;
  assign n538 = ( ~x66 & x184 ) | ( ~x66 & n341 ) | ( x184 & n341 ) ;
  assign n540 = n539 ^ n538 ^ n484 ;
  assign n541 = ( x216 & ~n537 ) | ( x216 & n540 ) | ( ~n537 & n540 ) ;
  assign n526 = x231 ^ x0 ^ 1'b0 ;
  assign n527 = n340 & n526 ;
  assign n528 = n527 ^ x138 ^ 1'b0 ;
  assign n529 = x163 & n528 ;
  assign n530 = n529 ^ n337 ^ x105 ;
  assign n531 = n530 ^ n323 ^ 1'b0 ;
  assign n532 = x12 & n531 ;
  assign n524 = ( x40 & ~n406 ) | ( x40 & n420 ) | ( ~n406 & n420 ) ;
  assign n523 = n402 ^ x172 ^ x140 ;
  assign n525 = n524 ^ n523 ^ x43 ;
  assign n533 = n532 ^ n525 ^ n487 ;
  assign n542 = n541 ^ n533 ^ n323 ;
  assign n548 = n547 ^ n542 ^ x26 ;
  assign n549 = n326 | n475 ;
  assign n550 = n457 | n549 ;
  assign n551 = ( x78 & x124 ) | ( x78 & ~x186 ) | ( x124 & ~x186 ) ;
  assign n552 = n551 ^ x70 ^ x46 ;
  assign n553 = x44 & ~n552 ;
  assign n554 = n553 ^ n273 ^ 1'b0 ;
  assign n555 = n400 ^ x59 ^ x5 ;
  assign n559 = n502 ^ x218 ^ x82 ;
  assign n556 = ( ~x183 & n272 ) | ( ~x183 & n391 ) | ( n272 & n391 ) ;
  assign n557 = n545 ^ x152 ^ x36 ;
  assign n558 = ( n414 & ~n556 ) | ( n414 & n557 ) | ( ~n556 & n557 ) ;
  assign n560 = n559 ^ n558 ^ n320 ;
  assign n563 = x144 ^ x114 ^ x33 ;
  assign n561 = n359 ^ x223 ^ x220 ;
  assign n562 = ( x108 & ~n364 ) | ( x108 & n561 ) | ( ~n364 & n561 ) ;
  assign n564 = n563 ^ n562 ^ 1'b0 ;
  assign n565 = n407 & ~n564 ;
  assign n566 = ( ~x153 & x209 ) | ( ~x153 & n387 ) | ( x209 & n387 ) ;
  assign n567 = x240 & ~n477 ;
  assign n568 = ( n565 & n566 ) | ( n565 & ~n567 ) | ( n566 & ~n567 ) ;
  assign n569 = n427 ^ x212 ^ x30 ;
  assign n570 = x189 ^ x173 ^ 1'b0 ;
  assign n571 = x182 & n570 ;
  assign n574 = ( ~x160 & x176 ) | ( ~x160 & n327 ) | ( x176 & n327 ) ;
  assign n572 = ( x43 & ~n317 ) | ( x43 & n505 ) | ( ~n317 & n505 ) ;
  assign n573 = x212 & ~n572 ;
  assign n575 = n574 ^ n573 ^ 1'b0 ;
  assign n576 = n571 & ~n575 ;
  assign n577 = ~n569 & n576 ;
  assign n578 = ( x1 & x57 ) | ( x1 & ~n332 ) | ( x57 & ~n332 ) ;
  assign n579 = n287 ^ x49 ^ 1'b0 ;
  assign n580 = ( n476 & ~n516 ) | ( n476 & n579 ) | ( ~n516 & n579 ) ;
  assign n581 = ( n294 & n337 ) | ( n294 & n580 ) | ( n337 & n580 ) ;
  assign n582 = ( n577 & n578 ) | ( n577 & ~n581 ) | ( n578 & ~n581 ) ;
  assign n583 = ( x20 & x113 ) | ( x20 & ~x141 ) | ( x113 & ~x141 ) ;
  assign n584 = n583 ^ x115 ^ x107 ;
  assign n585 = n584 ^ n319 ^ x111 ;
  assign n587 = n313 ^ n304 ^ x168 ;
  assign n586 = ~n323 & n568 ;
  assign n588 = n587 ^ n586 ^ 1'b0 ;
  assign n598 = n512 ^ n384 ^ n335 ;
  assign n591 = n361 ^ n256 ^ x138 ;
  assign n592 = n591 ^ n422 ^ 1'b0 ;
  assign n593 = n529 & ~n592 ;
  assign n594 = n343 ^ x203 ^ 1'b0 ;
  assign n595 = x165 & ~n594 ;
  assign n596 = n310 ^ x227 ^ x207 ;
  assign n597 = ( n593 & n595 ) | ( n593 & n596 ) | ( n595 & n596 ) ;
  assign n589 = ( x224 & n309 ) | ( x224 & ~n391 ) | ( n309 & ~n391 ) ;
  assign n590 = n589 ^ n577 ^ x95 ;
  assign n599 = n598 ^ n597 ^ n590 ;
  assign n603 = ( ~x98 & x237 ) | ( ~x98 & n546 ) | ( x237 & n546 ) ;
  assign n602 = ( x212 & x243 ) | ( x212 & n333 ) | ( x243 & n333 ) ;
  assign n600 = ( x118 & ~n284 ) | ( x118 & n416 ) | ( ~n284 & n416 ) ;
  assign n601 = ( x32 & ~x176 ) | ( x32 & n600 ) | ( ~x176 & n600 ) ;
  assign n604 = n603 ^ n602 ^ n601 ;
  assign n619 = ( ~x7 & x39 ) | ( ~x7 & x240 ) | ( x39 & x240 ) ;
  assign n607 = ( x116 & x150 ) | ( x116 & ~x201 ) | ( x150 & ~x201 ) ;
  assign n608 = x118 ^ x75 ^ x44 ;
  assign n609 = n608 ^ n301 ^ x190 ;
  assign n610 = n609 ^ x129 ^ x113 ;
  assign n611 = ( x40 & n506 ) | ( x40 & n610 ) | ( n506 & n610 ) ;
  assign n612 = ( x116 & x167 ) | ( x116 & ~x249 ) | ( x167 & ~x249 ) ;
  assign n613 = n612 ^ n469 ^ x194 ;
  assign n614 = ( x6 & x16 ) | ( x6 & ~n278 ) | ( x16 & ~n278 ) ;
  assign n615 = n317 ^ x29 ^ 1'b0 ;
  assign n616 = n614 & n615 ;
  assign n617 = ~n613 & n616 ;
  assign n618 = ( ~n607 & n611 ) | ( ~n607 & n617 ) | ( n611 & n617 ) ;
  assign n605 = x219 ^ x51 ^ x16 ;
  assign n606 = ( x16 & ~x41 ) | ( x16 & n605 ) | ( ~x41 & n605 ) ;
  assign n620 = n619 ^ n618 ^ n606 ;
  assign n621 = ( x47 & x121 ) | ( x47 & ~x150 ) | ( x121 & ~x150 ) ;
  assign n622 = ( n504 & n514 ) | ( n504 & n621 ) | ( n514 & n621 ) ;
  assign n623 = ( ~x137 & n620 ) | ( ~x137 & n622 ) | ( n620 & n622 ) ;
  assign n625 = n482 ^ x166 ^ x73 ;
  assign n624 = ( x93 & n429 ) | ( x93 & ~n431 ) | ( n429 & ~n431 ) ;
  assign n626 = n625 ^ n624 ^ x81 ;
  assign n627 = x47 ^ x18 ^ 1'b0 ;
  assign n628 = ( x111 & ~n414 ) | ( x111 & n627 ) | ( ~n414 & n627 ) ;
  assign n629 = n628 ^ n551 ^ n529 ;
  assign n630 = n407 & ~n629 ;
  assign n631 = ~n379 & n630 ;
  assign n632 = n631 ^ n433 ^ x84 ;
  assign n638 = ( ~x133 & x158 ) | ( ~x133 & x223 ) | ( x158 & x223 ) ;
  assign n633 = n417 ^ n322 ^ x180 ;
  assign n635 = ( x50 & n358 ) | ( x50 & n383 ) | ( n358 & n383 ) ;
  assign n634 = x6 & n513 ;
  assign n636 = n635 ^ n634 ^ 1'b0 ;
  assign n637 = ~n633 & n636 ;
  assign n639 = n638 ^ n637 ^ 1'b0 ;
  assign n657 = ( ~x9 & x136 ) | ( ~x9 & n352 ) | ( x136 & n352 ) ;
  assign n658 = n657 ^ x152 ^ x44 ;
  assign n659 = ( x183 & ~n388 ) | ( x183 & n658 ) | ( ~n388 & n658 ) ;
  assign n660 = ( x224 & ~x235 ) | ( x224 & n436 ) | ( ~x235 & n436 ) ;
  assign n662 = x200 ^ x194 ^ x96 ;
  assign n663 = n571 ^ x97 ^ x38 ;
  assign n664 = n663 ^ n427 ^ x104 ;
  assign n665 = ( x96 & n662 ) | ( x96 & ~n664 ) | ( n662 & ~n664 ) ;
  assign n661 = ( x151 & ~x237 ) | ( x151 & n298 ) | ( ~x237 & n298 ) ;
  assign n666 = n665 ^ n661 ^ x221 ;
  assign n667 = ( n659 & ~n660 ) | ( n659 & n666 ) | ( ~n660 & n666 ) ;
  assign n641 = ( x24 & ~n427 ) | ( x24 & n605 ) | ( ~n427 & n605 ) ;
  assign n640 = ( x35 & x123 ) | ( x35 & ~n332 ) | ( x123 & ~n332 ) ;
  assign n642 = n641 ^ n640 ^ x150 ;
  assign n643 = n518 ^ x212 ^ x19 ;
  assign n644 = ( x132 & n298 ) | ( x132 & ~n643 ) | ( n298 & ~n643 ) ;
  assign n645 = ( x170 & x194 ) | ( x170 & ~n263 ) | ( x194 & ~n263 ) ;
  assign n646 = ( n504 & n644 ) | ( n504 & n645 ) | ( n644 & n645 ) ;
  assign n651 = ( x7 & x194 ) | ( x7 & ~x244 ) | ( x194 & ~x244 ) ;
  assign n650 = n271 ^ x171 ^ x86 ;
  assign n648 = ( x110 & x173 ) | ( x110 & n318 ) | ( x173 & n318 ) ;
  assign n647 = n551 ^ n545 ^ x37 ;
  assign n649 = n648 ^ n647 ^ x157 ;
  assign n652 = n651 ^ n650 ^ n649 ;
  assign n653 = ( n495 & n646 ) | ( n495 & n652 ) | ( n646 & n652 ) ;
  assign n654 = n510 ^ n332 ^ x134 ;
  assign n655 = n654 ^ n617 ^ x244 ;
  assign n656 = ( n642 & ~n653 ) | ( n642 & n655 ) | ( ~n653 & n655 ) ;
  assign n668 = n667 ^ n656 ^ n361 ;
  assign n672 = x61 & x177 ;
  assign n673 = n378 & n672 ;
  assign n674 = n673 ^ n439 ^ n384 ;
  assign n675 = n674 ^ x254 ^ x167 ;
  assign n670 = x35 & x109 ;
  assign n671 = ~x69 & n670 ;
  assign n676 = n675 ^ n671 ^ n288 ;
  assign n678 = ( x181 & ~n439 ) | ( x181 & n676 ) | ( ~n439 & n676 ) ;
  assign n669 = x34 & ~n663 ;
  assign n677 = n676 ^ n669 ^ n465 ;
  assign n679 = n678 ^ n677 ^ n590 ;
  assign n680 = n673 ^ n587 ^ n305 ;
  assign n681 = n680 ^ n502 ^ x24 ;
  assign n682 = x142 ^ x128 ^ x111 ;
  assign n683 = ( x89 & n273 ) | ( x89 & ~n682 ) | ( n273 & ~n682 ) ;
  assign n684 = ( ~x161 & n681 ) | ( ~x161 & n683 ) | ( n681 & n683 ) ;
  assign n689 = n290 ^ n287 ^ x48 ;
  assign n690 = x233 & n689 ;
  assign n687 = n575 ^ n326 ^ n283 ;
  assign n685 = ( x187 & n410 ) | ( x187 & ~n494 ) | ( n410 & ~n494 ) ;
  assign n686 = ( ~x162 & n547 ) | ( ~x162 & n685 ) | ( n547 & n685 ) ;
  assign n688 = n687 ^ n686 ^ n638 ;
  assign n691 = n690 ^ n688 ^ x219 ;
  assign n700 = ( x43 & ~x67 ) | ( x43 & x202 ) | ( ~x67 & x202 ) ;
  assign n697 = n324 ^ n262 ^ 1'b0 ;
  assign n698 = x208 & ~n697 ;
  assign n695 = x9 & n355 ;
  assign n696 = n563 & n695 ;
  assign n694 = x192 ^ x76 ^ x33 ;
  assign n699 = n698 ^ n696 ^ n694 ;
  assign n692 = n516 ^ n420 ^ n266 ;
  assign n693 = ( x161 & n431 ) | ( x161 & n692 ) | ( n431 & n692 ) ;
  assign n701 = n700 ^ n699 ^ n693 ;
  assign n702 = n610 ^ n374 ^ x119 ;
  assign n703 = ( x75 & n277 ) | ( x75 & n702 ) | ( n277 & n702 ) ;
  assign n704 = x0 & x254 ;
  assign n705 = ( x211 & n298 ) | ( x211 & ~n404 ) | ( n298 & ~n404 ) ;
  assign n706 = ( x18 & ~x98 ) | ( x18 & n259 ) | ( ~x98 & n259 ) ;
  assign n707 = n706 ^ n561 ^ x185 ;
  assign n708 = n457 & n707 ;
  assign n709 = n705 & n708 ;
  assign n710 = ( n335 & n704 ) | ( n335 & n709 ) | ( n704 & n709 ) ;
  assign n711 = ( ~x13 & x14 ) | ( ~x13 & x20 ) | ( x14 & x20 ) ;
  assign n712 = x193 & n711 ;
  assign n713 = n712 ^ n327 ^ 1'b0 ;
  assign n714 = n713 ^ n470 ^ 1'b0 ;
  assign n715 = n422 | n714 ;
  assign n716 = ( x192 & ~x202 ) | ( x192 & n715 ) | ( ~x202 & n715 ) ;
  assign n719 = n414 ^ x60 ^ x29 ;
  assign n720 = ( n450 & n510 ) | ( n450 & ~n719 ) | ( n510 & ~n719 ) ;
  assign n721 = ( ~n667 & n694 ) | ( ~n667 & n720 ) | ( n694 & n720 ) ;
  assign n717 = ( ~x27 & n266 ) | ( ~x27 & n654 ) | ( n266 & n654 ) ;
  assign n718 = ( n283 & n295 ) | ( n283 & n717 ) | ( n295 & n717 ) ;
  assign n722 = n721 ^ n718 ^ n433 ;
  assign n726 = ( ~x109 & x240 ) | ( ~x109 & n284 ) | ( x240 & n284 ) ;
  assign n727 = ( n264 & ~n544 ) | ( n264 & n726 ) | ( ~n544 & n726 ) ;
  assign n723 = x199 & n491 ;
  assign n724 = ~x29 & n723 ;
  assign n725 = ( x184 & x239 ) | ( x184 & n724 ) | ( x239 & n724 ) ;
  assign n728 = n727 ^ n725 ^ 1'b0 ;
  assign n729 = n540 ^ x64 ^ 1'b0 ;
  assign n738 = ( x36 & ~n512 ) | ( x36 & n665 ) | ( ~n512 & n665 ) ;
  assign n735 = x221 & ~n319 ;
  assign n736 = n735 ^ x186 ^ 1'b0 ;
  assign n737 = n736 ^ n612 ^ n273 ;
  assign n730 = ( ~x66 & x121 ) | ( ~x66 & x136 ) | ( x121 & x136 ) ;
  assign n731 = x90 & x209 ;
  assign n732 = ~n730 & n731 ;
  assign n733 = ( ~x83 & n317 ) | ( ~x83 & n397 ) | ( n317 & n397 ) ;
  assign n734 = ( x119 & n732 ) | ( x119 & ~n733 ) | ( n732 & ~n733 ) ;
  assign n739 = n738 ^ n737 ^ n734 ;
  assign n740 = n739 ^ n359 ^ x208 ;
  assign n741 = ~n729 & n740 ;
  assign n742 = x148 & n741 ;
  assign n743 = ( ~x45 & n269 ) | ( ~x45 & n482 ) | ( n269 & n482 ) ;
  assign n744 = ( ~n357 & n571 ) | ( ~n357 & n651 ) | ( n571 & n651 ) ;
  assign n745 = ( ~x13 & x38 ) | ( ~x13 & x42 ) | ( x38 & x42 ) ;
  assign n746 = ( x172 & n644 ) | ( x172 & ~n745 ) | ( n644 & ~n745 ) ;
  assign n747 = n442 ^ n379 ^ x14 ;
  assign n748 = n746 | n747 ;
  assign n749 = n319 ^ x165 ^ 1'b0 ;
  assign n750 = x132 & ~n749 ;
  assign n751 = n750 ^ n674 ^ x9 ;
  assign n752 = ( x135 & n314 ) | ( x135 & n751 ) | ( n314 & n751 ) ;
  assign n756 = n619 ^ n324 ^ x47 ;
  assign n753 = x224 ^ x118 ^ x112 ;
  assign n754 = x95 & ~n506 ;
  assign n755 = n753 & n754 ;
  assign n757 = n756 ^ n755 ^ n354 ;
  assign n758 = ( x77 & ~n752 ) | ( x77 & n757 ) | ( ~n752 & n757 ) ;
  assign n759 = ( n744 & n748 ) | ( n744 & ~n758 ) | ( n748 & ~n758 ) ;
  assign n760 = x223 ^ x92 ^ x50 ;
  assign n761 = ( x30 & ~x168 ) | ( x30 & n760 ) | ( ~x168 & n760 ) ;
  assign n762 = ( x64 & x198 ) | ( x64 & n761 ) | ( x198 & n761 ) ;
  assign n763 = ( ~n607 & n759 ) | ( ~n607 & n762 ) | ( n759 & n762 ) ;
  assign n764 = x183 & x205 ;
  assign n765 = ~n763 & n764 ;
  assign n766 = ( ~n320 & n328 ) | ( ~n320 & n375 ) | ( n328 & n375 ) ;
  assign n767 = n628 ^ n496 ^ x77 ;
  assign n768 = ( n658 & ~n766 ) | ( n658 & n767 ) | ( ~n766 & n767 ) ;
  assign n770 = ( ~x183 & x186 ) | ( ~x183 & n440 ) | ( x186 & n440 ) ;
  assign n771 = n770 ^ x113 ^ 1'b0 ;
  assign n772 = n535 & ~n771 ;
  assign n773 = n772 ^ x111 ^ 1'b0 ;
  assign n769 = ( ~x64 & x82 ) | ( ~x64 & n507 ) | ( x82 & n507 ) ;
  assign n774 = n773 ^ n769 ^ x136 ;
  assign n782 = ( n336 & n579 ) | ( n336 & n709 ) | ( n579 & n709 ) ;
  assign n783 = ( ~x186 & n324 ) | ( ~x186 & n782 ) | ( n324 & n782 ) ;
  assign n775 = n652 ^ x209 ^ x14 ;
  assign n776 = n719 | n775 ;
  assign n777 = n776 ^ n341 ^ 1'b0 ;
  assign n778 = x177 & x235 ;
  assign n779 = ~n256 & n778 ;
  assign n780 = ( n477 & ~n622 ) | ( n477 & n779 ) | ( ~n622 & n779 ) ;
  assign n781 = ( n470 & n777 ) | ( n470 & n780 ) | ( n777 & n780 ) ;
  assign n784 = n783 ^ n781 ^ 1'b0 ;
  assign n785 = ( x60 & n264 ) | ( x60 & n286 ) | ( n264 & n286 ) ;
  assign n786 = ( ~x92 & n431 ) | ( ~x92 & n569 ) | ( n431 & n569 ) ;
  assign n787 = n786 ^ n391 ^ x210 ;
  assign n789 = ( ~x110 & x253 ) | ( ~x110 & n285 ) | ( x253 & n285 ) ;
  assign n790 = n694 | n789 ;
  assign n791 = x60 | n790 ;
  assign n792 = ( ~x204 & n552 ) | ( ~x204 & n791 ) | ( n552 & n791 ) ;
  assign n788 = n478 ^ n356 ^ x3 ;
  assign n793 = n792 ^ n788 ^ n357 ;
  assign n794 = ( ~n785 & n787 ) | ( ~n785 & n793 ) | ( n787 & n793 ) ;
  assign n806 = x141 ^ x98 ^ x67 ;
  assign n805 = n301 ^ x235 ^ x140 ;
  assign n804 = n650 ^ n293 ^ x245 ;
  assign n807 = n806 ^ n805 ^ n804 ;
  assign n798 = x225 ^ x40 ^ 1'b0 ;
  assign n799 = x58 & n798 ;
  assign n800 = ( x49 & n289 ) | ( x49 & ~n799 ) | ( n289 & ~n799 ) ;
  assign n801 = n800 ^ n430 ^ x40 ;
  assign n795 = n287 & n306 ;
  assign n796 = n350 & n795 ;
  assign n797 = n602 & ~n796 ;
  assign n802 = n801 ^ n797 ^ 1'b0 ;
  assign n803 = x58 & n802 ;
  assign n808 = n807 ^ n803 ^ 1'b0 ;
  assign n809 = n561 ^ x105 ^ x83 ;
  assign n810 = n698 ^ n608 ^ x211 ;
  assign n811 = ~n809 & n810 ;
  assign n812 = n811 ^ x191 ^ 1'b0 ;
  assign n813 = ( n349 & n401 ) | ( n349 & ~n548 ) | ( n401 & ~n548 ) ;
  assign n814 = ~x74 & n517 ;
  assign n815 = n814 ^ x206 ^ x3 ;
  assign n821 = n277 ^ x170 ^ x163 ;
  assign n822 = x249 & n472 ;
  assign n823 = ~n821 & n822 ;
  assign n816 = n574 ^ n379 ^ x207 ;
  assign n817 = ( x100 & x241 ) | ( x100 & n816 ) | ( x241 & n816 ) ;
  assign n818 = n495 ^ n281 ^ x223 ;
  assign n819 = ( x145 & ~n817 ) | ( x145 & n818 ) | ( ~n817 & n818 ) ;
  assign n820 = n819 ^ n709 ^ n700 ;
  assign n824 = n823 ^ n820 ^ x150 ;
  assign n825 = n598 ^ n571 ^ n494 ;
  assign n826 = n510 ^ n314 ^ x159 ;
  assign n827 = n826 ^ n733 ^ n665 ;
  assign n828 = ( x120 & ~n368 ) | ( x120 & n827 ) | ( ~n368 & n827 ) ;
  assign n829 = ( x53 & ~x141 ) | ( x53 & n828 ) | ( ~x141 & n828 ) ;
  assign n830 = n829 ^ n476 ^ n451 ;
  assign n831 = n557 ^ n293 ^ x147 ;
  assign n833 = n429 ^ x250 ^ x209 ;
  assign n834 = ( x38 & n433 ) | ( x38 & ~n833 ) | ( n433 & ~n833 ) ;
  assign n832 = ( x85 & x180 ) | ( x85 & ~n559 ) | ( x180 & ~n559 ) ;
  assign n835 = n834 ^ n832 ^ 1'b0 ;
  assign n836 = n384 ^ n375 ^ x14 ;
  assign n837 = x210 ^ x178 ^ x54 ;
  assign n838 = ( ~n298 & n416 ) | ( ~n298 & n469 ) | ( n416 & n469 ) ;
  assign n839 = ( n459 & n481 ) | ( n459 & ~n838 ) | ( n481 & ~n838 ) ;
  assign n845 = x3 & ~n271 ;
  assign n846 = ~x205 & n845 ;
  assign n847 = n846 ^ n401 ^ n263 ;
  assign n848 = ( n341 & n421 ) | ( n341 & n847 ) | ( n421 & n847 ) ;
  assign n840 = ( x57 & ~x190 ) | ( x57 & n479 ) | ( ~x190 & n479 ) ;
  assign n841 = ~n536 & n840 ;
  assign n842 = ~n403 & n841 ;
  assign n843 = ( x154 & x227 ) | ( x154 & n842 ) | ( x227 & n842 ) ;
  assign n844 = n819 & n843 ;
  assign n849 = n848 ^ n844 ^ 1'b0 ;
  assign n850 = ( n837 & ~n839 ) | ( n837 & n849 ) | ( ~n839 & n849 ) ;
  assign n851 = n656 ^ n402 ^ x61 ;
  assign n857 = ( x43 & x123 ) | ( x43 & n806 ) | ( x123 & n806 ) ;
  assign n856 = n479 ^ x108 ^ 1'b0 ;
  assign n852 = n569 ^ n328 ^ 1'b0 ;
  assign n853 = ( x27 & x163 ) | ( x27 & n852 ) | ( x163 & n852 ) ;
  assign n854 = ( ~n558 & n706 ) | ( ~n558 & n853 ) | ( n706 & n853 ) ;
  assign n855 = ( n273 & n624 ) | ( n273 & ~n854 ) | ( n624 & ~n854 ) ;
  assign n858 = n857 ^ n856 ^ n855 ;
  assign n859 = ( ~x244 & n435 ) | ( ~x244 & n460 ) | ( n435 & n460 ) ;
  assign n860 = n859 ^ n820 ^ x221 ;
  assign n870 = n361 ^ n262 ^ x224 ;
  assign n871 = n870 ^ n761 ^ x89 ;
  assign n861 = ~n418 & n551 ;
  assign n862 = n861 ^ n837 ^ 1'b0 ;
  assign n863 = ( n429 & n486 ) | ( n429 & ~n862 ) | ( n486 & ~n862 ) ;
  assign n865 = n662 ^ n308 ^ n295 ;
  assign n864 = x233 & n848 ;
  assign n866 = n865 ^ n864 ^ 1'b0 ;
  assign n867 = n713 ^ n633 ^ n401 ;
  assign n868 = ~n866 & n867 ;
  assign n869 = ( ~n863 & n866 ) | ( ~n863 & n868 ) | ( n866 & n868 ) ;
  assign n872 = n871 ^ n869 ^ n782 ;
  assign n876 = n477 ^ x103 ^ x80 ;
  assign n877 = ( x34 & ~x201 ) | ( x34 & n876 ) | ( ~x201 & n876 ) ;
  assign n873 = ( ~x100 & x127 ) | ( ~x100 & n424 ) | ( x127 & n424 ) ;
  assign n874 = ( n598 & n658 ) | ( n598 & n750 ) | ( n658 & n750 ) ;
  assign n875 = ( ~n557 & n873 ) | ( ~n557 & n874 ) | ( n873 & n874 ) ;
  assign n878 = n877 ^ n875 ^ n807 ;
  assign n879 = n400 ^ n357 ^ n291 ;
  assign n880 = n596 ^ n388 ^ x110 ;
  assign n881 = n544 ^ n389 ^ x140 ;
  assign n882 = n881 ^ n460 ^ x114 ;
  assign n884 = ( ~x73 & x113 ) | ( ~x73 & n498 ) | ( x113 & n498 ) ;
  assign n883 = n870 ^ n451 ^ x51 ;
  assign n885 = n884 ^ n883 ^ n298 ;
  assign n886 = ( n880 & n882 ) | ( n880 & n885 ) | ( n882 & n885 ) ;
  assign n887 = ( n590 & n785 ) | ( n590 & n886 ) | ( n785 & n886 ) ;
  assign n888 = ( ~n736 & n879 ) | ( ~n736 & n887 ) | ( n879 & n887 ) ;
  assign n898 = ( x111 & ~x217 ) | ( x111 & n862 ) | ( ~x217 & n862 ) ;
  assign n899 = n898 ^ n450 ^ n278 ;
  assign n900 = n658 & n899 ;
  assign n896 = ( x71 & ~x77 ) | ( x71 & n338 ) | ( ~x77 & n338 ) ;
  assign n890 = ( x166 & ~n469 ) | ( x166 & n481 ) | ( ~n469 & n481 ) ;
  assign n891 = x238 ^ x227 ^ x153 ;
  assign n892 = n890 & ~n891 ;
  assign n893 = n892 ^ x210 ^ 1'b0 ;
  assign n894 = ( ~n475 & n890 ) | ( ~n475 & n893 ) | ( n890 & n893 ) ;
  assign n895 = ( ~x7 & x155 ) | ( ~x7 & n894 ) | ( x155 & n894 ) ;
  assign n897 = n896 ^ n895 ^ n602 ;
  assign n901 = n900 ^ n897 ^ x36 ;
  assign n889 = ( n311 & n326 ) | ( n311 & ~n720 ) | ( n326 & ~n720 ) ;
  assign n902 = n901 ^ n889 ^ n611 ;
  assign n903 = ( x52 & n333 ) | ( x52 & ~n416 ) | ( n333 & ~n416 ) ;
  assign n904 = ( x124 & n294 ) | ( x124 & ~n903 ) | ( n294 & ~n903 ) ;
  assign n905 = n904 ^ x62 ^ 1'b0 ;
  assign n906 = n905 ^ n260 ^ x247 ;
  assign n907 = ( ~x27 & x110 ) | ( ~x27 & n355 ) | ( x110 & n355 ) ;
  assign n908 = ~n590 & n907 ;
  assign n909 = ~x35 & n908 ;
  assign n914 = n834 ^ n505 ^ n376 ;
  assign n910 = ( x106 & n460 ) | ( x106 & ~n862 ) | ( n460 & ~n862 ) ;
  assign n911 = n571 & ~n870 ;
  assign n912 = ~x254 & n911 ;
  assign n913 = n910 & ~n912 ;
  assign n915 = n914 ^ n913 ^ 1'b0 ;
  assign n916 = ( ~x189 & n909 ) | ( ~x189 & n915 ) | ( n909 & n915 ) ;
  assign n925 = n615 ^ n489 ^ n374 ;
  assign n923 = ( x2 & n361 ) | ( x2 & ~n609 ) | ( n361 & ~n609 ) ;
  assign n920 = x85 & x174 ;
  assign n921 = n920 ^ x91 ^ 1'b0 ;
  assign n922 = n921 ^ n442 ^ x178 ;
  assign n918 = ( n384 & n651 ) | ( n384 & n846 ) | ( n651 & n846 ) ;
  assign n917 = ( x253 & ~n274 ) | ( x253 & n312 ) | ( ~n274 & n312 ) ;
  assign n919 = n918 ^ n917 ^ n705 ;
  assign n924 = n923 ^ n922 ^ n919 ;
  assign n926 = n925 ^ n924 ^ 1'b0 ;
  assign n927 = ( x53 & ~n517 ) | ( x53 & n779 ) | ( ~n517 & n779 ) ;
  assign n928 = n689 ^ x109 ^ 1'b0 ;
  assign n929 = n927 | n928 ;
  assign n934 = x19 & x39 ;
  assign n930 = n546 ^ n423 ^ x193 ;
  assign n931 = n839 ^ x219 ^ x142 ;
  assign n932 = ( n583 & n930 ) | ( n583 & n931 ) | ( n930 & n931 ) ;
  assign n933 = ( x53 & n504 ) | ( x53 & ~n932 ) | ( n504 & ~n932 ) ;
  assign n935 = n934 ^ n933 ^ x244 ;
  assign n936 = n681 ^ x143 ^ x22 ;
  assign n937 = ( x39 & ~x189 ) | ( x39 & n598 ) | ( ~x189 & n598 ) ;
  assign n938 = n937 ^ n397 ^ x27 ;
  assign n966 = ( ~x139 & x150 ) | ( ~x139 & x227 ) | ( x150 & x227 ) ;
  assign n967 = n966 ^ x205 ^ x97 ;
  assign n968 = ( x160 & n273 ) | ( x160 & n967 ) | ( n273 & n967 ) ;
  assign n969 = ( x104 & ~n341 ) | ( x104 & n968 ) | ( ~n341 & n968 ) ;
  assign n970 = n321 ^ x121 ^ x47 ;
  assign n971 = ( n296 & n842 ) | ( n296 & n970 ) | ( n842 & n970 ) ;
  assign n972 = ( ~n280 & n969 ) | ( ~n280 & n971 ) | ( n969 & n971 ) ;
  assign n963 = n274 & n583 ;
  assign n964 = n963 ^ x61 ^ 1'b0 ;
  assign n942 = n449 ^ n428 ^ n335 ;
  assign n943 = n942 ^ n411 ^ 1'b0 ;
  assign n944 = x227 ^ x79 ^ x18 ;
  assign n945 = x218 | n944 ;
  assign n946 = n648 ^ n469 ^ x156 ;
  assign n947 = ( x10 & x228 ) | ( x10 & ~n512 ) | ( x228 & ~n512 ) ;
  assign n948 = n312 & n947 ;
  assign n949 = n948 ^ x230 ^ 1'b0 ;
  assign n950 = ( n661 & n946 ) | ( n661 & ~n949 ) | ( n946 & ~n949 ) ;
  assign n951 = n950 ^ x221 ^ x111 ;
  assign n952 = n951 ^ x64 ^ 1'b0 ;
  assign n953 = n945 & ~n952 ;
  assign n954 = ( ~x71 & x187 ) | ( ~x71 & n306 ) | ( x187 & n306 ) ;
  assign n955 = n954 ^ n434 ^ x4 ;
  assign n956 = n955 ^ n877 ^ n343 ;
  assign n957 = n956 ^ n497 ^ 1'b0 ;
  assign n958 = n957 ^ x79 ^ 1'b0 ;
  assign n959 = n953 & ~n958 ;
  assign n960 = ~n259 & n959 ;
  assign n961 = ~n943 & n960 ;
  assign n962 = ( x225 & n544 ) | ( x225 & ~n961 ) | ( n544 & ~n961 ) ;
  assign n965 = n964 ^ n962 ^ n410 ;
  assign n939 = ( n446 & ~n729 ) | ( n446 & n934 ) | ( ~n729 & n934 ) ;
  assign n940 = n558 & n939 ;
  assign n941 = ( x131 & x191 ) | ( x131 & ~n940 ) | ( x191 & ~n940 ) ;
  assign n973 = n972 ^ n965 ^ n941 ;
  assign n974 = ( ~x71 & n588 ) | ( ~x71 & n973 ) | ( n588 & n973 ) ;
  assign n975 = ( ~n285 & n938 ) | ( ~n285 & n974 ) | ( n938 & n974 ) ;
  assign n976 = x132 ^ x99 ^ 1'b0 ;
  assign n977 = n571 & n976 ;
  assign n978 = ( ~n327 & n415 ) | ( ~n327 & n977 ) | ( n415 & n977 ) ;
  assign n982 = n750 ^ n452 ^ n331 ;
  assign n983 = ( n420 & ~n783 ) | ( n420 & n982 ) | ( ~n783 & n982 ) ;
  assign n979 = ( ~x83 & x172 ) | ( ~x83 & n454 ) | ( x172 & n454 ) ;
  assign n980 = n979 ^ n659 ^ n360 ;
  assign n981 = ( ~x50 & n906 ) | ( ~x50 & n980 ) | ( n906 & n980 ) ;
  assign n984 = n983 ^ n981 ^ 1'b0 ;
  assign n1002 = ( x231 & n837 ) | ( x231 & ~n880 ) | ( n837 & ~n880 ) ;
  assign n991 = x2 & ~n805 ;
  assign n995 = n614 ^ n351 ^ x180 ;
  assign n992 = ( x49 & ~x220 ) | ( x49 & n364 ) | ( ~x220 & n364 ) ;
  assign n993 = ( n482 & n848 ) | ( n482 & ~n992 ) | ( n848 & ~n992 ) ;
  assign n994 = n322 & n993 ;
  assign n996 = n995 ^ n994 ^ 1'b0 ;
  assign n997 = n422 & n996 ;
  assign n998 = ( x233 & n499 ) | ( x233 & n997 ) | ( n499 & n997 ) ;
  assign n999 = ( n533 & ~n991 ) | ( n533 & n998 ) | ( ~n991 & n998 ) ;
  assign n1000 = n999 ^ n427 ^ x119 ;
  assign n987 = ( x189 & x191 ) | ( x189 & n449 ) | ( x191 & n449 ) ;
  assign n988 = ( x123 & n544 ) | ( x123 & ~n987 ) | ( n544 & ~n987 ) ;
  assign n985 = n450 ^ n413 ^ n341 ;
  assign n986 = n810 & n985 ;
  assign n989 = n988 ^ n986 ^ 1'b0 ;
  assign n990 = ( x153 & x209 ) | ( x153 & ~n989 ) | ( x209 & ~n989 ) ;
  assign n1001 = n1000 ^ n990 ^ x65 ;
  assign n1003 = n1002 ^ n1001 ^ n482 ;
  assign n1008 = n571 ^ x232 ^ x108 ;
  assign n1009 = ( n581 & n587 ) | ( n581 & ~n624 ) | ( n587 & ~n624 ) ;
  assign n1010 = n495 ^ n365 ^ x50 ;
  assign n1011 = ( ~n1008 & n1009 ) | ( ~n1008 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1004 = ( ~n287 & n593 ) | ( ~n287 & n917 ) | ( n593 & n917 ) ;
  assign n1005 = ( ~x87 & n309 ) | ( ~x87 & n1004 ) | ( n309 & n1004 ) ;
  assign n1006 = ( x217 & n800 ) | ( x217 & n1005 ) | ( n800 & n1005 ) ;
  assign n1007 = ( n422 & n652 ) | ( n422 & n1006 ) | ( n652 & n1006 ) ;
  assign n1012 = n1011 ^ n1007 ^ n302 ;
  assign n1024 = n859 ^ n399 ^ n359 ;
  assign n1025 = ( x97 & x117 ) | ( x97 & ~n613 ) | ( x117 & ~n613 ) ;
  assign n1026 = ( x203 & n964 ) | ( x203 & ~n1025 ) | ( n964 & ~n1025 ) ;
  assign n1027 = x84 & ~n572 ;
  assign n1028 = n1026 & n1027 ;
  assign n1029 = ( x56 & n1024 ) | ( x56 & ~n1028 ) | ( n1024 & ~n1028 ) ;
  assign n1013 = n378 ^ x177 ^ x173 ;
  assign n1014 = ( n282 & n491 ) | ( n282 & n1013 ) | ( n491 & n1013 ) ;
  assign n1015 = n877 ^ n598 ^ x234 ;
  assign n1016 = n617 ^ n615 ^ x123 ;
  assign n1017 = x155 & x189 ;
  assign n1018 = n1017 ^ n782 ^ 1'b0 ;
  assign n1019 = n1018 ^ n571 ^ n520 ;
  assign n1020 = n1019 ^ x80 ^ 1'b0 ;
  assign n1021 = x101 & ~n1020 ;
  assign n1022 = ( x16 & n1016 ) | ( x16 & ~n1021 ) | ( n1016 & ~n1021 ) ;
  assign n1023 = ( ~n1014 & n1015 ) | ( ~n1014 & n1022 ) | ( n1015 & n1022 ) ;
  assign n1030 = n1029 ^ n1023 ^ n990 ;
  assign n1039 = n1011 ^ n378 ^ n362 ;
  assign n1031 = n530 ^ x141 ^ 1'b0 ;
  assign n1032 = x185 & ~n1031 ;
  assign n1033 = ~n894 & n1032 ;
  assign n1034 = n1033 ^ n387 ^ x165 ;
  assign n1035 = n363 ^ x133 ^ x27 ;
  assign n1036 = n1035 ^ n389 ^ n370 ;
  assign n1037 = n715 | n1036 ;
  assign n1038 = n1034 & ~n1037 ;
  assign n1040 = n1039 ^ n1038 ^ 1'b0 ;
  assign n1041 = ~n860 & n1040 ;
  assign n1042 = n461 ^ n334 ^ x122 ;
  assign n1049 = n733 ^ n300 ^ x251 ;
  assign n1043 = x244 & n903 ;
  assign n1044 = n1043 ^ x47 ^ 1'b0 ;
  assign n1045 = n593 & ~n1044 ;
  assign n1046 = ~x198 & n1045 ;
  assign n1047 = n1046 ^ x140 ^ x73 ;
  assign n1048 = n1047 ^ n287 ^ x152 ;
  assign n1050 = n1049 ^ n1048 ^ n1026 ;
  assign n1051 = n1042 & ~n1050 ;
  assign n1052 = x127 | n386 ;
  assign n1053 = n1052 ^ n837 ^ n401 ;
  assign n1054 = n1053 ^ n769 ^ x122 ;
  assign n1061 = ( x149 & x225 ) | ( x149 & ~n707 ) | ( x225 & ~n707 ) ;
  assign n1055 = ( n565 & n786 ) | ( n565 & ~n817 ) | ( n786 & ~n817 ) ;
  assign n1057 = n625 ^ x77 ^ x16 ;
  assign n1056 = n853 ^ n511 ^ n410 ;
  assign n1058 = n1057 ^ n1056 ^ n580 ;
  assign n1059 = ( n883 & ~n1055 ) | ( n883 & n1058 ) | ( ~n1055 & n1058 ) ;
  assign n1060 = ( x76 & ~x141 ) | ( x76 & n1059 ) | ( ~x141 & n1059 ) ;
  assign n1062 = n1061 ^ n1060 ^ x73 ;
  assign n1063 = ( n625 & n1021 ) | ( n625 & ~n1062 ) | ( n1021 & ~n1062 ) ;
  assign n1064 = n1063 ^ x132 ^ x9 ;
  assign n1065 = n1064 ^ n545 ^ n305 ;
  assign n1081 = n288 ^ x153 ^ x93 ;
  assign n1082 = ( x105 & ~n847 ) | ( x105 & n1081 ) | ( ~n847 & n1081 ) ;
  assign n1066 = x186 & ~n713 ;
  assign n1067 = n625 & n1066 ;
  assign n1068 = n587 | n1067 ;
  assign n1069 = x4 | n1068 ;
  assign n1070 = n980 & n1069 ;
  assign n1071 = n468 & n1070 ;
  assign n1072 = x193 ^ x126 ^ x85 ;
  assign n1073 = n1072 ^ n536 ^ x218 ;
  assign n1074 = ( ~n628 & n874 ) | ( ~n628 & n1073 ) | ( n874 & n1073 ) ;
  assign n1075 = n1074 ^ n894 ^ n571 ;
  assign n1076 = ( x29 & n314 ) | ( x29 & ~n707 ) | ( n314 & ~n707 ) ;
  assign n1077 = n1076 ^ n372 ^ n360 ;
  assign n1078 = x192 ^ x175 ^ x84 ;
  assign n1079 = ( x190 & ~n1077 ) | ( x190 & n1078 ) | ( ~n1077 & n1078 ) ;
  assign n1080 = ( n1071 & n1075 ) | ( n1071 & ~n1079 ) | ( n1075 & ~n1079 ) ;
  assign n1083 = n1082 ^ n1080 ^ n454 ;
  assign n1084 = n640 ^ x154 ^ x44 ;
  assign n1085 = n1084 ^ n312 ^ x100 ;
  assign n1086 = ~n350 & n644 ;
  assign n1087 = ~n523 & n956 ;
  assign n1088 = n1086 & n1087 ;
  assign n1089 = ( ~x51 & x150 ) | ( ~x51 & x197 ) | ( x150 & x197 ) ;
  assign n1090 = ( x168 & x219 ) | ( x168 & ~n1089 ) | ( x219 & ~n1089 ) ;
  assign n1091 = n1090 ^ n508 ^ x69 ;
  assign n1092 = n1091 ^ n774 ^ n487 ;
  assign n1093 = ( ~n268 & n1088 ) | ( ~n268 & n1092 ) | ( n1088 & n1092 ) ;
  assign n1094 = n358 ^ x28 ^ 1'b0 ;
  assign n1095 = n476 ^ n273 ^ x107 ;
  assign n1096 = ( ~x28 & n568 ) | ( ~x28 & n1095 ) | ( n568 & n1095 ) ;
  assign n1097 = ( x39 & n339 ) | ( x39 & n773 ) | ( n339 & n773 ) ;
  assign n1098 = ( n423 & ~n623 ) | ( n423 & n809 ) | ( ~n623 & n809 ) ;
  assign n1099 = n1098 ^ n832 ^ x134 ;
  assign n1100 = n473 ^ x97 ^ x9 ;
  assign n1101 = ( n322 & n903 ) | ( n322 & ~n996 ) | ( n903 & ~n996 ) ;
  assign n1102 = ( n277 & n1100 ) | ( n277 & n1101 ) | ( n1100 & n1101 ) ;
  assign n1103 = ( x194 & n572 ) | ( x194 & n809 ) | ( n572 & n809 ) ;
  assign n1104 = ( ~n473 & n1102 ) | ( ~n473 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1105 = ( ~x119 & n283 ) | ( ~x119 & n386 ) | ( n283 & n386 ) ;
  assign n1106 = ( n511 & n905 ) | ( n511 & n1105 ) | ( n905 & n1105 ) ;
  assign n1107 = ( n657 & n921 ) | ( n657 & n1106 ) | ( n921 & n1106 ) ;
  assign n1108 = ( ~x236 & n266 ) | ( ~x236 & n1034 ) | ( n266 & n1034 ) ;
  assign n1109 = n1108 ^ n742 ^ x179 ;
  assign n1110 = x141 & n993 ;
  assign n1111 = ~n827 & n1110 ;
  assign n1112 = ( x169 & n904 ) | ( x169 & ~n953 ) | ( n904 & ~n953 ) ;
  assign n1113 = ( x204 & ~n1111 ) | ( x204 & n1112 ) | ( ~n1111 & n1112 ) ;
  assign n1114 = ( ~n391 & n773 ) | ( ~n391 & n1113 ) | ( n773 & n1113 ) ;
  assign n1115 = ( ~x44 & x168 ) | ( ~x44 & n505 ) | ( x168 & n505 ) ;
  assign n1116 = n1115 ^ n328 ^ x152 ;
  assign n1117 = x60 & ~n1116 ;
  assign n1122 = n946 ^ n721 ^ x110 ;
  assign n1123 = n1122 ^ n866 ^ x178 ;
  assign n1124 = n1123 ^ n762 ^ n620 ;
  assign n1118 = ( x52 & x240 ) | ( x52 & n424 ) | ( x240 & n424 ) ;
  assign n1119 = n1056 ^ n770 ^ x104 ;
  assign n1120 = ( x238 & ~n1014 ) | ( x238 & n1119 ) | ( ~n1014 & n1119 ) ;
  assign n1121 = ~n1118 & n1120 ;
  assign n1125 = n1124 ^ n1121 ^ n617 ;
  assign n1126 = n715 ^ x173 ^ 1'b0 ;
  assign n1127 = n487 & ~n1126 ;
  assign n1128 = x226 & n907 ;
  assign n1129 = ~x224 & n1128 ;
  assign n1130 = ( ~n319 & n527 ) | ( ~n319 & n806 ) | ( n527 & n806 ) ;
  assign n1131 = n1130 ^ x212 ^ x128 ;
  assign n1132 = n1131 ^ n290 ^ x229 ;
  assign n1133 = n1132 ^ n780 ^ x192 ;
  assign n1134 = ( ~n1127 & n1129 ) | ( ~n1127 & n1133 ) | ( n1129 & n1133 ) ;
  assign n1135 = n525 ^ n428 ^ n278 ;
  assign n1136 = ( x182 & n953 ) | ( x182 & ~n1135 ) | ( n953 & ~n1135 ) ;
  assign n1138 = n263 & n987 ;
  assign n1139 = n1138 ^ n985 ^ 1'b0 ;
  assign n1137 = n880 ^ n585 ^ n541 ;
  assign n1140 = n1139 ^ n1137 ^ 1'b0 ;
  assign n1141 = n1136 & n1140 ;
  assign n1142 = n619 ^ x183 ^ x168 ;
  assign n1143 = n1142 ^ n643 ^ x87 ;
  assign n1144 = n1143 ^ n326 ^ 1'b0 ;
  assign n1145 = x58 & ~n1144 ;
  assign n1146 = ( n607 & n618 ) | ( n607 & ~n1145 ) | ( n618 & ~n1145 ) ;
  assign n1147 = ( ~n363 & n1141 ) | ( ~n363 & n1146 ) | ( n1141 & n1146 ) ;
  assign n1148 = ( ~n701 & n748 ) | ( ~n701 & n840 ) | ( n748 & n840 ) ;
  assign n1151 = n661 ^ n417 ^ n342 ;
  assign n1152 = ( ~x107 & n602 ) | ( ~x107 & n1151 ) | ( n602 & n1151 ) ;
  assign n1149 = n482 ^ n308 ^ x72 ;
  assign n1150 = ( n295 & n1106 ) | ( n295 & n1149 ) | ( n1106 & n1149 ) ;
  assign n1153 = n1152 ^ n1150 ^ 1'b0 ;
  assign n1154 = n1132 ^ n293 ^ x12 ;
  assign n1155 = n1154 ^ x185 ^ 1'b0 ;
  assign n1156 = ( x47 & ~x130 ) | ( x47 & n1155 ) | ( ~x130 & n1155 ) ;
  assign n1157 = ~n1153 & n1156 ;
  assign n1158 = n931 ^ n914 ^ n382 ;
  assign n1159 = ( n431 & n729 ) | ( n431 & ~n1158 ) | ( n729 & ~n1158 ) ;
  assign n1160 = n1159 ^ n406 ^ x93 ;
  assign n1166 = ( n444 & n496 ) | ( n444 & ~n901 ) | ( n496 & ~n901 ) ;
  assign n1163 = n470 ^ n428 ^ 1'b0 ;
  assign n1164 = x160 & n1163 ;
  assign n1165 = n1164 ^ n876 ^ n551 ;
  assign n1161 = ( n393 & ~n867 ) | ( n393 & n1026 ) | ( ~n867 & n1026 ) ;
  assign n1162 = n563 | n1161 ;
  assign n1167 = n1166 ^ n1165 ^ n1162 ;
  assign n1168 = ~n755 & n1167 ;
  assign n1169 = ~n1160 & n1168 ;
  assign n1170 = ( x192 & x237 ) | ( x192 & ~n738 ) | ( x237 & ~n738 ) ;
  assign n1171 = x135 & ~n460 ;
  assign n1172 = ( n1062 & n1170 ) | ( n1062 & n1171 ) | ( n1170 & n1171 ) ;
  assign n1173 = n561 ^ n260 ^ x127 ;
  assign n1174 = ( ~n435 & n751 ) | ( ~n435 & n1173 ) | ( n751 & n1173 ) ;
  assign n1177 = x132 & ~n313 ;
  assign n1178 = n1177 ^ x118 ^ 1'b0 ;
  assign n1179 = n881 & ~n967 ;
  assign n1180 = n1178 & n1179 ;
  assign n1175 = n865 ^ n591 ^ n359 ;
  assign n1176 = ( ~x103 & n464 ) | ( ~x103 & n1175 ) | ( n464 & n1175 ) ;
  assign n1181 = n1180 ^ n1176 ^ x151 ;
  assign n1182 = n508 | n831 ;
  assign n1183 = ( x122 & ~n1181 ) | ( x122 & n1182 ) | ( ~n1181 & n1182 ) ;
  assign n1191 = n650 ^ x171 ^ x3 ;
  assign n1188 = n954 ^ x88 ^ x72 ;
  assign n1184 = n738 ^ n371 ^ n336 ;
  assign n1185 = x13 & x51 ;
  assign n1186 = ~n819 & n1185 ;
  assign n1187 = ( ~n642 & n1184 ) | ( ~n642 & n1186 ) | ( n1184 & n1186 ) ;
  assign n1189 = n1188 ^ n1187 ^ x41 ;
  assign n1190 = n524 | n1189 ;
  assign n1192 = n1191 ^ n1190 ^ 1'b0 ;
  assign n1193 = ( x100 & n349 ) | ( x100 & n730 ) | ( n349 & n730 ) ;
  assign n1194 = n1193 ^ n942 ^ n360 ;
  assign n1195 = n598 ^ x189 ^ x99 ;
  assign n1196 = n1131 ^ n650 ^ 1'b0 ;
  assign n1197 = n1171 ^ n643 ^ n309 ;
  assign n1198 = ( n1195 & n1196 ) | ( n1195 & ~n1197 ) | ( n1196 & ~n1197 ) ;
  assign n1199 = ( ~n356 & n686 ) | ( ~n356 & n874 ) | ( n686 & n874 ) ;
  assign n1200 = n1199 ^ n780 ^ 1'b0 ;
  assign n1201 = ( n1194 & ~n1198 ) | ( n1194 & n1200 ) | ( ~n1198 & n1200 ) ;
  assign n1205 = ( x46 & n256 ) | ( x46 & ~n491 ) | ( n256 & ~n491 ) ;
  assign n1204 = ( n490 & ~n840 ) | ( n490 & n983 ) | ( ~n840 & n983 ) ;
  assign n1202 = n450 | n814 ;
  assign n1203 = n574 | n1202 ;
  assign n1206 = n1205 ^ n1204 ^ n1203 ;
  assign n1207 = n518 ^ x60 ^ 1'b0 ;
  assign n1208 = ( ~x19 & x146 ) | ( ~x19 & n921 ) | ( x146 & n921 ) ;
  assign n1209 = n1208 ^ n724 ^ 1'b0 ;
  assign n1210 = n1209 ^ n1056 ^ n388 ;
  assign n1226 = n302 ^ n290 ^ x244 ;
  assign n1227 = n1226 ^ n947 ^ n614 ;
  assign n1224 = ( x37 & n580 ) | ( x37 & n760 ) | ( n580 & n760 ) ;
  assign n1222 = n427 ^ n414 ^ 1'b0 ;
  assign n1223 = n1222 ^ n877 ^ x12 ;
  assign n1225 = n1224 ^ n1223 ^ n987 ;
  assign n1228 = n1227 ^ n1225 ^ n1124 ;
  assign n1217 = ( x96 & ~n839 ) | ( x96 & n866 ) | ( ~n839 & n866 ) ;
  assign n1218 = ( ~n265 & n862 ) | ( ~n265 & n904 ) | ( n862 & n904 ) ;
  assign n1219 = n1218 ^ n597 ^ n263 ;
  assign n1220 = ( n317 & ~n1217 ) | ( n317 & n1219 ) | ( ~n1217 & n1219 ) ;
  assign n1213 = n427 ^ x145 ^ x109 ;
  assign n1214 = n1213 ^ n785 ^ n438 ;
  assign n1215 = ( x36 & ~n722 ) | ( x36 & n1214 ) | ( ~n722 & n1214 ) ;
  assign n1216 = n998 | n1215 ;
  assign n1221 = n1220 ^ n1216 ^ 1'b0 ;
  assign n1211 = n530 ^ n521 ^ x65 ;
  assign n1212 = ( n460 & n907 ) | ( n460 & ~n1211 ) | ( n907 & ~n1211 ) ;
  assign n1229 = n1228 ^ n1221 ^ n1212 ;
  assign n1230 = n1115 ^ n618 ^ x154 ;
  assign n1231 = n1230 ^ n1226 ^ x236 ;
  assign n1232 = ( x180 & n424 ) | ( x180 & ~n569 ) | ( n424 & ~n569 ) ;
  assign n1233 = n1232 ^ n782 ^ n567 ;
  assign n1234 = n1231 & n1233 ;
  assign n1235 = n1234 ^ n269 ^ 1'b0 ;
  assign n1236 = ( ~x71 & n583 ) | ( ~x71 & n1219 ) | ( n583 & n1219 ) ;
  assign n1237 = n640 & n917 ;
  assign n1238 = n1237 ^ n547 ^ 1'b0 ;
  assign n1239 = ( n865 & n1036 ) | ( n865 & n1238 ) | ( n1036 & n1238 ) ;
  assign n1240 = ( n998 & ~n1236 ) | ( n998 & n1239 ) | ( ~n1236 & n1239 ) ;
  assign n1245 = n394 ^ x186 ^ x54 ;
  assign n1244 = ( n338 & n396 ) | ( n338 & n561 ) | ( n396 & n561 ) ;
  assign n1246 = n1245 ^ n1244 ^ n921 ;
  assign n1241 = x209 & ~n979 ;
  assign n1242 = n1241 ^ n436 ^ 1'b0 ;
  assign n1243 = n1242 ^ n1132 ^ x237 ;
  assign n1247 = n1246 ^ n1243 ^ n813 ;
  assign n1256 = ( x60 & x190 ) | ( x60 & n467 ) | ( x190 & n467 ) ;
  assign n1257 = n1256 ^ n943 ^ n874 ;
  assign n1248 = ( x233 & x247 ) | ( x233 & ~n556 ) | ( x247 & ~n556 ) ;
  assign n1249 = ( x130 & x154 ) | ( x130 & ~x184 ) | ( x154 & ~x184 ) ;
  assign n1250 = n1249 ^ x173 ^ x37 ;
  assign n1251 = n1248 & ~n1250 ;
  assign n1252 = n370 & n1251 ;
  assign n1253 = x76 & n773 ;
  assign n1254 = n1252 & n1253 ;
  assign n1255 = ( n287 & n703 ) | ( n287 & n1254 ) | ( n703 & n1254 ) ;
  assign n1258 = n1257 ^ n1255 ^ n1078 ;
  assign n1259 = n895 ^ x157 ^ x4 ;
  assign n1260 = n1259 ^ x79 ^ 1'b0 ;
  assign n1270 = ( x229 & ~x244 ) | ( x229 & n883 ) | ( ~x244 & n883 ) ;
  assign n1264 = ( x101 & x189 ) | ( x101 & ~x233 ) | ( x189 & ~x233 ) ;
  assign n1265 = n1264 ^ n355 ^ x152 ;
  assign n1266 = n1265 ^ n1010 ^ n552 ;
  assign n1267 = n1266 ^ x37 ^ 1'b0 ;
  assign n1263 = n816 ^ n725 ^ n365 ;
  assign n1261 = n1250 ^ n698 ^ n372 ;
  assign n1262 = n1261 ^ n664 ^ n401 ;
  assign n1268 = n1267 ^ n1263 ^ n1262 ;
  assign n1269 = ( n424 & n1101 ) | ( n424 & n1268 ) | ( n1101 & n1268 ) ;
  assign n1271 = n1270 ^ n1269 ^ n323 ;
  assign n1272 = n739 & n1137 ;
  assign n1273 = x108 & ~n552 ;
  assign n1274 = ~n569 & n1273 ;
  assign n1275 = n890 ^ n457 ^ x132 ;
  assign n1279 = ( x91 & ~n266 ) | ( x91 & n370 ) | ( ~n266 & n370 ) ;
  assign n1276 = n791 ^ n534 ^ n347 ;
  assign n1277 = n1276 ^ n893 ^ x161 ;
  assign n1278 = n1277 ^ n1063 ^ n624 ;
  assign n1280 = n1279 ^ n1278 ^ n537 ;
  assign n1281 = ( n1274 & n1275 ) | ( n1274 & ~n1280 ) | ( n1275 & ~n1280 ) ;
  assign n1282 = n469 ^ x13 ^ x4 ;
  assign n1283 = ( x232 & ~n427 ) | ( x232 & n1195 ) | ( ~n427 & n1195 ) ;
  assign n1284 = n1283 ^ x101 ^ x29 ;
  assign n1285 = x83 ^ x30 ^ x25 ;
  assign n1286 = ( n1282 & n1284 ) | ( n1282 & n1285 ) | ( n1284 & n1285 ) ;
  assign n1287 = n1286 ^ n993 ^ x118 ;
  assign n1288 = ( n358 & ~n1131 ) | ( n358 & n1270 ) | ( ~n1131 & n1270 ) ;
  assign n1289 = x172 ^ x75 ^ x48 ;
  assign n1290 = ( n1016 & ~n1288 ) | ( n1016 & n1289 ) | ( ~n1288 & n1289 ) ;
  assign n1292 = n494 ^ x131 ^ x68 ;
  assign n1293 = n664 ^ x153 ^ x144 ;
  assign n1294 = ( x45 & ~n1292 ) | ( x45 & n1293 ) | ( ~n1292 & n1293 ) ;
  assign n1295 = ( n438 & n483 ) | ( n438 & ~n1294 ) | ( n483 & ~n1294 ) ;
  assign n1291 = n446 ^ n282 ^ x210 ;
  assign n1296 = n1295 ^ n1291 ^ n786 ;
  assign n1299 = ( n506 & ~n736 ) | ( n506 & n977 ) | ( ~n736 & n977 ) ;
  assign n1300 = n1299 ^ n883 ^ x115 ;
  assign n1297 = ( x8 & n437 ) | ( x8 & ~n1048 ) | ( n437 & ~n1048 ) ;
  assign n1298 = ( x94 & n924 ) | ( x94 & n1297 ) | ( n924 & n1297 ) ;
  assign n1301 = n1300 ^ n1298 ^ n965 ;
  assign n1302 = ( n652 & ~n1296 ) | ( n652 & n1301 ) | ( ~n1296 & n1301 ) ;
  assign n1303 = n1302 ^ n1105 ^ x87 ;
  assign n1308 = ( ~n391 & n415 ) | ( ~n391 & n618 ) | ( n415 & n618 ) ;
  assign n1309 = n1308 ^ n1193 ^ n457 ;
  assign n1310 = n1309 ^ n757 ^ 1'b0 ;
  assign n1307 = x184 & ~n627 ;
  assign n1311 = n1310 ^ n1307 ^ n513 ;
  assign n1304 = ( ~n611 & n649 ) | ( ~n611 & n834 ) | ( n649 & n834 ) ;
  assign n1305 = ( ~n870 & n1025 ) | ( ~n870 & n1304 ) | ( n1025 & n1304 ) ;
  assign n1306 = ( n648 & ~n819 ) | ( n648 & n1305 ) | ( ~n819 & n1305 ) ;
  assign n1312 = n1311 ^ n1306 ^ 1'b0 ;
  assign n1322 = ( x69 & ~x149 ) | ( x69 & x162 ) | ( ~x149 & x162 ) ;
  assign n1323 = ( n275 & n426 ) | ( n275 & n1322 ) | ( n426 & n1322 ) ;
  assign n1324 = ( n277 & n400 ) | ( n277 & n1323 ) | ( n400 & n1323 ) ;
  assign n1319 = n345 ^ n306 ^ x242 ;
  assign n1320 = ( x131 & ~n687 ) | ( x131 & n1319 ) | ( ~n687 & n1319 ) ;
  assign n1321 = n1320 ^ n909 ^ n707 ;
  assign n1325 = n1324 ^ n1321 ^ n657 ;
  assign n1317 = x226 ^ x209 ^ x171 ;
  assign n1318 = n1317 ^ n1277 ^ n1073 ;
  assign n1314 = ( x164 & n833 ) | ( x164 & n1218 ) | ( n833 & n1218 ) ;
  assign n1313 = n669 ^ n417 ^ 1'b0 ;
  assign n1315 = n1314 ^ n1313 ^ n1136 ;
  assign n1316 = n1315 ^ n978 ^ n635 ;
  assign n1326 = n1325 ^ n1318 ^ n1316 ;
  assign n1327 = ( n774 & ~n1051 ) | ( n774 & n1326 ) | ( ~n1051 & n1326 ) ;
  assign n1330 = ( n534 & ~n721 ) | ( n534 & n838 ) | ( ~n721 & n838 ) ;
  assign n1331 = n1330 ^ n750 ^ 1'b0 ;
  assign n1332 = x152 & ~n1331 ;
  assign n1333 = ( n765 & ~n1151 ) | ( n765 & n1332 ) | ( ~n1151 & n1332 ) ;
  assign n1329 = n809 ^ n707 ^ n256 ;
  assign n1328 = ( ~x118 & n266 ) | ( ~x118 & n789 ) | ( n266 & n789 ) ;
  assign n1334 = n1333 ^ n1329 ^ n1328 ;
  assign n1335 = n1334 ^ n983 ^ n625 ;
  assign n1336 = n848 ^ n337 ^ x186 ;
  assign n1337 = ( n304 & n725 ) | ( n304 & ~n1336 ) | ( n725 & ~n1336 ) ;
  assign n1338 = ( ~n886 & n1142 ) | ( ~n886 & n1337 ) | ( n1142 & n1337 ) ;
  assign n1339 = n1338 ^ n372 ^ x241 ;
  assign n1340 = n1098 ^ n512 ^ x153 ;
  assign n1341 = ~n938 & n1340 ;
  assign n1342 = ( x4 & x99 ) | ( x4 & ~n799 ) | ( x99 & ~n799 ) ;
  assign n1343 = ( ~n261 & n560 ) | ( ~n261 & n1132 ) | ( n560 & n1132 ) ;
  assign n1344 = ( n748 & n1342 ) | ( n748 & n1343 ) | ( n1342 & n1343 ) ;
  assign n1345 = n717 ^ x211 ^ 1'b0 ;
  assign n1346 = n1345 ^ n342 ^ x116 ;
  assign n1347 = n1344 & n1346 ;
  assign n1348 = ( x128 & ~x166 ) | ( x128 & n286 ) | ( ~x166 & n286 ) ;
  assign n1349 = ( x124 & n277 ) | ( x124 & ~n1055 ) | ( n277 & ~n1055 ) ;
  assign n1350 = ( n1220 & n1348 ) | ( n1220 & ~n1349 ) | ( n1348 & ~n1349 ) ;
  assign n1351 = ( n677 & ~n742 ) | ( n677 & n1350 ) | ( ~n742 & n1350 ) ;
  assign n1352 = ( n1014 & n1289 ) | ( n1014 & ~n1351 ) | ( n1289 & ~n1351 ) ;
  assign n1353 = n527 & ~n1352 ;
  assign n1354 = n1353 ^ n1141 ^ 1'b0 ;
  assign n1355 = ( n1000 & ~n1046 ) | ( n1000 & n1354 ) | ( ~n1046 & n1354 ) ;
  assign n1358 = n880 ^ n499 ^ x151 ;
  assign n1359 = n1358 ^ n900 ^ n375 ;
  assign n1356 = n261 & ~n589 ;
  assign n1357 = n1356 ^ n720 ^ x13 ;
  assign n1360 = n1359 ^ n1357 ^ x144 ;
  assign n1361 = ( n665 & n1086 ) | ( n665 & n1343 ) | ( n1086 & n1343 ) ;
  assign n1362 = n1361 ^ n767 ^ n548 ;
  assign n1363 = n1362 ^ n991 ^ x202 ;
  assign n1364 = n1363 ^ n319 ^ 1'b0 ;
  assign n1365 = x115 & ~x197 ;
  assign n1366 = n464 & n937 ;
  assign n1367 = ~x129 & n1366 ;
  assign n1368 = ( n393 & n1291 ) | ( n393 & ~n1367 ) | ( n1291 & ~n1367 ) ;
  assign n1369 = n643 ^ x3 ^ 1'b0 ;
  assign n1370 = n433 & n1369 ;
  assign n1371 = ~n609 & n1370 ;
  assign n1372 = n1368 & n1371 ;
  assign n1373 = ( ~n865 & n1365 ) | ( ~n865 & n1372 ) | ( n1365 & n1372 ) ;
  assign n1374 = ( ~x107 & n569 ) | ( ~x107 & n1048 ) | ( n569 & n1048 ) ;
  assign n1375 = ( x239 & n1373 ) | ( x239 & ~n1374 ) | ( n1373 & ~n1374 ) ;
  assign n1385 = n739 ^ n259 ^ 1'b0 ;
  assign n1386 = n772 ^ n554 ^ 1'b0 ;
  assign n1387 = n1385 & n1386 ;
  assign n1388 = n1387 ^ n311 ^ x218 ;
  assign n1377 = n646 ^ x247 ^ x163 ;
  assign n1376 = ( ~x119 & x136 ) | ( ~x119 & x230 ) | ( x136 & x230 ) ;
  assign n1378 = n1377 ^ n1376 ^ x213 ;
  assign n1379 = ( n899 & ~n1145 ) | ( n899 & n1378 ) | ( ~n1145 & n1378 ) ;
  assign n1380 = n1379 ^ x240 ^ x154 ;
  assign n1381 = n961 ^ n423 ^ n406 ;
  assign n1382 = n1013 ^ n966 ^ n873 ;
  assign n1383 = n1382 ^ n1145 ^ x127 ;
  assign n1384 = ( n1380 & ~n1381 ) | ( n1380 & n1383 ) | ( ~n1381 & n1383 ) ;
  assign n1389 = n1388 ^ n1384 ^ x136 ;
  assign n1397 = n936 ^ n923 ^ n433 ;
  assign n1392 = ( x198 & ~n853 ) | ( x198 & n992 ) | ( ~n853 & n992 ) ;
  assign n1393 = n1392 ^ n420 ^ x186 ;
  assign n1394 = ( ~n565 & n1336 ) | ( ~n565 & n1393 ) | ( n1336 & n1393 ) ;
  assign n1395 = ( ~x252 & n1294 ) | ( ~x252 & n1394 ) | ( n1294 & n1394 ) ;
  assign n1396 = n1395 ^ n673 ^ 1'b0 ;
  assign n1390 = ( n311 & n617 ) | ( n311 & n1245 ) | ( n617 & n1245 ) ;
  assign n1391 = ( n1006 & n1131 ) | ( n1006 & ~n1390 ) | ( n1131 & ~n1390 ) ;
  assign n1398 = n1397 ^ n1396 ^ n1391 ;
  assign n1399 = ( x124 & n1094 ) | ( x124 & ~n1292 ) | ( n1094 & ~n1292 ) ;
  assign n1403 = ( x54 & x110 ) | ( x54 & n1171 ) | ( x110 & n1171 ) ;
  assign n1400 = x243 & ~n343 ;
  assign n1401 = ~n345 & n1400 ;
  assign n1402 = n1401 ^ x79 ^ 1'b0 ;
  assign n1404 = n1403 ^ n1402 ^ n272 ;
  assign n1405 = n556 ^ x190 ^ x17 ;
  assign n1406 = n1385 ^ n924 ^ n271 ;
  assign n1407 = ( n724 & n1405 ) | ( n724 & ~n1406 ) | ( n1405 & ~n1406 ) ;
  assign n1413 = n706 ^ n305 ^ 1'b0 ;
  assign n1414 = ( x181 & n1323 ) | ( x181 & ~n1413 ) | ( n1323 & ~n1413 ) ;
  assign n1415 = n1414 ^ x216 ^ x103 ;
  assign n1416 = ( n287 & n782 ) | ( n287 & n1415 ) | ( n782 & n1415 ) ;
  assign n1411 = n745 ^ n339 ^ x59 ;
  assign n1408 = n1264 ^ n853 ^ n617 ;
  assign n1409 = n1408 ^ n890 ^ n457 ;
  assign n1410 = n1409 ^ x177 ^ 1'b0 ;
  assign n1412 = n1411 ^ n1410 ^ n990 ;
  assign n1417 = n1416 ^ n1412 ^ n1078 ;
  assign n1423 = n1365 ^ n802 ^ n671 ;
  assign n1418 = ( x169 & n391 ) | ( x169 & n469 ) | ( n391 & n469 ) ;
  assign n1419 = n595 & ~n1418 ;
  assign n1420 = ( n437 & n752 ) | ( n437 & n1419 ) | ( n752 & n1419 ) ;
  assign n1421 = ( ~n498 & n650 ) | ( ~n498 & n1420 ) | ( n650 & n1420 ) ;
  assign n1422 = ( x9 & n669 ) | ( x9 & ~n1421 ) | ( n669 & ~n1421 ) ;
  assign n1424 = n1423 ^ n1422 ^ n1267 ;
  assign n1425 = ( ~x76 & n1417 ) | ( ~x76 & n1424 ) | ( n1417 & n1424 ) ;
  assign n1440 = ( n341 & n363 ) | ( n341 & n499 ) | ( n363 & n499 ) ;
  assign n1441 = x238 ^ x105 ^ 1'b0 ;
  assign n1442 = n374 & n1441 ;
  assign n1436 = ( n292 & n496 ) | ( n292 & ~n625 ) | ( n496 & ~n625 ) ;
  assign n1437 = n1436 ^ n1028 ^ n551 ;
  assign n1443 = n1442 ^ n1437 ^ n817 ;
  assign n1444 = n1443 ^ n1406 ^ 1'b0 ;
  assign n1445 = n365 & n1444 ;
  assign n1446 = ( n825 & n1440 ) | ( n825 & n1445 ) | ( n1440 & n1445 ) ;
  assign n1429 = x201 & n627 ;
  assign n1430 = n1429 ^ x103 ^ 1'b0 ;
  assign n1431 = ( x134 & ~n947 ) | ( x134 & n1430 ) | ( ~n947 & n1430 ) ;
  assign n1432 = ( x138 & n940 ) | ( x138 & n1431 ) | ( n940 & n1431 ) ;
  assign n1433 = x148 ^ x45 ^ x42 ;
  assign n1434 = ( ~x87 & n1432 ) | ( ~x87 & n1433 ) | ( n1432 & n1433 ) ;
  assign n1435 = n1434 ^ n650 ^ n302 ;
  assign n1438 = n490 & n1437 ;
  assign n1439 = n1435 & n1438 ;
  assign n1426 = n612 ^ n495 ^ x32 ;
  assign n1427 = ( n783 & n1131 ) | ( n783 & n1426 ) | ( n1131 & n1426 ) ;
  assign n1428 = ( n465 & n1198 ) | ( n465 & n1427 ) | ( n1198 & n1427 ) ;
  assign n1447 = n1446 ^ n1439 ^ n1428 ;
  assign n1448 = ( ~x181 & n402 ) | ( ~x181 & n1122 ) | ( n402 & n1122 ) ;
  assign n1449 = ( n341 & n874 ) | ( n341 & n1448 ) | ( n874 & n1448 ) ;
  assign n1450 = n361 ^ x240 ^ x69 ;
  assign n1451 = ( n436 & n471 ) | ( n436 & n953 ) | ( n471 & n953 ) ;
  assign n1452 = ( n375 & n807 ) | ( n375 & ~n1451 ) | ( n807 & ~n1451 ) ;
  assign n1453 = n265 & n1452 ;
  assign n1454 = ~n521 & n1453 ;
  assign n1455 = n1450 & ~n1454 ;
  assign n1456 = ~n752 & n1455 ;
  assign n1459 = ( x139 & n615 ) | ( x139 & n1367 ) | ( n615 & n1367 ) ;
  assign n1460 = n1459 ^ n668 ^ 1'b0 ;
  assign n1457 = n542 ^ n369 ^ x189 ;
  assign n1458 = n1457 ^ n972 ^ n940 ;
  assign n1461 = n1460 ^ n1458 ^ n833 ;
  assign n1462 = n1461 ^ n545 ^ 1'b0 ;
  assign n1463 = n1178 | n1462 ;
  assign n1464 = ( n310 & ~n334 ) | ( n310 & n578 ) | ( ~n334 & n578 ) ;
  assign n1465 = n1464 ^ n1284 ^ n430 ;
  assign n1466 = n1078 ^ x9 ^ 1'b0 ;
  assign n1467 = n1465 & ~n1466 ;
  assign n1468 = n540 ^ n428 ^ n371 ;
  assign n1469 = ( n901 & ~n1397 ) | ( n901 & n1468 ) | ( ~n1397 & n1468 ) ;
  assign n1470 = n1467 & n1469 ;
  assign n1473 = ( x196 & n346 ) | ( x196 & n411 ) | ( n346 & n411 ) ;
  assign n1474 = ( n907 & n1067 ) | ( n907 & ~n1473 ) | ( n1067 & ~n1473 ) ;
  assign n1475 = n1474 ^ n1209 ^ x70 ;
  assign n1471 = n1074 ^ n763 ^ x194 ;
  assign n1472 = n1471 ^ n1248 ^ n547 ;
  assign n1476 = n1475 ^ n1472 ^ n257 ;
  assign n1489 = ( x231 & n324 ) | ( x231 & ~n363 ) | ( n324 & ~n363 ) ;
  assign n1484 = ( ~x130 & x213 ) | ( ~x130 & n625 ) | ( x213 & n625 ) ;
  assign n1485 = n1484 ^ x89 ^ 1'b0 ;
  assign n1486 = n1085 & ~n1485 ;
  assign n1487 = n1486 ^ n772 ^ 1'b0 ;
  assign n1477 = n891 ^ n726 ^ 1'b0 ;
  assign n1478 = ( n464 & n1067 ) | ( n464 & n1173 ) | ( n1067 & n1173 ) ;
  assign n1479 = n1478 ^ n1358 ^ n1171 ;
  assign n1480 = n890 & ~n1479 ;
  assign n1481 = ~n1282 & n1480 ;
  assign n1482 = ( n825 & n1477 ) | ( n825 & ~n1481 ) | ( n1477 & ~n1481 ) ;
  assign n1483 = n1325 & n1482 ;
  assign n1488 = n1487 ^ n1483 ^ 1'b0 ;
  assign n1490 = n1489 ^ n1488 ^ x196 ;
  assign n1491 = ( x62 & n562 ) | ( x62 & n736 ) | ( n562 & n736 ) ;
  assign n1492 = ( ~n941 & n1490 ) | ( ~n941 & n1491 ) | ( n1490 & n1491 ) ;
  assign n1493 = n807 & ~n971 ;
  assign n1494 = n930 & n1493 ;
  assign n1495 = n1494 ^ n684 ^ x235 ;
  assign n1503 = ( n292 & ~n439 ) | ( n292 & n673 ) | ( ~n439 & n673 ) ;
  assign n1502 = ( x113 & n660 ) | ( x113 & n1184 ) | ( n660 & n1184 ) ;
  assign n1504 = n1503 ^ n1502 ^ x214 ;
  assign n1501 = ( ~x23 & n261 ) | ( ~x23 & n319 ) | ( n261 & n319 ) ;
  assign n1505 = n1504 ^ n1501 ^ x31 ;
  assign n1506 = n1505 ^ n510 ^ x208 ;
  assign n1496 = n988 ^ n680 ^ n593 ;
  assign n1497 = n360 ^ x248 ^ 1'b0 ;
  assign n1498 = n1497 ^ n1485 ^ n379 ;
  assign n1499 = ( x108 & n1496 ) | ( x108 & ~n1498 ) | ( n1496 & ~n1498 ) ;
  assign n1500 = n1499 ^ n1039 ^ n449 ;
  assign n1507 = n1506 ^ n1500 ^ n1044 ;
  assign n1508 = x233 ^ x143 ^ 1'b0 ;
  assign n1509 = x201 & n1508 ;
  assign n1510 = ( n812 & n1293 ) | ( n812 & ~n1509 ) | ( n1293 & ~n1509 ) ;
  assign n1511 = ( n311 & ~n833 ) | ( n311 & n946 ) | ( ~n833 & n946 ) ;
  assign n1512 = n727 ^ n256 ^ x104 ;
  assign n1513 = n1291 & ~n1512 ;
  assign n1514 = n1511 & n1513 ;
  assign n1515 = ( n1024 & ~n1394 ) | ( n1024 & n1477 ) | ( ~n1394 & n1477 ) ;
  assign n1518 = ( x59 & n532 ) | ( x59 & n1142 ) | ( n532 & n1142 ) ;
  assign n1519 = n1518 ^ n1368 ^ x28 ;
  assign n1516 = n298 | n371 ;
  assign n1517 = n1516 ^ n1512 ^ 1'b0 ;
  assign n1520 = n1519 ^ n1517 ^ 1'b0 ;
  assign n1521 = ~n1515 & n1520 ;
  assign n1522 = n1184 ^ n401 ^ x115 ;
  assign n1523 = ( n922 & n931 ) | ( n922 & ~n1522 ) | ( n931 & ~n1522 ) ;
  assign n1524 = ( ~x45 & n571 ) | ( ~x45 & n578 ) | ( n571 & n578 ) ;
  assign n1525 = ~n1523 & n1524 ;
  assign n1526 = n466 & n1525 ;
  assign n1527 = ( x50 & ~n621 ) | ( x50 & n1085 ) | ( ~n621 & n1085 ) ;
  assign n1528 = ( n1521 & n1526 ) | ( n1521 & ~n1527 ) | ( n1526 & ~n1527 ) ;
  assign n1529 = ( n887 & n1514 ) | ( n887 & ~n1528 ) | ( n1514 & ~n1528 ) ;
  assign n1539 = n638 ^ n322 ^ n277 ;
  assign n1536 = ( ~x74 & n627 ) | ( ~x74 & n932 ) | ( n627 & n932 ) ;
  assign n1537 = x252 ^ x134 ^ x50 ;
  assign n1538 = ( ~n674 & n1536 ) | ( ~n674 & n1537 ) | ( n1536 & n1537 ) ;
  assign n1535 = n953 ^ x29 ^ x16 ;
  assign n1540 = n1539 ^ n1538 ^ n1535 ;
  assign n1530 = ( n264 & n442 ) | ( n264 & ~n863 ) | ( n442 & ~n863 ) ;
  assign n1531 = n1299 ^ n982 ^ n577 ;
  assign n1532 = n1531 ^ n1248 ^ n561 ;
  assign n1533 = n931 ^ n915 ^ x240 ;
  assign n1534 = ( ~n1530 & n1532 ) | ( ~n1530 & n1533 ) | ( n1532 & n1533 ) ;
  assign n1541 = n1540 ^ n1534 ^ n1416 ;
  assign n1542 = n434 ^ x89 ^ 1'b0 ;
  assign n1543 = ( x109 & n934 ) | ( x109 & ~n1542 ) | ( n934 & ~n1542 ) ;
  assign n1544 = ( x198 & n800 ) | ( x198 & ~n959 ) | ( n800 & ~n959 ) ;
  assign n1545 = ( x45 & ~n1543 ) | ( x45 & n1544 ) | ( ~n1543 & n1544 ) ;
  assign n1546 = n1545 ^ n1115 ^ n435 ;
  assign n1547 = n905 ^ n617 ^ x29 ;
  assign n1548 = ( ~n269 & n989 ) | ( ~n269 & n1547 ) | ( n989 & n1547 ) ;
  assign n1549 = ( n671 & n901 ) | ( n671 & ~n1496 ) | ( n901 & ~n1496 ) ;
  assign n1550 = n1549 ^ n1443 ^ n334 ;
  assign n1551 = ( ~x201 & x226 ) | ( ~x201 & n1025 ) | ( x226 & n1025 ) ;
  assign n1552 = n1437 ^ n1370 ^ x64 ;
  assign n1553 = ( x42 & n1551 ) | ( x42 & n1552 ) | ( n1551 & n1552 ) ;
  assign n1555 = n650 ^ n530 ^ n340 ;
  assign n1556 = n1035 ^ n643 ^ 1'b0 ;
  assign n1557 = n1556 ^ n817 ^ n628 ;
  assign n1558 = ( n848 & ~n1014 ) | ( n848 & n1557 ) | ( ~n1014 & n1557 ) ;
  assign n1559 = ( n488 & n1555 ) | ( n488 & ~n1558 ) | ( n1555 & ~n1558 ) ;
  assign n1560 = n1559 ^ n1089 ^ n957 ;
  assign n1554 = x228 & ~n1427 ;
  assign n1561 = n1560 ^ n1554 ^ 1'b0 ;
  assign n1562 = n1553 | n1561 ;
  assign n1581 = n847 ^ n651 ^ x37 ;
  assign n1582 = ( x42 & n264 ) | ( x42 & n765 ) | ( n264 & n765 ) ;
  assign n1583 = ( n1048 & n1277 ) | ( n1048 & ~n1582 ) | ( n1277 & ~n1582 ) ;
  assign n1584 = ( ~n277 & n1581 ) | ( ~n277 & n1583 ) | ( n1581 & n1583 ) ;
  assign n1563 = n561 ^ x232 ^ x170 ;
  assign n1564 = n1563 ^ n1013 ^ 1'b0 ;
  assign n1565 = x51 | n921 ;
  assign n1566 = ~n1055 & n1194 ;
  assign n1567 = n1566 ^ n1010 ^ n801 ;
  assign n1568 = n1159 ^ n709 ^ 1'b0 ;
  assign n1569 = n624 & n1568 ;
  assign n1570 = ( n1244 & n1567 ) | ( n1244 & ~n1569 ) | ( n1567 & ~n1569 ) ;
  assign n1571 = ( n1564 & n1565 ) | ( n1564 & ~n1570 ) | ( n1565 & ~n1570 ) ;
  assign n1572 = n609 ^ n414 ^ n299 ;
  assign n1573 = ( x84 & n613 ) | ( x84 & n1572 ) | ( n613 & n1572 ) ;
  assign n1574 = n785 & ~n1573 ;
  assign n1575 = n1274 ^ x107 ^ 1'b0 ;
  assign n1576 = n1575 ^ n1367 ^ n599 ;
  assign n1577 = n1576 ^ x110 ^ 1'b0 ;
  assign n1578 = n1577 ^ n1403 ^ n914 ;
  assign n1579 = n1578 ^ n897 ^ n379 ;
  assign n1580 = ( n1571 & n1574 ) | ( n1571 & n1579 ) | ( n1574 & n1579 ) ;
  assign n1585 = n1584 ^ n1580 ^ 1'b0 ;
  assign n1587 = ( n426 & ~n927 ) | ( n426 & n1250 ) | ( ~n927 & n1250 ) ;
  assign n1586 = ( ~x160 & n351 ) | ( ~x160 & n378 ) | ( n351 & n378 ) ;
  assign n1588 = n1587 ^ n1586 ^ n371 ;
  assign n1593 = ( ~x75 & x136 ) | ( ~x75 & n360 ) | ( x136 & n360 ) ;
  assign n1591 = n799 ^ n619 ^ x134 ;
  assign n1589 = n1345 ^ n1314 ^ n734 ;
  assign n1590 = n866 | n1589 ;
  assign n1592 = n1591 ^ n1590 ^ n1154 ;
  assign n1594 = n1593 ^ n1592 ^ n831 ;
  assign n1595 = n730 ^ n715 ^ n602 ;
  assign n1596 = n1595 ^ n983 ^ n633 ;
  assign n1597 = ( n1072 & n1314 ) | ( n1072 & n1596 ) | ( n1314 & n1596 ) ;
  assign n1598 = ( ~n297 & n1594 ) | ( ~n297 & n1597 ) | ( n1594 & n1597 ) ;
  assign n1600 = ( x77 & ~n428 ) | ( x77 & n544 ) | ( ~n428 & n544 ) ;
  assign n1601 = n1600 ^ n730 ^ x104 ;
  assign n1602 = ( n1028 & n1053 ) | ( n1028 & ~n1601 ) | ( n1053 & ~n1601 ) ;
  assign n1599 = ( x78 & x232 ) | ( x78 & ~n925 ) | ( x232 & ~n925 ) ;
  assign n1603 = n1602 ^ n1599 ^ n437 ;
  assign n1604 = n545 | n909 ;
  assign n1605 = n985 | n1604 ;
  assign n1607 = ( n757 & n1047 ) | ( n757 & ~n1173 ) | ( n1047 & ~n1173 ) ;
  assign n1606 = n1376 ^ n1325 ^ x119 ;
  assign n1608 = n1607 ^ n1606 ^ n530 ;
  assign n1609 = ( n354 & ~n1531 ) | ( n354 & n1608 ) | ( ~n1531 & n1608 ) ;
  assign n1610 = n1609 ^ n427 ^ x205 ;
  assign n1611 = ( ~x137 & n1605 ) | ( ~x137 & n1610 ) | ( n1605 & n1610 ) ;
  assign n1614 = n588 ^ n383 ^ x190 ;
  assign n1612 = n1060 ^ n416 ^ x197 ;
  assign n1613 = ( n654 & n871 ) | ( n654 & n1612 ) | ( n871 & n1612 ) ;
  assign n1615 = n1614 ^ n1613 ^ n379 ;
  assign n1616 = n1615 ^ x250 ^ 1'b0 ;
  assign n1617 = ~n358 & n1616 ;
  assign n1628 = ( x26 & ~x53 ) | ( x26 & n552 ) | ( ~x53 & n552 ) ;
  assign n1629 = n1628 ^ n949 ^ x133 ;
  assign n1618 = n1289 ^ n1056 ^ n499 ;
  assign n1619 = n371 ^ x191 ^ x71 ;
  assign n1620 = n502 ^ n263 ^ x247 ;
  assign n1621 = ( x61 & ~n831 ) | ( x61 & n1620 ) | ( ~n831 & n1620 ) ;
  assign n1622 = ( x12 & ~n1619 ) | ( x12 & n1621 ) | ( ~n1619 & n1621 ) ;
  assign n1623 = ( ~x62 & x121 ) | ( ~x62 & n1622 ) | ( x121 & n1622 ) ;
  assign n1624 = n737 ^ n273 ^ 1'b0 ;
  assign n1625 = n1624 ^ n877 ^ 1'b0 ;
  assign n1626 = n830 & ~n1625 ;
  assign n1627 = ( n1618 & n1623 ) | ( n1618 & ~n1626 ) | ( n1623 & ~n1626 ) ;
  assign n1630 = n1629 ^ n1627 ^ n1443 ;
  assign n1631 = n932 ^ x72 ^ 1'b0 ;
  assign n1632 = n1631 ^ n1271 ^ n298 ;
  assign n1633 = n546 ^ n457 ^ n294 ;
  assign n1634 = n1633 ^ n527 ^ n362 ;
  assign n1635 = n1634 ^ n937 ^ 1'b0 ;
  assign n1636 = n1632 | n1635 ;
  assign n1637 = n1033 ^ n1005 ^ x36 ;
  assign n1638 = n971 ^ n869 ^ n384 ;
  assign n1639 = ( n1030 & n1637 ) | ( n1030 & n1638 ) | ( n1637 & n1638 ) ;
  assign n1640 = ( x247 & ~n665 ) | ( x247 & n1274 ) | ( ~n665 & n1274 ) ;
  assign n1641 = n1640 ^ n919 ^ n423 ;
  assign n1642 = x67 & n728 ;
  assign n1643 = ~n1641 & n1642 ;
  assign n1644 = ~x86 & n1450 ;
  assign n1645 = n1644 ^ n1227 ^ n1123 ;
  assign n1648 = n306 ^ x173 ^ x118 ;
  assign n1646 = n422 ^ n333 ^ n310 ;
  assign n1647 = ( n411 & n603 ) | ( n411 & ~n1646 ) | ( n603 & ~n1646 ) ;
  assign n1649 = n1648 ^ n1647 ^ n1382 ;
  assign n1650 = n1649 ^ n1137 ^ n686 ;
  assign n1651 = ( n874 & n1645 ) | ( n874 & ~n1650 ) | ( n1645 & ~n1650 ) ;
  assign n1652 = ~n1643 & n1651 ;
  assign n1653 = n399 ^ x162 ^ x143 ;
  assign n1654 = ( n678 & ~n1446 ) | ( n678 & n1653 ) | ( ~n1446 & n1653 ) ;
  assign n1655 = ( ~n961 & n1410 ) | ( ~n961 & n1654 ) | ( n1410 & n1654 ) ;
  assign n1656 = ( x50 & n885 ) | ( x50 & n1595 ) | ( n885 & n1595 ) ;
  assign n1657 = n1656 ^ n1547 ^ n393 ;
  assign n1658 = ( n964 & n1014 ) | ( n964 & ~n1657 ) | ( n1014 & ~n1657 ) ;
  assign n1659 = n1658 ^ n404 ^ n313 ;
  assign n1660 = n456 ^ x228 ^ x6 ;
  assign n1661 = ( x209 & ~n1035 ) | ( x209 & n1660 ) | ( ~n1035 & n1660 ) ;
  assign n1662 = n1661 ^ n1337 ^ n831 ;
  assign n1663 = n1662 ^ n618 ^ n507 ;
  assign n1664 = n1659 | n1663 ;
  assign n1665 = n950 ^ n302 ^ x244 ;
  assign n1666 = ( x12 & ~n1414 ) | ( x12 & n1665 ) | ( ~n1414 & n1665 ) ;
  assign n1667 = ( x183 & n748 ) | ( x183 & ~n973 ) | ( n748 & ~n973 ) ;
  assign n1668 = ( ~x249 & n451 ) | ( ~x249 & n1593 ) | ( n451 & n1593 ) ;
  assign n1669 = n547 | n1668 ;
  assign n1670 = n1669 ^ n1538 ^ 1'b0 ;
  assign n1671 = ( x241 & n1290 ) | ( x241 & ~n1670 ) | ( n1290 & ~n1670 ) ;
  assign n1672 = ( n1666 & n1667 ) | ( n1666 & n1671 ) | ( n1667 & n1671 ) ;
  assign n1675 = n551 & ~n775 ;
  assign n1676 = ~n698 & n1675 ;
  assign n1677 = n1676 ^ n618 ^ n340 ;
  assign n1673 = n542 ^ n462 ^ 1'b0 ;
  assign n1674 = n1673 ^ n258 ^ x223 ;
  assign n1678 = n1677 ^ n1674 ^ n1242 ;
  assign n1679 = n806 | n1269 ;
  assign n1680 = n1679 ^ n1645 ^ 1'b0 ;
  assign n1681 = ( n1396 & n1678 ) | ( n1396 & n1680 ) | ( n1678 & n1680 ) ;
  assign n1682 = n909 ^ n728 ^ x249 ;
  assign n1683 = n983 ^ x199 ^ x172 ;
  assign n1684 = n1367 ^ n559 ^ n421 ;
  assign n1685 = n527 & n1684 ;
  assign n1686 = ~n1683 & n1685 ;
  assign n1687 = ( ~x105 & n388 ) | ( ~x105 & n1686 ) | ( n388 & n1686 ) ;
  assign n1688 = n660 ^ n452 ^ n324 ;
  assign n1689 = ( ~n418 & n1271 ) | ( ~n418 & n1688 ) | ( n1271 & n1688 ) ;
  assign n1690 = ( n326 & ~n426 ) | ( n326 & n905 ) | ( ~n426 & n905 ) ;
  assign n1691 = ( ~n1235 & n1426 ) | ( ~n1235 & n1690 ) | ( n1426 & n1690 ) ;
  assign n1700 = n1587 ^ n1264 ^ x170 ;
  assign n1694 = n420 ^ n354 ^ x41 ;
  assign n1695 = n1694 ^ n595 ^ n579 ;
  assign n1692 = n834 ^ x15 ^ 1'b0 ;
  assign n1693 = n554 & n1692 ;
  assign n1696 = n1695 ^ n1693 ^ n947 ;
  assign n1697 = ( n329 & n337 ) | ( n329 & ~n956 ) | ( n337 & ~n956 ) ;
  assign n1698 = n1697 ^ n653 ^ n593 ;
  assign n1699 = n1696 & n1698 ;
  assign n1701 = n1700 ^ n1699 ^ 1'b0 ;
  assign n1712 = n423 & ~n1618 ;
  assign n1713 = n547 ^ x127 ^ 1'b0 ;
  assign n1714 = n646 | n1713 ;
  assign n1715 = x193 & ~n386 ;
  assign n1716 = ~x43 & n1715 ;
  assign n1717 = n1716 ^ n766 ^ n317 ;
  assign n1718 = ( n383 & n1714 ) | ( n383 & n1717 ) | ( n1714 & n1717 ) ;
  assign n1720 = x99 ^ x70 ^ x39 ;
  assign n1719 = ( ~x36 & n288 ) | ( ~x36 & n807 ) | ( n288 & n807 ) ;
  assign n1721 = n1720 ^ n1719 ^ 1'b0 ;
  assign n1722 = x138 & n1721 ;
  assign n1723 = ~n849 & n1722 ;
  assign n1724 = ~x106 & n1723 ;
  assign n1725 = ( n1712 & ~n1718 ) | ( n1712 & n1724 ) | ( ~n1718 & n1724 ) ;
  assign n1726 = n1725 ^ n852 ^ n643 ;
  assign n1702 = n682 ^ n449 ^ x153 ;
  assign n1703 = n1012 & ~n1702 ;
  assign n1704 = n378 & n1703 ;
  assign n1705 = n516 ^ n506 ^ n343 ;
  assign n1707 = ( n765 & n985 ) | ( n765 & ~n1622 ) | ( n985 & ~n1622 ) ;
  assign n1706 = ( x49 & n438 ) | ( x49 & ~n1349 ) | ( n438 & ~n1349 ) ;
  assign n1708 = n1707 ^ n1706 ^ n1135 ;
  assign n1709 = ( n1242 & ~n1705 ) | ( n1242 & n1708 ) | ( ~n1705 & n1708 ) ;
  assign n1710 = ( n647 & n1704 ) | ( n647 & ~n1709 ) | ( n1704 & ~n1709 ) ;
  assign n1711 = n1710 ^ n1537 ^ n734 ;
  assign n1727 = n1726 ^ n1711 ^ x173 ;
  assign n1732 = ( x174 & n868 ) | ( x174 & ~n1275 ) | ( n868 & ~n1275 ) ;
  assign n1733 = ( x114 & n1431 ) | ( x114 & n1732 ) | ( n1431 & n1732 ) ;
  assign n1730 = n862 ^ n561 ^ n271 ;
  assign n1728 = n324 ^ x31 ^ 1'b0 ;
  assign n1729 = ~n1005 & n1728 ;
  assign n1731 = n1730 ^ n1729 ^ n775 ;
  assign n1734 = n1733 ^ n1731 ^ n1133 ;
  assign n1735 = ( x39 & ~n391 ) | ( x39 & n692 ) | ( ~n391 & n692 ) ;
  assign n1736 = x104 & ~n1735 ;
  assign n1737 = n678 & n1736 ;
  assign n1751 = n343 ^ x196 ^ x60 ;
  assign n1752 = ( n343 & ~n437 ) | ( n343 & n1751 ) | ( ~n437 & n1751 ) ;
  assign n1753 = n1752 ^ n1720 ^ 1'b0 ;
  assign n1754 = n884 | n1753 ;
  assign n1738 = n945 ^ n400 ^ x42 ;
  assign n1739 = n1738 ^ n1236 ^ n444 ;
  assign n1740 = n1358 ^ n991 ^ n787 ;
  assign n1741 = ( n340 & ~n1479 ) | ( n340 & n1740 ) | ( ~n1479 & n1740 ) ;
  assign n1742 = ( n301 & n1739 ) | ( n301 & n1741 ) | ( n1739 & n1741 ) ;
  assign n1743 = ~n921 & n1638 ;
  assign n1744 = n1743 ^ n853 ^ 1'b0 ;
  assign n1745 = ( n1243 & ~n1381 ) | ( n1243 & n1744 ) | ( ~n1381 & n1744 ) ;
  assign n1746 = n479 ^ n355 ^ n294 ;
  assign n1747 = ( ~x123 & x216 ) | ( ~x123 & n512 ) | ( x216 & n512 ) ;
  assign n1748 = n1747 ^ n566 ^ n379 ;
  assign n1749 = ( n1059 & n1746 ) | ( n1059 & ~n1748 ) | ( n1746 & ~n1748 ) ;
  assign n1750 = ( ~n1742 & n1745 ) | ( ~n1742 & n1749 ) | ( n1745 & n1749 ) ;
  assign n1755 = n1754 ^ n1750 ^ 1'b0 ;
  assign n1756 = ( ~n629 & n1737 ) | ( ~n629 & n1755 ) | ( n1737 & n1755 ) ;
  assign n1758 = ( x28 & ~x135 ) | ( x28 & x143 ) | ( ~x135 & x143 ) ;
  assign n1757 = n1747 ^ n428 ^ x37 ;
  assign n1759 = n1758 ^ n1757 ^ n1308 ;
  assign n1760 = n1759 ^ n1505 ^ x69 ;
  assign n1765 = n356 & ~n1279 ;
  assign n1766 = n1765 ^ x148 ^ 1'b0 ;
  assign n1761 = ( x174 & ~n291 ) | ( x174 & n358 ) | ( ~n291 & n358 ) ;
  assign n1762 = n404 ^ n370 ^ x36 ;
  assign n1763 = ( n660 & n1761 ) | ( n660 & ~n1762 ) | ( n1761 & ~n1762 ) ;
  assign n1764 = ( x167 & n1602 ) | ( x167 & n1763 ) | ( n1602 & n1763 ) ;
  assign n1767 = n1766 ^ n1764 ^ n781 ;
  assign n1768 = n1767 ^ n1746 ^ n1432 ;
  assign n1777 = n756 ^ n585 ^ x254 ;
  assign n1769 = x105 & ~n313 ;
  assign n1770 = ~x44 & n1769 ;
  assign n1771 = n1770 ^ n1530 ^ n548 ;
  assign n1772 = n1771 ^ n882 ^ n659 ;
  assign n1773 = x200 & n296 ;
  assign n1774 = ~n1297 & n1773 ;
  assign n1775 = n1052 ^ n721 ^ n595 ;
  assign n1776 = ( n1772 & ~n1774 ) | ( n1772 & n1775 ) | ( ~n1774 & n1775 ) ;
  assign n1778 = n1777 ^ n1776 ^ n1526 ;
  assign n1779 = ( n969 & n1614 ) | ( n969 & n1778 ) | ( n1614 & n1778 ) ;
  assign n1780 = ( ~n1760 & n1768 ) | ( ~n1760 & n1779 ) | ( n1768 & n1779 ) ;
  assign n1781 = ( n880 & n1137 ) | ( n880 & n1381 ) | ( n1137 & n1381 ) ;
  assign n1782 = n1172 ^ n709 ^ 1'b0 ;
  assign n1783 = ~n1415 & n1782 ;
  assign n1784 = ( ~n1322 & n1781 ) | ( ~n1322 & n1783 ) | ( n1781 & n1783 ) ;
  assign n1785 = ( n287 & n504 ) | ( n287 & n837 ) | ( n504 & n837 ) ;
  assign n1786 = n461 ^ n423 ^ x5 ;
  assign n1787 = ( n383 & ~n546 ) | ( n383 & n1786 ) | ( ~n546 & n1786 ) ;
  assign n1788 = ( n1431 & ~n1785 ) | ( n1431 & n1787 ) | ( ~n1785 & n1787 ) ;
  assign n1789 = n1788 ^ n1661 ^ n1510 ;
  assign n1794 = ~n805 & n946 ;
  assign n1790 = n1496 ^ n862 ^ n597 ;
  assign n1791 = n1790 ^ n1684 ^ 1'b0 ;
  assign n1792 = n1018 & n1791 ;
  assign n1793 = ( ~n1063 & n1073 ) | ( ~n1063 & n1792 ) | ( n1073 & n1792 ) ;
  assign n1795 = n1794 ^ n1793 ^ n1178 ;
  assign n1803 = n1297 ^ n444 ^ x251 ;
  assign n1800 = ( n736 & n985 ) | ( n736 & n995 ) | ( n985 & n995 ) ;
  assign n1801 = n1593 & ~n1800 ;
  assign n1802 = n1801 ^ n439 ^ x206 ;
  assign n1796 = ( ~n633 & n1409 ) | ( ~n633 & n1512 ) | ( n1409 & n1512 ) ;
  assign n1797 = ( ~x135 & n311 ) | ( ~x135 & n1796 ) | ( n311 & n1796 ) ;
  assign n1798 = n1797 ^ n1378 ^ 1'b0 ;
  assign n1799 = ~n370 & n1798 ;
  assign n1804 = n1803 ^ n1802 ^ n1799 ;
  assign n1805 = ( x220 & n1321 ) | ( x220 & ~n1351 ) | ( n1321 & ~n1351 ) ;
  assign n1806 = n1501 ^ n514 ^ x165 ;
  assign n1807 = ( x1 & n1751 ) | ( x1 & ~n1806 ) | ( n1751 & ~n1806 ) ;
  assign n1808 = n1807 ^ n400 ^ x234 ;
  assign n1809 = n1062 ^ n752 ^ n376 ;
  assign n1810 = x201 ^ x197 ^ 1'b0 ;
  assign n1811 = ( ~n1282 & n1809 ) | ( ~n1282 & n1810 ) | ( n1809 & n1810 ) ;
  assign n1812 = n1811 ^ n1448 ^ n520 ;
  assign n1813 = ( n345 & n815 ) | ( n345 & n1180 ) | ( n815 & n1180 ) ;
  assign n1822 = n1751 ^ n870 ^ n540 ;
  assign n1823 = n1822 ^ n937 ^ x189 ;
  assign n1820 = n525 | n582 ;
  assign n1821 = x227 | n1820 ;
  assign n1817 = n1593 ^ x79 ^ 1'b0 ;
  assign n1814 = ( x70 & n587 ) | ( x70 & n910 ) | ( n587 & n910 ) ;
  assign n1815 = n537 & n1814 ;
  assign n1816 = n1815 ^ n1300 ^ 1'b0 ;
  assign n1818 = n1817 ^ n1816 ^ n1230 ;
  assign n1819 = n745 & ~n1818 ;
  assign n1824 = n1823 ^ n1821 ^ n1819 ;
  assign n1826 = x17 & ~n423 ;
  assign n1827 = n1826 ^ n643 ^ 1'b0 ;
  assign n1825 = ( ~n545 & n1115 ) | ( ~n545 & n1665 ) | ( n1115 & n1665 ) ;
  assign n1828 = n1827 ^ n1825 ^ x239 ;
  assign n1829 = n1828 ^ n1587 ^ n483 ;
  assign n1830 = n1829 ^ x185 ^ x83 ;
  assign n1831 = n1161 ^ n619 ^ n324 ;
  assign n1832 = n1831 ^ x7 ^ 1'b0 ;
  assign n1833 = n993 & ~n1832 ;
  assign n1834 = ( ~n659 & n1830 ) | ( ~n659 & n1833 ) | ( n1830 & n1833 ) ;
  assign n1836 = ( ~x25 & n529 ) | ( ~x25 & n791 ) | ( n529 & n791 ) ;
  assign n1835 = n1474 ^ n955 ^ n725 ;
  assign n1837 = n1836 ^ n1835 ^ n1262 ;
  assign n1838 = ( n667 & n964 ) | ( n667 & ~n1600 ) | ( n964 & ~n1600 ) ;
  assign n1839 = n1838 ^ n700 ^ x168 ;
  assign n1840 = ( n1239 & n1837 ) | ( n1239 & ~n1839 ) | ( n1837 & ~n1839 ) ;
  assign n1841 = n581 ^ x93 ^ x33 ;
  assign n1842 = n1841 ^ n834 ^ n556 ;
  assign n1843 = n740 ^ n568 ^ n325 ;
  assign n1844 = n1843 ^ n342 ^ x155 ;
  assign n1845 = ( x128 & n956 ) | ( x128 & ~n1844 ) | ( n956 & ~n1844 ) ;
  assign n1846 = n1845 ^ n309 ^ x193 ;
  assign n1847 = ( n1188 & ~n1842 ) | ( n1188 & n1846 ) | ( ~n1842 & n1846 ) ;
  assign n1848 = n1847 ^ n1061 ^ n979 ;
  assign n1850 = n674 ^ n512 ^ x34 ;
  assign n1849 = n1300 ^ x138 ^ x23 ;
  assign n1851 = n1850 ^ n1849 ^ x25 ;
  assign n1852 = ( x155 & ~n1848 ) | ( x155 & n1851 ) | ( ~n1848 & n1851 ) ;
  assign n1853 = ( ~n537 & n666 ) | ( ~n537 & n1496 ) | ( n666 & n1496 ) ;
  assign n1861 = n1572 ^ x239 ^ 1'b0 ;
  assign n1862 = n1861 ^ n1460 ^ n505 ;
  assign n1863 = n1862 ^ n1226 ^ n1137 ;
  assign n1854 = ~n420 & n1001 ;
  assign n1855 = n446 & n1854 ;
  assign n1856 = n1082 ^ n858 ^ n372 ;
  assign n1857 = x190 ^ x134 ^ 1'b0 ;
  assign n1858 = ~n1856 & n1857 ;
  assign n1859 = ( ~n624 & n1855 ) | ( ~n624 & n1858 ) | ( n1855 & n1858 ) ;
  assign n1860 = x242 & ~n1859 ;
  assign n1864 = n1863 ^ n1860 ^ 1'b0 ;
  assign n1866 = n449 ^ n256 ^ x100 ;
  assign n1867 = n1511 & n1866 ;
  assign n1868 = ~n1761 & n1867 ;
  assign n1865 = ( n533 & n689 ) | ( n533 & n1707 ) | ( n689 & n1707 ) ;
  assign n1869 = n1868 ^ n1865 ^ x234 ;
  assign n1870 = n1802 ^ n1614 ^ n486 ;
  assign n1871 = n1869 | n1870 ;
  assign n1872 = n1871 ^ n1464 ^ 1'b0 ;
  assign n1873 = x201 & ~n1872 ;
  assign n1874 = n859 ^ n816 ^ n410 ;
  assign n1875 = n391 | n1874 ;
  assign n1876 = ~n546 & n1875 ;
  assign n1877 = ~n835 & n1876 ;
  assign n1878 = n1877 ^ n1704 ^ 1'b0 ;
  assign n1879 = n785 & n1878 ;
  assign n1880 = n1645 ^ n1211 ^ x216 ;
  assign n1881 = n1761 ^ n658 ^ x201 ;
  assign n1882 = n1022 ^ n934 ^ 1'b0 ;
  assign n1883 = n1881 & n1882 ;
  assign n1884 = n1883 ^ n1640 ^ n753 ;
  assign n1885 = n352 & ~n1884 ;
  assign n1886 = n1885 ^ n1555 ^ 1'b0 ;
  assign n1887 = n997 ^ x167 ^ 1'b0 ;
  assign n1888 = ( x179 & n806 ) | ( x179 & n1887 ) | ( n806 & n1887 ) ;
  assign n1889 = ( n1880 & ~n1886 ) | ( n1880 & n1888 ) | ( ~n1886 & n1888 ) ;
  assign n1890 = x43 & n434 ;
  assign n1891 = n1890 ^ n487 ^ 1'b0 ;
  assign n1892 = n1891 ^ n259 ^ 1'b0 ;
  assign n1893 = n541 ^ n507 ^ n311 ;
  assign n1894 = n559 | n891 ;
  assign n1895 = n1894 ^ n350 ^ x48 ;
  assign n1896 = ( n336 & n1893 ) | ( n336 & n1895 ) | ( n1893 & n1895 ) ;
  assign n1897 = n444 ^ x244 ^ x9 ;
  assign n1898 = ( ~n620 & n653 ) | ( ~n620 & n1897 ) | ( n653 & n1897 ) ;
  assign n1899 = ( n785 & n1041 ) | ( n785 & ~n1898 ) | ( n1041 & ~n1898 ) ;
  assign n1900 = ( n1892 & ~n1896 ) | ( n1892 & n1899 ) | ( ~n1896 & n1899 ) ;
  assign n1901 = ( x98 & ~x130 ) | ( x98 & n605 ) | ( ~x130 & n605 ) ;
  assign n1902 = ( ~x164 & n393 ) | ( ~x164 & n1901 ) | ( n393 & n1901 ) ;
  assign n1903 = ( x231 & x237 ) | ( x231 & n1902 ) | ( x237 & n1902 ) ;
  assign n1904 = n1903 ^ n775 ^ 1'b0 ;
  assign n1905 = n1904 ^ n1489 ^ n1248 ;
  assign n1906 = ( ~n1889 & n1900 ) | ( ~n1889 & n1905 ) | ( n1900 & n1905 ) ;
  assign n1907 = n406 | n814 ;
  assign n1908 = x82 & n890 ;
  assign n1909 = ~n638 & n1908 ;
  assign n1910 = ( n546 & n706 ) | ( n546 & ~n1909 ) | ( n706 & ~n1909 ) ;
  assign n1911 = ~n768 & n1405 ;
  assign n1912 = n1911 ^ n1887 ^ n833 ;
  assign n1924 = ( x179 & n646 ) | ( x179 & ~n946 ) | ( n646 & ~n946 ) ;
  assign n1925 = ( n338 & ~n1436 ) | ( n338 & n1512 ) | ( ~n1436 & n1512 ) ;
  assign n1926 = n1925 ^ n1897 ^ n970 ;
  assign n1927 = ( x59 & n817 ) | ( x59 & n1031 ) | ( n817 & n1031 ) ;
  assign n1928 = x116 & ~n1927 ;
  assign n1929 = n1928 ^ n1415 ^ n409 ;
  assign n1930 = ( n1924 & ~n1926 ) | ( n1924 & n1929 ) | ( ~n1926 & n1929 ) ;
  assign n1913 = x186 & ~n277 ;
  assign n1914 = n1913 ^ n925 ^ 1'b0 ;
  assign n1915 = ( x45 & ~x57 ) | ( x45 & n784 ) | ( ~x57 & n784 ) ;
  assign n1916 = n1915 ^ n879 ^ 1'b0 ;
  assign n1917 = ~n1914 & n1916 ;
  assign n1918 = ~n659 & n1803 ;
  assign n1919 = n692 & n1918 ;
  assign n1920 = n1919 ^ x14 ^ 1'b0 ;
  assign n1921 = n722 & ~n1920 ;
  assign n1922 = n1921 ^ n1846 ^ x113 ;
  assign n1923 = n1917 & ~n1922 ;
  assign n1931 = n1930 ^ n1923 ^ 1'b0 ;
  assign n1932 = ( ~n964 & n1912 ) | ( ~n964 & n1931 ) | ( n1912 & n1931 ) ;
  assign n1933 = ( ~n968 & n1910 ) | ( ~n968 & n1932 ) | ( n1910 & n1932 ) ;
  assign n1934 = ( ~n698 & n1539 ) | ( ~n698 & n1763 ) | ( n1539 & n1763 ) ;
  assign n1936 = ( ~n818 & n987 ) | ( ~n818 & n1292 ) | ( n987 & n1292 ) ;
  assign n1935 = n1279 ^ n1189 ^ 1'b0 ;
  assign n1937 = n1936 ^ n1935 ^ n508 ;
  assign n1938 = ( x134 & n655 ) | ( x134 & n1937 ) | ( n655 & n1937 ) ;
  assign n1941 = n1299 ^ n659 ^ n274 ;
  assign n1942 = n1205 & ~n1941 ;
  assign n1943 = n1942 ^ n1850 ^ x158 ;
  assign n1939 = n1801 ^ n659 ^ x19 ;
  assign n1940 = n1449 | n1939 ;
  assign n1944 = n1943 ^ n1940 ^ n256 ;
  assign n1945 = n365 & n719 ;
  assign n1947 = n383 ^ x217 ^ x36 ;
  assign n1946 = ( n1746 & n1764 ) | ( n1746 & n1794 ) | ( n1764 & n1794 ) ;
  assign n1948 = n1947 ^ n1946 ^ n748 ;
  assign n1949 = ( ~n538 & n1160 ) | ( ~n538 & n1948 ) | ( n1160 & n1948 ) ;
  assign n1950 = n580 ^ n491 ^ n426 ;
  assign n1951 = x17 & n1950 ;
  assign n1952 = n1951 ^ n1195 ^ 1'b0 ;
  assign n1959 = n418 ^ x141 ^ x111 ;
  assign n1960 = n1959 ^ n853 ^ n772 ;
  assign n1961 = ( n823 & n1477 ) | ( n823 & ~n1960 ) | ( n1477 & ~n1960 ) ;
  assign n1953 = n374 ^ n339 ^ x12 ;
  assign n1954 = n1796 ^ x241 ^ 1'b0 ;
  assign n1955 = ( n583 & n1953 ) | ( n583 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1956 = ( ~x248 & n1086 ) | ( ~x248 & n1955 ) | ( n1086 & n1955 ) ;
  assign n1957 = ( n329 & n1214 ) | ( n329 & ~n1956 ) | ( n1214 & ~n1956 ) ;
  assign n1958 = ( ~n317 & n910 ) | ( ~n317 & n1957 ) | ( n910 & n1957 ) ;
  assign n1962 = n1961 ^ n1958 ^ n1744 ;
  assign n1963 = ( x26 & n291 ) | ( x26 & ~n500 ) | ( n291 & ~n500 ) ;
  assign n1964 = ( ~n467 & n1962 ) | ( ~n467 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1965 = ( x214 & ~n1952 ) | ( x214 & n1964 ) | ( ~n1952 & n1964 ) ;
  assign n1966 = n1697 ^ x58 ^ 1'b0 ;
  assign n1967 = ( ~x116 & n877 ) | ( ~x116 & n1966 ) | ( n877 & n1966 ) ;
  assign n1969 = ( ~n584 & n762 ) | ( ~n584 & n1484 ) | ( n762 & n1484 ) ;
  assign n1968 = ( n959 & ~n1019 ) | ( n959 & n1284 ) | ( ~n1019 & n1284 ) ;
  assign n1970 = n1969 ^ n1968 ^ n1254 ;
  assign n1971 = n1283 ^ n349 ^ 1'b0 ;
  assign n1972 = ( ~n1967 & n1970 ) | ( ~n1967 & n1971 ) | ( n1970 & n1971 ) ;
  assign n1973 = ( x34 & n912 ) | ( x34 & n1022 ) | ( n912 & n1022 ) ;
  assign n1974 = n1973 ^ n1142 ^ x123 ;
  assign n1975 = n1593 & n1974 ;
  assign n1976 = n1975 ^ n1893 ^ n997 ;
  assign n1977 = ( n832 & n1233 ) | ( n832 & ~n1361 ) | ( n1233 & ~n1361 ) ;
  assign n1978 = n780 ^ n444 ^ 1'b0 ;
  assign n1979 = n1977 & n1978 ;
  assign n1980 = ( n456 & n482 ) | ( n456 & ~n1077 ) | ( n482 & ~n1077 ) ;
  assign n1981 = n1980 ^ x173 ^ 1'b0 ;
  assign n1982 = ( ~n1235 & n1979 ) | ( ~n1235 & n1981 ) | ( n1979 & n1981 ) ;
  assign n1983 = x148 & ~n362 ;
  assign n1984 = ( n1139 & ~n1196 ) | ( n1139 & n1983 ) | ( ~n1196 & n1983 ) ;
  assign n1985 = n1172 & n1984 ;
  assign n1986 = n1985 ^ n1915 ^ n1450 ;
  assign n1987 = ( n321 & ~n640 ) | ( n321 & n1895 ) | ( ~n640 & n1895 ) ;
  assign n1988 = ( n389 & n1411 ) | ( n389 & ~n1464 ) | ( n1411 & ~n1464 ) ;
  assign n1989 = n1988 ^ n467 ^ x37 ;
  assign n1990 = ( ~n1698 & n1915 ) | ( ~n1698 & n1989 ) | ( n1915 & n1989 ) ;
  assign n1991 = ~n597 & n613 ;
  assign n1992 = ( n673 & ~n838 ) | ( n673 & n1991 ) | ( ~n838 & n1991 ) ;
  assign n1993 = n1992 ^ n1720 ^ n905 ;
  assign n1994 = ( x182 & ~n481 ) | ( x182 & n1633 ) | ( ~n481 & n1633 ) ;
  assign n1995 = n1468 ^ n675 ^ 1'b0 ;
  assign n1996 = n1994 & ~n1995 ;
  assign n1997 = ( ~n740 & n1418 ) | ( ~n740 & n1996 ) | ( n1418 & n1996 ) ;
  assign n1998 = ( n1133 & ~n1993 ) | ( n1133 & n1997 ) | ( ~n1993 & n1997 ) ;
  assign n1999 = n1990 & n1998 ;
  assign n2000 = ~n941 & n1999 ;
  assign n2006 = ( ~x182 & n569 ) | ( ~x182 & n817 ) | ( n569 & n817 ) ;
  assign n2007 = n2006 ^ n1509 ^ x107 ;
  assign n2008 = n2007 ^ n1602 ^ 1'b0 ;
  assign n2009 = ~n1189 & n2008 ;
  assign n2001 = n580 ^ x230 ^ x6 ;
  assign n2002 = n1401 ^ n571 ^ n519 ;
  assign n2003 = ( n522 & n1085 ) | ( n522 & ~n2002 ) | ( n1085 & ~n2002 ) ;
  assign n2004 = n2003 ^ n857 ^ x101 ;
  assign n2005 = n2001 | n2004 ;
  assign n2010 = n2009 ^ n2005 ^ 1'b0 ;
  assign n2019 = ( x17 & n502 ) | ( x17 & n1485 ) | ( n502 & n1485 ) ;
  assign n2020 = ( n580 & n642 ) | ( n580 & n1368 ) | ( n642 & n1368 ) ;
  assign n2021 = n2020 ^ n746 ^ n649 ;
  assign n2022 = n2021 ^ n1915 ^ n987 ;
  assign n2023 = ( x97 & n431 ) | ( x97 & ~n2022 ) | ( n431 & ~n2022 ) ;
  assign n2024 = n1275 | n2023 ;
  assign n2025 = n2019 & ~n2024 ;
  assign n2016 = ( n284 & n744 ) | ( n284 & ~n1295 ) | ( n744 & ~n1295 ) ;
  assign n2017 = n2016 ^ n1897 ^ n446 ;
  assign n2011 = ( ~n439 & n1244 ) | ( ~n439 & n1269 ) | ( n1244 & n1269 ) ;
  assign n2012 = ( x66 & x226 ) | ( x66 & n2011 ) | ( x226 & n2011 ) ;
  assign n2013 = n1686 ^ n660 ^ x31 ;
  assign n2014 = ( x170 & n2012 ) | ( x170 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2015 = n2014 ^ n788 ^ 1'b0 ;
  assign n2018 = n2017 ^ n2015 ^ n1644 ;
  assign n2026 = n2025 ^ n2018 ^ x252 ;
  assign n2028 = ( x25 & ~n298 ) | ( x25 & n466 ) | ( ~n298 & n466 ) ;
  assign n2027 = n1670 ^ n1035 ^ n324 ;
  assign n2029 = n2028 ^ n2027 ^ n1197 ;
  assign n2030 = ~n453 & n1220 ;
  assign n2031 = n2030 ^ n1213 ^ 1'b0 ;
  assign n2032 = n1624 ^ n896 ^ 1'b0 ;
  assign n2033 = n391 & n2032 ;
  assign n2034 = n2033 ^ n1929 ^ n881 ;
  assign n2035 = ( n863 & ~n2031 ) | ( n863 & n2034 ) | ( ~n2031 & n2034 ) ;
  assign n2039 = ( n263 & ~n816 ) | ( n263 & n1067 ) | ( ~n816 & n1067 ) ;
  assign n2040 = x148 & n2039 ;
  assign n2041 = ~n1102 & n2040 ;
  assign n2036 = ( ~n287 & n349 ) | ( ~n287 & n1320 ) | ( n349 & n1320 ) ;
  assign n2037 = n2036 ^ n1300 ^ n628 ;
  assign n2038 = n2037 ^ n1055 ^ n495 ;
  assign n2042 = n2041 ^ n2038 ^ n1709 ;
  assign n2046 = x142 & ~n605 ;
  assign n2043 = ( ~n343 & n756 ) | ( ~n343 & n787 ) | ( n756 & n787 ) ;
  assign n2044 = ( x44 & ~n1947 ) | ( x44 & n2043 ) | ( ~n1947 & n2043 ) ;
  assign n2045 = ( ~n1469 & n1796 ) | ( ~n1469 & n2044 ) | ( n1796 & n2044 ) ;
  assign n2047 = n2046 ^ n2045 ^ n1733 ;
  assign n2048 = n588 & ~n691 ;
  assign n2049 = ~n1264 & n2048 ;
  assign n2050 = ( n436 & n1966 ) | ( n436 & ~n1970 ) | ( n1966 & ~n1970 ) ;
  assign n2051 = n2050 ^ n1010 ^ n679 ;
  assign n2052 = ( ~n367 & n2049 ) | ( ~n367 & n2051 ) | ( n2049 & n2051 ) ;
  assign n2053 = n2052 ^ n1370 ^ x160 ;
  assign n2054 = n2053 ^ n1252 ^ x239 ;
  assign n2055 = ( n2042 & n2047 ) | ( n2042 & ~n2054 ) | ( n2047 & ~n2054 ) ;
  assign n2056 = n1764 ^ n1573 ^ n1321 ;
  assign n2057 = n1204 | n1379 ;
  assign n2058 = n2057 ^ n1268 ^ 1'b0 ;
  assign n2059 = ( n1596 & ~n1925 ) | ( n1596 & n2058 ) | ( ~n1925 & n2058 ) ;
  assign n2060 = n1060 ^ n350 ^ n301 ;
  assign n2061 = ( n2056 & ~n2059 ) | ( n2056 & n2060 ) | ( ~n2059 & n2060 ) ;
  assign n2062 = ( n625 & n966 ) | ( n625 & ~n1026 ) | ( n966 & ~n1026 ) ;
  assign n2063 = ( n272 & n1003 ) | ( n272 & ~n2046 ) | ( n1003 & ~n2046 ) ;
  assign n2064 = ( n508 & n2062 ) | ( n508 & ~n2063 ) | ( n2062 & ~n2063 ) ;
  assign n2071 = n1955 ^ n901 ^ n869 ;
  assign n2072 = ( ~n1535 & n1601 ) | ( ~n1535 & n2071 ) | ( n1601 & n2071 ) ;
  assign n2065 = ( n499 & n627 ) | ( n499 & n1590 ) | ( n627 & n1590 ) ;
  assign n2068 = ( x88 & n577 ) | ( x88 & n870 ) | ( n577 & n870 ) ;
  assign n2066 = n1422 ^ n688 ^ n686 ;
  assign n2067 = ( x161 & n1262 ) | ( x161 & ~n2066 ) | ( n1262 & ~n2066 ) ;
  assign n2069 = n2068 ^ n2067 ^ n1275 ;
  assign n2070 = ~n2065 & n2069 ;
  assign n2073 = n2072 ^ n2070 ^ n1147 ;
  assign n2074 = ( ~n513 & n827 ) | ( ~n513 & n2073 ) | ( n827 & n2073 ) ;
  assign n2075 = x226 & n1942 ;
  assign n2076 = ~n666 & n2075 ;
  assign n2077 = n1842 | n2076 ;
  assign n2078 = ( x133 & ~x139 ) | ( x133 & n1953 ) | ( ~x139 & n1953 ) ;
  assign n2079 = x95 & n308 ;
  assign n2080 = n2079 ^ x248 ^ 1'b0 ;
  assign n2081 = ( ~x77 & n326 ) | ( ~x77 & n1836 ) | ( n326 & n1836 ) ;
  assign n2082 = ( n1142 & n1676 ) | ( n1142 & ~n2081 ) | ( n1676 & ~n2081 ) ;
  assign n2083 = n1243 ^ n816 ^ 1'b0 ;
  assign n2084 = ~n2082 & n2083 ;
  assign n2085 = ( ~n750 & n1739 ) | ( ~n750 & n2084 ) | ( n1739 & n2084 ) ;
  assign n2086 = ( n2078 & n2080 ) | ( n2078 & ~n2085 ) | ( n2080 & ~n2085 ) ;
  assign n2087 = x16 & ~n2086 ;
  assign n2088 = x134 & ~n569 ;
  assign n2089 = ( n454 & ~n468 ) | ( n454 & n1431 ) | ( ~n468 & n1431 ) ;
  assign n2090 = x204 & ~n2089 ;
  assign n2091 = n2090 ^ n1504 ^ 1'b0 ;
  assign n2092 = n1712 ^ n275 ^ 1'b0 ;
  assign n2093 = ~n1637 & n2092 ;
  assign n2094 = ( n2088 & ~n2091 ) | ( n2088 & n2093 ) | ( ~n2091 & n2093 ) ;
  assign n2095 = x114 & n987 ;
  assign n2096 = n2094 & n2095 ;
  assign n2097 = n1503 ^ n1002 ^ n287 ;
  assign n2098 = n1075 ^ n601 ^ n557 ;
  assign n2099 = n2098 ^ n2097 ^ n325 ;
  assign n2100 = ( ~n1130 & n2097 ) | ( ~n1130 & n2099 ) | ( n2097 & n2099 ) ;
  assign n2101 = n2100 ^ n1594 ^ 1'b0 ;
  assign n2102 = n1921 ^ n1030 ^ n335 ;
  assign n2103 = ( n755 & n1912 ) | ( n755 & n2102 ) | ( n1912 & n2102 ) ;
  assign n2104 = ( n2096 & n2101 ) | ( n2096 & n2103 ) | ( n2101 & n2103 ) ;
  assign n2117 = n2091 ^ n1016 ^ n836 ;
  assign n2118 = ( ~n362 & n1238 ) | ( ~n362 & n2117 ) | ( n1238 & n2117 ) ;
  assign n2119 = n2118 ^ n305 ^ x82 ;
  assign n2120 = n1113 & n1371 ;
  assign n2121 = n2119 & n2120 ;
  assign n2122 = n2121 ^ n1222 ^ n866 ;
  assign n2108 = n827 ^ n662 ^ n386 ;
  assign n2109 = ~n806 & n1145 ;
  assign n2110 = n2109 ^ n849 ^ 1'b0 ;
  assign n2111 = ~n984 & n2110 ;
  assign n2112 = n2108 & n2111 ;
  assign n2113 = ( n893 & ~n1650 ) | ( n893 & n1827 ) | ( ~n1650 & n1827 ) ;
  assign n2114 = ( n311 & n2112 ) | ( n311 & ~n2113 ) | ( n2112 & ~n2113 ) ;
  assign n2105 = n463 ^ n343 ^ x186 ;
  assign n2106 = ( n846 & n1161 ) | ( n846 & ~n2105 ) | ( n1161 & ~n2105 ) ;
  assign n2107 = n2106 ^ n560 ^ n540 ;
  assign n2115 = n2114 ^ n2107 ^ n1637 ;
  assign n2116 = ( n597 & ~n1894 ) | ( n597 & n2115 ) | ( ~n1894 & n2115 ) ;
  assign n2123 = n2122 ^ n2116 ^ 1'b0 ;
  assign n2124 = n651 & ~n2123 ;
  assign n2127 = n1297 ^ n932 ^ n665 ;
  assign n2128 = ( n323 & n896 ) | ( n323 & n2127 ) | ( n896 & n2127 ) ;
  assign n2125 = n1371 ^ n514 ^ n406 ;
  assign n2126 = ( ~n635 & n1522 ) | ( ~n635 & n2125 ) | ( n1522 & n2125 ) ;
  assign n2129 = n2128 ^ n2126 ^ n2009 ;
  assign n2130 = ( n1019 & ~n1167 ) | ( n1019 & n1624 ) | ( ~n1167 & n1624 ) ;
  assign n2133 = ( ~x31 & x149 ) | ( ~x31 & x191 ) | ( x149 & x191 ) ;
  assign n2131 = ( x250 & n376 ) | ( x250 & n593 ) | ( n376 & n593 ) ;
  assign n2132 = ~n1191 & n2131 ;
  assign n2134 = n2133 ^ n2132 ^ 1'b0 ;
  assign n2138 = ( n463 & ~n556 ) | ( n463 & n1294 ) | ( ~n556 & n1294 ) ;
  assign n2135 = n424 | n489 ;
  assign n2136 = n694 & ~n2135 ;
  assign n2137 = n2136 ^ n1836 ^ n1201 ;
  assign n2139 = n2138 ^ n2137 ^ n876 ;
  assign n2147 = n587 ^ n483 ^ n319 ;
  assign n2145 = ( x250 & ~n287 ) | ( x250 & n950 ) | ( ~n287 & n950 ) ;
  assign n2146 = n2145 ^ n1222 ^ x240 ;
  assign n2142 = x219 & ~n1719 ;
  assign n2143 = n2142 ^ n1503 ^ 1'b0 ;
  assign n2140 = n1941 ^ n1595 ^ x60 ;
  assign n2141 = ( x105 & ~n1159 ) | ( x105 & n2140 ) | ( ~n1159 & n2140 ) ;
  assign n2144 = n2143 ^ n2141 ^ n534 ;
  assign n2148 = n2147 ^ n2146 ^ n2144 ;
  assign n2149 = x88 & x124 ;
  assign n2150 = ~x232 & n2149 ;
  assign n2151 = n2150 ^ n565 ^ n473 ;
  assign n2152 = n2136 ^ n1925 ^ 1'b0 ;
  assign n2153 = n1275 ^ n662 ^ n584 ;
  assign n2154 = ~n1946 & n2153 ;
  assign n2155 = ( n264 & n954 ) | ( n264 & ~n2154 ) | ( n954 & ~n2154 ) ;
  assign n2156 = n1752 ^ n304 ^ x100 ;
  assign n2157 = n2156 ^ n1219 ^ n1158 ;
  assign n2158 = ( ~n343 & n547 ) | ( ~n343 & n635 ) | ( n547 & n635 ) ;
  assign n2159 = ( n575 & n1566 ) | ( n575 & ~n2158 ) | ( n1566 & ~n2158 ) ;
  assign n2160 = ( n1330 & n1757 ) | ( n1330 & n2159 ) | ( n1757 & n2159 ) ;
  assign n2161 = n2160 ^ n1917 ^ 1'b0 ;
  assign n2162 = n1763 | n2161 ;
  assign n2163 = ( ~n1638 & n2157 ) | ( ~n1638 & n2162 ) | ( n2157 & n2162 ) ;
  assign n2164 = ( n2152 & n2155 ) | ( n2152 & n2163 ) | ( n2155 & n2163 ) ;
  assign n2165 = ( n2100 & n2151 ) | ( n2100 & ~n2164 ) | ( n2151 & ~n2164 ) ;
  assign n2166 = ( n605 & n2148 ) | ( n605 & ~n2165 ) | ( n2148 & ~n2165 ) ;
  assign n2167 = n448 ^ n271 ^ x157 ;
  assign n2175 = ( ~x253 & n273 ) | ( ~x253 & n819 ) | ( n273 & n819 ) ;
  assign n2169 = n2088 ^ n1342 ^ x74 ;
  assign n2170 = n520 ^ x73 ^ 1'b0 ;
  assign n2171 = n345 & n2170 ;
  assign n2172 = ( n545 & n2147 ) | ( n545 & n2171 ) | ( n2147 & n2171 ) ;
  assign n2173 = ( n1372 & n1866 ) | ( n1372 & n2172 ) | ( n1866 & n2172 ) ;
  assign n2174 = ( n2031 & n2169 ) | ( n2031 & n2173 ) | ( n2169 & n2173 ) ;
  assign n2168 = n1634 ^ n1263 ^ n1060 ;
  assign n2176 = n2175 ^ n2174 ^ n2168 ;
  assign n2177 = n1719 | n1830 ;
  assign n2178 = n2177 ^ n1310 ^ 1'b0 ;
  assign n2179 = ( n357 & ~n1129 ) | ( n357 & n1797 ) | ( ~n1129 & n1797 ) ;
  assign n2180 = n965 ^ n396 ^ n309 ;
  assign n2181 = n1319 ^ n628 ^ n484 ;
  assign n2182 = n2181 ^ n604 ^ 1'b0 ;
  assign n2183 = n1276 & n2182 ;
  assign n2184 = ( n681 & ~n1052 ) | ( n681 & n2183 ) | ( ~n1052 & n2183 ) ;
  assign n2185 = n2184 ^ n1363 ^ n1120 ;
  assign n2186 = ( n738 & n1545 ) | ( n738 & n2185 ) | ( n1545 & n2185 ) ;
  assign n2187 = n2180 & n2186 ;
  assign n2188 = n2187 ^ x160 ^ 1'b0 ;
  assign n2189 = n2188 ^ n1896 ^ n1361 ;
  assign n2190 = n2189 ^ n863 ^ x241 ;
  assign n2222 = ( x59 & x197 ) | ( x59 & n814 ) | ( x197 & n814 ) ;
  assign n2208 = n1294 ^ n614 ^ 1'b0 ;
  assign n2209 = n482 & n2208 ;
  assign n2206 = n419 ^ n289 ^ x126 ;
  assign n2207 = ( n420 & n1953 ) | ( n420 & ~n2206 ) | ( n1953 & ~n2206 ) ;
  assign n2210 = n2209 ^ n2207 ^ n1478 ;
  assign n2204 = n1988 ^ n1527 ^ x236 ;
  assign n2205 = n2204 ^ n1645 ^ n789 ;
  assign n2201 = n1661 ^ n1214 ^ n1053 ;
  assign n2202 = ( ~n740 & n930 ) | ( ~n740 & n2201 ) | ( n930 & n2201 ) ;
  assign n2199 = ( n1123 & n1887 ) | ( n1123 & n1983 ) | ( n1887 & n1983 ) ;
  assign n2198 = n1761 ^ n1220 ^ n868 ;
  assign n2197 = ( x40 & n693 ) | ( x40 & n1077 ) | ( n693 & n1077 ) ;
  assign n2200 = n2199 ^ n2198 ^ n2197 ;
  assign n2192 = n572 ^ n305 ^ x55 ;
  assign n2191 = x99 & n1213 ;
  assign n2193 = n2192 ^ n2191 ^ 1'b0 ;
  assign n2194 = n725 & ~n1648 ;
  assign n2195 = n2193 & n2194 ;
  assign n2196 = n2195 ^ n973 ^ n965 ;
  assign n2203 = n2202 ^ n2200 ^ n2196 ;
  assign n2211 = n2210 ^ n2205 ^ n2203 ;
  assign n2216 = ~x239 & n799 ;
  assign n2217 = n2216 ^ n1810 ^ n851 ;
  assign n2218 = ( ~n584 & n1726 ) | ( ~n584 & n2217 ) | ( n1726 & n2217 ) ;
  assign n2212 = ( n471 & n1532 ) | ( n471 & ~n2192 ) | ( n1532 & ~n2192 ) ;
  assign n2213 = n658 ^ n417 ^ 1'b0 ;
  assign n2214 = n2213 ^ n848 ^ n482 ;
  assign n2215 = n2212 & n2214 ;
  assign n2219 = n2218 ^ n2215 ^ 1'b0 ;
  assign n2220 = ( ~n1362 & n2211 ) | ( ~n1362 & n2219 ) | ( n2211 & n2219 ) ;
  assign n2221 = ~n1042 & n2220 ;
  assign n2223 = n2222 ^ n2221 ^ n949 ;
  assign n2241 = n696 | n1801 ;
  assign n2237 = n511 | n983 ;
  assign n2238 = n1194 ^ n502 ^ n359 ;
  assign n2239 = ( n310 & n2237 ) | ( n310 & ~n2238 ) | ( n2237 & ~n2238 ) ;
  assign n2234 = ( x81 & n371 ) | ( x81 & n1338 ) | ( n371 & n1338 ) ;
  assign n2235 = n2234 ^ n1426 ^ n1135 ;
  assign n2232 = x14 & x22 ;
  assign n2233 = n2232 ^ x210 ^ 1'b0 ;
  assign n2224 = ( n645 & n772 ) | ( n645 & n891 ) | ( n772 & n891 ) ;
  assign n2225 = n2002 ^ n1176 ^ x193 ;
  assign n2226 = n2225 ^ n1217 ^ n810 ;
  assign n2228 = x167 ^ x63 ^ 1'b0 ;
  assign n2227 = x209 & x223 ;
  assign n2229 = n2228 ^ n2227 ^ 1'b0 ;
  assign n2230 = ( ~n633 & n1633 ) | ( ~n633 & n2229 ) | ( n1633 & n2229 ) ;
  assign n2231 = ( n2224 & ~n2226 ) | ( n2224 & n2230 ) | ( ~n2226 & n2230 ) ;
  assign n2236 = n2235 ^ n2233 ^ n2231 ;
  assign n2240 = n2239 ^ n2236 ^ n1722 ;
  assign n2242 = n2241 ^ n2240 ^ n1311 ;
  assign n2243 = n2242 ^ n1121 ^ n821 ;
  assign n2244 = n2243 ^ n839 ^ x237 ;
  assign n2246 = ( n327 & n343 ) | ( n327 & ~n389 ) | ( n343 & ~n389 ) ;
  assign n2247 = n2246 ^ n1838 ^ x143 ;
  assign n2245 = ( n409 & n1309 ) | ( n409 & ~n1313 ) | ( n1309 & ~n1313 ) ;
  assign n2248 = n2247 ^ n2245 ^ n1822 ;
  assign n2249 = ( ~n587 & n2035 ) | ( ~n587 & n2248 ) | ( n2035 & n2248 ) ;
  assign n2250 = ( n685 & n951 ) | ( n685 & ~n1055 ) | ( n951 & ~n1055 ) ;
  assign n2257 = n1902 ^ n322 ^ x142 ;
  assign n2258 = ( x8 & n313 ) | ( x8 & n2257 ) | ( n313 & n2257 ) ;
  assign n2255 = n720 ^ x150 ^ x66 ;
  assign n2256 = n2255 ^ n827 ^ n572 ;
  assign n2259 = n2258 ^ n2256 ^ x77 ;
  assign n2260 = n2259 ^ n1255 ^ x106 ;
  assign n2252 = ( x9 & ~x82 ) | ( x9 & n537 ) | ( ~x82 & n537 ) ;
  assign n2251 = n1021 ^ n597 ^ n459 ;
  assign n2253 = n2252 ^ n2251 ^ 1'b0 ;
  assign n2254 = n2253 ^ n743 ^ n317 ;
  assign n2261 = n2260 ^ n2254 ^ n1133 ;
  assign n2262 = ( n2038 & ~n2250 ) | ( n2038 & n2261 ) | ( ~n2250 & n2261 ) ;
  assign n2263 = ( ~n294 & n295 ) | ( ~n294 & n442 ) | ( n295 & n442 ) ;
  assign n2264 = n2263 ^ x172 ^ 1'b0 ;
  assign n2265 = ( n835 & ~n1409 ) | ( n835 & n1504 ) | ( ~n1409 & n1504 ) ;
  assign n2266 = x250 ^ x25 ^ 1'b0 ;
  assign n2267 = x103 & n2266 ;
  assign n2268 = n2267 ^ n898 ^ n496 ;
  assign n2269 = ( n1262 & n2265 ) | ( n1262 & ~n2268 ) | ( n2265 & ~n2268 ) ;
  assign n2303 = ( n817 & n1283 ) | ( n817 & ~n1450 ) | ( n1283 & ~n1450 ) ;
  assign n2299 = ( x248 & n358 ) | ( x248 & ~n1071 ) | ( n358 & ~n1071 ) ;
  assign n2300 = ( x33 & ~n2158 ) | ( x33 & n2181 ) | ( ~n2158 & n2181 ) ;
  assign n2301 = n2300 ^ n698 ^ 1'b0 ;
  assign n2302 = n2299 & n2301 ;
  assign n2304 = n2303 ^ n2302 ^ x245 ;
  assign n2305 = ( n614 & n1382 ) | ( n614 & ~n1570 ) | ( n1382 & ~n1570 ) ;
  assign n2306 = ( x161 & n2304 ) | ( x161 & ~n2305 ) | ( n2304 & ~n2305 ) ;
  assign n2292 = n574 ^ x208 ^ x16 ;
  assign n2293 = n753 | n1874 ;
  assign n2294 = n380 | n2293 ;
  assign n2295 = n2294 ^ n1345 ^ 1'b0 ;
  assign n2296 = n2295 ^ n671 ^ n287 ;
  assign n2297 = n337 & n2296 ;
  assign n2298 = n2292 & n2297 ;
  assign n2270 = n1573 ^ n1566 ^ n597 ;
  assign n2271 = n1980 ^ n1219 ^ x231 ;
  assign n2272 = ( ~n668 & n2270 ) | ( ~n668 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2277 = ( ~n511 & n934 ) | ( ~n511 & n1966 ) | ( n934 & n1966 ) ;
  assign n2278 = ( n534 & n1767 ) | ( n534 & n2277 ) | ( n1767 & n2277 ) ;
  assign n2273 = n661 ^ n574 ^ x133 ;
  assign n2274 = ~n871 & n2273 ;
  assign n2275 = n2192 ^ n2039 ^ 1'b0 ;
  assign n2276 = n2274 & ~n2275 ;
  assign n2279 = n2278 ^ n2276 ^ 1'b0 ;
  assign n2287 = n1026 ^ n589 ^ x253 ;
  assign n2285 = n462 & ~n1515 ;
  assign n2286 = ~n2250 & n2285 ;
  assign n2284 = ( x180 & n452 ) | ( x180 & n878 ) | ( n452 & n878 ) ;
  assign n2288 = n2287 ^ n2286 ^ n2284 ;
  assign n2289 = ~n1824 & n2288 ;
  assign n2280 = n1925 ^ n1028 ^ n1014 ;
  assign n2281 = n1970 & ~n2280 ;
  assign n2282 = ~n2183 & n2281 ;
  assign n2283 = n1593 | n2282 ;
  assign n2290 = n2289 ^ n2283 ^ 1'b0 ;
  assign n2291 = ( n2272 & n2279 ) | ( n2272 & ~n2290 ) | ( n2279 & ~n2290 ) ;
  assign n2307 = n2306 ^ n2298 ^ n2291 ;
  assign n2309 = ( x191 & ~n275 ) | ( x191 & n839 ) | ( ~n275 & n839 ) ;
  assign n2310 = n2309 ^ n619 ^ n370 ;
  assign n2308 = ( n692 & n1137 ) | ( n692 & n2224 ) | ( n1137 & n2224 ) ;
  assign n2311 = n2310 ^ n2308 ^ n657 ;
  assign n2313 = n382 | n682 ;
  assign n2314 = n297 | n2313 ;
  assign n2312 = n1422 ^ n1097 ^ n800 ;
  assign n2315 = n2314 ^ n2312 ^ 1'b0 ;
  assign n2316 = n1135 & ~n2315 ;
  assign n2317 = n1838 ^ n1057 ^ x107 ;
  assign n2318 = n995 ^ n336 ^ 1'b0 ;
  assign n2319 = n1771 ^ n1770 ^ n1706 ;
  assign n2320 = ( ~n650 & n2318 ) | ( ~n650 & n2319 ) | ( n2318 & n2319 ) ;
  assign n2321 = ~n2317 & n2320 ;
  assign n2322 = n2321 ^ n2098 ^ 1'b0 ;
  assign n2323 = ( n2311 & n2316 ) | ( n2311 & n2322 ) | ( n2316 & n2322 ) ;
  assign n2324 = x133 & ~n2171 ;
  assign n2325 = ( n694 & n1235 ) | ( n694 & n2324 ) | ( n1235 & n2324 ) ;
  assign n2326 = ( x212 & n568 ) | ( x212 & ~n2267 ) | ( n568 & ~n2267 ) ;
  assign n2327 = ( ~n961 & n1797 ) | ( ~n961 & n2326 ) | ( n1797 & n2326 ) ;
  assign n2346 = x3 & x24 ;
  assign n2336 = n1288 ^ n688 ^ n601 ;
  assign n2337 = n2336 ^ n1814 ^ n1184 ;
  assign n2338 = x19 & n1055 ;
  assign n2340 = ( x133 & ~n800 ) | ( x133 & n2002 ) | ( ~n800 & n2002 ) ;
  assign n2339 = x70 & n1063 ;
  assign n2341 = n2340 ^ n2339 ^ 1'b0 ;
  assign n2342 = ( x133 & n2338 ) | ( x133 & ~n2341 ) | ( n2338 & ~n2341 ) ;
  assign n2343 = n2337 | n2342 ;
  assign n2344 = n434 | n2343 ;
  assign n2331 = n962 & ~n2268 ;
  assign n2332 = n2331 ^ n2036 ^ x196 ;
  assign n2333 = n710 ^ x227 ^ x53 ;
  assign n2334 = n2333 ^ n1730 ^ n537 ;
  assign n2335 = ( ~n2099 & n2332 ) | ( ~n2099 & n2334 ) | ( n2332 & n2334 ) ;
  assign n2329 = n1504 ^ n1242 ^ n556 ;
  assign n2328 = n1248 ^ n1230 ^ n461 ;
  assign n2330 = n2329 ^ n2328 ^ x45 ;
  assign n2345 = n2344 ^ n2335 ^ n2330 ;
  assign n2347 = n2346 ^ n2345 ^ n1426 ;
  assign n2348 = ( ~x92 & n2327 ) | ( ~x92 & n2347 ) | ( n2327 & n2347 ) ;
  assign n2349 = n1479 ^ n1318 ^ n1194 ;
  assign n2350 = n2150 ^ n736 ^ x148 ;
  assign n2351 = n2350 ^ n1761 ^ n947 ;
  assign n2352 = n2351 ^ n2311 ^ 1'b0 ;
  assign n2353 = n1749 & n2352 ;
  assign n2354 = n1385 & n2353 ;
  assign n2355 = n2349 & n2354 ;
  assign n2357 = n1034 ^ x59 ^ 1'b0 ;
  assign n2358 = n1081 & ~n2357 ;
  assign n2356 = ( x249 & n852 ) | ( x249 & n1956 ) | ( n852 & n1956 ) ;
  assign n2359 = n2358 ^ n2356 ^ x28 ;
  assign n2361 = n423 ^ x95 ^ 1'b0 ;
  assign n2362 = x123 & ~n2361 ;
  assign n2360 = ( ~n325 & n1442 ) | ( ~n325 & n1865 ) | ( n1442 & n1865 ) ;
  assign n2363 = n2362 ^ n2360 ^ n2317 ;
  assign n2364 = n2252 ^ n1060 ^ n977 ;
  assign n2365 = ( x239 & ~n351 ) | ( x239 & n389 ) | ( ~n351 & n389 ) ;
  assign n2366 = n2365 ^ n2108 ^ x163 ;
  assign n2367 = n2366 ^ n438 ^ 1'b0 ;
  assign n2368 = n1295 ^ n818 ^ 1'b0 ;
  assign n2369 = n2368 ^ n1802 ^ x28 ;
  assign n2370 = ( n2364 & ~n2367 ) | ( n2364 & n2369 ) | ( ~n2367 & n2369 ) ;
  assign n2371 = n1330 ^ n1029 ^ n949 ;
  assign n2372 = ( ~n1484 & n2366 ) | ( ~n1484 & n2371 ) | ( n2366 & n2371 ) ;
  assign n2373 = ( x54 & n273 ) | ( x54 & n1582 ) | ( n273 & n1582 ) ;
  assign n2374 = n696 ^ n548 ^ x42 ;
  assign n2382 = n753 ^ n566 ^ x2 ;
  assign n2383 = ( n516 & n2299 ) | ( n516 & n2382 ) | ( n2299 & n2382 ) ;
  assign n2381 = ( ~n335 & n571 ) | ( ~n335 & n1751 ) | ( n571 & n1751 ) ;
  assign n2379 = ( n922 & n1738 ) | ( n922 & n1845 ) | ( n1738 & n1845 ) ;
  assign n2375 = ( x41 & n620 ) | ( x41 & n1282 ) | ( n620 & n1282 ) ;
  assign n2376 = n2375 ^ n815 ^ n360 ;
  assign n2377 = n2376 ^ n640 ^ 1'b0 ;
  assign n2378 = n1717 & ~n2377 ;
  assign n2380 = n2379 ^ n2378 ^ n1057 ;
  assign n2384 = n2383 ^ n2381 ^ n2380 ;
  assign n2385 = ( n312 & n2374 ) | ( n312 & ~n2384 ) | ( n2374 & ~n2384 ) ;
  assign n2386 = ( n1142 & ~n2373 ) | ( n1142 & n2385 ) | ( ~n2373 & n2385 ) ;
  assign n2387 = ( n2370 & n2372 ) | ( n2370 & n2386 ) | ( n2372 & n2386 ) ;
  assign n2388 = ( n2359 & n2363 ) | ( n2359 & n2387 ) | ( n2363 & n2387 ) ;
  assign n2389 = n1891 ^ n365 ^ 1'b0 ;
  assign n2390 = n617 ^ n257 ^ x2 ;
  assign n2391 = n431 ^ n400 ^ 1'b0 ;
  assign n2392 = ( n2389 & n2390 ) | ( n2389 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = ( n371 & n559 ) | ( n371 & n1006 ) | ( n559 & n1006 ) ;
  assign n2394 = ( n515 & n873 ) | ( n515 & n2393 ) | ( n873 & n2393 ) ;
  assign n2395 = ( n1105 & ~n1171 ) | ( n1105 & n2394 ) | ( ~n1171 & n2394 ) ;
  assign n2396 = ( n662 & n1522 ) | ( n662 & ~n2395 ) | ( n1522 & ~n2395 ) ;
  assign n2397 = n2396 ^ n1595 ^ 1'b0 ;
  assign n2398 = ( n464 & n943 ) | ( n464 & ~n2228 ) | ( n943 & ~n2228 ) ;
  assign n2399 = n2398 ^ n2225 ^ n1170 ;
  assign n2400 = ( ~x241 & n1372 ) | ( ~x241 & n1806 ) | ( n1372 & n1806 ) ;
  assign n2401 = n2036 ^ n1415 ^ 1'b0 ;
  assign n2402 = n2401 ^ n1927 ^ n507 ;
  assign n2403 = ( n418 & n512 ) | ( n418 & n580 ) | ( n512 & n580 ) ;
  assign n2404 = n1647 ^ x60 ^ 1'b0 ;
  assign n2405 = x203 & n2404 ;
  assign n2406 = ( x119 & ~n2403 ) | ( x119 & n2405 ) | ( ~n2403 & n2405 ) ;
  assign n2407 = ( ~n2400 & n2402 ) | ( ~n2400 & n2406 ) | ( n2402 & n2406 ) ;
  assign n2408 = ( n2397 & n2399 ) | ( n2397 & ~n2407 ) | ( n2399 & ~n2407 ) ;
  assign n2411 = n1188 ^ n738 ^ n258 ;
  assign n2409 = x37 & n1833 ;
  assign n2410 = n2409 ^ n1346 ^ 1'b0 ;
  assign n2412 = n2411 ^ n2410 ^ n781 ;
  assign n2413 = n1239 ^ n1000 ^ 1'b0 ;
  assign n2414 = n2413 ^ n456 ^ 1'b0 ;
  assign n2415 = n2256 | n2414 ;
  assign n2416 = ( n323 & n846 ) | ( n323 & n1077 ) | ( n846 & n1077 ) ;
  assign n2417 = ( n783 & n1211 ) | ( n783 & n2416 ) | ( n1211 & n2416 ) ;
  assign n2418 = ( ~n513 & n1546 ) | ( ~n513 & n2417 ) | ( n1546 & n2417 ) ;
  assign n2420 = ( ~n525 & n783 ) | ( ~n525 & n1047 ) | ( n783 & n1047 ) ;
  assign n2419 = n1532 & n2295 ;
  assign n2421 = n2420 ^ n2419 ^ 1'b0 ;
  assign n2422 = ( n1142 & n1555 ) | ( n1142 & n2421 ) | ( n1555 & n2421 ) ;
  assign n2423 = n2422 ^ n904 ^ x94 ;
  assign n2424 = n2311 ^ n1301 ^ n1013 ;
  assign n2425 = n1029 & n2424 ;
  assign n2426 = ( n2418 & ~n2423 ) | ( n2418 & n2425 ) | ( ~n2423 & n2425 ) ;
  assign n2432 = ( ~n1370 & n1481 ) | ( ~n1370 & n1845 ) | ( n1481 & n1845 ) ;
  assign n2433 = n2432 ^ n1436 ^ 1'b0 ;
  assign n2430 = ( ~x48 & x83 ) | ( ~x48 & n470 ) | ( x83 & n470 ) ;
  assign n2428 = n541 ^ x114 ^ x95 ;
  assign n2429 = n2428 ^ n1226 ^ n524 ;
  assign n2427 = n1741 ^ n1127 ^ n1005 ;
  assign n2431 = n2430 ^ n2429 ^ n2427 ;
  assign n2434 = n2433 ^ n2431 ^ n1221 ;
  assign n2438 = ( n323 & n1039 ) | ( n323 & n1539 ) | ( n1039 & n1539 ) ;
  assign n2439 = n2438 ^ n2091 ^ n1794 ;
  assign n2436 = ( n466 & ~n604 ) | ( n466 & n2226 ) | ( ~n604 & n2226 ) ;
  assign n2435 = ( n644 & n2027 ) | ( n644 & n2395 ) | ( n2027 & n2395 ) ;
  assign n2437 = n2436 ^ n2435 ^ n1149 ;
  assign n2440 = n2439 ^ n2437 ^ n386 ;
  assign n2441 = n2028 ^ n454 ^ x184 ;
  assign n2442 = ~n277 & n2441 ;
  assign n2443 = ~n1605 & n2442 ;
  assign n2444 = n1730 ^ n835 ^ n277 ;
  assign n2445 = n1562 ^ n1416 ^ n1193 ;
  assign n2446 = n2444 & n2445 ;
  assign n2447 = n2446 ^ n912 ^ 1'b0 ;
  assign n2448 = ( n538 & n627 ) | ( n538 & n2447 ) | ( n627 & n2447 ) ;
  assign n2449 = n2152 ^ n1310 ^ n765 ;
  assign n2450 = n2449 ^ n2150 ^ n1244 ;
  assign n2452 = n1474 ^ n1452 ^ n411 ;
  assign n2451 = ( n274 & ~n1482 ) | ( n274 & n1838 ) | ( ~n1482 & n1838 ) ;
  assign n2453 = n2452 ^ n2451 ^ n624 ;
  assign n2454 = ~n2450 & n2453 ;
  assign n2455 = n657 ^ x251 ^ 1'b0 ;
  assign n2457 = ~n912 & n996 ;
  assign n2458 = ( n1414 & n2304 ) | ( n1414 & n2457 ) | ( n2304 & n2457 ) ;
  assign n2456 = n1197 ^ n1080 ^ n565 ;
  assign n2459 = n2458 ^ n2456 ^ x210 ;
  assign n2460 = n2459 ^ n368 ^ 1'b0 ;
  assign n2461 = n2455 & ~n2460 ;
  assign n2462 = ( n932 & ~n1018 ) | ( n932 & n1777 ) | ( ~n1018 & n1777 ) ;
  assign n2463 = n2462 ^ n1731 ^ n652 ;
  assign n2464 = ( n1497 & ~n1603 ) | ( n1497 & n2463 ) | ( ~n1603 & n2463 ) ;
  assign n2465 = n1226 & n2464 ;
  assign n2466 = ~n1396 & n2465 ;
  assign n2467 = ( x134 & n1363 ) | ( x134 & n2255 ) | ( n1363 & n2255 ) ;
  assign n2468 = n1419 ^ n575 ^ x42 ;
  assign n2469 = ( x14 & n852 ) | ( x14 & ~n2468 ) | ( n852 & ~n2468 ) ;
  assign n2470 = n688 ^ x252 ^ 1'b0 ;
  assign n2471 = n2470 ^ n709 ^ n423 ;
  assign n2472 = ~n1055 & n2471 ;
  assign n2473 = n2472 ^ n1744 ^ 1'b0 ;
  assign n2474 = ( ~n831 & n996 ) | ( ~n831 & n2473 ) | ( n996 & n2473 ) ;
  assign n2475 = ( n675 & ~n2469 ) | ( n675 & n2474 ) | ( ~n2469 & n2474 ) ;
  assign n2477 = ( x143 & n792 ) | ( x143 & ~n925 ) | ( n792 & ~n925 ) ;
  assign n2478 = n2477 ^ n540 ^ n520 ;
  assign n2476 = x54 & n1330 ;
  assign n2479 = n2478 ^ n2476 ^ n1069 ;
  assign n2480 = n2198 ^ n1922 ^ 1'b0 ;
  assign n2481 = n1618 ^ n1227 ^ 1'b0 ;
  assign n2482 = ~n2160 & n2481 ;
  assign n2483 = ~n2169 & n2482 ;
  assign n2484 = ( x63 & n2162 ) | ( x63 & ~n2483 ) | ( n2162 & ~n2483 ) ;
  assign n2485 = ( n1515 & ~n2480 ) | ( n1515 & n2484 ) | ( ~n2480 & n2484 ) ;
  assign n2492 = n1740 ^ n1442 ^ n1300 ;
  assign n2493 = ( n333 & ~n396 ) | ( n333 & n2303 ) | ( ~n396 & n2303 ) ;
  assign n2494 = ( n588 & n2492 ) | ( n588 & n2493 ) | ( n2492 & n2493 ) ;
  assign n2488 = ( ~x110 & n467 ) | ( ~x110 & n483 ) | ( n467 & n483 ) ;
  assign n2489 = n2488 ^ n2468 ^ n2020 ;
  assign n2486 = ( n287 & n816 ) | ( n287 & n1730 ) | ( n816 & n1730 ) ;
  assign n2487 = ( n689 & n1488 ) | ( n689 & ~n2486 ) | ( n1488 & ~n2486 ) ;
  assign n2490 = n2489 ^ n2487 ^ 1'b0 ;
  assign n2491 = ~n1289 & n2490 ;
  assign n2495 = n2494 ^ n2491 ^ n1119 ;
  assign n2496 = n2485 & ~n2495 ;
  assign n2497 = n2479 & n2496 ;
  assign n2498 = ( n1417 & n1899 ) | ( n1417 & ~n2497 ) | ( n1899 & ~n2497 ) ;
  assign n2499 = ( x171 & ~n588 ) | ( x171 & n653 ) | ( ~n588 & n653 ) ;
  assign n2500 = n2499 ^ n2026 ^ n1823 ;
  assign n2501 = n2305 ^ n1539 ^ 1'b0 ;
  assign n2502 = ~n567 & n2501 ;
  assign n2506 = ( ~x180 & x220 ) | ( ~x180 & n1089 ) | ( x220 & n1089 ) ;
  assign n2503 = n1434 ^ n943 ^ 1'b0 ;
  assign n2504 = n2006 & ~n2503 ;
  assign n2505 = ~n1021 & n2504 ;
  assign n2507 = n2506 ^ n2505 ^ x202 ;
  assign n2508 = ( x140 & n955 ) | ( x140 & n1162 ) | ( n955 & n1162 ) ;
  assign n2509 = ( n1071 & n1339 ) | ( n1071 & n2508 ) | ( n1339 & n2508 ) ;
  assign n2510 = x205 & n396 ;
  assign n2511 = ( x172 & n968 ) | ( x172 & n1013 ) | ( n968 & n1013 ) ;
  assign n2512 = ( n361 & ~n2510 ) | ( n361 & n2511 ) | ( ~n2510 & n2511 ) ;
  assign n2513 = n2509 & ~n2512 ;
  assign n2514 = n2241 ^ n1605 ^ n1503 ;
  assign n2515 = ( n876 & n1337 ) | ( n876 & n2514 ) | ( n1337 & n2514 ) ;
  assign n2516 = n2515 ^ n1336 ^ n404 ;
  assign n2517 = n1307 ^ n1264 ^ 1'b0 ;
  assign n2518 = n2517 ^ n1937 ^ 1'b0 ;
  assign n2519 = ( n1408 & ~n1503 ) | ( n1408 & n1809 ) | ( ~n1503 & n1809 ) ;
  assign n2520 = ~n437 & n2258 ;
  assign n2521 = ~n2519 & n2520 ;
  assign n2522 = n491 & ~n2521 ;
  assign n2523 = n2522 ^ n959 ^ 1'b0 ;
  assign n2524 = n2523 ^ n484 ^ 1'b0 ;
  assign n2535 = ( n530 & n896 ) | ( n530 & n1478 ) | ( n896 & n1478 ) ;
  assign n2536 = n1720 ^ n1323 ^ n523 ;
  assign n2537 = ( x216 & n1628 ) | ( x216 & ~n2536 ) | ( n1628 & ~n2536 ) ;
  assign n2538 = ~x132 & x197 ;
  assign n2539 = ( ~n2535 & n2537 ) | ( ~n2535 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2525 = n1270 & ~n1960 ;
  assign n2526 = n1000 & n2525 ;
  assign n2527 = ( x129 & x214 ) | ( x129 & n2526 ) | ( x214 & n2526 ) ;
  assign n2528 = n2527 ^ n2097 ^ n1069 ;
  assign n2529 = ( x138 & x195 ) | ( x138 & ~n430 ) | ( x195 & ~n430 ) ;
  assign n2530 = ( ~x138 & n706 ) | ( ~x138 & n2529 ) | ( n706 & n2529 ) ;
  assign n2531 = n314 | n2530 ;
  assign n2532 = n2531 ^ n947 ^ 1'b0 ;
  assign n2533 = ( n375 & ~n2528 ) | ( n375 & n2532 ) | ( ~n2528 & n2532 ) ;
  assign n2534 = n2533 ^ n1983 ^ n1774 ;
  assign n2540 = n2539 ^ n2534 ^ n1566 ;
  assign n2542 = ( n536 & ~n829 ) | ( n536 & n1350 ) | ( ~n829 & n1350 ) ;
  assign n2543 = n1323 ^ n1137 ^ n819 ;
  assign n2544 = ( n690 & n726 ) | ( n690 & ~n1678 ) | ( n726 & ~n1678 ) ;
  assign n2545 = ( ~x237 & n2046 ) | ( ~x237 & n2544 ) | ( n2046 & n2544 ) ;
  assign n2546 = ( ~n2542 & n2543 ) | ( ~n2542 & n2545 ) | ( n2543 & n2545 ) ;
  assign n2547 = n666 & ~n781 ;
  assign n2548 = n2547 ^ n675 ^ 1'b0 ;
  assign n2549 = ( n2199 & n2546 ) | ( n2199 & ~n2548 ) | ( n2546 & ~n2548 ) ;
  assign n2541 = ( n296 & n431 ) | ( n296 & ~n1874 ) | ( n431 & ~n1874 ) ;
  assign n2550 = n2549 ^ n2541 ^ 1'b0 ;
  assign n2562 = x244 & n626 ;
  assign n2551 = n1928 ^ n1628 ^ n839 ;
  assign n2552 = n603 ^ n388 ^ n386 ;
  assign n2553 = ( x163 & n535 ) | ( x163 & n1036 ) | ( n535 & n1036 ) ;
  assign n2554 = n485 | n1034 ;
  assign n2555 = n2554 ^ x1 ^ 1'b0 ;
  assign n2556 = ( n2141 & n2553 ) | ( n2141 & ~n2555 ) | ( n2553 & ~n2555 ) ;
  assign n2557 = ( n1700 & n2552 ) | ( n1700 & ~n2556 ) | ( n2552 & ~n2556 ) ;
  assign n2558 = x184 & ~n2557 ;
  assign n2559 = ~n2551 & n2558 ;
  assign n2560 = x76 & ~n2559 ;
  assign n2561 = n1470 & n2560 ;
  assign n2563 = n2562 ^ n2561 ^ x31 ;
  assign n2564 = n1101 ^ n750 ^ n596 ;
  assign n2565 = n2564 ^ n949 ^ n610 ;
  assign n2566 = n2565 ^ n800 ^ x96 ;
  assign n2576 = n2370 ^ n2073 ^ n619 ;
  assign n2567 = ( x133 & n314 ) | ( x133 & ~n582 ) | ( n314 & ~n582 ) ;
  assign n2568 = ( ~n355 & n1471 ) | ( ~n355 & n2567 ) | ( n1471 & n2567 ) ;
  assign n2569 = n2568 ^ n837 ^ n815 ;
  assign n2570 = ( x169 & n1111 ) | ( x169 & ~n2569 ) | ( n1111 & ~n2569 ) ;
  assign n2571 = n1823 ^ n660 ^ 1'b0 ;
  assign n2572 = ( n843 & n946 ) | ( n843 & n2571 ) | ( n946 & n2571 ) ;
  assign n2573 = ( n1141 & n1827 ) | ( n1141 & ~n2050 ) | ( n1827 & ~n2050 ) ;
  assign n2574 = n2572 & n2573 ;
  assign n2575 = n2570 & n2574 ;
  assign n2577 = n2576 ^ n2575 ^ n1807 ;
  assign n2578 = n1385 ^ n773 ^ x252 ;
  assign n2579 = ( n615 & n673 ) | ( n615 & ~n2578 ) | ( n673 & ~n2578 ) ;
  assign n2580 = ( ~n415 & n683 ) | ( ~n415 & n1289 ) | ( n683 & n1289 ) ;
  assign n2581 = n993 ^ n693 ^ 1'b0 ;
  assign n2582 = n2580 | n2581 ;
  assign n2583 = ( ~n984 & n2579 ) | ( ~n984 & n2582 ) | ( n2579 & n2582 ) ;
  assign n2584 = ( n1991 & n2510 ) | ( n1991 & n2583 ) | ( n2510 & n2583 ) ;
  assign n2586 = n718 ^ n617 ^ n497 ;
  assign n2587 = ( ~n1498 & n1901 ) | ( ~n1498 & n2586 ) | ( n1901 & n2586 ) ;
  assign n2585 = n2133 ^ n1239 ^ n1077 ;
  assign n2588 = n2587 ^ n2585 ^ x220 ;
  assign n2589 = ( n1542 & n1881 ) | ( n1542 & ~n2319 ) | ( n1881 & ~n2319 ) ;
  assign n2590 = ( n618 & n1684 ) | ( n618 & n2589 ) | ( n1684 & n2589 ) ;
  assign n2591 = n2590 ^ n1099 ^ x246 ;
  assign n2592 = x9 & n2591 ;
  assign n2593 = n2592 ^ n766 ^ 1'b0 ;
  assign n2594 = ( n590 & n1792 ) | ( n590 & ~n2478 ) | ( n1792 & ~n2478 ) ;
  assign n2595 = n2594 ^ n724 ^ 1'b0 ;
  assign n2596 = ( x199 & ~n1970 ) | ( x199 & n2340 ) | ( ~n1970 & n2340 ) ;
  assign n2597 = n1647 ^ n1414 ^ 1'b0 ;
  assign n2598 = n1184 ^ n479 ^ x72 ;
  assign n2599 = ( n870 & ~n1774 ) | ( n870 & n2598 ) | ( ~n1774 & n2598 ) ;
  assign n2600 = ( n2596 & ~n2597 ) | ( n2596 & n2599 ) | ( ~n2597 & n2599 ) ;
  assign n2601 = n1118 ^ n831 ^ x32 ;
  assign n2602 = n1266 ^ n653 ^ x156 ;
  assign n2603 = n1224 ^ n1127 ^ x166 ;
  assign n2604 = n2602 | n2603 ;
  assign n2605 = n2601 & ~n2604 ;
  assign n2606 = ( x244 & n2600 ) | ( x244 & ~n2605 ) | ( n2600 & ~n2605 ) ;
  assign n2607 = ( ~n2289 & n2595 ) | ( ~n2289 & n2606 ) | ( n2595 & n2606 ) ;
  assign n2608 = n973 ^ x8 ^ 1'b0 ;
  assign n2609 = ( x251 & ~n2494 ) | ( x251 & n2608 ) | ( ~n2494 & n2608 ) ;
  assign n2610 = n1992 ^ n818 ^ 1'b0 ;
  assign n2611 = n1033 | n2610 ;
  assign n2612 = n2611 ^ n1475 ^ n1201 ;
  assign n2613 = n2612 ^ n2376 ^ x157 ;
  assign n2614 = n2242 & n2471 ;
  assign n2615 = n2614 ^ n351 ^ x6 ;
  assign n2616 = ( ~n1141 & n2613 ) | ( ~n1141 & n2615 ) | ( n2613 & n2615 ) ;
  assign n2627 = ( x78 & n264 ) | ( x78 & n521 ) | ( n264 & n521 ) ;
  assign n2628 = n2627 ^ n1288 ^ x3 ;
  assign n2629 = x170 & n640 ;
  assign n2630 = ( ~n800 & n2628 ) | ( ~n800 & n2629 ) | ( n2628 & n2629 ) ;
  assign n2624 = n580 & ~n2336 ;
  assign n2625 = ( ~x242 & n668 ) | ( ~x242 & n2624 ) | ( n668 & n2624 ) ;
  assign n2620 = ( ~n605 & n1419 ) | ( ~n605 & n1522 ) | ( n1419 & n1522 ) ;
  assign n2621 = ( n511 & n1042 ) | ( n511 & ~n2620 ) | ( n1042 & ~n2620 ) ;
  assign n2617 = n2579 ^ n1122 ^ n297 ;
  assign n2618 = ( x178 & ~n1704 ) | ( x178 & n2031 ) | ( ~n1704 & n2031 ) ;
  assign n2619 = ( n448 & ~n2617 ) | ( n448 & n2618 ) | ( ~n2617 & n2618 ) ;
  assign n2622 = n2621 ^ n2619 ^ x47 ;
  assign n2623 = ( n851 & n1578 ) | ( n851 & n2622 ) | ( n1578 & n2622 ) ;
  assign n2626 = n2625 ^ n2623 ^ n1502 ;
  assign n2631 = n2630 ^ n2626 ^ n429 ;
  assign n2635 = n2091 ^ n1469 ^ n751 ;
  assign n2632 = n1730 ^ n1351 ^ 1'b0 ;
  assign n2633 = ~n875 & n2632 ;
  assign n2634 = ( ~n799 & n2094 ) | ( ~n799 & n2633 ) | ( n2094 & n2633 ) ;
  assign n2636 = n2635 ^ n2634 ^ n1280 ;
  assign n2637 = n2159 ^ n1249 ^ n567 ;
  assign n2638 = n1897 ^ n973 ^ x140 ;
  assign n2639 = n2638 ^ n1739 ^ x223 ;
  assign n2640 = ( x0 & n2151 ) | ( x0 & n2639 ) | ( n2151 & n2639 ) ;
  assign n2641 = ( n1148 & ~n2637 ) | ( n1148 & n2640 ) | ( ~n2637 & n2640 ) ;
  assign n2642 = ~n449 & n1504 ;
  assign n2643 = ( x192 & n584 ) | ( x192 & ~n1423 ) | ( n584 & ~n1423 ) ;
  assign n2644 = ( ~x151 & n1152 ) | ( ~x151 & n2643 ) | ( n1152 & n2643 ) ;
  assign n2645 = ( ~n434 & n2642 ) | ( ~n434 & n2644 ) | ( n2642 & n2644 ) ;
  assign n2650 = ~n298 & n1351 ;
  assign n2651 = n2650 ^ n1231 ^ 1'b0 ;
  assign n2652 = n2651 ^ n1695 ^ x251 ;
  assign n2646 = x239 | n2088 ;
  assign n2647 = n2314 ^ n1368 ^ n809 ;
  assign n2648 = n2647 ^ n680 ^ 1'b0 ;
  assign n2649 = n2646 & ~n2648 ;
  assign n2653 = n2652 ^ n2649 ^ n260 ;
  assign n2654 = n1593 ^ n1067 ^ n274 ;
  assign n2655 = ( n1368 & ~n1620 ) | ( n1368 & n2654 ) | ( ~n1620 & n2654 ) ;
  assign n2656 = n2263 ^ n310 ^ x171 ;
  assign n2657 = n2656 ^ n2020 ^ x244 ;
  assign n2658 = ( n1268 & n1536 ) | ( n1268 & n2657 ) | ( n1536 & n2657 ) ;
  assign n2659 = ( n1547 & ~n2216 ) | ( n1547 & n2658 ) | ( ~n2216 & n2658 ) ;
  assign n2660 = n2655 | n2659 ;
  assign n2661 = n1754 & ~n2660 ;
  assign n2662 = ( x249 & n770 ) | ( x249 & ~n1960 ) | ( n770 & ~n1960 ) ;
  assign n2663 = n2615 & n2662 ;
  assign n2664 = n2661 & n2663 ;
  assign n2667 = ( n786 & n1915 ) | ( n786 & ~n2304 ) | ( n1915 & ~n2304 ) ;
  assign n2668 = n598 ^ x245 ^ x198 ;
  assign n2669 = ( n299 & n2667 ) | ( n299 & ~n2668 ) | ( n2667 & ~n2668 ) ;
  assign n2670 = ( ~n1612 & n2067 ) | ( ~n1612 & n2669 ) | ( n2067 & n2669 ) ;
  assign n2665 = x144 & n1225 ;
  assign n2666 = ~n2452 & n2665 ;
  assign n2671 = n2670 ^ n2666 ^ x242 ;
  assign n2672 = n2511 ^ n1219 ^ n310 ;
  assign n2673 = n2672 ^ n1526 ^ n1186 ;
  assign n2674 = n2673 ^ n821 ^ x28 ;
  assign n2675 = ( n283 & n1809 ) | ( n283 & n2674 ) | ( n1809 & n2674 ) ;
  assign n2680 = n567 & ~n605 ;
  assign n2681 = ( n1717 & n1775 ) | ( n1717 & n2680 ) | ( n1775 & n2680 ) ;
  assign n2676 = x156 & n1564 ;
  assign n2677 = n649 & n2676 ;
  assign n2678 = n2677 ^ n2572 ^ x90 ;
  assign n2679 = n2678 ^ n1490 ^ n483 ;
  assign n2682 = n2681 ^ n2679 ^ n1000 ;
  assign n2683 = ( n1044 & ~n2675 ) | ( n1044 & n2682 ) | ( ~n2675 & n2682 ) ;
  assign n2684 = ~n1416 & n2683 ;
  assign n2685 = n646 ^ x109 ^ 1'b0 ;
  assign n2687 = n1935 ^ n919 ^ n760 ;
  assign n2686 = n2252 ^ n651 ^ x171 ;
  assign n2688 = n2687 ^ n2686 ^ n1069 ;
  assign n2695 = n1395 ^ x234 ^ x158 ;
  assign n2696 = ( ~n561 & n2530 ) | ( ~n561 & n2695 ) | ( n2530 & n2695 ) ;
  assign n2689 = ( x166 & n904 ) | ( x166 & ~n1106 ) | ( n904 & ~n1106 ) ;
  assign n2690 = n2689 ^ n1758 ^ n1091 ;
  assign n2692 = ~n258 & n992 ;
  assign n2691 = ( n666 & n826 ) | ( n666 & n1064 ) | ( n826 & n1064 ) ;
  assign n2693 = n2692 ^ n2691 ^ n1550 ;
  assign n2694 = ( n2015 & n2690 ) | ( n2015 & n2693 ) | ( n2690 & n2693 ) ;
  assign n2697 = n2696 ^ n2694 ^ n755 ;
  assign n2698 = n1481 ^ n1246 ^ n377 ;
  assign n2699 = ( x233 & ~n1209 ) | ( x233 & n2698 ) | ( ~n1209 & n2698 ) ;
  assign n2700 = ( ~n1031 & n2066 ) | ( ~n1031 & n2293 ) | ( n2066 & n2293 ) ;
  assign n2701 = n2700 ^ n1109 ^ x209 ;
  assign n2702 = n857 ^ n826 ^ n298 ;
  assign n2703 = n2318 ^ n1365 ^ n1019 ;
  assign n2704 = ( n596 & n2702 ) | ( n596 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2705 = ( ~n2699 & n2701 ) | ( ~n2699 & n2704 ) | ( n2701 & n2704 ) ;
  assign n2706 = ( n382 & n2337 ) | ( n382 & n2705 ) | ( n2337 & n2705 ) ;
  assign n2707 = n1222 | n1415 ;
  assign n2708 = n2706 & ~n2707 ;
  assign n2709 = ( ~n1115 & n2067 ) | ( ~n1115 & n2085 ) | ( n2067 & n2085 ) ;
  assign n2710 = n2709 ^ n884 ^ 1'b0 ;
  assign n2711 = n1637 ^ n1373 ^ n620 ;
  assign n2712 = ( ~x176 & n2710 ) | ( ~x176 & n2711 ) | ( n2710 & n2711 ) ;
  assign n2727 = n2701 ^ n1204 ^ n688 ;
  assign n2720 = n1738 ^ n1100 ^ n493 ;
  assign n2723 = ( x103 & n501 ) | ( x103 & n804 ) | ( n501 & n804 ) ;
  assign n2721 = ( ~x98 & x160 ) | ( ~x98 & n1503 ) | ( x160 & n1503 ) ;
  assign n2722 = ( x40 & ~n374 ) | ( x40 & n2721 ) | ( ~n374 & n2721 ) ;
  assign n2724 = n2723 ^ n2722 ^ x79 ;
  assign n2725 = ( ~x14 & n2720 ) | ( ~x14 & n2724 ) | ( n2720 & n2724 ) ;
  assign n2726 = ~n758 & n2725 ;
  assign n2728 = n2727 ^ n2726 ^ 1'b0 ;
  assign n2718 = n631 ^ x244 ^ x199 ;
  assign n2719 = ( n1225 & n2421 ) | ( n1225 & n2718 ) | ( n2421 & n2718 ) ;
  assign n2713 = ( n1411 & n2438 ) | ( n1411 & ~n2703 ) | ( n2438 & ~n2703 ) ;
  assign n2714 = ( ~n523 & n2591 ) | ( ~n523 & n2713 ) | ( n2591 & n2713 ) ;
  assign n2715 = n2714 ^ n1377 ^ 1'b0 ;
  assign n2716 = ( x66 & n343 ) | ( x66 & ~n1859 ) | ( n343 & ~n1859 ) ;
  assign n2717 = ( n2308 & n2715 ) | ( n2308 & ~n2716 ) | ( n2715 & ~n2716 ) ;
  assign n2729 = n2728 ^ n2719 ^ n2717 ;
  assign n2751 = n584 ^ n538 ^ x166 ;
  assign n2752 = ( ~n2416 & n2640 ) | ( ~n2416 & n2751 ) | ( n2640 & n2751 ) ;
  assign n2742 = n675 ^ x7 ^ 1'b0 ;
  assign n2743 = ( ~n1082 & n2338 ) | ( ~n1082 & n2742 ) | ( n2338 & n2742 ) ;
  assign n2744 = ( x40 & n840 ) | ( x40 & n891 ) | ( n840 & n891 ) ;
  assign n2745 = n1310 ^ n1188 ^ n629 ;
  assign n2746 = n2745 ^ n2724 ^ 1'b0 ;
  assign n2747 = n2744 & n2746 ;
  assign n2748 = n2747 ^ n2539 ^ x167 ;
  assign n2749 = ( ~n2013 & n2743 ) | ( ~n2013 & n2748 ) | ( n2743 & n2748 ) ;
  assign n2730 = n2308 ^ n1494 ^ n1151 ;
  assign n2731 = ( x12 & n893 ) | ( x12 & n1777 ) | ( n893 & n1777 ) ;
  assign n2734 = x174 & n1249 ;
  assign n2735 = n663 & n2734 ;
  assign n2732 = n1601 ^ n1593 ^ x116 ;
  assign n2733 = n2732 ^ n399 ^ x156 ;
  assign n2736 = n2735 ^ n2733 ^ n943 ;
  assign n2737 = ( n929 & n2731 ) | ( n929 & n2736 ) | ( n2731 & n2736 ) ;
  assign n2738 = ( n746 & n2730 ) | ( n746 & ~n2737 ) | ( n2730 & ~n2737 ) ;
  assign n2739 = n2544 & ~n2738 ;
  assign n2740 = n2739 ^ x193 ^ 1'b0 ;
  assign n2741 = x107 & ~n2740 ;
  assign n2750 = n2749 ^ n2741 ^ n1581 ;
  assign n2753 = n2752 ^ n2750 ^ n2733 ;
  assign n2754 = ( n806 & n829 ) | ( n806 & n2153 ) | ( n829 & n2153 ) ;
  assign n2755 = n2754 ^ n343 ^ n290 ;
  assign n2756 = n2755 ^ n2269 ^ 1'b0 ;
  assign n2757 = ( ~n391 & n1336 ) | ( ~n391 & n2263 ) | ( n1336 & n2263 ) ;
  assign n2758 = n2247 ^ n2068 ^ n521 ;
  assign n2759 = n1171 ^ n938 ^ n440 ;
  assign n2760 = ( n2757 & n2758 ) | ( n2757 & ~n2759 ) | ( n2758 & ~n2759 ) ;
  assign n2761 = n2760 ^ n1100 ^ n460 ;
  assign n2762 = n1991 ^ n820 ^ n767 ;
  assign n2763 = n2762 ^ n304 ^ 1'b0 ;
  assign n2764 = n2761 | n2763 ;
  assign n2766 = ( n453 & n719 ) | ( n453 & ~n737 ) | ( n719 & ~n737 ) ;
  assign n2765 = n2723 ^ n452 ^ x159 ;
  assign n2767 = n2766 ^ n2765 ^ n580 ;
  assign n2768 = ( n1843 & n1865 ) | ( n1843 & n1875 ) | ( n1865 & n1875 ) ;
  assign n2769 = ( ~n276 & n1229 ) | ( ~n276 & n1527 ) | ( n1229 & n1527 ) ;
  assign n2770 = n1246 ^ n681 ^ x101 ;
  assign n2771 = ( n1023 & ~n2769 ) | ( n1023 & n2770 ) | ( ~n2769 & n2770 ) ;
  assign n2772 = n738 & ~n2771 ;
  assign n2773 = n2768 & n2772 ;
  assign n2775 = n2529 ^ n691 ^ x1 ;
  assign n2774 = n2108 ^ n1063 ^ x197 ;
  assign n2776 = n2775 ^ n2774 ^ n401 ;
  assign n2777 = n2776 ^ n1884 ^ 1'b0 ;
  assign n2778 = ( n2767 & ~n2773 ) | ( n2767 & n2777 ) | ( ~n2773 & n2777 ) ;
  assign n2786 = ( n1076 & n1089 ) | ( n1076 & ~n1424 ) | ( n1089 & ~n1424 ) ;
  assign n2783 = n1055 ^ n473 ^ 1'b0 ;
  assign n2781 = n662 ^ n259 ^ x140 ;
  assign n2782 = ( ~n679 & n2222 ) | ( ~n679 & n2781 ) | ( n2222 & n2781 ) ;
  assign n2779 = n400 ^ x124 ^ 1'b0 ;
  assign n2780 = ~n468 & n2779 ;
  assign n2784 = n2783 ^ n2782 ^ n2780 ;
  assign n2785 = n2784 ^ n2762 ^ n1264 ;
  assign n2787 = n2786 ^ n2785 ^ n2022 ;
  assign n2788 = n523 & ~n1415 ;
  assign n2789 = n274 & n598 ;
  assign n2790 = n882 & n2789 ;
  assign n2791 = n2790 ^ n272 ^ 1'b0 ;
  assign n2805 = x96 | n1440 ;
  assign n2803 = n1026 ^ x204 ^ 1'b0 ;
  assign n2804 = ( n1714 & n2371 ) | ( n1714 & ~n2803 ) | ( n2371 & ~n2803 ) ;
  assign n2796 = n393 ^ x195 ^ x161 ;
  assign n2794 = x50 & x169 ;
  assign n2795 = n396 & n2794 ;
  assign n2797 = n2796 ^ n2795 ^ n2097 ;
  assign n2798 = ~n662 & n2797 ;
  assign n2799 = n2798 ^ x186 ^ 1'b0 ;
  assign n2800 = n2799 ^ n2212 ^ n985 ;
  assign n2801 = ( n403 & n2238 ) | ( n403 & ~n2800 ) | ( n2238 & ~n2800 ) ;
  assign n2792 = n297 & n580 ;
  assign n2793 = n1772 & n2792 ;
  assign n2802 = n2801 ^ n2793 ^ n1151 ;
  assign n2806 = n2805 ^ n2804 ^ n2802 ;
  assign n2807 = n1362 ^ n601 ^ 1'b0 ;
  assign n2808 = ( n1356 & n1458 ) | ( n1356 & n2807 ) | ( n1458 & n2807 ) ;
  assign n2809 = n1809 ^ n445 ^ n437 ;
  assign n2810 = n902 ^ x169 ^ 1'b0 ;
  assign n2811 = x200 & ~n2810 ;
  assign n2812 = n1807 & n2811 ;
  assign n2813 = ~n2809 & n2812 ;
  assign n2814 = ( n2410 & n2505 ) | ( n2410 & n2813 ) | ( n2505 & n2813 ) ;
  assign n2819 = ( n904 & ~n2034 ) | ( n904 & n2195 ) | ( ~n2034 & n2195 ) ;
  assign n2815 = n1271 ^ n377 ^ x144 ;
  assign n2816 = x203 & n2815 ;
  assign n2817 = ~n1224 & n2816 ;
  assign n2818 = n2817 ^ n801 ^ n613 ;
  assign n2820 = n2819 ^ n2818 ^ x170 ;
  assign n2839 = n1861 ^ n1103 ^ x98 ;
  assign n2821 = ( n1531 & n1532 ) | ( n1531 & n1842 ) | ( n1532 & n1842 ) ;
  assign n2822 = n2821 ^ n1850 ^ n1423 ;
  assign n2830 = ~n1227 & n2627 ;
  assign n2831 = n2830 ^ n1522 ^ 1'b0 ;
  assign n2832 = n1319 ^ n787 ^ x77 ;
  assign n2833 = ( n530 & n666 ) | ( n530 & n998 ) | ( n666 & n998 ) ;
  assign n2834 = ( x77 & ~n2832 ) | ( x77 & n2833 ) | ( ~n2832 & n2833 ) ;
  assign n2835 = ( x102 & n2831 ) | ( x102 & n2834 ) | ( n2831 & n2834 ) ;
  assign n2836 = ( x135 & n2435 ) | ( x135 & ~n2835 ) | ( n2435 & ~n2835 ) ;
  assign n2825 = ( ~n999 & n1511 ) | ( ~n999 & n2781 ) | ( n1511 & n2781 ) ;
  assign n2826 = n2825 ^ n1186 ^ x189 ;
  assign n2827 = n2826 ^ n760 ^ n351 ;
  assign n2828 = ( n962 & n1393 ) | ( n962 & ~n2827 ) | ( n1393 & ~n2827 ) ;
  assign n2829 = ( n1407 & n1633 ) | ( n1407 & n2828 ) | ( n1633 & n2828 ) ;
  assign n2823 = ( n349 & n751 ) | ( n349 & ~n942 ) | ( n751 & ~n942 ) ;
  assign n2824 = ( x199 & ~n1895 ) | ( x199 & n2823 ) | ( ~n1895 & n2823 ) ;
  assign n2837 = n2836 ^ n2829 ^ n2824 ;
  assign n2838 = ( n2721 & n2822 ) | ( n2721 & n2837 ) | ( n2822 & n2837 ) ;
  assign n2840 = n2839 ^ n2838 ^ x56 ;
  assign n2841 = n2840 ^ n1644 ^ n1417 ;
  assign n2842 = ( ~x37 & n955 ) | ( ~x37 & n1276 ) | ( n955 & n1276 ) ;
  assign n2843 = n2842 ^ n1637 ^ n1445 ;
  assign n2844 = n653 ^ x217 ^ 1'b0 ;
  assign n2845 = n2844 ^ n2136 ^ n1154 ;
  assign n2846 = ( n1094 & ~n2843 ) | ( n1094 & n2845 ) | ( ~n2843 & n2845 ) ;
  assign n2847 = ( n799 & n1286 ) | ( n799 & ~n2458 ) | ( n1286 & ~n2458 ) ;
  assign n2848 = n1924 | n2847 ;
  assign n2849 = n2848 ^ x210 ^ 1'b0 ;
  assign n2850 = n1095 ^ n406 ^ x115 ;
  assign n2851 = ( n604 & ~n2100 ) | ( n604 & n2850 ) | ( ~n2100 & n2850 ) ;
  assign n2852 = ~n2849 & n2851 ;
  assign n2853 = ( n1180 & n1868 ) | ( n1180 & n1875 ) | ( n1868 & n1875 ) ;
  assign n2854 = n2273 ^ n2251 ^ n1274 ;
  assign n2855 = ( n632 & ~n2620 ) | ( n632 & n2854 ) | ( ~n2620 & n2854 ) ;
  assign n2856 = n2855 ^ n636 ^ 1'b0 ;
  assign n2857 = ( x38 & n2853 ) | ( x38 & n2856 ) | ( n2853 & n2856 ) ;
  assign n2858 = n1305 ^ n898 ^ 1'b0 ;
  assign n2859 = n2858 ^ n2052 ^ x41 ;
  assign n2860 = ( ~n544 & n1010 ) | ( ~n544 & n1187 ) | ( n1010 & n1187 ) ;
  assign n2861 = n2860 ^ n2576 ^ n814 ;
  assign n2862 = ( n551 & ~n785 ) | ( n551 & n2359 ) | ( ~n785 & n2359 ) ;
  assign n2864 = n726 | n1504 ;
  assign n2863 = n1631 ^ n655 ^ n315 ;
  assign n2865 = n2864 ^ n2863 ^ n1166 ;
  assign n2866 = ( x165 & n2862 ) | ( x165 & n2865 ) | ( n2862 & n2865 ) ;
  assign n2867 = ( ~n941 & n2861 ) | ( ~n941 & n2866 ) | ( n2861 & n2866 ) ;
  assign n2868 = n2867 ^ n2484 ^ n370 ;
  assign n2885 = ( ~n772 & n817 ) | ( ~n772 & n956 ) | ( n817 & n956 ) ;
  assign n2886 = n2885 ^ n580 ^ n398 ;
  assign n2869 = n1308 ^ n1272 ^ n595 ;
  assign n2870 = n596 ^ n363 ^ x74 ;
  assign n2871 = ~n1351 & n2870 ;
  assign n2881 = ( n554 & n590 ) | ( n554 & n1807 ) | ( n590 & n1807 ) ;
  assign n2878 = ( n718 & n852 ) | ( n718 & ~n1716 ) | ( n852 & ~n1716 ) ;
  assign n2877 = n2651 ^ n1695 ^ n1322 ;
  assign n2879 = n2878 ^ n2877 ^ n1507 ;
  assign n2872 = n1930 ^ n1502 ^ n1069 ;
  assign n2873 = n772 & ~n2031 ;
  assign n2874 = n2873 ^ n681 ^ 1'b0 ;
  assign n2875 = ( ~n1706 & n2183 ) | ( ~n1706 & n2874 ) | ( n2183 & n2874 ) ;
  assign n2876 = n2872 & n2875 ;
  assign n2880 = n2879 ^ n2876 ^ 1'b0 ;
  assign n2882 = n2881 ^ n2880 ^ 1'b0 ;
  assign n2883 = n1089 & n2882 ;
  assign n2884 = ( ~n2869 & n2871 ) | ( ~n2869 & n2883 ) | ( n2871 & n2883 ) ;
  assign n2887 = n2886 ^ n2884 ^ n571 ;
  assign n2888 = ( ~x34 & x173 ) | ( ~x34 & n677 ) | ( x173 & n677 ) ;
  assign n2889 = ( x75 & n1637 ) | ( x75 & ~n2888 ) | ( n1637 & ~n2888 ) ;
  assign n2890 = n2889 ^ n313 ^ n295 ;
  assign n2891 = ( ~n600 & n785 ) | ( ~n600 & n801 ) | ( n785 & n801 ) ;
  assign n2892 = n1620 ^ n821 ^ 1'b0 ;
  assign n2893 = n2184 | n2892 ;
  assign n2894 = ( x253 & n666 ) | ( x253 & ~n2893 ) | ( n666 & ~n2893 ) ;
  assign n2895 = ( ~x97 & n2891 ) | ( ~x97 & n2894 ) | ( n2891 & n2894 ) ;
  assign n2896 = ~n2890 & n2895 ;
  assign n2897 = n2896 ^ n282 ^ 1'b0 ;
  assign n2898 = ( x114 & ~n1298 ) | ( x114 & n2056 ) | ( ~n1298 & n2056 ) ;
  assign n2899 = n2898 ^ n2185 ^ n1165 ;
  assign n2900 = n2680 ^ n2613 ^ n1182 ;
  assign n2901 = n2899 & ~n2900 ;
  assign n2904 = n1855 ^ n462 ^ 1'b0 ;
  assign n2905 = n1729 & ~n2904 ;
  assign n2906 = ~n1801 & n2864 ;
  assign n2907 = ~n2905 & n2906 ;
  assign n2902 = n856 ^ n506 ^ x45 ;
  assign n2903 = n1206 & n2902 ;
  assign n2908 = n2907 ^ n2903 ^ 1'b0 ;
  assign n2909 = ( ~n1395 & n2275 ) | ( ~n1395 & n2908 ) | ( n2275 & n2908 ) ;
  assign n2917 = n2375 ^ n918 ^ n566 ;
  assign n2910 = n686 ^ n439 ^ x4 ;
  assign n2911 = ( n278 & n1540 ) | ( n278 & ~n2691 ) | ( n1540 & ~n2691 ) ;
  assign n2912 = n2910 & ~n2911 ;
  assign n2913 = n1825 ^ n312 ^ x250 ;
  assign n2914 = n1785 ^ n1333 ^ n740 ;
  assign n2915 = ( ~n1877 & n2913 ) | ( ~n1877 & n2914 ) | ( n2913 & n2914 ) ;
  assign n2916 = ( n1088 & ~n2912 ) | ( n1088 & n2915 ) | ( ~n2912 & n2915 ) ;
  assign n2918 = n2917 ^ n2916 ^ n2617 ;
  assign n2919 = ( n1236 & n1394 ) | ( n1236 & ~n2181 ) | ( n1394 & ~n2181 ) ;
  assign n2920 = n2919 ^ n1823 ^ n882 ;
  assign n2921 = ( ~n1356 & n2752 ) | ( ~n1356 & n2920 ) | ( n2752 & n2920 ) ;
  assign n2922 = ~n1424 & n2921 ;
  assign n2923 = ( n1996 & n2130 ) | ( n1996 & ~n2922 ) | ( n2130 & ~n2922 ) ;
  assign n2930 = n1102 ^ n863 ^ n499 ;
  assign n2931 = n2930 ^ n1362 ^ 1'b0 ;
  assign n2932 = n1036 | n2931 ;
  assign n2924 = ~n1257 & n2311 ;
  assign n2925 = ~n615 & n2924 ;
  assign n2926 = n2603 ^ n2365 ^ n2349 ;
  assign n2927 = n2926 ^ n2117 ^ n1534 ;
  assign n2928 = n2927 ^ n1638 ^ 1'b0 ;
  assign n2929 = n2925 | n2928 ;
  assign n2933 = n2932 ^ n2929 ^ n1680 ;
  assign n2937 = ( x145 & x195 ) | ( x145 & ~n368 ) | ( x195 & ~n368 ) ;
  assign n2935 = ( ~x195 & n286 ) | ( ~x195 & n1509 ) | ( n286 & n1509 ) ;
  assign n2934 = ( n876 & ~n1569 ) | ( n876 & n1631 ) | ( ~n1569 & n1631 ) ;
  assign n2936 = n2935 ^ n2934 ^ n2723 ;
  assign n2938 = n2937 ^ n2936 ^ n2368 ;
  assign n2939 = x171 & n559 ;
  assign n2940 = n2939 ^ n1567 ^ 1'b0 ;
  assign n2943 = n1479 ^ n1424 ^ n339 ;
  assign n2941 = n1907 ^ n1777 ^ n1409 ;
  assign n2942 = ( ~n1147 & n1787 ) | ( ~n1147 & n2941 ) | ( n1787 & n2941 ) ;
  assign n2944 = n2943 ^ n2942 ^ n1409 ;
  assign n2945 = ( n1660 & ~n2940 ) | ( n1660 & n2944 ) | ( ~n2940 & n2944 ) ;
  assign n2946 = n2945 ^ n814 ^ 1'b0 ;
  assign n2947 = ~n2938 & n2946 ;
  assign n2948 = n2807 ^ n2643 ^ n1901 ;
  assign n2951 = n2031 ^ n1517 ^ n683 ;
  assign n2952 = n2951 ^ n2668 ^ n2657 ;
  assign n2949 = ( n299 & ~n1644 ) | ( n299 & n1796 ) | ( ~n1644 & n1796 ) ;
  assign n2950 = n1001 & ~n2949 ;
  assign n2953 = n2952 ^ n2950 ^ 1'b0 ;
  assign n2954 = ( x29 & ~n1464 ) | ( x29 & n2953 ) | ( ~n1464 & n2953 ) ;
  assign n2960 = n1724 ^ n1165 ^ n332 ;
  assign n2961 = n2960 ^ n2031 ^ 1'b0 ;
  assign n2962 = n2402 & ~n2961 ;
  assign n2958 = n1909 ^ n653 ^ n404 ;
  assign n2956 = ( x109 & ~n866 ) | ( x109 & n2703 ) | ( ~n866 & n2703 ) ;
  assign n2955 = ( n365 & n882 ) | ( n365 & n1806 ) | ( n882 & n1806 ) ;
  assign n2957 = n2956 ^ n2955 ^ x227 ;
  assign n2959 = n2958 ^ n2957 ^ n2186 ;
  assign n2963 = n2962 ^ n2959 ^ n1639 ;
  assign n2964 = ( n399 & n1848 ) | ( n399 & ~n2963 ) | ( n1848 & ~n2963 ) ;
  assign n2965 = ( n1052 & n1975 ) | ( n1052 & n2290 ) | ( n1975 & n2290 ) ;
  assign n2969 = n821 | n1267 ;
  assign n2966 = n453 ^ x116 ^ x115 ;
  assign n2967 = ( ~x214 & n308 ) | ( ~x214 & n2966 ) | ( n308 & n2966 ) ;
  assign n2968 = n2967 ^ n2124 ^ n940 ;
  assign n2970 = n2969 ^ n2968 ^ x216 ;
  assign n2973 = n499 | n1725 ;
  assign n2974 = n2973 ^ n1121 ^ 1'b0 ;
  assign n2975 = ( x8 & n2774 ) | ( x8 & n2974 ) | ( n2774 & n2974 ) ;
  assign n2971 = n1536 ^ n874 ^ n362 ;
  assign n2972 = ( n1537 & ~n1969 ) | ( n1537 & n2971 ) | ( ~n1969 & n2971 ) ;
  assign n2976 = n2975 ^ n2972 ^ n599 ;
  assign n2985 = n969 ^ n967 ^ n738 ;
  assign n2984 = n1924 ^ n1817 ^ n1094 ;
  assign n2979 = ( ~x55 & n456 ) | ( ~x55 & n891 ) | ( n456 & n891 ) ;
  assign n2977 = ( n324 & n423 ) | ( n324 & ~n1367 ) | ( n423 & ~n1367 ) ;
  assign n2978 = n2977 ^ n2329 ^ n1098 ;
  assign n2980 = n2979 ^ n2978 ^ n2216 ;
  assign n2981 = n2980 ^ n760 ^ n732 ;
  assign n2982 = ( ~n304 & n2529 ) | ( ~n304 & n2981 ) | ( n2529 & n2981 ) ;
  assign n2983 = n2982 ^ n1318 ^ n544 ;
  assign n2986 = n2985 ^ n2984 ^ n2983 ;
  assign n2987 = ( ~x159 & n435 ) | ( ~x159 & n1301 ) | ( n435 & n1301 ) ;
  assign n2988 = n1392 & ~n2987 ;
  assign n2989 = n2988 ^ n2486 ^ 1'b0 ;
  assign n2990 = ( n457 & ~n835 ) | ( n457 & n2989 ) | ( ~n835 & n2989 ) ;
  assign n2991 = n2990 ^ n1628 ^ n1158 ;
  assign n2992 = n1861 ^ n1626 ^ n895 ;
  assign n2993 = n2992 ^ n1069 ^ x69 ;
  assign n2994 = ( ~n2145 & n2400 ) | ( ~n2145 & n2993 ) | ( n2400 & n2993 ) ;
  assign n2995 = n2700 ^ n2268 ^ n1592 ;
  assign n2996 = ( ~n661 & n663 ) | ( ~n661 & n2995 ) | ( n663 & n2995 ) ;
  assign n2997 = ( n826 & n2994 ) | ( n826 & ~n2996 ) | ( n2994 & ~n2996 ) ;
  assign n2998 = ( ~x239 & n654 ) | ( ~x239 & n2997 ) | ( n654 & n2997 ) ;
  assign n2999 = ( n2160 & n2991 ) | ( n2160 & ~n2998 ) | ( n2991 & ~n2998 ) ;
  assign n3000 = n2499 ^ n2247 ^ 1'b0 ;
  assign n3001 = n2207 ^ n1517 ^ 1'b0 ;
  assign n3002 = ~n3000 & n3001 ;
  assign n3003 = n3002 ^ n2043 ^ n1657 ;
  assign n3006 = ( x30 & x211 ) | ( x30 & n713 ) | ( x211 & n713 ) ;
  assign n3007 = ( x68 & n666 ) | ( x68 & ~n3006 ) | ( n666 & ~n3006 ) ;
  assign n3008 = ( x166 & n2603 ) | ( x166 & ~n3007 ) | ( n2603 & ~n3007 ) ;
  assign n3004 = ( x156 & x205 ) | ( x156 & ~x215 ) | ( x205 & ~x215 ) ;
  assign n3005 = n3004 ^ n1191 ^ n945 ;
  assign n3009 = n3008 ^ n3005 ^ n848 ;
  assign n3010 = n1276 & n3009 ;
  assign n3011 = ~n726 & n3010 ;
  assign n3012 = n3011 ^ n2548 ^ n1053 ;
  assign n3013 = n693 ^ n579 ^ x92 ;
  assign n3014 = n660 | n1101 ;
  assign n3015 = ( n2913 & n3013 ) | ( n2913 & ~n3014 ) | ( n3013 & ~n3014 ) ;
  assign n3016 = n2239 ^ n356 ^ x189 ;
  assign n3017 = n759 & ~n3016 ;
  assign n3018 = n3015 & n3017 ;
  assign n3019 = n3012 & ~n3018 ;
  assign n3020 = ( n2567 & ~n3003 ) | ( n2567 & n3019 ) | ( ~n3003 & n3019 ) ;
  assign n3021 = n1348 & n3004 ;
  assign n3022 = ~n1696 & n3021 ;
  assign n3023 = n3022 ^ n2211 ^ x185 ;
  assign n3024 = n2205 ^ n1154 ^ x22 ;
  assign n3025 = ( n460 & ~n1459 ) | ( n460 & n2819 ) | ( ~n1459 & n2819 ) ;
  assign n3026 = n3025 ^ n563 ^ 1'b0 ;
  assign n3027 = ~n3024 & n3026 ;
  assign n3028 = n1582 & n3027 ;
  assign n3029 = n3023 | n3028 ;
  assign n3030 = n1208 & ~n3029 ;
  assign n3031 = n2147 ^ n2143 ^ n335 ;
  assign n3032 = n3031 ^ n1161 ^ 1'b0 ;
  assign n3038 = n1720 ^ n1349 ^ 1'b0 ;
  assign n3033 = ~n301 & n669 ;
  assign n3034 = ~x228 & n3033 ;
  assign n3035 = n915 ^ n384 ^ x53 ;
  assign n3036 = n3035 ^ n2140 ^ n388 ;
  assign n3037 = ( ~n2190 & n3034 ) | ( ~n2190 & n3036 ) | ( n3034 & n3036 ) ;
  assign n3039 = n3038 ^ n3037 ^ 1'b0 ;
  assign n3049 = n660 & ~n774 ;
  assign n3045 = ( x129 & n1325 ) | ( x129 & ~n1915 ) | ( n1325 & ~n1915 ) ;
  assign n3046 = n3045 ^ n1887 ^ 1'b0 ;
  assign n3047 = n2823 | n3046 ;
  assign n3043 = n819 & ~n1158 ;
  assign n3040 = ( x40 & n953 ) | ( x40 & ~n2760 ) | ( n953 & ~n2760 ) ;
  assign n3041 = ~n362 & n3040 ;
  assign n3042 = n1948 & n3041 ;
  assign n3044 = n3043 ^ n3042 ^ n2203 ;
  assign n3048 = n3047 ^ n3044 ^ n3042 ;
  assign n3050 = n3049 ^ n3048 ^ n2224 ;
  assign n3051 = n666 ^ n508 ^ n303 ;
  assign n3052 = ( x229 & ~n516 ) | ( x229 & n1072 ) | ( ~n516 & n1072 ) ;
  assign n3053 = ( n269 & n613 ) | ( n269 & n2089 ) | ( n613 & n2089 ) ;
  assign n3054 = ( n2590 & ~n3052 ) | ( n2590 & n3053 ) | ( ~n3052 & n3053 ) ;
  assign n3055 = n3051 | n3054 ;
  assign n3056 = n3055 ^ n2229 ^ 1'b0 ;
  assign n3057 = n3056 ^ n378 ^ 1'b0 ;
  assign n3058 = n3057 ^ n1552 ^ 1'b0 ;
  assign n3059 = n3058 ^ n711 ^ 1'b0 ;
  assign n3067 = n2769 ^ n1476 ^ n1111 ;
  assign n3065 = ( n273 & ~n1014 ) | ( n273 & n2971 ) | ( ~n1014 & n2971 ) ;
  assign n3062 = ( x215 & ~n1015 ) | ( x215 & n1029 ) | ( ~n1015 & n1029 ) ;
  assign n3063 = n3062 ^ n609 ^ n403 ;
  assign n3060 = n450 | n2790 ;
  assign n3061 = n3060 ^ n843 ^ 1'b0 ;
  assign n3064 = n3063 ^ n3061 ^ 1'b0 ;
  assign n3066 = n3065 ^ n3064 ^ n2133 ;
  assign n3068 = n3067 ^ n3066 ^ n1510 ;
  assign n3069 = n1960 ^ n1593 ^ x65 ;
  assign n3070 = n3069 ^ n721 ^ n533 ;
  assign n3071 = ( n1164 & ~n1362 ) | ( n1164 & n1775 ) | ( ~n1362 & n1775 ) ;
  assign n3072 = ( n287 & n1375 ) | ( n287 & ~n3071 ) | ( n1375 & ~n3071 ) ;
  assign n3073 = ( n2698 & n3070 ) | ( n2698 & n3072 ) | ( n3070 & n3072 ) ;
  assign n3074 = n3073 ^ x171 ^ x104 ;
  assign n3075 = n3074 ^ n1469 ^ n739 ;
  assign n3076 = n676 | n2892 ;
  assign n3077 = n3076 ^ n1211 ^ 1'b0 ;
  assign n3078 = n2341 & n3077 ;
  assign n3079 = ( x175 & n341 ) | ( x175 & ~n1958 ) | ( n341 & ~n1958 ) ;
  assign n3080 = ( n954 & n1192 ) | ( n954 & n1779 ) | ( n1192 & n1779 ) ;
  assign n3081 = n3080 ^ n1401 ^ 1'b0 ;
  assign n3084 = ( n1521 & n2521 ) | ( n1521 & n2602 ) | ( n2521 & n2602 ) ;
  assign n3082 = ( ~x121 & n2411 ) | ( ~x121 & n2515 ) | ( n2411 & n2515 ) ;
  assign n3083 = n3082 ^ n1451 ^ n916 ;
  assign n3085 = n3084 ^ n3083 ^ n1257 ;
  assign n3086 = ( n2236 & n3081 ) | ( n2236 & n3085 ) | ( n3081 & n3085 ) ;
  assign n3087 = ( ~n1058 & n3079 ) | ( ~n1058 & n3086 ) | ( n3079 & n3086 ) ;
  assign n3092 = ( ~n702 & n1219 ) | ( ~n702 & n1401 ) | ( n1219 & n1401 ) ;
  assign n3089 = n1409 ^ n1265 ^ x102 ;
  assign n3090 = n3089 ^ n1325 ^ n886 ;
  assign n3091 = ( n897 & n1730 ) | ( n897 & n3090 ) | ( n1730 & n3090 ) ;
  assign n3088 = n1812 ^ n469 ^ x92 ;
  assign n3093 = n3092 ^ n3091 ^ n3088 ;
  assign n3102 = n653 ^ n552 ^ n551 ;
  assign n3103 = n3102 ^ n2171 ^ n1567 ;
  assign n3099 = ~n1159 & n1432 ;
  assign n3100 = ~n1657 & n3099 ;
  assign n3098 = ( n515 & n802 ) | ( n515 & ~n965 ) | ( n802 & ~n965 ) ;
  assign n3094 = n1991 ^ n1014 ^ x211 ;
  assign n3095 = n3094 ^ n2342 ^ n1028 ;
  assign n3096 = n943 & ~n3095 ;
  assign n3097 = ~n257 & n3096 ;
  assign n3101 = n3100 ^ n3098 ^ n3097 ;
  assign n3104 = n3103 ^ n3101 ^ n2101 ;
  assign n3106 = n1269 ^ n1125 ^ x231 ;
  assign n3105 = ( n1942 & n2201 ) | ( n1942 & ~n2358 ) | ( n2201 & ~n2358 ) ;
  assign n3107 = n3106 ^ n3105 ^ 1'b0 ;
  assign n3108 = ( n619 & n728 ) | ( n619 & ~n1143 ) | ( n728 & ~n1143 ) ;
  assign n3109 = ( ~x90 & n1656 ) | ( ~x90 & n1666 ) | ( n1656 & n1666 ) ;
  assign n3110 = ( ~n1638 & n1670 ) | ( ~n1638 & n3109 ) | ( n1670 & n3109 ) ;
  assign n3111 = n3108 & n3110 ;
  assign n3112 = ~x252 & n3111 ;
  assign n3113 = n3112 ^ n1019 ^ 1'b0 ;
  assign n3114 = x57 & n3113 ;
  assign n3115 = n1894 ^ n889 ^ 1'b0 ;
  assign n3116 = n762 ^ x154 ^ x41 ;
  assign n3117 = n3116 ^ n3008 ^ n2825 ;
  assign n3118 = ( ~n782 & n3115 ) | ( ~n782 & n3117 ) | ( n3115 & n3117 ) ;
  assign n3119 = ( ~x106 & n681 ) | ( ~x106 & n2199 ) | ( n681 & n2199 ) ;
  assign n3120 = ( n1518 & n2282 ) | ( n1518 & ~n3119 ) | ( n2282 & ~n3119 ) ;
  assign n3121 = n3120 ^ n2606 ^ n1501 ;
  assign n3122 = x87 & x141 ;
  assign n3123 = n3122 ^ x192 ^ 1'b0 ;
  assign n3124 = ( x8 & n848 ) | ( x8 & n1668 ) | ( n848 & n1668 ) ;
  assign n3125 = ( n1317 & n1473 ) | ( n1317 & ~n3124 ) | ( n1473 & ~n3124 ) ;
  assign n3126 = n3123 & ~n3125 ;
  assign n3127 = n529 & n1332 ;
  assign n3128 = ~n3126 & n3127 ;
  assign n3129 = n1868 & n3128 ;
  assign n3130 = ( n631 & n2744 ) | ( n631 & ~n3094 ) | ( n2744 & ~n3094 ) ;
  assign n3131 = n3130 ^ n810 ^ n673 ;
  assign n3132 = n2197 ^ x89 ^ x88 ;
  assign n3133 = ( n2822 & n3131 ) | ( n2822 & ~n3132 ) | ( n3131 & ~n3132 ) ;
  assign n3134 = ( x160 & n1794 ) | ( x160 & n2169 ) | ( n1794 & n2169 ) ;
  assign n3135 = ( ~x194 & n3133 ) | ( ~x194 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3136 = n3092 & n3135 ;
  assign n3137 = n3079 & n3136 ;
  assign n3145 = n813 & n2854 ;
  assign n3146 = n3145 ^ n1576 ^ 1'b0 ;
  assign n3147 = ( ~n372 & n1551 ) | ( ~n372 & n2949 ) | ( n1551 & n2949 ) ;
  assign n3148 = ~n326 & n1361 ;
  assign n3149 = ( ~n3146 & n3147 ) | ( ~n3146 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3142 = n1145 ^ n304 ^ x34 ;
  assign n3139 = ( n687 & n1305 ) | ( n687 & n1868 ) | ( n1305 & n1868 ) ;
  assign n3138 = ( n577 & n2127 ) | ( n577 & ~n2655 ) | ( n2127 & ~n2655 ) ;
  assign n3140 = n3139 ^ n3138 ^ n306 ;
  assign n3141 = n3140 ^ n1649 ^ n365 ;
  assign n3143 = n3142 ^ n3141 ^ n3014 ;
  assign n3144 = n3032 & ~n3143 ;
  assign n3150 = n3149 ^ n3144 ^ 1'b0 ;
  assign n3151 = n753 ^ n729 ^ n328 ;
  assign n3152 = ( ~n411 & n607 ) | ( ~n411 & n3151 ) | ( n607 & n3151 ) ;
  assign n3153 = n3152 ^ n2241 ^ n1704 ;
  assign n3154 = n3153 ^ n2902 ^ x63 ;
  assign n3155 = ( n292 & ~n894 ) | ( n292 & n3154 ) | ( ~n894 & n3154 ) ;
  assign n3157 = ( n1143 & n2037 ) | ( n1143 & n2156 ) | ( n2037 & n2156 ) ;
  assign n3156 = ( x89 & ~n418 ) | ( x89 & n789 ) | ( ~n418 & n789 ) ;
  assign n3158 = n3157 ^ n3156 ^ n1341 ;
  assign n3159 = n471 & n1903 ;
  assign n3160 = ( x179 & ~n1898 ) | ( x179 & n3159 ) | ( ~n1898 & n3159 ) ;
  assign n3161 = n1683 ^ n610 ^ 1'b0 ;
  assign n3162 = n2711 & n3161 ;
  assign n3166 = n260 & ~n1478 ;
  assign n3167 = n3166 ^ x167 ^ 1'b0 ;
  assign n3165 = ( n256 & n1230 ) | ( n256 & ~n1317 ) | ( n1230 & ~n1317 ) ;
  assign n3164 = n2196 ^ n1050 ^ 1'b0 ;
  assign n3168 = n3167 ^ n3165 ^ n3164 ;
  assign n3163 = n651 & ~n3116 ;
  assign n3169 = n3168 ^ n3163 ^ 1'b0 ;
  assign n3170 = ( n3142 & ~n3162 ) | ( n3142 & n3169 ) | ( ~n3162 & n3169 ) ;
  assign n3180 = ( x49 & n277 ) | ( x49 & ~n838 ) | ( n277 & ~n838 ) ;
  assign n3181 = ( x59 & n2969 ) | ( x59 & ~n3180 ) | ( n2969 & ~n3180 ) ;
  assign n3171 = n726 ^ n495 ^ n333 ;
  assign n3172 = n789 ^ n699 ^ n411 ;
  assign n3173 = ( ~n464 & n2405 ) | ( ~n464 & n3172 ) | ( n2405 & n3172 ) ;
  assign n3174 = n1133 ^ n720 ^ n277 ;
  assign n3175 = n3174 ^ n2456 ^ n513 ;
  assign n3176 = ( n3171 & n3173 ) | ( n3171 & ~n3175 ) | ( n3173 & ~n3175 ) ;
  assign n3177 = n2536 ^ n1157 ^ n378 ;
  assign n3178 = n3177 ^ n2431 ^ n977 ;
  assign n3179 = ~n3176 & n3178 ;
  assign n3182 = n3181 ^ n3179 ^ 1'b0 ;
  assign n3186 = ~n572 & n1697 ;
  assign n3187 = n3186 ^ n3043 ^ 1'b0 ;
  assign n3188 = ~n2210 & n3187 ;
  assign n3184 = ( x78 & ~n1403 ) | ( x78 & n1660 ) | ( ~n1403 & n1660 ) ;
  assign n3183 = n3073 ^ n2492 ^ x150 ;
  assign n3185 = n3184 ^ n3183 ^ n1726 ;
  assign n3189 = n3188 ^ n3185 ^ n2980 ;
  assign n3190 = n1289 ^ n1007 ^ 1'b0 ;
  assign n3191 = n774 | n3190 ;
  assign n3192 = n3138 ^ n2822 ^ n1260 ;
  assign n3193 = n3192 ^ n2239 ^ 1'b0 ;
  assign n3194 = n739 & ~n3193 ;
  assign n3195 = n3194 ^ n880 ^ 1'b0 ;
  assign n3196 = ( n949 & n3191 ) | ( n949 & n3195 ) | ( n3191 & n3195 ) ;
  assign n3197 = n3196 ^ n1311 ^ n924 ;
  assign n3198 = ( n2272 & ~n2481 ) | ( n2272 & n2579 ) | ( ~n2481 & n2579 ) ;
  assign n3199 = ( n1599 & n1942 ) | ( n1599 & n2256 ) | ( n1942 & n2256 ) ;
  assign n3200 = n1665 ^ n1316 ^ n275 ;
  assign n3201 = ( n645 & ~n652 ) | ( n645 & n862 ) | ( ~n652 & n862 ) ;
  assign n3202 = n3201 ^ n1275 ^ x49 ;
  assign n3203 = n1823 ^ n329 ^ x182 ;
  assign n3204 = n3203 ^ x150 ^ x139 ;
  assign n3205 = ( n3200 & ~n3202 ) | ( n3200 & n3204 ) | ( ~n3202 & n3204 ) ;
  assign n3206 = ( n1309 & ~n3199 ) | ( n1309 & n3205 ) | ( ~n3199 & n3205 ) ;
  assign n3207 = ( ~x82 & n1957 ) | ( ~x82 & n3206 ) | ( n1957 & n3206 ) ;
  assign n3208 = n3198 | n3207 ;
  assign n3209 = n3208 ^ x199 ^ 1'b0 ;
  assign n3212 = ( n545 & n1448 ) | ( n545 & n2571 ) | ( n1448 & n2571 ) ;
  assign n3213 = ( x39 & ~n1074 ) | ( x39 & n3212 ) | ( ~n1074 & n3212 ) ;
  assign n3210 = n1801 ^ n1544 ^ n1212 ;
  assign n3211 = n3210 ^ x164 ^ x71 ;
  assign n3214 = n3213 ^ n3211 ^ n3173 ;
  assign n3215 = ~n1716 & n3214 ;
  assign n3224 = ( ~x122 & n1252 ) | ( ~x122 & n1437 ) | ( n1252 & n1437 ) ;
  assign n3222 = n3005 ^ n662 ^ n502 ;
  assign n3219 = n2181 ^ n1696 ^ n1448 ;
  assign n3220 = n3219 ^ n1301 ^ n826 ;
  assign n3218 = n2891 ^ n2669 ^ n719 ;
  assign n3216 = ~x183 & n593 ;
  assign n3217 = n3216 ^ n1440 ^ n1391 ;
  assign n3221 = n3220 ^ n3218 ^ n3217 ;
  assign n3223 = n3222 ^ n3221 ^ n2470 ;
  assign n3225 = n3224 ^ n3223 ^ n2268 ;
  assign n3226 = n3225 ^ n850 ^ 1'b0 ;
  assign n3227 = n2787 & n3226 ;
  assign n3228 = ( x18 & n1171 ) | ( x18 & ~n1957 ) | ( n1171 & ~n1957 ) ;
  assign n3229 = n3228 ^ n2593 ^ 1'b0 ;
  assign n3231 = ~n459 & n1249 ;
  assign n3232 = ~x89 & n3231 ;
  assign n3230 = ~x14 & x92 ;
  assign n3233 = n3232 ^ n3230 ^ n625 ;
  assign n3234 = n1774 ^ n1705 ^ x4 ;
  assign n3235 = ( x176 & ~n1537 ) | ( x176 & n1557 ) | ( ~n1537 & n1557 ) ;
  assign n3236 = ~n3234 & n3235 ;
  assign n3237 = n2718 ^ n395 ^ 1'b0 ;
  assign n3238 = ( n3233 & n3236 ) | ( n3233 & ~n3237 ) | ( n3236 & ~n3237 ) ;
  assign n3239 = n3238 ^ n1953 ^ n1010 ;
  assign n3240 = n2299 ^ n1208 ^ x109 ;
  assign n3241 = n3240 ^ n2329 ^ 1'b0 ;
  assign n3249 = n1322 ^ n1211 ^ n1046 ;
  assign n3250 = n876 | n1132 ;
  assign n3251 = n3250 ^ n2994 ^ n668 ;
  assign n3252 = ( n457 & ~n3249 ) | ( n457 & n3251 ) | ( ~n3249 & n3251 ) ;
  assign n3247 = ( n700 & n759 ) | ( n700 & n1556 ) | ( n759 & n1556 ) ;
  assign n3244 = ( x76 & n272 ) | ( x76 & ~n393 ) | ( n272 & ~n393 ) ;
  assign n3245 = ( ~n1256 & n1370 ) | ( ~n1256 & n3244 ) | ( n1370 & n3244 ) ;
  assign n3246 = n3245 ^ n1601 ^ n805 ;
  assign n3248 = n3247 ^ n3246 ^ x80 ;
  assign n3242 = n2853 ^ n2207 ^ n506 ;
  assign n3243 = n3242 ^ n1695 ^ n894 ;
  assign n3253 = n3252 ^ n3248 ^ n3243 ;
  assign n3254 = n2892 ^ n821 ^ n431 ;
  assign n3255 = n1502 ^ n1220 ^ n760 ;
  assign n3256 = ( ~x144 & n2775 ) | ( ~x144 & n3255 ) | ( n2775 & n3255 ) ;
  assign n3257 = n3256 ^ n3036 ^ n1059 ;
  assign n3258 = n650 ^ n476 ^ 1'b0 ;
  assign n3259 = n355 & ~n3258 ;
  assign n3260 = ( ~x28 & n758 ) | ( ~x28 & n3259 ) | ( n758 & n3259 ) ;
  assign n3261 = n3260 ^ n774 ^ n627 ;
  assign n3262 = ( n716 & n1047 ) | ( n716 & ~n3261 ) | ( n1047 & ~n3261 ) ;
  assign n3263 = n3262 ^ n1898 ^ 1'b0 ;
  assign n3264 = ( n277 & ~n765 ) | ( n277 & n1551 ) | ( ~n765 & n1551 ) ;
  assign n3265 = ( n1367 & ~n3115 ) | ( n1367 & n3264 ) | ( ~n3115 & n3264 ) ;
  assign n3266 = ( n936 & n3263 ) | ( n936 & ~n3265 ) | ( n3263 & ~n3265 ) ;
  assign n3267 = n2185 & n3266 ;
  assign n3268 = n1555 ^ n510 ^ 1'b0 ;
  assign n3269 = n596 & n3268 ;
  assign n3270 = ( ~x20 & n2864 ) | ( ~x20 & n3269 ) | ( n2864 & n3269 ) ;
  assign n3271 = n3270 ^ n1612 ^ n898 ;
  assign n3272 = n1080 ^ n777 ^ n391 ;
  assign n3273 = ( x195 & n2535 ) | ( x195 & n3272 ) | ( n2535 & n3272 ) ;
  assign n3274 = n3273 ^ n698 ^ 1'b0 ;
  assign n3276 = n1143 ^ n599 ^ n358 ;
  assign n3275 = n1937 | n2672 ;
  assign n3277 = n3276 ^ n3275 ^ n782 ;
  assign n3278 = n1249 & n3277 ;
  assign n3279 = n2654 ^ n2643 ^ n256 ;
  assign n3280 = ~n2972 & n3279 ;
  assign n3281 = ~n1812 & n3280 ;
  assign n3290 = ( ~x69 & n1343 ) | ( ~x69 & n2499 ) | ( n1343 & n2499 ) ;
  assign n3284 = ( n524 & n753 ) | ( n524 & n881 ) | ( n753 & n881 ) ;
  assign n3282 = ( n461 & n713 ) | ( n461 & n772 ) | ( n713 & n772 ) ;
  assign n3283 = n3282 ^ n1142 ^ n364 ;
  assign n3285 = n3284 ^ n3283 ^ n2344 ;
  assign n3286 = n1250 ^ n1079 ^ n718 ;
  assign n3287 = n3286 ^ n607 ^ x197 ;
  assign n3288 = n3287 ^ n3072 ^ n1351 ;
  assign n3289 = n3285 & ~n3288 ;
  assign n3291 = n3290 ^ n3289 ^ 1'b0 ;
  assign n3297 = n1925 ^ n799 ^ n753 ;
  assign n3292 = ( ~n1863 & n2250 ) | ( ~n1863 & n2668 ) | ( n2250 & n2668 ) ;
  assign n3293 = ( n1295 & n1619 ) | ( n1295 & n3123 ) | ( n1619 & n3123 ) ;
  assign n3294 = n3293 ^ n614 ^ 1'b0 ;
  assign n3295 = n617 | n3294 ;
  assign n3296 = n3292 & ~n3295 ;
  assign n3298 = n3297 ^ n3296 ^ n1301 ;
  assign n3299 = x223 & n763 ;
  assign n3300 = n1188 & n3299 ;
  assign n3301 = x154 & ~n1173 ;
  assign n3302 = n3301 ^ n1457 ^ 1'b0 ;
  assign n3303 = n3302 ^ n657 ^ n409 ;
  assign n3304 = ( ~n497 & n2110 ) | ( ~n497 & n3303 ) | ( n2110 & n3303 ) ;
  assign n3305 = ( n322 & n461 ) | ( n322 & n814 ) | ( n461 & n814 ) ;
  assign n3307 = n1192 ^ n978 ^ x246 ;
  assign n3306 = ( x154 & n314 ) | ( x154 & ~n2612 ) | ( n314 & ~n2612 ) ;
  assign n3308 = n3307 ^ n3306 ^ n2605 ;
  assign n3309 = ( n889 & n3202 ) | ( n889 & ~n3308 ) | ( n3202 & ~n3308 ) ;
  assign n3310 = ( ~n2579 & n3305 ) | ( ~n2579 & n3309 ) | ( n3305 & n3309 ) ;
  assign n3311 = ( ~n2265 & n3304 ) | ( ~n2265 & n3310 ) | ( n3304 & n3310 ) ;
  assign n3312 = ( n2613 & n3300 ) | ( n2613 & ~n3311 ) | ( n3300 & ~n3311 ) ;
  assign n3313 = n3312 ^ n2899 ^ n1981 ;
  assign n3317 = ( ~n1130 & n1304 ) | ( ~n1130 & n1309 ) | ( n1304 & n1309 ) ;
  assign n3314 = ( n1709 & ~n1861 ) | ( n1709 & n2181 ) | ( ~n1861 & n2181 ) ;
  assign n3315 = n1097 & n3314 ;
  assign n3316 = n1577 & n3315 ;
  assign n3318 = n3317 ^ n3316 ^ n1474 ;
  assign n3319 = n1267 ^ n610 ^ 1'b0 ;
  assign n3322 = n2211 ^ n546 ^ 1'b0 ;
  assign n3320 = ( n696 & ~n1533 ) | ( n696 & n1844 ) | ( ~n1533 & n1844 ) ;
  assign n3321 = n1408 & n3320 ;
  assign n3323 = n3322 ^ n3321 ^ 1'b0 ;
  assign n3324 = n3319 | n3323 ;
  assign n3325 = n3324 ^ n1371 ^ 1'b0 ;
  assign n3326 = n3325 ^ n700 ^ x183 ;
  assign n3327 = ( n2481 & ~n3318 ) | ( n2481 & n3326 ) | ( ~n3318 & n3326 ) ;
  assign n3328 = n2393 ^ n1408 ^ n1330 ;
  assign n3329 = n2723 ^ n1003 ^ x97 ;
  assign n3330 = n2667 & n3199 ;
  assign n3331 = n3329 & n3330 ;
  assign n3332 = n3331 ^ n2796 ^ n759 ;
  assign n3333 = ( ~n568 & n2216 ) | ( ~n568 & n3332 ) | ( n2216 & n3332 ) ;
  assign n3334 = ( n2236 & n3328 ) | ( n2236 & n3333 ) | ( n3328 & n3333 ) ;
  assign n3341 = ~n268 & n1700 ;
  assign n3342 = n3341 ^ n1061 ^ 1'b0 ;
  assign n3343 = n3342 ^ n2834 ^ n852 ;
  assign n3338 = n2552 ^ n1501 ^ n1051 ;
  assign n3339 = n3338 ^ n1285 ^ n1062 ;
  assign n3340 = n3339 ^ n1822 ^ n1403 ;
  assign n3335 = ( n1670 & n2174 ) | ( n1670 & ~n2755 ) | ( n2174 & ~n2755 ) ;
  assign n3336 = ( n362 & n907 ) | ( n362 & ~n1831 ) | ( n907 & ~n1831 ) ;
  assign n3337 = ( n382 & ~n3335 ) | ( n382 & n3336 ) | ( ~n3335 & n3336 ) ;
  assign n3344 = n3343 ^ n3340 ^ n3337 ;
  assign n3345 = n577 ^ x188 ^ x24 ;
  assign n3346 = ( n1395 & ~n2745 ) | ( n1395 & n3345 ) | ( ~n2745 & n3345 ) ;
  assign n3347 = n1994 ^ n751 ^ 1'b0 ;
  assign n3348 = n3347 ^ n1693 ^ n1150 ;
  assign n3349 = n3346 | n3348 ;
  assign n3352 = ( n940 & ~n1329 ) | ( n940 & n3142 ) | ( ~n1329 & n3142 ) ;
  assign n3350 = ( ~x113 & n2255 ) | ( ~x113 & n2509 ) | ( n2255 & n2509 ) ;
  assign n3351 = n1109 & ~n3350 ;
  assign n3353 = n3352 ^ n3351 ^ 1'b0 ;
  assign n3354 = n3353 ^ n2804 ^ x0 ;
  assign n3355 = ( n1201 & ~n2113 ) | ( n1201 & n2370 ) | ( ~n2113 & n2370 ) ;
  assign n3356 = n1030 & n3355 ;
  assign n3357 = ( ~x36 & n471 ) | ( ~x36 & n1317 ) | ( n471 & n1317 ) ;
  assign n3358 = ( n2233 & ~n2335 ) | ( n2233 & n3357 ) | ( ~n2335 & n3357 ) ;
  assign n3359 = n3358 ^ n2261 ^ 1'b0 ;
  assign n3360 = ( n2588 & n3356 ) | ( n2588 & ~n3359 ) | ( n3356 & ~n3359 ) ;
  assign n3361 = n3360 ^ n2778 ^ n502 ;
  assign n3364 = x50 & ~n692 ;
  assign n3365 = ~x181 & n3364 ;
  assign n3362 = n1437 & n2153 ;
  assign n3363 = n3362 ^ n2273 ^ 1'b0 ;
  assign n3366 = n3365 ^ n3363 ^ n2618 ;
  assign n3367 = ( n1154 & n1481 ) | ( n1154 & n3366 ) | ( n1481 & n3366 ) ;
  assign n3368 = n2955 ^ n2699 ^ n1205 ;
  assign n3369 = ( x214 & n780 ) | ( x214 & n3368 ) | ( n780 & n3368 ) ;
  assign n3370 = ( n3212 & ~n3367 ) | ( n3212 & n3369 ) | ( ~n3367 & n3369 ) ;
  assign n3371 = ( n2049 & ~n2440 ) | ( n2049 & n3112 ) | ( ~n2440 & n3112 ) ;
  assign n3372 = ( n1111 & n1309 ) | ( n1111 & n1646 ) | ( n1309 & n1646 ) ;
  assign n3373 = n1039 ^ n1035 ^ n983 ;
  assign n3374 = ( n840 & ~n2569 ) | ( n840 & n3373 ) | ( ~n2569 & n3373 ) ;
  assign n3375 = ( n851 & n2967 ) | ( n851 & ~n3374 ) | ( n2967 & ~n3374 ) ;
  assign n3376 = ( n462 & n828 ) | ( n462 & ~n3375 ) | ( n828 & ~n3375 ) ;
  assign n3377 = n3376 ^ n2590 ^ 1'b0 ;
  assign n3378 = ~n3372 & n3377 ;
  assign n3379 = n3378 ^ n2410 ^ n1217 ;
  assign n3380 = n2432 | n3379 ;
  assign n3382 = n1164 ^ n973 ^ n740 ;
  assign n3383 = n2201 ^ n652 ^ 1'b0 ;
  assign n3384 = ( n3056 & ~n3382 ) | ( n3056 & n3383 ) | ( ~n3382 & n3383 ) ;
  assign n3381 = n3259 ^ n1803 ^ n1109 ;
  assign n3385 = n3384 ^ n3381 ^ n1637 ;
  assign n3386 = n3385 ^ n1435 ^ 1'b0 ;
  assign n3390 = ( ~n359 & n442 ) | ( ~n359 & n2172 ) | ( n442 & n2172 ) ;
  assign n3387 = n2689 ^ n761 ^ 1'b0 ;
  assign n3388 = n3213 & ~n3387 ;
  assign n3389 = n3388 ^ n2344 ^ 1'b0 ;
  assign n3391 = n3390 ^ n3389 ^ n2249 ;
  assign n3392 = n3391 ^ n3091 ^ n1792 ;
  assign n3398 = n2687 ^ n2602 ^ n1343 ;
  assign n3393 = ( x42 & n1304 ) | ( x42 & n2598 ) | ( n1304 & n2598 ) ;
  assign n3394 = ~n687 & n2078 ;
  assign n3395 = ~n3151 & n3394 ;
  assign n3396 = ( ~n655 & n1392 ) | ( ~n655 & n3395 ) | ( n1392 & n3395 ) ;
  assign n3397 = n3393 & n3396 ;
  assign n3399 = n3398 ^ n3397 ^ 1'b0 ;
  assign n3400 = n2396 ^ n536 ^ x113 ;
  assign n3401 = ( n587 & ~n2300 ) | ( n587 & n3400 ) | ( ~n2300 & n3400 ) ;
  assign n3402 = n3401 ^ n1581 ^ n1114 ;
  assign n3403 = ( n2326 & ~n2430 ) | ( n2326 & n3402 ) | ( ~n2430 & n3402 ) ;
  assign n3404 = x90 & n3127 ;
  assign n3405 = n2499 ^ n640 ^ x63 ;
  assign n3406 = n1660 ^ n1227 ^ x180 ;
  assign n3407 = ( ~n2274 & n3405 ) | ( ~n2274 & n3406 ) | ( n3405 & n3406 ) ;
  assign n3408 = n3407 ^ n2697 ^ n2247 ;
  assign n3409 = ( n3051 & n3404 ) | ( n3051 & n3408 ) | ( n3404 & n3408 ) ;
  assign n3414 = n875 ^ n694 ^ n337 ;
  assign n3415 = ( n1221 & ~n3300 ) | ( n1221 & n3414 ) | ( ~n3300 & n3414 ) ;
  assign n3411 = n3357 ^ x132 ^ 1'b0 ;
  assign n3412 = n602 & ~n3411 ;
  assign n3413 = n3412 ^ n2350 ^ n2289 ;
  assign n3410 = n3242 ^ n2529 ^ x147 ;
  assign n3416 = n3415 ^ n3413 ^ n3410 ;
  assign n3417 = n1077 ^ n459 ^ n388 ;
  assign n3418 = n3417 ^ n2042 ^ 1'b0 ;
  assign n3419 = ~n2333 & n3418 ;
  assign n3420 = n3419 ^ n3172 ^ n2605 ;
  assign n3421 = n585 | n3054 ;
  assign n3422 = n3421 ^ n535 ^ 1'b0 ;
  assign n3423 = ( n750 & ~n2633 ) | ( n750 & n2782 ) | ( ~n2633 & n2782 ) ;
  assign n3424 = n3423 ^ x94 ^ x44 ;
  assign n3425 = ( n835 & ~n3422 ) | ( n835 & n3424 ) | ( ~n3422 & n3424 ) ;
  assign n3426 = ( n756 & ~n2011 ) | ( n756 & n3425 ) | ( ~n2011 & n3425 ) ;
  assign n3427 = ( x206 & n3420 ) | ( x206 & ~n3426 ) | ( n3420 & ~n3426 ) ;
  assign n3428 = n1232 & n1292 ;
  assign n3429 = n2328 ^ n914 ^ x72 ;
  assign n3430 = n2702 ^ n596 ^ n262 ;
  assign n3431 = ( n3428 & n3429 ) | ( n3428 & ~n3430 ) | ( n3429 & ~n3430 ) ;
  assign n3432 = ( x39 & n775 ) | ( x39 & n856 ) | ( n775 & n856 ) ;
  assign n3433 = n3432 ^ n1896 ^ n1547 ;
  assign n3436 = n2776 ^ n1870 ^ n805 ;
  assign n3434 = n2766 ^ x237 ^ 1'b0 ;
  assign n3435 = n360 | n3434 ;
  assign n3437 = n3436 ^ n3435 ^ n3076 ;
  assign n3438 = n3433 & ~n3437 ;
  assign n3439 = ~n3431 & n3438 ;
  assign n3440 = n603 ^ n437 ^ 1'b0 ;
  assign n3449 = ( ~n893 & n2207 ) | ( ~n893 & n2258 ) | ( n2207 & n2258 ) ;
  assign n3443 = n2732 ^ n2477 ^ 1'b0 ;
  assign n3444 = n643 & ~n884 ;
  assign n3445 = ~n820 & n3444 ;
  assign n3446 = ( n606 & n705 ) | ( n606 & n1006 ) | ( n705 & n1006 ) ;
  assign n3447 = n3445 | n3446 ;
  assign n3448 = n3443 & ~n3447 ;
  assign n3441 = n1557 ^ n1445 ^ n633 ;
  assign n3442 = n3441 ^ n3184 ^ n804 ;
  assign n3450 = n3449 ^ n3448 ^ n3442 ;
  assign n3454 = n3368 ^ n1181 ^ n520 ;
  assign n3451 = ( n296 & n434 ) | ( n296 & ~n2620 ) | ( n434 & ~n2620 ) ;
  assign n3452 = n3451 ^ n1473 ^ 1'b0 ;
  assign n3453 = n3452 ^ n1954 ^ x98 ;
  assign n3455 = n3454 ^ n3453 ^ n1039 ;
  assign n3456 = n3455 ^ n379 ^ x136 ;
  assign n3470 = ( x118 & ~n993 ) | ( x118 & n1803 ) | ( ~n993 & n1803 ) ;
  assign n3471 = ( n360 & n1898 ) | ( n360 & n3470 ) | ( n1898 & n3470 ) ;
  assign n3472 = ( n1121 & ~n3084 ) | ( n1121 & n3471 ) | ( ~n3084 & n3471 ) ;
  assign n3463 = ( ~n336 & n351 ) | ( ~n336 & n376 ) | ( n351 & n376 ) ;
  assign n3464 = n1442 ^ n629 ^ n276 ;
  assign n3465 = n3463 | n3464 ;
  assign n3466 = n2612 ^ n623 ^ 1'b0 ;
  assign n3467 = ( ~n684 & n3465 ) | ( ~n684 & n3466 ) | ( n3465 & n3466 ) ;
  assign n3460 = n1539 ^ n1496 ^ n1073 ;
  assign n3461 = n3460 ^ n700 ^ x67 ;
  assign n3462 = ( ~n1081 & n1263 ) | ( ~n1081 & n3461 ) | ( n1263 & n3461 ) ;
  assign n3468 = n3467 ^ n3462 ^ n584 ;
  assign n3457 = ( n883 & ~n1063 ) | ( n883 & n2800 ) | ( ~n1063 & n2800 ) ;
  assign n3458 = ( n1611 & ~n3272 ) | ( n1611 & n3457 ) | ( ~n3272 & n3457 ) ;
  assign n3459 = n1451 & n3458 ;
  assign n3469 = n3468 ^ n3459 ^ 1'b0 ;
  assign n3473 = n3472 ^ n3469 ^ n1990 ;
  assign n3474 = ( n816 & n1402 ) | ( n816 & n3355 ) | ( n1402 & n3355 ) ;
  assign n3475 = n3474 ^ n2128 ^ 1'b0 ;
  assign n3476 = ( n860 & ~n2136 ) | ( n860 & n3475 ) | ( ~n2136 & n3475 ) ;
  assign n3477 = n3185 ^ n2284 ^ n1547 ;
  assign n3488 = ( x7 & x50 ) | ( x7 & ~n1264 ) | ( x50 & ~n1264 ) ;
  assign n3489 = n3488 ^ n3302 ^ n742 ;
  assign n3485 = ~n1572 & n2300 ;
  assign n3486 = n3485 ^ n609 ^ 1'b0 ;
  assign n3483 = n1637 ^ n1542 ^ n1248 ;
  assign n3484 = n3483 ^ n1895 ^ n736 ;
  assign n3481 = n2382 ^ n1062 ^ x109 ;
  assign n3478 = n2293 ^ n1390 ^ n1145 ;
  assign n3479 = ( x80 & ~n2341 ) | ( x80 & n3478 ) | ( ~n2341 & n3478 ) ;
  assign n3480 = n3479 ^ n312 ^ 1'b0 ;
  assign n3482 = n3481 ^ n3480 ^ n313 ;
  assign n3487 = n3486 ^ n3484 ^ n3482 ;
  assign n3490 = n3489 ^ n3487 ^ x35 ;
  assign n3491 = ( n2012 & n3477 ) | ( n2012 & n3490 ) | ( n3477 & n3490 ) ;
  assign n3492 = n3491 ^ n1083 ^ x241 ;
  assign n3493 = n3492 ^ n1379 ^ n437 ;
  assign n3494 = n2497 ^ n739 ^ 1'b0 ;
  assign n3495 = n3494 ^ n1657 ^ n726 ;
  assign n3496 = ( ~n662 & n761 ) | ( ~n662 & n943 ) | ( n761 & n943 ) ;
  assign n3497 = ( ~n333 & n1839 ) | ( ~n333 & n2268 ) | ( n1839 & n2268 ) ;
  assign n3498 = ( n2677 & n3496 ) | ( n2677 & n3497 ) | ( n3496 & n3497 ) ;
  assign n3499 = ( n2063 & n3288 ) | ( n2063 & ~n3498 ) | ( n3288 & ~n3498 ) ;
  assign n3502 = ( x95 & ~n889 ) | ( x95 & n1365 ) | ( ~n889 & n1365 ) ;
  assign n3503 = ( ~n943 & n1300 ) | ( ~n943 & n3502 ) | ( n1300 & n3502 ) ;
  assign n3501 = ( ~n756 & n896 ) | ( ~n756 & n3222 ) | ( n896 & n3222 ) ;
  assign n3504 = n3503 ^ n3501 ^ n1235 ;
  assign n3500 = ~n427 & n2793 ;
  assign n3505 = n3504 ^ n3500 ^ 1'b0 ;
  assign n3506 = n3310 ^ n2861 ^ n2739 ;
  assign n3507 = n1513 & n1974 ;
  assign n3508 = n1245 ^ n1074 ^ n949 ;
  assign n3509 = ( n837 & n2724 ) | ( n837 & ~n3508 ) | ( n2724 & ~n3508 ) ;
  assign n3510 = x206 | n3509 ;
  assign n3518 = n2131 ^ n1102 ^ n975 ;
  assign n3519 = n3518 ^ n998 ^ n786 ;
  assign n3515 = n1952 ^ n1950 ^ n1451 ;
  assign n3516 = n3515 ^ n1181 ^ n578 ;
  assign n3513 = n2844 ^ n703 ^ x149 ;
  assign n3514 = n3513 ^ n1502 ^ x19 ;
  assign n3511 = ( n467 & n869 ) | ( n467 & ~n1800 ) | ( n869 & ~n1800 ) ;
  assign n3512 = n3511 ^ n1811 ^ n741 ;
  assign n3517 = n3516 ^ n3514 ^ n3512 ;
  assign n3520 = n3519 ^ n3517 ^ 1'b0 ;
  assign n3521 = n3520 ^ n2045 ^ n1320 ;
  assign n3522 = n799 ^ n725 ^ x27 ;
  assign n3523 = n1577 & ~n3522 ;
  assign n3524 = ( x131 & n269 ) | ( x131 & ~n769 ) | ( n269 & ~n769 ) ;
  assign n3525 = n2375 ^ n1083 ^ 1'b0 ;
  assign n3526 = ( n289 & n3524 ) | ( n289 & ~n3525 ) | ( n3524 & ~n3525 ) ;
  assign n3527 = ( n2069 & n3523 ) | ( n2069 & ~n3526 ) | ( n3523 & ~n3526 ) ;
  assign n3528 = ( n1226 & ~n2459 ) | ( n1226 & n3527 ) | ( ~n2459 & n3527 ) ;
  assign n3541 = ( n284 & n555 ) | ( n284 & n1662 ) | ( n555 & n1662 ) ;
  assign n3542 = ( ~x16 & n1793 ) | ( ~x16 & n3541 ) | ( n1793 & n3541 ) ;
  assign n3543 = ( n1013 & n3002 ) | ( n1013 & n3542 ) | ( n3002 & n3542 ) ;
  assign n3544 = ( ~x143 & n1581 ) | ( ~x143 & n3543 ) | ( n1581 & n3543 ) ;
  assign n3532 = n507 ^ n305 ^ 1'b0 ;
  assign n3534 = ( n1320 & ~n1640 ) | ( n1320 & n3034 ) | ( ~n1640 & n3034 ) ;
  assign n3533 = ( n451 & ~n568 ) | ( n451 & n2225 ) | ( ~n568 & n2225 ) ;
  assign n3535 = n3534 ^ n3533 ^ n1005 ;
  assign n3536 = n3535 ^ n688 ^ 1'b0 ;
  assign n3537 = n2943 | n3536 ;
  assign n3538 = n377 | n3537 ;
  assign n3539 = ( n887 & ~n3532 ) | ( n887 & n3538 ) | ( ~n3532 & n3538 ) ;
  assign n3529 = ~n618 & n2267 ;
  assign n3530 = n3529 ^ n1167 ^ 1'b0 ;
  assign n3531 = n3530 ^ n3296 ^ n2888 ;
  assign n3540 = n3539 ^ n3531 ^ n1744 ;
  assign n3545 = n3544 ^ n3540 ^ n906 ;
  assign n3546 = n3350 ^ n3184 ^ n1807 ;
  assign n3547 = n2195 ^ n970 ^ n687 ;
  assign n3548 = n3547 ^ n2856 ^ n2356 ;
  assign n3549 = ( x61 & n3546 ) | ( x61 & n3548 ) | ( n3546 & n3548 ) ;
  assign n3552 = n1430 ^ n898 ^ n293 ;
  assign n3553 = ( ~n431 & n802 ) | ( ~n431 & n3552 ) | ( n802 & n3552 ) ;
  assign n3550 = n2870 ^ n1775 ^ n1073 ;
  assign n3551 = n2228 & n3550 ;
  assign n3554 = n3553 ^ n3551 ^ 1'b0 ;
  assign n3555 = ( n487 & ~n1731 ) | ( n487 & n3554 ) | ( ~n1731 & n3554 ) ;
  assign n3556 = n2912 ^ n1822 ^ 1'b0 ;
  assign n3557 = ~n1116 & n3556 ;
  assign n3558 = ( x132 & n1240 ) | ( x132 & n2552 ) | ( n1240 & n2552 ) ;
  assign n3559 = n1489 ^ n1018 ^ n437 ;
  assign n3560 = ( n1157 & n1645 ) | ( n1157 & n1992 ) | ( n1645 & n1992 ) ;
  assign n3561 = ( n320 & n3559 ) | ( n320 & n3560 ) | ( n3559 & n3560 ) ;
  assign n3562 = ( n1358 & n3558 ) | ( n1358 & n3561 ) | ( n3558 & n3561 ) ;
  assign n3563 = n2209 ^ x206 ^ 1'b0 ;
  assign n3564 = ~n1105 & n3563 ;
  assign n3565 = n3564 ^ n2381 ^ n1401 ;
  assign n3566 = ( n802 & n2317 ) | ( n802 & n2956 ) | ( n2317 & n2956 ) ;
  assign n3567 = n3566 ^ n437 ^ x14 ;
  assign n3568 = ( n926 & n3565 ) | ( n926 & n3567 ) | ( n3565 & n3567 ) ;
  assign n3575 = ( x97 & n1180 ) | ( x97 & n1265 ) | ( n1180 & n1265 ) ;
  assign n3576 = ( x197 & n989 ) | ( x197 & n2306 ) | ( n989 & n2306 ) ;
  assign n3577 = ( n1031 & n1484 ) | ( n1031 & n3576 ) | ( n1484 & n3576 ) ;
  assign n3579 = ( ~n548 & n975 ) | ( ~n548 & n1129 ) | ( n975 & n1129 ) ;
  assign n3578 = n1989 ^ n600 ^ x80 ;
  assign n3580 = n3579 ^ n3578 ^ n1022 ;
  assign n3581 = ( n3575 & n3577 ) | ( n3575 & ~n3580 ) | ( n3577 & ~n3580 ) ;
  assign n3569 = n2428 ^ n1621 ^ n1581 ;
  assign n3570 = n3569 ^ n1534 ^ n814 ;
  assign n3571 = ( n1078 & ~n1875 ) | ( n1078 & n3570 ) | ( ~n1875 & n3570 ) ;
  assign n3572 = ( x251 & ~n821 ) | ( x251 & n1661 ) | ( ~n821 & n1661 ) ;
  assign n3573 = ( n1200 & n3489 ) | ( n1200 & ~n3572 ) | ( n3489 & ~n3572 ) ;
  assign n3574 = n3571 | n3573 ;
  assign n3582 = n3581 ^ n3574 ^ 1'b0 ;
  assign n3583 = x15 & ~n1519 ;
  assign n3584 = n3583 ^ n2571 ^ 1'b0 ;
  assign n3585 = ( n1754 & ~n2877 ) | ( n1754 & n3584 ) | ( ~n2877 & n3584 ) ;
  assign n3586 = n3585 ^ n3463 ^ n1593 ;
  assign n3587 = n3586 ^ n3517 ^ 1'b0 ;
  assign n3589 = ( n1540 & n2956 ) | ( n1540 & n3558 ) | ( n2956 & n3558 ) ;
  assign n3590 = n1247 | n3589 ;
  assign n3588 = n2186 ^ n541 ^ 1'b0 ;
  assign n3591 = n3590 ^ n3588 ^ n2974 ;
  assign n3594 = x80 & ~n413 ;
  assign n3595 = n3594 ^ n2979 ^ n872 ;
  assign n3596 = ( x207 & ~n1647 ) | ( x207 & n3595 ) | ( ~n1647 & n3595 ) ;
  assign n3592 = ( ~x139 & x174 ) | ( ~x139 & n755 ) | ( x174 & n755 ) ;
  assign n3593 = ( n465 & n997 ) | ( n465 & ~n3592 ) | ( n997 & ~n3592 ) ;
  assign n3597 = n3596 ^ n3593 ^ n1652 ;
  assign n3598 = n537 ^ x158 ^ x44 ;
  assign n3599 = ~n1800 & n2247 ;
  assign n3600 = n3599 ^ n1825 ^ 1'b0 ;
  assign n3601 = ( n791 & n3598 ) | ( n791 & n3600 ) | ( n3598 & n3600 ) ;
  assign n3602 = n3601 ^ n1484 ^ n1376 ;
  assign n3603 = x207 ^ x7 ^ 1'b0 ;
  assign n3604 = n1283 & n3603 ;
  assign n3605 = ( n2545 & ~n2782 ) | ( n2545 & n3604 ) | ( ~n2782 & n3604 ) ;
  assign n3606 = n1593 | n3605 ;
  assign n3607 = n3602 & ~n3606 ;
  assign n3608 = ( ~n1003 & n2893 ) | ( ~n1003 & n3092 ) | ( n2893 & n3092 ) ;
  assign n3609 = ~n696 & n1732 ;
  assign n3610 = ~x105 & n3609 ;
  assign n3620 = ( ~n517 & n1880 ) | ( ~n517 & n2826 ) | ( n1880 & n2826 ) ;
  assign n3618 = n438 & n445 ;
  assign n3616 = ( n1829 & ~n2718 ) | ( n1829 & n2853 ) | ( ~n2718 & n2853 ) ;
  assign n3617 = n3616 ^ n1529 ^ n478 ;
  assign n3619 = n3618 ^ n3617 ^ x85 ;
  assign n3611 = n2229 ^ n505 ^ 1'b0 ;
  assign n3612 = ~n1956 & n3611 ;
  assign n3613 = n3612 ^ n748 ^ n332 ;
  assign n3614 = ( ~n562 & n1075 ) | ( ~n562 & n3613 ) | ( n1075 & n3613 ) ;
  assign n3615 = n3614 ^ n2598 ^ n1410 ;
  assign n3621 = n3620 ^ n3619 ^ n3615 ;
  assign n3622 = n3621 ^ n2103 ^ n740 ;
  assign n3623 = ( x125 & n491 ) | ( x125 & ~n2720 ) | ( n491 & ~n2720 ) ;
  assign n3624 = ~n1925 & n3623 ;
  assign n3634 = ( ~n860 & n1289 ) | ( ~n860 & n2678 ) | ( n1289 & n2678 ) ;
  assign n3633 = ~n885 & n2259 ;
  assign n3635 = n3634 ^ n3633 ^ 1'b0 ;
  assign n3625 = n3445 ^ n1188 ^ n1053 ;
  assign n3626 = n1220 ^ x232 ^ 1'b0 ;
  assign n3627 = ~n383 & n3626 ;
  assign n3628 = ( ~n368 & n1208 ) | ( ~n368 & n3627 ) | ( n1208 & n3627 ) ;
  assign n3629 = n1097 & ~n1419 ;
  assign n3630 = n3628 & n3629 ;
  assign n3631 = n3625 | n3630 ;
  assign n3632 = n3631 ^ n2553 ^ n2441 ;
  assign n3636 = n3635 ^ n3632 ^ n3053 ;
  assign n3637 = n3636 ^ n313 ^ n309 ;
  assign n3639 = ( n632 & n1292 ) | ( n632 & ~n2169 ) | ( n1292 & ~n2169 ) ;
  assign n3640 = ~n665 & n3639 ;
  assign n3641 = ( n436 & n1969 ) | ( n436 & n3640 ) | ( n1969 & n3640 ) ;
  assign n3638 = ( n1005 & n1638 ) | ( n1005 & n3074 ) | ( n1638 & n3074 ) ;
  assign n3642 = n3641 ^ n3638 ^ n1488 ;
  assign n3656 = ( x193 & ~n1002 ) | ( x193 & n2703 ) | ( ~n1002 & n2703 ) ;
  assign n3657 = n3656 ^ n2255 ^ n457 ;
  assign n3658 = ( n818 & ~n1101 ) | ( n818 & n1282 ) | ( ~n1101 & n1282 ) ;
  assign n3659 = n3658 ^ n1565 ^ n1380 ;
  assign n3660 = n3659 ^ n938 ^ 1'b0 ;
  assign n3661 = n2911 & ~n3660 ;
  assign n3662 = n3657 & n3661 ;
  assign n3663 = n3662 ^ n2659 ^ 1'b0 ;
  assign n3664 = n3663 ^ n2130 ^ n1899 ;
  assign n3650 = ( n2140 & n2160 ) | ( n2140 & n2299 ) | ( n2160 & n2299 ) ;
  assign n3651 = n3650 ^ n2800 ^ n2168 ;
  assign n3649 = ~n1762 & n2705 ;
  assign n3652 = n3651 ^ n3649 ^ n2243 ;
  assign n3653 = n3652 ^ n1848 ^ n533 ;
  assign n3643 = ( n619 & n747 ) | ( n619 & ~n1414 ) | ( n747 & ~n1414 ) ;
  assign n3644 = ~n2317 & n3643 ;
  assign n3645 = n548 & n3644 ;
  assign n3646 = ( ~n2870 & n3559 ) | ( ~n2870 & n3645 ) | ( n3559 & n3645 ) ;
  assign n3647 = n3598 | n3646 ;
  assign n3648 = n297 | n3647 ;
  assign n3654 = n3653 ^ n3648 ^ n3202 ;
  assign n3655 = ( n2413 & n3076 ) | ( n2413 & ~n3654 ) | ( n3076 & ~n3654 ) ;
  assign n3665 = n3664 ^ n3655 ^ 1'b0 ;
  assign n3666 = n3487 ^ n2110 ^ 1'b0 ;
  assign n3667 = n2093 ^ n1025 ^ 1'b0 ;
  assign n3668 = n3667 ^ n1061 ^ n987 ;
  assign n3669 = n580 ^ x59 ^ 1'b0 ;
  assign n3670 = ( n1761 & n1802 ) | ( n1761 & ~n3669 ) | ( n1802 & ~n3669 ) ;
  assign n3671 = ( ~n2114 & n3285 ) | ( ~n2114 & n3670 ) | ( n3285 & n3670 ) ;
  assign n3672 = ( n560 & n2033 ) | ( n560 & n3331 ) | ( n2033 & n3331 ) ;
  assign n3673 = ( n3668 & ~n3671 ) | ( n3668 & n3672 ) | ( ~n3671 & n3672 ) ;
  assign n3674 = ( n1393 & n2001 ) | ( n1393 & ~n2282 ) | ( n2001 & ~n2282 ) ;
  assign n3675 = ( n501 & n3673 ) | ( n501 & n3674 ) | ( n3673 & n3674 ) ;
  assign n3677 = n701 ^ x117 ^ 1'b0 ;
  assign n3678 = n1902 | n3677 ;
  assign n3679 = n3678 ^ n3429 ^ 1'b0 ;
  assign n3676 = n2033 ^ n786 ^ n457 ;
  assign n3680 = n3679 ^ n3676 ^ n740 ;
  assign n3681 = ( n3666 & ~n3675 ) | ( n3666 & n3680 ) | ( ~n3675 & n3680 ) ;
  assign n3682 = n3519 ^ n2295 ^ 1'b0 ;
  assign n3683 = ( n1764 & n3325 ) | ( n1764 & n3682 ) | ( n3325 & n3682 ) ;
  assign n3684 = n967 | n3230 ;
  assign n3685 = x180 | n3684 ;
  assign n3686 = n2310 ^ n1473 ^ n334 ;
  assign n3687 = ( x189 & ~n2471 ) | ( x189 & n3686 ) | ( ~n2471 & n3686 ) ;
  assign n3688 = ( x176 & n3685 ) | ( x176 & n3687 ) | ( n3685 & n3687 ) ;
  assign n3689 = ~n3516 & n3688 ;
  assign n3690 = n3689 ^ n3164 ^ n2477 ;
  assign n3736 = n1058 ^ n1016 ^ n442 ;
  assign n3734 = ( n759 & n1660 ) | ( n759 & n2375 ) | ( n1660 & n2375 ) ;
  assign n3735 = n3734 ^ n1220 ^ x15 ;
  assign n3726 = n744 ^ n363 ^ x10 ;
  assign n3727 = n2338 ^ n1079 ^ x115 ;
  assign n3728 = ( n361 & n791 ) | ( n361 & ~n1152 ) | ( n791 & ~n1152 ) ;
  assign n3729 = n3728 ^ x169 ^ x92 ;
  assign n3730 = n3729 ^ n1479 ^ n1116 ;
  assign n3731 = n3730 ^ n2755 ^ n1495 ;
  assign n3732 = ( ~n1189 & n3727 ) | ( ~n1189 & n3731 ) | ( n3727 & n3731 ) ;
  assign n3733 = ( n1653 & n3726 ) | ( n1653 & ~n3732 ) | ( n3726 & ~n3732 ) ;
  assign n3737 = n3736 ^ n3735 ^ n3733 ;
  assign n3718 = ( x197 & n925 ) | ( x197 & ~n2143 ) | ( n925 & ~n2143 ) ;
  assign n3719 = n3718 ^ n715 ^ n517 ;
  assign n3720 = ( n518 & ~n980 ) | ( n518 & n1947 ) | ( ~n980 & n1947 ) ;
  assign n3721 = ( n1200 & n1589 ) | ( n1200 & n2277 ) | ( n1589 & n2277 ) ;
  assign n3722 = n2766 | n3721 ;
  assign n3723 = n3720 & ~n3722 ;
  assign n3724 = ( n1363 & n3719 ) | ( n1363 & ~n3723 ) | ( n3719 & ~n3723 ) ;
  assign n3715 = n520 ^ n310 ^ n291 ;
  assign n3716 = n3715 ^ n624 ^ x195 ;
  assign n3713 = ( x215 & n718 ) | ( x215 & ~n1283 ) | ( n718 & ~n1283 ) ;
  assign n3714 = ( ~x147 & n2210 ) | ( ~x147 & n3713 ) | ( n2210 & n3713 ) ;
  assign n3703 = n471 ^ n345 ^ x109 ;
  assign n3704 = n3703 ^ n1154 ^ 1'b0 ;
  assign n3705 = n1928 | n3704 ;
  assign n3706 = n3705 ^ n1176 ^ n1093 ;
  assign n3707 = n863 | n1634 ;
  assign n3708 = n1931 & ~n3707 ;
  assign n3709 = ( n1398 & n3706 ) | ( n1398 & n3708 ) | ( n3706 & n3708 ) ;
  assign n3710 = n2956 ^ n2548 ^ n1149 ;
  assign n3711 = n3710 ^ n3052 ^ 1'b0 ;
  assign n3712 = ( n2733 & ~n3709 ) | ( n2733 & n3711 ) | ( ~n3709 & n3711 ) ;
  assign n3717 = n3716 ^ n3714 ^ n3712 ;
  assign n3693 = n2138 ^ n1289 ^ n1024 ;
  assign n3694 = ( n417 & n1772 ) | ( n417 & n3693 ) | ( n1772 & n3693 ) ;
  assign n3695 = n1069 ^ n895 ^ n781 ;
  assign n3696 = n3695 ^ n3417 ^ n2689 ;
  assign n3697 = ( n729 & n828 ) | ( n729 & ~n882 ) | ( n828 & ~n882 ) ;
  assign n3698 = ( x244 & n1807 ) | ( x244 & n3630 ) | ( n1807 & n3630 ) ;
  assign n3699 = ( n3269 & n3697 ) | ( n3269 & ~n3698 ) | ( n3697 & ~n3698 ) ;
  assign n3700 = ( ~n1549 & n3696 ) | ( ~n1549 & n3699 ) | ( n3696 & n3699 ) ;
  assign n3701 = n3700 ^ n2786 ^ n2687 ;
  assign n3702 = ( n2766 & ~n3694 ) | ( n2766 & n3701 ) | ( ~n3694 & n3701 ) ;
  assign n3725 = n3724 ^ n3717 ^ n3702 ;
  assign n3691 = n1960 ^ n1143 ^ x104 ;
  assign n3692 = n3691 ^ n3039 ^ n2429 ;
  assign n3738 = n3737 ^ n3725 ^ n3692 ;
  assign n3739 = ( n1540 & ~n2885 ) | ( n1540 & n3533 ) | ( ~n2885 & n3533 ) ;
  assign n3740 = n3739 ^ n1598 ^ n1142 ;
  assign n3741 = n3740 ^ n1152 ^ n659 ;
  assign n3780 = n2011 ^ n1402 ^ n1370 ;
  assign n3781 = ( n1165 & n1427 ) | ( n1165 & n3780 ) | ( n1427 & n3780 ) ;
  assign n3782 = n3781 ^ n636 ^ x142 ;
  assign n3775 = x245 & n1771 ;
  assign n3776 = n3775 ^ x85 ^ 1'b0 ;
  assign n3777 = n3776 ^ n3576 ^ n1667 ;
  assign n3778 = x161 & n3777 ;
  assign n3779 = n1336 & n3778 ;
  assign n3783 = n3782 ^ n3779 ^ n3661 ;
  assign n3742 = n3716 ^ n3317 ^ n1911 ;
  assign n3743 = ( n650 & ~n1259 ) | ( n650 & n1587 ) | ( ~n1259 & n1587 ) ;
  assign n3744 = ( n529 & ~n2228 ) | ( n529 & n3743 ) | ( ~n2228 & n3743 ) ;
  assign n3745 = n1060 & n3744 ;
  assign n3746 = n3745 ^ n2006 ^ 1'b0 ;
  assign n3747 = n772 & n3490 ;
  assign n3748 = n3746 & n3747 ;
  assign n3749 = n2382 ^ n1349 ^ x68 ;
  assign n3750 = ( n589 & n885 ) | ( n589 & n3749 ) | ( n885 & n3749 ) ;
  assign n3751 = ( ~n786 & n884 ) | ( ~n786 & n1458 ) | ( n884 & n1458 ) ;
  assign n3752 = n2318 ^ n717 ^ n448 ;
  assign n3753 = ( n2594 & n3751 ) | ( n2594 & n3752 ) | ( n3751 & n3752 ) ;
  assign n3754 = n3753 ^ n3212 ^ 1'b0 ;
  assign n3755 = n1980 & ~n3754 ;
  assign n3756 = n2506 ^ n1105 ^ 1'b0 ;
  assign n3757 = n3756 ^ n1296 ^ 1'b0 ;
  assign n3759 = n866 & n1345 ;
  assign n3758 = n2949 ^ n2403 ^ n2186 ;
  assign n3760 = n3759 ^ n3758 ^ n2424 ;
  assign n3761 = ( n3630 & n3757 ) | ( n3630 & ~n3760 ) | ( n3757 & ~n3760 ) ;
  assign n3762 = ( n3750 & n3755 ) | ( n3750 & n3761 ) | ( n3755 & n3761 ) ;
  assign n3763 = ( ~n1112 & n3748 ) | ( ~n1112 & n3762 ) | ( n3748 & n3762 ) ;
  assign n3764 = ( n3352 & n3742 ) | ( n3352 & n3763 ) | ( n3742 & n3763 ) ;
  assign n3765 = n3764 ^ x66 ^ x17 ;
  assign n3769 = x80 & x120 ;
  assign n3770 = n3769 ^ x176 ^ 1'b0 ;
  assign n3771 = n3770 ^ n962 ^ n713 ;
  assign n3772 = ( ~n2378 & n3480 ) | ( ~n2378 & n3771 ) | ( n3480 & n3771 ) ;
  assign n3766 = x168 & n2246 ;
  assign n3767 = ( n2113 & n3268 ) | ( n2113 & n3766 ) | ( n3268 & n3766 ) ;
  assign n3768 = ( ~n2485 & n3250 ) | ( ~n2485 & n3767 ) | ( n3250 & n3767 ) ;
  assign n3773 = n3772 ^ n3768 ^ n3615 ;
  assign n3774 = n3765 & ~n3773 ;
  assign n3784 = n3783 ^ n3774 ^ 1'b0 ;
  assign n3785 = n3594 ^ n1123 ^ x42 ;
  assign n3786 = n3785 ^ n3234 ^ n725 ;
  assign n3787 = n3786 ^ n1125 ^ 1'b0 ;
  assign n3797 = ( n287 & n1422 ) | ( n287 & ~n1666 ) | ( n1422 & ~n1666 ) ;
  assign n3796 = ( ~x145 & n1748 ) | ( ~x145 & n2393 ) | ( n1748 & n2393 ) ;
  assign n3794 = n2280 ^ n1990 ^ n1347 ;
  assign n3795 = n3794 ^ n938 ^ x183 ;
  assign n3798 = n3797 ^ n3796 ^ n3795 ;
  assign n3789 = n875 ^ n555 ^ n434 ;
  assign n3788 = ( x63 & n653 ) | ( x63 & n1838 ) | ( n653 & n1838 ) ;
  assign n3790 = n3789 ^ n3788 ^ 1'b0 ;
  assign n3791 = n3790 ^ n3376 ^ n365 ;
  assign n3792 = ( n673 & n1399 ) | ( n673 & n1698 ) | ( n1399 & n1698 ) ;
  assign n3793 = n3791 & ~n3792 ;
  assign n3799 = n3798 ^ n3793 ^ n1650 ;
  assign n3800 = ( n1459 & n2953 ) | ( n1459 & ~n3799 ) | ( n2953 & ~n3799 ) ;
  assign n3807 = n1802 ^ n1478 ^ x194 ;
  assign n3804 = n2293 ^ n872 ^ n404 ;
  assign n3803 = n1505 | n3732 ;
  assign n3805 = n3804 ^ n3803 ^ n824 ;
  assign n3801 = ( n1010 & n1012 ) | ( n1010 & ~n2299 ) | ( n1012 & ~n2299 ) ;
  assign n3802 = n3801 ^ n3109 ^ n2637 ;
  assign n3806 = n3805 ^ n3802 ^ n819 ;
  assign n3808 = n3807 ^ n3806 ^ n522 ;
  assign n3819 = n1485 ^ n1218 ^ n337 ;
  assign n3822 = n2760 ^ n467 ^ x164 ;
  assign n3820 = ( n1261 & n1909 ) | ( n1261 & ~n2781 ) | ( n1909 & ~n2781 ) ;
  assign n3821 = n2692 | n3820 ;
  assign n3823 = n3822 ^ n3821 ^ 1'b0 ;
  assign n3824 = ~n3350 & n3823 ;
  assign n3825 = n3824 ^ n2693 ^ 1'b0 ;
  assign n3826 = ( n1840 & n3819 ) | ( n1840 & n3825 ) | ( n3819 & n3825 ) ;
  assign n3815 = ( ~n1207 & n1214 ) | ( ~n1207 & n1296 ) | ( n1214 & n1296 ) ;
  assign n3816 = n1774 & ~n3815 ;
  assign n3817 = n3816 ^ n3657 ^ 1'b0 ;
  assign n3818 = n1102 & ~n3817 ;
  assign n3809 = ( ~n977 & n989 ) | ( ~n977 & n2969 ) | ( n989 & n2969 ) ;
  assign n3810 = n1193 ^ n1192 ^ n743 ;
  assign n3811 = ( ~n921 & n3008 ) | ( ~n921 & n3810 ) | ( n3008 & n3810 ) ;
  assign n3812 = ( n1537 & n3002 ) | ( n1537 & ~n3811 ) | ( n3002 & ~n3811 ) ;
  assign n3813 = ( x204 & ~n1035 ) | ( x204 & n3054 ) | ( ~n1035 & n3054 ) ;
  assign n3814 = ( ~n3809 & n3812 ) | ( ~n3809 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3827 = n3826 ^ n3818 ^ n3814 ;
  assign n3832 = ( n2119 & n2491 ) | ( n2119 & ~n3382 ) | ( n2491 & ~n3382 ) ;
  assign n3828 = ~n269 & n1542 ;
  assign n3829 = n3828 ^ n3228 ^ n1565 ;
  assign n3830 = n2728 ^ n2311 ^ n1030 ;
  assign n3831 = ( x66 & ~n3829 ) | ( x66 & n3830 ) | ( ~n3829 & n3830 ) ;
  assign n3833 = n3832 ^ n3831 ^ n1447 ;
  assign n3834 = n3294 ^ n2042 ^ n1209 ;
  assign n3835 = n2317 ^ n1002 ^ n364 ;
  assign n3836 = ( n2478 & n3183 ) | ( n2478 & ~n3835 ) | ( n3183 & ~n3835 ) ;
  assign n3837 = ( n1544 & ~n3834 ) | ( n1544 & n3836 ) | ( ~n3834 & n3836 ) ;
  assign n3841 = ( ~n538 & n806 ) | ( ~n538 & n1969 ) | ( n806 & n1969 ) ;
  assign n3838 = ( n336 & n2647 ) | ( n336 & ~n2889 ) | ( n2647 & ~n2889 ) ;
  assign n3839 = n624 & n2551 ;
  assign n3840 = ~n3838 & n3839 ;
  assign n3842 = n3841 ^ n3840 ^ n580 ;
  assign n3843 = ( n862 & n1974 ) | ( n862 & ~n3842 ) | ( n1974 & ~n3842 ) ;
  assign n3844 = ( n1132 & n1334 ) | ( n1132 & n3843 ) | ( n1334 & n3843 ) ;
  assign n3845 = ( n1443 & ~n3837 ) | ( n1443 & n3844 ) | ( ~n3837 & n3844 ) ;
  assign n3846 = ( x122 & ~n894 ) | ( x122 & n2041 ) | ( ~n894 & n2041 ) ;
  assign n3847 = ( x171 & n1868 ) | ( x171 & ~n2674 ) | ( n1868 & ~n2674 ) ;
  assign n3850 = n1578 ^ n979 ^ n857 ;
  assign n3852 = ( n384 & n541 ) | ( n384 & ~n866 ) | ( n541 & ~n866 ) ;
  assign n3851 = ( x11 & ~n288 ) | ( x11 & n1094 ) | ( ~n288 & n1094 ) ;
  assign n3853 = n3852 ^ n3851 ^ n3156 ;
  assign n3854 = ( n2340 & ~n3850 ) | ( n2340 & n3853 ) | ( ~n3850 & n3853 ) ;
  assign n3849 = ( n287 & n806 ) | ( n287 & ~n2398 ) | ( n806 & ~n2398 ) ;
  assign n3848 = n2768 ^ n1551 ^ 1'b0 ;
  assign n3855 = n3854 ^ n3849 ^ n3848 ;
  assign n3856 = ( x127 & n1272 ) | ( x127 & ~n1381 ) | ( n1272 & ~n1381 ) ;
  assign n3857 = n365 & ~n2519 ;
  assign n3858 = ( x31 & n393 ) | ( x31 & n3857 ) | ( n393 & n3857 ) ;
  assign n3859 = n3858 ^ n1160 ^ n1057 ;
  assign n3860 = ( n2175 & n3856 ) | ( n2175 & ~n3859 ) | ( n3856 & ~n3859 ) ;
  assign n3866 = n1503 ^ n1338 ^ n818 ;
  assign n3862 = ( n584 & ~n1141 ) | ( n584 & n1816 ) | ( ~n1141 & n1816 ) ;
  assign n3863 = ( n1764 & ~n2602 ) | ( n1764 & n3862 ) | ( ~n2602 & n3862 ) ;
  assign n3864 = n3863 ^ n767 ^ x57 ;
  assign n3861 = ( ~n750 & n2193 ) | ( ~n750 & n3553 ) | ( n2193 & n3553 ) ;
  assign n3865 = n3864 ^ n3861 ^ n3729 ;
  assign n3867 = n3866 ^ n3865 ^ n3483 ;
  assign n3868 = ( ~n1262 & n3036 ) | ( ~n1262 & n3480 ) | ( n3036 & n3480 ) ;
  assign n3869 = ( n587 & n752 ) | ( n587 & n1814 ) | ( n752 & n1814 ) ;
  assign n3870 = ( ~x159 & n1606 ) | ( ~x159 & n1612 ) | ( n1606 & n1612 ) ;
  assign n3871 = ( n2545 & n3869 ) | ( n2545 & n3870 ) | ( n3869 & n3870 ) ;
  assign n3872 = ( n1132 & ~n1812 ) | ( n1132 & n3871 ) | ( ~n1812 & n3871 ) ;
  assign n3873 = n3872 ^ n1482 ^ n1183 ;
  assign n3876 = n2775 ^ n1955 ^ 1'b0 ;
  assign n3877 = n593 & n3876 ;
  assign n3874 = ( n364 & ~n739 ) | ( n364 & n1823 ) | ( ~n739 & n1823 ) ;
  assign n3875 = ~n3577 & n3874 ;
  assign n3878 = n3877 ^ n3875 ^ 1'b0 ;
  assign n3879 = ( ~n871 & n1213 ) | ( ~n871 & n3878 ) | ( n1213 & n3878 ) ;
  assign n3880 = ( ~x252 & n2279 ) | ( ~x252 & n3879 ) | ( n2279 & n3879 ) ;
  assign n3881 = ( n478 & ~n1899 ) | ( n478 & n3880 ) | ( ~n1899 & n3880 ) ;
  assign n3882 = n3881 ^ n2225 ^ 1'b0 ;
  assign n3883 = n3194 | n3882 ;
  assign n3884 = n1633 ^ n1142 ^ 1'b0 ;
  assign n3885 = x140 & n3884 ;
  assign n3886 = ( n827 & n872 ) | ( n827 & ~n3885 ) | ( n872 & ~n3885 ) ;
  assign n3887 = n1348 ^ n989 ^ n970 ;
  assign n3888 = ( x61 & n1086 ) | ( x61 & ~n3887 ) | ( n1086 & ~n3887 ) ;
  assign n3889 = ( n834 & n3012 ) | ( n834 & ~n3888 ) | ( n3012 & ~n3888 ) ;
  assign n3890 = ( n1115 & n3886 ) | ( n1115 & ~n3889 ) | ( n3886 & ~n3889 ) ;
  assign n3897 = ( ~n866 & n1367 ) | ( ~n866 & n1901 ) | ( n1367 & n1901 ) ;
  assign n3892 = ( n645 & ~n1319 ) | ( n645 & n1739 ) | ( ~n1319 & n1739 ) ;
  assign n3893 = n3892 ^ n1248 ^ x121 ;
  assign n3891 = n1332 ^ n1059 ^ x14 ;
  assign n3894 = n3893 ^ n3891 ^ n418 ;
  assign n3895 = n3894 ^ n2888 ^ n1236 ;
  assign n3896 = ( n1463 & n3066 ) | ( n1463 & ~n3895 ) | ( n3066 & ~n3895 ) ;
  assign n3898 = n3897 ^ n3896 ^ n943 ;
  assign n3899 = ( n883 & n927 ) | ( n883 & ~n2286 ) | ( n927 & ~n2286 ) ;
  assign n3900 = x192 ^ x132 ^ x73 ;
  assign n3901 = ( x1 & n1589 ) | ( x1 & ~n3900 ) | ( n1589 & ~n3900 ) ;
  assign n3902 = ( n2179 & n2595 ) | ( n2179 & ~n3525 ) | ( n2595 & ~n3525 ) ;
  assign n3903 = ( n2750 & n3901 ) | ( n2750 & n3902 ) | ( n3901 & n3902 ) ;
  assign n3904 = ( ~n396 & n415 ) | ( ~n396 & n1105 ) | ( n415 & n1105 ) ;
  assign n3905 = n3904 ^ n1690 ^ n277 ;
  assign n3906 = ( n3899 & ~n3903 ) | ( n3899 & n3905 ) | ( ~n3903 & n3905 ) ;
  assign n3907 = n914 ^ n661 ^ n599 ;
  assign n3908 = n3907 ^ n1796 ^ x209 ;
  assign n3914 = ( x188 & ~n1825 ) | ( x188 & n3864 ) | ( ~n1825 & n3864 ) ;
  assign n3909 = n310 & n1652 ;
  assign n3910 = ~n818 & n3909 ;
  assign n3911 = n3910 ^ n1521 ^ n1006 ;
  assign n3912 = ( x249 & ~n430 ) | ( x249 & n3911 ) | ( ~n430 & n3911 ) ;
  assign n3913 = n1821 & n3912 ;
  assign n3915 = n3914 ^ n3913 ^ 1'b0 ;
  assign n3916 = ( n2056 & n3908 ) | ( n2056 & ~n3915 ) | ( n3908 & ~n3915 ) ;
  assign n3917 = ( n423 & n1218 ) | ( n423 & ~n1904 ) | ( n1218 & ~n1904 ) ;
  assign n3918 = x162 & ~n2082 ;
  assign n3919 = n3918 ^ n1134 ^ 1'b0 ;
  assign n3920 = ( n550 & ~n557 ) | ( n550 & n610 ) | ( ~n557 & n610 ) ;
  assign n3921 = ( n725 & n3919 ) | ( n725 & ~n3920 ) | ( n3919 & ~n3920 ) ;
  assign n3922 = x43 & n3921 ;
  assign n3923 = n3917 | n3922 ;
  assign n3924 = ( n2062 & ~n2942 ) | ( n2062 & n3923 ) | ( ~n2942 & n3923 ) ;
  assign n3925 = n3924 ^ n3008 ^ n2169 ;
  assign n3926 = ( n1977 & n2843 ) | ( n1977 & n3925 ) | ( n2843 & n3925 ) ;
  assign n3927 = n327 & ~n3443 ;
  assign n3928 = n2964 ^ n2697 ^ n600 ;
  assign n3929 = ( ~n274 & n3927 ) | ( ~n274 & n3928 ) | ( n3927 & n3928 ) ;
  assign n3930 = n3656 ^ n1786 ^ n1550 ;
  assign n3931 = n2202 ^ n2147 ^ 1'b0 ;
  assign n3932 = ~n3003 & n3931 ;
  assign n3933 = ( x134 & ~n1467 ) | ( x134 & n2099 ) | ( ~n1467 & n2099 ) ;
  assign n3934 = ( n1256 & n3932 ) | ( n1256 & ~n3933 ) | ( n3932 & ~n3933 ) ;
  assign n3935 = n3934 ^ n3879 ^ n1398 ;
  assign n3936 = n3935 ^ n3130 ^ 1'b0 ;
  assign n3937 = n3930 & n3936 ;
  assign n3938 = n2021 ^ x93 ^ 1'b0 ;
  assign n3939 = n3938 ^ n3123 ^ n1724 ;
  assign n3965 = ( n1800 & ~n2741 ) | ( n1800 & n3396 ) | ( ~n2741 & n3396 ) ;
  assign n3962 = n1513 ^ x127 ^ 1'b0 ;
  assign n3960 = ( n261 & n1072 ) | ( n261 & n1382 ) | ( n1072 & n1382 ) ;
  assign n3961 = n1975 & n3960 ;
  assign n3963 = n3962 ^ n3961 ^ 1'b0 ;
  assign n3964 = n3963 ^ n2775 ^ n2022 ;
  assign n3955 = n863 ^ x72 ^ 1'b0 ;
  assign n3956 = x77 & ~n3955 ;
  assign n3950 = ( x136 & x224 ) | ( x136 & ~n2411 ) | ( x224 & ~n2411 ) ;
  assign n3951 = n3110 ^ n2781 ^ n1189 ;
  assign n3952 = n3950 & n3951 ;
  assign n3953 = n3286 ^ n662 ^ 1'b0 ;
  assign n3954 = ~n3952 & n3953 ;
  assign n3949 = ( ~x141 & n2396 ) | ( ~x141 & n3795 ) | ( n2396 & n3795 ) ;
  assign n3957 = n3956 ^ n3954 ^ n3949 ;
  assign n3947 = ( ~n821 & n945 ) | ( ~n821 & n1467 ) | ( n945 & n1467 ) ;
  assign n3948 = ( n2510 & ~n3287 ) | ( n2510 & n3947 ) | ( ~n3287 & n3947 ) ;
  assign n3958 = n3957 ^ n3948 ^ n2336 ;
  assign n3943 = ( x239 & n1405 ) | ( x239 & n1619 ) | ( n1405 & n1619 ) ;
  assign n3940 = n1230 | n1770 ;
  assign n3941 = n3940 ^ n597 ^ 1'b0 ;
  assign n3942 = n3941 ^ n702 ^ x54 ;
  assign n3944 = n3943 ^ n3942 ^ n601 ;
  assign n3945 = ( ~n351 & n1411 ) | ( ~n351 & n3138 ) | ( n1411 & n3138 ) ;
  assign n3946 = n3944 & ~n3945 ;
  assign n3959 = n3958 ^ n3946 ^ 1'b0 ;
  assign n3966 = n3965 ^ n3964 ^ n3959 ;
  assign n3974 = ( n929 & n1379 ) | ( n929 & n2084 ) | ( n1379 & n2084 ) ;
  assign n3975 = n3974 ^ n2736 ^ n1077 ;
  assign n3976 = ( n620 & ~n734 ) | ( n620 & n1408 ) | ( ~n734 & n1408 ) ;
  assign n3977 = ( n1108 & ~n2703 ) | ( n1108 & n3976 ) | ( ~n2703 & n3976 ) ;
  assign n3978 = n1828 ^ n1171 ^ 1'b0 ;
  assign n3979 = n1660 | n3978 ;
  assign n3980 = ( n283 & n973 ) | ( n283 & ~n2186 ) | ( n973 & ~n2186 ) ;
  assign n3981 = ( n3977 & ~n3979 ) | ( n3977 & n3980 ) | ( ~n3979 & n3980 ) ;
  assign n3982 = ( n1602 & n3975 ) | ( n1602 & ~n3981 ) | ( n3975 & ~n3981 ) ;
  assign n3967 = x153 & ~n1481 ;
  assign n3968 = ~x133 & n3967 ;
  assign n3969 = n1993 ^ n722 ^ x175 ;
  assign n3970 = n1362 & ~n3969 ;
  assign n3971 = n3968 & n3970 ;
  assign n3972 = ( ~n264 & n419 ) | ( ~n264 & n2890 ) | ( n419 & n2890 ) ;
  assign n3973 = n3971 | n3972 ;
  assign n3983 = n3982 ^ n3973 ^ 1'b0 ;
  assign n3984 = n1266 ^ n931 ^ x216 ;
  assign n3985 = n1286 ^ n1028 ^ 1'b0 ;
  assign n3986 = n3984 & n3985 ;
  assign n3987 = ( x183 & n755 ) | ( x183 & ~n3986 ) | ( n755 & ~n3986 ) ;
  assign n3991 = n2796 ^ n1505 ^ x201 ;
  assign n3992 = n3991 ^ n658 ^ x33 ;
  assign n3993 = n823 | n3992 ;
  assign n3994 = n269 & ~n3993 ;
  assign n3995 = n1063 & n3994 ;
  assign n3988 = n2038 ^ n1519 ^ n1109 ;
  assign n3989 = n3988 ^ n2730 ^ n1440 ;
  assign n3990 = ( ~n1556 & n1930 ) | ( ~n1556 & n3989 ) | ( n1930 & n3989 ) ;
  assign n3996 = n3995 ^ n3990 ^ n3554 ;
  assign n3997 = ( x98 & n1323 ) | ( x98 & n3252 ) | ( n1323 & n3252 ) ;
  assign n3998 = ( n1895 & ~n2335 ) | ( n1895 & n3997 ) | ( ~n2335 & n3997 ) ;
  assign n3999 = n3406 ^ n1738 ^ n369 ;
  assign n4000 = ( n2171 & n3998 ) | ( n2171 & n3999 ) | ( n3998 & n3999 ) ;
  assign n4001 = n3346 ^ n2143 ^ x78 ;
  assign n4002 = n4001 ^ n2831 ^ n451 ;
  assign n4003 = n3152 & n4002 ;
  assign n4004 = n1868 ^ n1573 ^ 1'b0 ;
  assign n4005 = n2114 & ~n4004 ;
  assign n4006 = ~n1585 & n4005 ;
  assign n4007 = ~n4003 & n4006 ;
  assign n4008 = ( n2625 & n3065 ) | ( n2625 & ~n4007 ) | ( n3065 & ~n4007 ) ;
  assign n4019 = n3141 ^ n2011 ^ n1266 ;
  assign n4017 = n1931 | n2761 ;
  assign n4018 = n1082 | n4017 ;
  assign n4009 = n2069 ^ n1895 ^ n1106 ;
  assign n4010 = ( ~x138 & n2206 ) | ( ~x138 & n3092 ) | ( n2206 & n3092 ) ;
  assign n4011 = ( x230 & ~n873 ) | ( x230 & n1478 ) | ( ~n873 & n1478 ) ;
  assign n4012 = ( n265 & n468 ) | ( n265 & ~n4011 ) | ( n468 & ~n4011 ) ;
  assign n4013 = ( n278 & ~n1012 ) | ( n278 & n1026 ) | ( ~n1012 & n1026 ) ;
  assign n4014 = n4012 | n4013 ;
  assign n4015 = n4010 | n4014 ;
  assign n4016 = ( ~n635 & n4009 ) | ( ~n635 & n4015 ) | ( n4009 & n4015 ) ;
  assign n4020 = n4019 ^ n4018 ^ n4016 ;
  assign n4021 = n4020 ^ n2429 ^ n1838 ;
  assign n4022 = ( x135 & n924 ) | ( x135 & n3950 ) | ( n924 & n3950 ) ;
  assign n4023 = n4022 ^ n2094 ^ n1271 ;
  assign n4024 = ( x118 & ~n281 ) | ( x118 & n462 ) | ( ~n281 & n462 ) ;
  assign n4025 = n4024 ^ n1676 ^ n1428 ;
  assign n4026 = n1917 & n1935 ;
  assign n4027 = n4025 & n4026 ;
  assign n4028 = ( x140 & n4023 ) | ( x140 & ~n4027 ) | ( n4023 & ~n4027 ) ;
  assign n4030 = n2452 & ~n3659 ;
  assign n4031 = n4030 ^ x165 ^ 1'b0 ;
  assign n4029 = n2002 ^ n420 ^ n290 ;
  assign n4032 = n4031 ^ n4029 ^ n671 ;
  assign n4033 = ( ~n1006 & n1627 ) | ( ~n1006 & n4032 ) | ( n1627 & n4032 ) ;
  assign n4034 = ( ~n2345 & n2594 ) | ( ~n2345 & n3616 ) | ( n2594 & n3616 ) ;
  assign n4040 = n3600 ^ n379 ^ x63 ;
  assign n4035 = n3564 ^ n827 ^ 1'b0 ;
  assign n4036 = n1120 & n4035 ;
  assign n4037 = n4036 ^ n3986 ^ n403 ;
  assign n4038 = ( ~n575 & n1937 ) | ( ~n575 & n4037 ) | ( n1937 & n4037 ) ;
  assign n4039 = n4038 ^ n1551 ^ 1'b0 ;
  assign n4041 = n4040 ^ n4039 ^ x213 ;
  assign n4042 = n3002 ^ n1473 ^ n781 ;
  assign n4043 = n3576 ^ n1072 ^ 1'b0 ;
  assign n4044 = n4042 & ~n4043 ;
  assign n4045 = ~n4041 & n4044 ;
  assign n4046 = n2510 | n4045 ;
  assign n4047 = n4034 | n4046 ;
  assign n4074 = n1953 ^ n1049 ^ n752 ;
  assign n4075 = ( ~n2002 & n2580 ) | ( ~n2002 & n4074 ) | ( n2580 & n4074 ) ;
  assign n4076 = n1505 & ~n3785 ;
  assign n4077 = ~n4075 & n4076 ;
  assign n4072 = ~n2886 & n3008 ;
  assign n4069 = ( ~x47 & n1260 ) | ( ~x47 & n2850 ) | ( n1260 & n2850 ) ;
  assign n4070 = ( n411 & n1374 ) | ( n411 & ~n4069 ) | ( n1374 & ~n4069 ) ;
  assign n4071 = n4070 ^ n2662 ^ n1818 ;
  assign n4073 = n4072 ^ n4071 ^ n3174 ;
  assign n4049 = ( ~n1030 & n1113 ) | ( ~n1030 & n3230 ) | ( n1113 & n3230 ) ;
  assign n4050 = n4049 ^ n3002 ^ x190 ;
  assign n4051 = n4050 ^ n3405 ^ n533 ;
  assign n4048 = n3653 ^ n3352 ^ n1862 ;
  assign n4052 = n4051 ^ n4048 ^ n1275 ;
  assign n4056 = n1595 ^ n309 ^ 1'b0 ;
  assign n4054 = n2383 ^ n1121 ^ n608 ;
  assign n4053 = n3669 ^ n2479 ^ n860 ;
  assign n4055 = n4054 ^ n4053 ^ n618 ;
  assign n4057 = n4056 ^ n4055 ^ 1'b0 ;
  assign n4058 = ( n975 & ~n1476 ) | ( n975 & n3677 ) | ( ~n1476 & n3677 ) ;
  assign n4059 = n1684 & n4058 ;
  assign n4060 = ~n578 & n4059 ;
  assign n4061 = n4060 ^ n3340 ^ n1075 ;
  assign n4062 = n4057 & ~n4061 ;
  assign n4063 = n4062 ^ n1059 ^ 1'b0 ;
  assign n4064 = n1937 ^ n652 ^ n464 ;
  assign n4065 = ( n1057 & ~n1930 ) | ( n1057 & n3596 ) | ( ~n1930 & n3596 ) ;
  assign n4066 = n4065 ^ n1416 ^ 1'b0 ;
  assign n4067 = n4064 & ~n4066 ;
  assign n4068 = ( n4052 & n4063 ) | ( n4052 & n4067 ) | ( n4063 & n4067 ) ;
  assign n4078 = n4077 ^ n4073 ^ n4068 ;
  assign n4079 = n2742 ^ n2329 ^ n568 ;
  assign n4080 = n4079 ^ n2274 ^ n759 ;
  assign n4081 = ~n1198 & n4080 ;
  assign n4082 = ~n1803 & n4081 ;
  assign n4083 = ( n2251 & n2842 ) | ( n2251 & ~n4082 ) | ( n2842 & ~n4082 ) ;
  assign n4084 = n625 | n1406 ;
  assign n4085 = n1443 & ~n4084 ;
  assign n4086 = ( ~n310 & n2701 ) | ( ~n310 & n4085 ) | ( n2701 & n4085 ) ;
  assign n4090 = n2767 ^ n1139 ^ n673 ;
  assign n4087 = ( ~x165 & n1897 ) | ( ~x165 & n2368 ) | ( n1897 & n2368 ) ;
  assign n4088 = n4087 ^ n1388 ^ x36 ;
  assign n4089 = ~n2128 & n4088 ;
  assign n4091 = n4090 ^ n4089 ^ 1'b0 ;
  assign n4092 = ( n4083 & n4086 ) | ( n4083 & ~n4091 ) | ( n4086 & ~n4091 ) ;
  assign n4100 = ( n2157 & n2336 ) | ( n2157 & n3643 ) | ( n2336 & n3643 ) ;
  assign n4101 = n4100 ^ n1383 ^ n1152 ;
  assign n4093 = n3186 ^ n882 ^ 1'b0 ;
  assign n4096 = n3369 ^ n2192 ^ n2037 ;
  assign n4097 = ( ~n3006 & n3350 ) | ( ~n3006 & n4096 ) | ( n3350 & n4096 ) ;
  assign n4094 = ( ~n760 & n1390 ) | ( ~n760 & n1474 ) | ( n1390 & n1474 ) ;
  assign n4095 = n4094 ^ n2081 ^ n846 ;
  assign n4098 = n4097 ^ n4095 ^ 1'b0 ;
  assign n4099 = ( x173 & n4093 ) | ( x173 & ~n4098 ) | ( n4093 & ~n4098 ) ;
  assign n4102 = n4101 ^ n4099 ^ n1595 ;
  assign n4103 = ( ~n866 & n4092 ) | ( ~n866 & n4102 ) | ( n4092 & n4102 ) ;
  assign n4112 = n3807 ^ n2509 ^ n2328 ;
  assign n4108 = ~n525 & n827 ;
  assign n4109 = n4108 ^ n3259 ^ 1'b0 ;
  assign n4110 = n4109 ^ n729 ^ n535 ;
  assign n4111 = ( ~n2687 & n3016 ) | ( ~n2687 & n4110 ) | ( n3016 & n4110 ) ;
  assign n4113 = n4112 ^ n4111 ^ n4065 ;
  assign n4114 = n914 | n1227 ;
  assign n4115 = n4114 ^ n608 ^ 1'b0 ;
  assign n4116 = ( x32 & ~n2235 ) | ( x32 & n3065 ) | ( ~n2235 & n3065 ) ;
  assign n4117 = n3804 ^ n2781 ^ n334 ;
  assign n4118 = ~n4116 & n4117 ;
  assign n4119 = ( n2516 & n4115 ) | ( n2516 & ~n4118 ) | ( n4115 & ~n4118 ) ;
  assign n4120 = ( n3616 & ~n4113 ) | ( n3616 & n4119 ) | ( ~n4113 & n4119 ) ;
  assign n4121 = ( n1838 & n2862 ) | ( n1838 & n4120 ) | ( n2862 & n4120 ) ;
  assign n4104 = ( ~n387 & n2198 ) | ( ~n387 & n3089 ) | ( n2198 & n3089 ) ;
  assign n4105 = ( n2275 & n2714 ) | ( n2275 & n4104 ) | ( n2714 & n4104 ) ;
  assign n4106 = n2679 & n4105 ;
  assign n4107 = n780 & n4106 ;
  assign n4122 = n4121 ^ n4107 ^ n3564 ;
  assign n4123 = ( n488 & n2652 ) | ( n488 & n3451 ) | ( n2652 & n3451 ) ;
  assign n4124 = n651 & n4123 ;
  assign n4125 = n2172 & n4124 ;
  assign n4133 = n1650 ^ n449 ^ x1 ;
  assign n4134 = ( x193 & ~n3357 ) | ( x193 & n4133 ) | ( ~n3357 & n4133 ) ;
  assign n4132 = ( n855 & n1436 ) | ( n855 & n2499 ) | ( n1436 & n2499 ) ;
  assign n4128 = ( n542 & n598 ) | ( n542 & ~n3726 ) | ( n598 & ~n3726 ) ;
  assign n4126 = n2553 ^ n1389 ^ n971 ;
  assign n4127 = ( n1533 & ~n1645 ) | ( n1533 & n4126 ) | ( ~n1645 & n4126 ) ;
  assign n4129 = n4128 ^ n4127 ^ n1235 ;
  assign n4130 = n3409 | n4129 ;
  assign n4131 = n978 | n4130 ;
  assign n4135 = n4134 ^ n4132 ^ n4131 ;
  assign n4136 = ( ~x186 & n1181 ) | ( ~x186 & n3165 ) | ( n1181 & n3165 ) ;
  assign n4137 = n4136 ^ n1527 ^ 1'b0 ;
  assign n4140 = ( x171 & n625 ) | ( x171 & n1297 ) | ( n625 & n1297 ) ;
  assign n4141 = n4140 ^ n2899 ^ 1'b0 ;
  assign n4138 = n2499 ^ n1888 ^ 1'b0 ;
  assign n4139 = x103 & n4138 ;
  assign n4142 = n4141 ^ n4139 ^ n2169 ;
  assign n4148 = ( ~n305 & n312 ) | ( ~n305 & n1010 ) | ( n312 & n1010 ) ;
  assign n4149 = n4148 ^ n334 ^ x41 ;
  assign n4147 = n3921 ^ n1745 ^ x25 ;
  assign n4150 = n4149 ^ n4147 ^ n895 ;
  assign n4144 = n1292 ^ n859 ^ n846 ;
  assign n4143 = n2659 ^ x72 ^ 1'b0 ;
  assign n4145 = n4144 ^ n4143 ^ n1752 ;
  assign n4146 = ~n3302 & n4145 ;
  assign n4151 = n4150 ^ n4146 ^ 1'b0 ;
  assign n4152 = n3923 ^ n1169 ^ n846 ;
  assign n4153 = ( n3540 & n4151 ) | ( n3540 & ~n4152 ) | ( n4151 & ~n4152 ) ;
  assign n4154 = ( ~n471 & n1061 ) | ( ~n471 & n1288 ) | ( n1061 & n1288 ) ;
  assign n4155 = n4154 ^ n3917 ^ n541 ;
  assign n4156 = n2902 ^ n1511 ^ 1'b0 ;
  assign n4157 = ( n1055 & n1307 ) | ( n1055 & n4156 ) | ( n1307 & n4156 ) ;
  assign n4158 = n529 ^ n511 ^ 1'b0 ;
  assign n4159 = n912 ^ n710 ^ 1'b0 ;
  assign n4160 = ( n2523 & n4158 ) | ( n2523 & n4159 ) | ( n4158 & n4159 ) ;
  assign n4161 = n3653 ^ n2296 ^ n1271 ;
  assign n4162 = n400 & ~n1307 ;
  assign n4163 = ~n2257 & n4162 ;
  assign n4164 = n4163 ^ n1900 ^ 1'b0 ;
  assign n4165 = ( n629 & n1141 ) | ( n629 & n4164 ) | ( n1141 & n4164 ) ;
  assign n4166 = ( n4160 & n4161 ) | ( n4160 & ~n4165 ) | ( n4161 & ~n4165 ) ;
  assign n4181 = ( ~n1270 & n1309 ) | ( ~n1270 & n1563 ) | ( n1309 & n1563 ) ;
  assign n4182 = n4181 ^ n1440 ^ n583 ;
  assign n4183 = n1973 ^ n1297 ^ 1'b0 ;
  assign n4184 = ~n4182 & n4183 ;
  assign n4176 = ( x53 & ~n627 ) | ( x53 & n2066 ) | ( ~n627 & n2066 ) ;
  assign n4177 = ( n372 & ~n2085 ) | ( n372 & n4176 ) | ( ~n2085 & n4176 ) ;
  assign n4174 = n1348 ^ n583 ^ x173 ;
  assign n4175 = x202 & ~n4174 ;
  assign n4178 = n4177 ^ n4175 ^ 1'b0 ;
  assign n4171 = ( n614 & ~n1219 ) | ( n614 & n2536 ) | ( ~n1219 & n2536 ) ;
  assign n4172 = ( n488 & n1668 ) | ( n488 & ~n4171 ) | ( n1668 & ~n4171 ) ;
  assign n4173 = ( ~n575 & n1958 ) | ( ~n575 & n4172 ) | ( n1958 & n4172 ) ;
  assign n4179 = n4178 ^ n4173 ^ 1'b0 ;
  assign n4180 = ~n1985 & n4179 ;
  assign n4167 = ( x125 & ~n1941 ) | ( x125 & n3382 ) | ( ~n1941 & n3382 ) ;
  assign n4168 = n2378 ^ n1613 ^ n857 ;
  assign n4169 = ( n745 & n1718 ) | ( n745 & n1827 ) | ( n1718 & n1827 ) ;
  assign n4170 = ( n4167 & ~n4168 ) | ( n4167 & n4169 ) | ( ~n4168 & n4169 ) ;
  assign n4185 = n4184 ^ n4180 ^ n4170 ;
  assign n4201 = n3103 ^ n1589 ^ x67 ;
  assign n4186 = n1423 ^ n597 ^ 1'b0 ;
  assign n4187 = n733 | n4186 ;
  assign n4198 = n2222 ^ n589 ^ x61 ;
  assign n4196 = n1829 ^ n981 ^ n548 ;
  assign n4190 = n817 & ~n1757 ;
  assign n4191 = n4190 ^ n2656 ^ 1'b0 ;
  assign n4192 = ( n727 & ~n1377 ) | ( n727 & n4191 ) | ( ~n1377 & n4191 ) ;
  assign n4193 = ~n4177 & n4192 ;
  assign n4194 = ~n2662 & n4193 ;
  assign n4195 = n4194 ^ n1031 ^ 1'b0 ;
  assign n4188 = x179 & ~n2831 ;
  assign n4189 = n2292 & n4188 ;
  assign n4197 = n4196 ^ n4195 ^ n4189 ;
  assign n4199 = n4198 ^ n4197 ^ x135 ;
  assign n4200 = n4187 | n4199 ;
  assign n4202 = n4201 ^ n4200 ^ 1'b0 ;
  assign n4203 = ( ~n418 & n2237 ) | ( ~n418 & n4202 ) | ( n2237 & n4202 ) ;
  assign n4204 = n968 ^ n813 ^ x49 ;
  assign n4205 = n3412 & ~n3788 ;
  assign n4206 = ( x52 & ~n332 ) | ( x52 & n4205 ) | ( ~n332 & n4205 ) ;
  assign n4207 = ( n1452 & n4204 ) | ( n1452 & ~n4206 ) | ( n4204 & ~n4206 ) ;
  assign n4210 = ( n260 & ~n1217 ) | ( n260 & n2337 ) | ( ~n1217 & n2337 ) ;
  assign n4209 = n1617 ^ n1238 ^ 1'b0 ;
  assign n4208 = ( x82 & ~n266 ) | ( x82 & n1244 ) | ( ~n266 & n1244 ) ;
  assign n4211 = n4210 ^ n4209 ^ n4208 ;
  assign n4212 = ( ~n1300 & n1557 ) | ( ~n1300 & n3862 ) | ( n1557 & n3862 ) ;
  assign n4213 = n4212 ^ n3064 ^ 1'b0 ;
  assign n4219 = ( ~n2200 & n2844 ) | ( ~n2200 & n3650 ) | ( n2844 & n3650 ) ;
  assign n4214 = ( n305 & n1063 ) | ( n305 & n2282 ) | ( n1063 & n2282 ) ;
  assign n4215 = ( x177 & ~n1206 ) | ( x177 & n2261 ) | ( ~n1206 & n2261 ) ;
  assign n4216 = ( n4094 & n4214 ) | ( n4094 & ~n4215 ) | ( n4214 & ~n4215 ) ;
  assign n4217 = ( ~n266 & n1154 ) | ( ~n266 & n1423 ) | ( n1154 & n1423 ) ;
  assign n4218 = ( ~n2801 & n4216 ) | ( ~n2801 & n4217 ) | ( n4216 & n4217 ) ;
  assign n4220 = n4219 ^ n4218 ^ 1'b0 ;
  assign n4221 = ( n3720 & n4213 ) | ( n3720 & n4220 ) | ( n4213 & n4220 ) ;
  assign n4225 = x110 & ~n519 ;
  assign n4226 = ~n4087 & n4225 ;
  assign n4224 = ( ~x200 & n1478 ) | ( ~x200 & n2760 ) | ( n1478 & n2760 ) ;
  assign n4227 = n4226 ^ n4224 ^ n1877 ;
  assign n4228 = n4227 ^ n3997 ^ x247 ;
  assign n4222 = ( x165 & n424 ) | ( x165 & ~n1897 ) | ( n424 & ~n1897 ) ;
  assign n4223 = n310 & ~n4222 ;
  assign n4229 = n4228 ^ n4223 ^ n2385 ;
  assign n4230 = n1673 ^ n730 ^ x25 ;
  assign n4234 = n2651 ^ n1645 ^ 1'b0 ;
  assign n4235 = n4234 ^ n1121 ^ x189 ;
  assign n4232 = n1365 ^ n1100 ^ n1088 ;
  assign n4233 = ( n2533 & ~n3084 ) | ( n2533 & n4232 ) | ( ~n3084 & n4232 ) ;
  assign n4231 = n2669 ^ n1695 ^ n1115 ;
  assign n4236 = n4235 ^ n4233 ^ n4231 ;
  assign n4237 = n257 & ~n4236 ;
  assign n4238 = n2877 ^ n1233 ^ n628 ;
  assign n4239 = n4085 ^ n3338 ^ n728 ;
  assign n4240 = n4239 ^ n2874 ^ n2617 ;
  assign n4241 = ( ~n1194 & n4238 ) | ( ~n1194 & n4240 ) | ( n4238 & n4240 ) ;
  assign n4242 = ( ~n479 & n1751 ) | ( ~n479 & n4241 ) | ( n1751 & n4241 ) ;
  assign n4243 = ( n4230 & n4237 ) | ( n4230 & ~n4242 ) | ( n4237 & ~n4242 ) ;
  assign n4244 = ( n452 & n1191 ) | ( n452 & ~n2510 ) | ( n1191 & ~n2510 ) ;
  assign n4245 = ( ~n430 & n1771 ) | ( ~n430 & n3119 ) | ( n1771 & n3119 ) ;
  assign n4246 = ( ~n1506 & n2278 ) | ( ~n1506 & n4245 ) | ( n2278 & n4245 ) ;
  assign n4247 = n4246 ^ n4145 ^ n1457 ;
  assign n4248 = ( n2257 & n4244 ) | ( n2257 & ~n4247 ) | ( n4244 & ~n4247 ) ;
  assign n4249 = n554 & n1145 ;
  assign n4250 = n4249 ^ n2085 ^ 1'b0 ;
  assign n4251 = ~n2557 & n4250 ;
  assign n4252 = ~n640 & n4251 ;
  assign n4253 = n326 | n4252 ;
  assign n4254 = n4248 | n4253 ;
  assign n4255 = n4083 & n4254 ;
  assign n4256 = n4255 ^ n2217 ^ 1'b0 ;
  assign n4260 = n3165 ^ n1509 ^ n602 ;
  assign n4261 = ( n3534 & n3897 ) | ( n3534 & ~n4260 ) | ( n3897 & ~n4260 ) ;
  assign n4258 = n768 ^ n466 ^ 1'b0 ;
  assign n4257 = n3486 ^ n1123 ^ x126 ;
  assign n4259 = n4258 ^ n4257 ^ n2148 ;
  assign n4262 = n4261 ^ n4259 ^ n2358 ;
  assign n4263 = n4262 ^ n1323 ^ n660 ;
  assign n4264 = ( n1471 & ~n2600 ) | ( n1471 & n4263 ) | ( ~n2600 & n4263 ) ;
  assign n4266 = ~n300 & n520 ;
  assign n4265 = n3432 ^ n1549 ^ n512 ;
  assign n4267 = n4266 ^ n4265 ^ n3524 ;
  assign n4268 = n4264 & ~n4267 ;
  assign n4269 = ~n2099 & n4268 ;
  assign n4270 = n610 ^ n386 ^ 1'b0 ;
  assign n4271 = n3070 | n4270 ;
  assign n4272 = n1543 & ~n4271 ;
  assign n4273 = n4272 ^ n2172 ^ 1'b0 ;
  assign n4274 = ( ~n386 & n2668 ) | ( ~n386 & n4273 ) | ( n2668 & n4273 ) ;
  assign n4275 = ( n1667 & ~n2877 ) | ( n1667 & n3598 ) | ( ~n2877 & n3598 ) ;
  assign n4276 = n337 & n4275 ;
  assign n4277 = ~x217 & n4276 ;
  assign n4278 = n4277 ^ n2987 ^ n775 ;
  assign n4279 = n4278 ^ n3957 ^ n1977 ;
  assign n4280 = n1811 ^ n884 ^ 1'b0 ;
  assign n4281 = ~n1529 & n4280 ;
  assign n4282 = ( n2041 & n2386 ) | ( n2041 & n4281 ) | ( n2386 & n4281 ) ;
  assign n4283 = ~n2223 & n4282 ;
  assign n4284 = ( n1264 & n2771 ) | ( n1264 & ~n3308 ) | ( n2771 & ~n3308 ) ;
  assign n4285 = n3744 ^ n1737 ^ n1133 ;
  assign n4286 = ( n984 & n1943 ) | ( n984 & n4285 ) | ( n1943 & n4285 ) ;
  assign n4287 = n4286 ^ n3675 ^ n1903 ;
  assign n4288 = n3436 ^ n983 ^ x24 ;
  assign n4289 = ( n4284 & ~n4287 ) | ( n4284 & n4288 ) | ( ~n4287 & n4288 ) ;
  assign n4290 = n4283 & n4289 ;
  assign n4304 = ( n831 & n1472 ) | ( n831 & ~n1714 ) | ( n1472 & ~n1714 ) ;
  assign n4302 = ( ~x239 & n601 ) | ( ~x239 & n1929 ) | ( n601 & n1929 ) ;
  assign n4303 = ( n2732 & n3771 ) | ( n2732 & n4302 ) | ( n3771 & n4302 ) ;
  assign n4291 = ( n262 & n2152 ) | ( n262 & n2784 ) | ( n2152 & n2784 ) ;
  assign n4292 = ( n3205 & n3841 ) | ( n3205 & n4291 ) | ( n3841 & n4291 ) ;
  assign n4293 = ( n534 & ~n1225 ) | ( n534 & n3461 ) | ( ~n1225 & n3461 ) ;
  assign n4294 = ( x101 & ~n853 ) | ( x101 & n2952 ) | ( ~n853 & n2952 ) ;
  assign n4295 = ( ~n923 & n2381 ) | ( ~n923 & n4294 ) | ( n2381 & n4294 ) ;
  assign n4296 = n1864 | n4295 ;
  assign n4297 = n2287 & ~n4296 ;
  assign n4298 = ( ~n3687 & n4293 ) | ( ~n3687 & n4297 ) | ( n4293 & n4297 ) ;
  assign n4299 = ( ~n915 & n1576 ) | ( ~n915 & n3002 ) | ( n1576 & n3002 ) ;
  assign n4300 = ( n1175 & ~n4298 ) | ( n1175 & n4299 ) | ( ~n4298 & n4299 ) ;
  assign n4301 = n4292 | n4300 ;
  assign n4305 = n4304 ^ n4303 ^ n4301 ;
  assign n4306 = n1696 ^ n1507 ^ x15 ;
  assign n4307 = n4306 ^ x197 ^ x151 ;
  assign n4308 = n2303 ^ n1313 ^ n367 ;
  assign n4309 = n4308 ^ n2735 ^ n985 ;
  assign n4310 = n4309 ^ n3138 ^ n828 ;
  assign n4311 = ~n4307 & n4310 ;
  assign n4312 = n4311 ^ n3068 ^ 1'b0 ;
  assign n4313 = x200 & n2860 ;
  assign n4314 = n4313 ^ n690 ^ 1'b0 ;
  assign n4315 = ( ~n990 & n2886 ) | ( ~n990 & n4314 ) | ( n2886 & n4314 ) ;
  assign n4316 = n1785 ^ n1129 ^ n843 ;
  assign n4317 = ( n350 & n2359 ) | ( n350 & ~n4316 ) | ( n2359 & ~n4316 ) ;
  assign n4318 = n4043 | n4317 ;
  assign n4326 = n2620 ^ n883 ^ n686 ;
  assign n4319 = ( ~n857 & n2825 ) | ( ~n857 & n3780 ) | ( n2825 & n3780 ) ;
  assign n4320 = ( x36 & n729 ) | ( x36 & n758 ) | ( n729 & n758 ) ;
  assign n4321 = ( n683 & n743 ) | ( n683 & n2984 ) | ( n743 & n2984 ) ;
  assign n4322 = n1141 ^ n745 ^ x132 ;
  assign n4323 = n4322 ^ n1671 ^ n507 ;
  assign n4324 = ( n4320 & n4321 ) | ( n4320 & ~n4323 ) | ( n4321 & ~n4323 ) ;
  assign n4325 = ~n4319 & n4324 ;
  assign n4327 = n4326 ^ n4325 ^ 1'b0 ;
  assign n4329 = ( n691 & ~n899 ) | ( n691 & n1542 ) | ( ~n899 & n1542 ) ;
  assign n4330 = x163 & ~n3406 ;
  assign n4331 = n4329 & n4330 ;
  assign n4332 = n4331 ^ n2679 ^ n848 ;
  assign n4328 = n685 & n3465 ;
  assign n4333 = n4332 ^ n4328 ^ 1'b0 ;
  assign n4334 = ( n918 & n3114 ) | ( n918 & n4333 ) | ( n3114 & n4333 ) ;
  assign n4335 = ( n2933 & ~n3368 ) | ( n2933 & n4334 ) | ( ~n3368 & n4334 ) ;
  assign n4336 = n2735 ^ n1188 ^ n338 ;
  assign n4337 = ( n1288 & n2014 ) | ( n1288 & ~n4336 ) | ( n2014 & ~n4336 ) ;
  assign n4338 = n2545 ^ n1579 ^ x11 ;
  assign n4339 = ( ~n1257 & n4337 ) | ( ~n1257 & n4338 ) | ( n4337 & n4338 ) ;
  assign n4340 = ( ~n302 & n869 ) | ( ~n302 & n1485 ) | ( n869 & n1485 ) ;
  assign n4341 = ( n463 & n3703 ) | ( n463 & ~n4340 ) | ( n3703 & ~n4340 ) ;
  assign n4342 = ( n740 & ~n3376 ) | ( n740 & n4341 ) | ( ~n3376 & n4341 ) ;
  assign n4343 = n4342 ^ n1861 ^ n1266 ;
  assign n4344 = n3991 ^ n3356 ^ x250 ;
  assign n4345 = n4344 ^ n4266 ^ n2952 ;
  assign n4346 = n1297 & ~n4345 ;
  assign n4347 = n1244 ^ n1060 ^ n688 ;
  assign n4350 = n1573 ^ n1474 ^ n805 ;
  assign n4351 = ( n1794 & ~n3532 ) | ( n1794 & n4350 ) | ( ~n3532 & n4350 ) ;
  assign n4348 = n2907 ^ n2702 ^ 1'b0 ;
  assign n4349 = n324 & ~n4348 ;
  assign n4352 = n4351 ^ n4349 ^ n1847 ;
  assign n4353 = ( n1428 & n4347 ) | ( n1428 & n4352 ) | ( n4347 & n4352 ) ;
  assign n4354 = n3432 ^ n1254 ^ n1165 ;
  assign n4355 = ( n2930 & ~n3348 ) | ( n2930 & n4354 ) | ( ~n3348 & n4354 ) ;
  assign n4356 = ( n1839 & ~n4353 ) | ( n1839 & n4355 ) | ( ~n4353 & n4355 ) ;
  assign n4357 = n1336 ^ n700 ^ n311 ;
  assign n4358 = ( n1585 & n2398 ) | ( n1585 & n4357 ) | ( n2398 & n4357 ) ;
  assign n4359 = n1797 | n4358 ;
  assign n4360 = n4052 ^ n2001 ^ n473 ;
  assign n4361 = ( n352 & ~n462 ) | ( n352 & n4360 ) | ( ~n462 & n4360 ) ;
  assign n4362 = ( n3218 & n4359 ) | ( n3218 & n4361 ) | ( n4359 & n4361 ) ;
  assign n4363 = ( ~n1135 & n3525 ) | ( ~n1135 & n4362 ) | ( n3525 & n4362 ) ;
  assign n4364 = ( n326 & n1268 ) | ( n326 & ~n1328 ) | ( n1268 & ~n1328 ) ;
  assign n4365 = n3414 | n4364 ;
  assign n4366 = n4365 ^ n2724 ^ 1'b0 ;
  assign n4367 = n4366 ^ n3641 ^ n312 ;
  assign n4368 = n4367 ^ n3383 ^ 1'b0 ;
  assign n4369 = ( x39 & n261 ) | ( x39 & n4368 ) | ( n261 & n4368 ) ;
  assign n4370 = ( ~x153 & x204 ) | ( ~x153 & n2199 ) | ( x204 & n2199 ) ;
  assign n4371 = n2233 ^ n1761 ^ n1098 ;
  assign n4372 = ~n1245 & n2072 ;
  assign n4373 = n4372 ^ n3305 ^ 1'b0 ;
  assign n4374 = ( n4370 & ~n4371 ) | ( n4370 & n4373 ) | ( ~n4371 & n4373 ) ;
  assign n4376 = n2492 ^ n1574 ^ n1356 ;
  assign n4377 = ( n1146 & n1442 ) | ( n1146 & ~n4376 ) | ( n1442 & ~n4376 ) ;
  assign n4375 = ( n930 & n1118 ) | ( n930 & ~n2303 ) | ( n1118 & ~n2303 ) ;
  assign n4378 = n4377 ^ n4375 ^ n1714 ;
  assign n4379 = n4378 ^ n329 ^ 1'b0 ;
  assign n4380 = ( n269 & n673 ) | ( n269 & n4126 ) | ( n673 & n4126 ) ;
  assign n4381 = n4048 ^ n2620 ^ n2028 ;
  assign n4382 = ( n709 & n3382 ) | ( n709 & ~n4381 ) | ( n3382 & ~n4381 ) ;
  assign n4383 = ( x113 & n4380 ) | ( x113 & n4382 ) | ( n4380 & n4382 ) ;
  assign n4384 = ( n465 & n3182 ) | ( n465 & n4383 ) | ( n3182 & n4383 ) ;
  assign n4385 = n2601 ^ n271 ^ x104 ;
  assign n4386 = ( n1119 & ~n2423 ) | ( n1119 & n4385 ) | ( ~n2423 & n4385 ) ;
  assign n4390 = ( n789 & ~n1152 ) | ( n789 & n1292 ) | ( ~n1152 & n1292 ) ;
  assign n4391 = ( n1194 & n2515 ) | ( n1194 & ~n4390 ) | ( n2515 & ~n4390 ) ;
  assign n4393 = n1029 ^ n906 ^ n269 ;
  assign n4394 = n4393 ^ n2727 ^ n1377 ;
  assign n4395 = n4394 ^ n767 ^ n751 ;
  assign n4392 = n2536 & n3535 ;
  assign n4396 = n4395 ^ n4392 ^ 1'b0 ;
  assign n4397 = n1147 ^ n605 ^ 1'b0 ;
  assign n4398 = ~n4085 & n4397 ;
  assign n4399 = n4398 ^ n653 ^ n477 ;
  assign n4400 = n4399 ^ n1973 ^ n1228 ;
  assign n4401 = ( ~n4391 & n4396 ) | ( ~n4391 & n4400 ) | ( n4396 & n4400 ) ;
  assign n4404 = n2140 ^ n979 ^ 1'b0 ;
  assign n4402 = n2429 ^ n1293 ^ n680 ;
  assign n4403 = ( x235 & n1334 ) | ( x235 & ~n4402 ) | ( n1334 & ~n4402 ) ;
  assign n4405 = n4404 ^ n4403 ^ n2941 ;
  assign n4406 = ( n1367 & n4401 ) | ( n1367 & ~n4405 ) | ( n4401 & ~n4405 ) ;
  assign n4387 = n601 ^ n582 ^ x2 ;
  assign n4388 = n3559 ^ n2674 ^ 1'b0 ;
  assign n4389 = n4387 | n4388 ;
  assign n4407 = n4406 ^ n4389 ^ n973 ;
  assign n4408 = ~n729 & n1024 ;
  assign n4409 = n759 & ~n1002 ;
  assign n4410 = n4409 ^ n648 ^ 1'b0 ;
  assign n4411 = ( n2047 & ~n3763 ) | ( n2047 & n4410 ) | ( ~n3763 & n4410 ) ;
  assign n4412 = n1559 ^ n1349 ^ n1191 ;
  assign n4413 = ( ~n2454 & n2777 ) | ( ~n2454 & n4412 ) | ( n2777 & n4412 ) ;
  assign n4414 = ( ~n4408 & n4411 ) | ( ~n4408 & n4413 ) | ( n4411 & n4413 ) ;
  assign n4424 = n1629 ^ n1619 ^ n1427 ;
  assign n4421 = x41 & ~n988 ;
  assign n4422 = n2002 & n4421 ;
  assign n4419 = n3743 ^ n1634 ^ 1'b0 ;
  assign n4420 = n4419 ^ n3098 ^ n2508 ;
  assign n4423 = n4422 ^ n4420 ^ n1272 ;
  assign n4417 = ( ~x134 & x215 ) | ( ~x134 & n741 ) | ( x215 & n741 ) ;
  assign n4415 = n656 ^ n321 ^ 1'b0 ;
  assign n4416 = ( ~x24 & n1966 ) | ( ~x24 & n4415 ) | ( n1966 & n4415 ) ;
  assign n4418 = n4417 ^ n4416 ^ n938 ;
  assign n4425 = n4424 ^ n4423 ^ n4418 ;
  assign n4433 = n2578 ^ n2206 ^ 1'b0 ;
  assign n4434 = n4433 ^ n1478 ^ n1030 ;
  assign n4426 = n3639 ^ n2205 ^ n1371 ;
  assign n4427 = ( ~n846 & n2914 ) | ( ~n846 & n4426 ) | ( n2914 & n4426 ) ;
  assign n4428 = n4427 ^ x24 ^ 1'b0 ;
  assign n4429 = n759 & n3798 ;
  assign n4430 = n4429 ^ n3661 ^ n2093 ;
  assign n4431 = n4430 ^ n3891 ^ n3282 ;
  assign n4432 = ~n4428 & n4431 ;
  assign n4435 = n4434 ^ n4432 ^ 1'b0 ;
  assign n4436 = n1513 ^ n1049 ^ x68 ;
  assign n4437 = ( n2744 & n4051 ) | ( n2744 & ~n4436 ) | ( n4051 & ~n4436 ) ;
  assign n4439 = ( ~x151 & x156 ) | ( ~x151 & n513 ) | ( x156 & n513 ) ;
  assign n4440 = n3488 ^ n3035 ^ n710 ;
  assign n4441 = ( n1524 & n4439 ) | ( n1524 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4438 = n608 & n759 ;
  assign n4442 = n4441 ^ n4438 ^ n3462 ;
  assign n4443 = ( n975 & n1667 ) | ( n975 & n2611 ) | ( n1667 & n2611 ) ;
  assign n4444 = ( ~n1212 & n2218 ) | ( ~n1212 & n4443 ) | ( n2218 & n4443 ) ;
  assign n4460 = ( n510 & ~n859 ) | ( n510 & n1787 ) | ( ~n859 & n1787 ) ;
  assign n4461 = x67 & n4460 ;
  assign n4462 = n4461 ^ n286 ^ 1'b0 ;
  assign n4459 = n519 | n639 ;
  assign n4463 = n4462 ^ n4459 ^ n1346 ;
  assign n4456 = ( x38 & ~n1232 ) | ( x38 & n2195 ) | ( ~n1232 & n2195 ) ;
  assign n4457 = n518 & n2420 ;
  assign n4458 = ( n1801 & n4456 ) | ( n1801 & n4457 ) | ( n4456 & n4457 ) ;
  assign n4464 = n4463 ^ n4458 ^ n1909 ;
  assign n4454 = x145 & n3640 ;
  assign n4455 = n4454 ^ n821 ^ n716 ;
  assign n4450 = n1605 & ~n3286 ;
  assign n4451 = n918 & n4450 ;
  assign n4452 = n4451 ^ n2811 ^ 1'b0 ;
  assign n4453 = n4452 ^ n2159 ^ n1059 ;
  assign n4465 = n4464 ^ n4455 ^ n4453 ;
  assign n4445 = n3643 ^ n471 ^ x17 ;
  assign n4446 = n4445 ^ n2303 ^ n1580 ;
  assign n4447 = n2557 ^ n1902 ^ x156 ;
  assign n4448 = ( n1548 & n2121 ) | ( n1548 & ~n4447 ) | ( n2121 & ~n4447 ) ;
  assign n4449 = ( n314 & ~n4446 ) | ( n314 & n4448 ) | ( ~n4446 & n4448 ) ;
  assign n4466 = n4465 ^ n4449 ^ n3384 ;
  assign n4467 = n600 & n2316 ;
  assign n4468 = ( x27 & x242 ) | ( x27 & ~n1077 ) | ( x242 & ~n1077 ) ;
  assign n4469 = n4316 ^ n673 ^ x208 ;
  assign n4470 = ( n2150 & n4468 ) | ( n2150 & ~n4469 ) | ( n4468 & ~n4469 ) ;
  assign n4475 = ~n1347 & n1428 ;
  assign n4473 = n636 ^ n274 ^ 1'b0 ;
  assign n4471 = ( n591 & ~n1337 ) | ( n591 & n1802 ) | ( ~n1337 & n1802 ) ;
  assign n4472 = ( ~n1396 & n4302 ) | ( ~n1396 & n4471 ) | ( n4302 & n4471 ) ;
  assign n4474 = n4473 ^ n4472 ^ n1236 ;
  assign n4476 = n4475 ^ n4474 ^ n3276 ;
  assign n4477 = ( n4467 & n4470 ) | ( n4467 & n4476 ) | ( n4470 & n4476 ) ;
  assign n4478 = ( n4444 & n4466 ) | ( n4444 & n4477 ) | ( n4466 & n4477 ) ;
  assign n4495 = ( x47 & n2476 ) | ( x47 & ~n3100 ) | ( n2476 & ~n3100 ) ;
  assign n4496 = n2826 ^ n2314 ^ n1755 ;
  assign n4497 = n4496 ^ n1632 ^ 1'b0 ;
  assign n4498 = ( ~n2756 & n4495 ) | ( ~n2756 & n4497 ) | ( n4495 & n4497 ) ;
  assign n4491 = n1856 ^ n1210 ^ 1'b0 ;
  assign n4492 = ~n719 & n4491 ;
  assign n4493 = n4492 ^ n1592 ^ n640 ;
  assign n4486 = n917 & n1322 ;
  assign n4487 = n1198 & n4486 ;
  assign n4484 = ( n724 & ~n889 ) | ( n724 & n1856 ) | ( ~n889 & n1856 ) ;
  assign n4485 = ( n1335 & n3203 ) | ( n1335 & ~n4484 ) | ( n3203 & ~n4484 ) ;
  assign n4479 = n2127 ^ n1330 ^ 1'b0 ;
  assign n4480 = x43 & n4479 ;
  assign n4481 = ( n2310 & n4275 ) | ( n2310 & ~n4480 ) | ( n4275 & ~n4480 ) ;
  assign n4482 = ( n1187 & n2063 ) | ( n1187 & ~n2690 ) | ( n2063 & ~n2690 ) ;
  assign n4483 = n4481 | n4482 ;
  assign n4488 = n4487 ^ n4485 ^ n4483 ;
  assign n4489 = n4488 ^ n1755 ^ 1'b0 ;
  assign n4490 = n3461 & ~n4489 ;
  assign n4494 = n4493 ^ n4490 ^ x172 ;
  assign n4499 = n4498 ^ n4494 ^ n4148 ;
  assign n4502 = x6 | n1035 ;
  assign n4503 = n1582 | n4502 ;
  assign n4504 = ( n838 & n2458 ) | ( n838 & ~n4503 ) | ( n2458 & ~n4503 ) ;
  assign n4500 = n2657 ^ n1385 ^ n685 ;
  assign n4501 = n4500 ^ n3387 ^ n1787 ;
  assign n4505 = n4504 ^ n4501 ^ x253 ;
  assign n4506 = n4505 ^ n3846 ^ n362 ;
  assign n4509 = n4314 ^ n2842 ^ n1708 ;
  assign n4507 = x211 & ~n2813 ;
  assign n4508 = ( n1235 & ~n2006 ) | ( n1235 & n4507 ) | ( ~n2006 & n4507 ) ;
  assign n4510 = n4509 ^ n4508 ^ n1586 ;
  assign n4511 = n2822 ^ n1959 ^ n1259 ;
  assign n4512 = n4510 & n4511 ;
  assign n4513 = n2751 & n4512 ;
  assign n4514 = n4140 ^ n2373 ^ n2333 ;
  assign n4515 = n4514 ^ n4492 ^ n326 ;
  assign n4516 = n2221 ^ n256 ^ x115 ;
  assign n4518 = n1330 ^ n1211 ^ x249 ;
  assign n4517 = n4376 ^ n3332 ^ 1'b0 ;
  assign n4519 = n4518 ^ n4517 ^ n4473 ;
  assign n4520 = n3464 ^ n2206 ^ n1341 ;
  assign n4528 = ( n416 & ~n1035 ) | ( n416 & n1622 ) | ( ~n1035 & n1622 ) ;
  assign n4524 = n3539 | n4037 ;
  assign n4525 = n4524 ^ n1286 ^ 1'b0 ;
  assign n4526 = ( ~n1589 & n1653 ) | ( ~n1589 & n4525 ) | ( n1653 & n4525 ) ;
  assign n4522 = ( x121 & n1261 ) | ( x121 & ~n1277 ) | ( n1261 & ~n1277 ) ;
  assign n4521 = ( n498 & ~n2058 ) | ( n498 & n2226 ) | ( ~n2058 & n2226 ) ;
  assign n4523 = n4522 ^ n4521 ^ n4111 ;
  assign n4527 = n4526 ^ n4523 ^ x242 ;
  assign n4529 = n4528 ^ n4527 ^ n870 ;
  assign n4530 = n4529 ^ x8 ^ 1'b0 ;
  assign n4531 = n4520 | n4530 ;
  assign n4532 = ( n836 & ~n1893 ) | ( n836 & n3088 ) | ( ~n1893 & n3088 ) ;
  assign n4533 = ( ~x224 & n1093 ) | ( ~x224 & n1947 ) | ( n1093 & n1947 ) ;
  assign n4534 = ( n1712 & ~n2591 ) | ( n1712 & n4533 ) | ( ~n2591 & n4533 ) ;
  assign n4535 = n2687 ^ n2047 ^ n912 ;
  assign n4541 = n2338 ^ n1233 ^ 1'b0 ;
  assign n4542 = n3838 & ~n4541 ;
  assign n4540 = n4501 ^ n1388 ^ n261 ;
  assign n4543 = n4542 ^ n4540 ^ n2096 ;
  assign n4544 = ( n796 & ~n2428 ) | ( n796 & n3656 ) | ( ~n2428 & n3656 ) ;
  assign n4545 = ( n3533 & n4503 ) | ( n3533 & ~n4544 ) | ( n4503 & ~n4544 ) ;
  assign n4546 = n4545 ^ n535 ^ 1'b0 ;
  assign n4547 = ~n4543 & n4546 ;
  assign n4536 = n4332 ^ n2364 ^ n367 ;
  assign n4537 = n929 | n4536 ;
  assign n4538 = n3831 | n4537 ;
  assign n4539 = ( n514 & ~n2362 ) | ( n514 & n4538 ) | ( ~n2362 & n4538 ) ;
  assign n4548 = n4547 ^ n4539 ^ n1858 ;
  assign n4549 = ( n1152 & n1750 ) | ( n1152 & n2369 ) | ( n1750 & n2369 ) ;
  assign n4556 = ( n2013 & n2234 ) | ( n2013 & n3342 ) | ( n2234 & n3342 ) ;
  assign n4554 = ( n403 & ~n655 ) | ( n403 & n3125 ) | ( ~n655 & n3125 ) ;
  assign n4555 = ~n2709 & n4554 ;
  assign n4550 = x189 & ~n4297 ;
  assign n4551 = n1785 & n4550 ;
  assign n4552 = n2840 | n3763 ;
  assign n4553 = n4551 & ~n4552 ;
  assign n4557 = n4556 ^ n4555 ^ n4553 ;
  assign n4558 = ( n3012 & n4549 ) | ( n3012 & ~n4557 ) | ( n4549 & ~n4557 ) ;
  assign n4559 = n3759 ^ n1802 ^ n1778 ;
  assign n4566 = ( ~n781 & n3974 ) | ( ~n781 & n4364 ) | ( n3974 & n4364 ) ;
  assign n4560 = n3541 ^ n2338 ^ n1917 ;
  assign n4561 = ~n2119 & n4391 ;
  assign n4562 = n1019 & n4561 ;
  assign n4563 = ( ~n423 & n534 ) | ( ~n423 & n2336 ) | ( n534 & n2336 ) ;
  assign n4564 = ( n4560 & n4562 ) | ( n4560 & ~n4563 ) | ( n4562 & ~n4563 ) ;
  assign n4565 = ( n2879 & ~n3518 ) | ( n2879 & n4564 ) | ( ~n3518 & n4564 ) ;
  assign n4567 = n4566 ^ n4565 ^ n2156 ;
  assign n4568 = n4567 ^ n2915 ^ n494 ;
  assign n4569 = ( n2516 & n4559 ) | ( n2516 & ~n4568 ) | ( n4559 & ~n4568 ) ;
  assign n4578 = ( ~n743 & n2537 ) | ( ~n743 & n3232 ) | ( n2537 & n3232 ) ;
  assign n4579 = ( n1527 & ~n2910 ) | ( n1527 & n4578 ) | ( ~n2910 & n4578 ) ;
  assign n4580 = ( n1030 & n1433 ) | ( n1030 & ~n1716 ) | ( n1433 & ~n1716 ) ;
  assign n4581 = n4580 ^ n1974 ^ n781 ;
  assign n4582 = n2603 ^ n1970 ^ n834 ;
  assign n4583 = n4582 ^ n3217 ^ n2969 ;
  assign n4584 = ( n661 & ~n4581 ) | ( n661 & n4583 ) | ( ~n4581 & n4583 ) ;
  assign n4585 = ( ~n420 & n4579 ) | ( ~n420 & n4584 ) | ( n4579 & n4584 ) ;
  assign n4586 = n4585 ^ n4127 ^ n858 ;
  assign n4570 = ( x164 & ~n601 ) | ( x164 & n809 ) | ( ~n601 & n809 ) ;
  assign n4571 = ( n2687 & n3385 ) | ( n2687 & n4570 ) | ( n3385 & n4570 ) ;
  assign n4573 = ( x86 & n501 ) | ( x86 & ~n3702 ) | ( n501 & ~n3702 ) ;
  assign n4572 = n345 & ~n891 ;
  assign n4574 = n4573 ^ n4572 ^ 1'b0 ;
  assign n4575 = n2633 ^ n2532 ^ n1609 ;
  assign n4576 = n4575 ^ n1755 ^ n1733 ;
  assign n4577 = ( ~n4571 & n4574 ) | ( ~n4571 & n4576 ) | ( n4574 & n4576 ) ;
  assign n4587 = n4586 ^ n4577 ^ n3013 ;
  assign n4588 = ( n1362 & n1720 ) | ( n1362 & n1785 ) | ( n1720 & n1785 ) ;
  assign n4589 = n4588 ^ n3014 ^ n1063 ;
  assign n4590 = n807 & n3670 ;
  assign n4591 = n4590 ^ x231 ^ 1'b0 ;
  assign n4592 = ( n4422 & n4589 ) | ( n4422 & n4591 ) | ( n4589 & n4591 ) ;
  assign n4593 = ( n1115 & n1811 ) | ( n1115 & n2273 ) | ( n1811 & n2273 ) ;
  assign n4594 = ~n835 & n1114 ;
  assign n4595 = n4594 ^ n1801 ^ n900 ;
  assign n4596 = ~n1470 & n4595 ;
  assign n4597 = n4596 ^ n1757 ^ 1'b0 ;
  assign n4598 = n3464 ^ n2212 ^ n938 ;
  assign n4599 = n3696 ^ n2932 ^ n1001 ;
  assign n4600 = ( ~n3975 & n4598 ) | ( ~n3975 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4601 = n3350 ^ n1289 ^ 1'b0 ;
  assign n4602 = ~n4600 & n4601 ;
  assign n4603 = ( n4593 & ~n4597 ) | ( n4593 & n4602 ) | ( ~n4597 & n4602 ) ;
  assign n4604 = n1969 ^ n574 ^ x201 ;
  assign n4605 = ( n1319 & n2754 ) | ( n1319 & ~n4604 ) | ( n2754 & ~n4604 ) ;
  assign n4606 = n4605 ^ n2519 ^ n517 ;
  assign n4607 = n4606 ^ n2757 ^ n837 ;
  assign n4616 = x203 & n1505 ;
  assign n4617 = n4616 ^ n2164 ^ n665 ;
  assign n4615 = n2436 ^ n2035 ^ n1784 ;
  assign n4610 = ~n1722 & n3320 ;
  assign n4611 = ( n579 & n1653 ) | ( n579 & ~n4610 ) | ( n1653 & ~n4610 ) ;
  assign n4612 = n4611 ^ n1828 ^ n777 ;
  assign n4608 = n3047 ^ n2220 ^ n1754 ;
  assign n4609 = n4608 ^ n736 ^ n674 ;
  assign n4613 = n4612 ^ n4609 ^ 1'b0 ;
  assign n4614 = n4248 & ~n4613 ;
  assign n4618 = n4617 ^ n4615 ^ n4614 ;
  assign n4619 = ( n1272 & ~n2141 ) | ( n1272 & n3550 ) | ( ~n2141 & n3550 ) ;
  assign n4620 = n3188 ^ n1589 ^ n1484 ;
  assign n4621 = ( n683 & ~n1141 ) | ( n683 & n1345 ) | ( ~n1141 & n1345 ) ;
  assign n4622 = n2644 ^ n1671 ^ 1'b0 ;
  assign n4623 = ( ~n1044 & n4621 ) | ( ~n1044 & n4622 ) | ( n4621 & n4622 ) ;
  assign n4624 = n585 | n1494 ;
  assign n4625 = n4624 ^ n2080 ^ 1'b0 ;
  assign n4626 = n937 & ~n4222 ;
  assign n4627 = n4267 & n4626 ;
  assign n4628 = n943 & ~n4627 ;
  assign n4629 = n4625 & n4628 ;
  assign n4630 = n4629 ^ n2803 ^ n1396 ;
  assign n4631 = ( ~n4620 & n4623 ) | ( ~n4620 & n4630 ) | ( n4623 & n4630 ) ;
  assign n4637 = n2390 ^ n406 ^ x153 ;
  assign n4636 = x234 & n1336 ;
  assign n4638 = n4637 ^ n4636 ^ n2720 ;
  assign n4634 = n2827 ^ n821 ^ 1'b0 ;
  assign n4635 = ~n1591 & n4634 ;
  assign n4639 = n4638 ^ n4635 ^ n1701 ;
  assign n4632 = ( ~n2258 & n3627 ) | ( ~n2258 & n3904 ) | ( n3627 & n3904 ) ;
  assign n4633 = n4632 ^ n4449 ^ n2795 ;
  assign n4640 = n4639 ^ n4633 ^ n2607 ;
  assign n4641 = n4631 & n4640 ;
  assign n4642 = n4619 & n4641 ;
  assign n4643 = n1607 ^ n1443 ^ n1081 ;
  assign n4644 = n3502 ^ n2844 ^ n554 ;
  assign n4645 = n3224 ^ n1364 ^ n898 ;
  assign n4646 = n1424 & n1674 ;
  assign n4647 = ( n839 & n1735 ) | ( n839 & ~n3194 ) | ( n1735 & ~n3194 ) ;
  assign n4648 = n996 ^ n819 ^ x52 ;
  assign n4649 = ( n4646 & n4647 ) | ( n4646 & n4648 ) | ( n4647 & n4648 ) ;
  assign n4650 = ( ~n4644 & n4645 ) | ( ~n4644 & n4649 ) | ( n4645 & n4649 ) ;
  assign n4651 = ( ~n4113 & n4643 ) | ( ~n4113 & n4650 ) | ( n4643 & n4650 ) ;
  assign n4652 = n4651 ^ n2631 ^ n2429 ;
  assign n4653 = n4652 ^ n2452 ^ 1'b0 ;
  assign n4654 = ( n489 & n747 ) | ( n489 & ~n4012 ) | ( n747 & ~n4012 ) ;
  assign n4655 = ( x42 & n967 ) | ( x42 & ~n4654 ) | ( n967 & ~n4654 ) ;
  assign n4656 = n2340 ^ n1811 ^ n266 ;
  assign n4657 = n4656 ^ n3146 ^ n2583 ;
  assign n4660 = n3515 ^ n1745 ^ n1021 ;
  assign n4658 = ( ~n1014 & n2038 ) | ( ~n1014 & n3475 ) | ( n2038 & n3475 ) ;
  assign n4659 = n4658 ^ n2373 ^ n561 ;
  assign n4661 = n4660 ^ n4659 ^ 1'b0 ;
  assign n4662 = ( n4655 & n4657 ) | ( n4655 & ~n4661 ) | ( n4657 & ~n4661 ) ;
  assign n4663 = ( n1288 & n2628 ) | ( n1288 & n2690 ) | ( n2628 & n2690 ) ;
  assign n4672 = n2559 ^ n943 ^ x185 ;
  assign n4670 = ( x183 & n338 ) | ( x183 & ~n1771 ) | ( n338 & ~n1771 ) ;
  assign n4668 = n2370 ^ n1352 ^ n1009 ;
  assign n4669 = ( ~n1257 & n1668 ) | ( ~n1257 & n4668 ) | ( n1668 & n4668 ) ;
  assign n4664 = ~n2147 & n3005 ;
  assign n4665 = n4664 ^ n3173 ^ 1'b0 ;
  assign n4666 = ~n2730 & n4665 ;
  assign n4667 = ~n1282 & n4666 ;
  assign n4671 = n4670 ^ n4669 ^ n4667 ;
  assign n4673 = n4672 ^ n4671 ^ n2965 ;
  assign n4674 = ( ~n4316 & n4663 ) | ( ~n4316 & n4673 ) | ( n4663 & n4673 ) ;
  assign n4678 = ( n818 & n1470 ) | ( n818 & n3328 ) | ( n1470 & n3328 ) ;
  assign n4679 = n4678 ^ n1659 ^ n1637 ;
  assign n4680 = n4679 ^ n3497 ^ n2124 ;
  assign n4681 = n4680 ^ n2324 ^ 1'b0 ;
  assign n4676 = n2089 ^ n1851 ^ x13 ;
  assign n4677 = n4676 ^ n2506 ^ n2351 ;
  assign n4675 = ( n285 & ~n635 ) | ( n285 & n2870 ) | ( ~n635 & n2870 ) ;
  assign n4682 = n4681 ^ n4677 ^ n4675 ;
  assign n4683 = ~n4646 & n4682 ;
  assign n4684 = ( x78 & n957 ) | ( x78 & n2238 ) | ( n957 & n2238 ) ;
  assign n4690 = n1694 ^ n624 ^ x154 ;
  assign n4691 = ( n2230 & ~n2402 ) | ( n2230 & n3734 ) | ( ~n2402 & n3734 ) ;
  assign n4692 = ( n969 & n4690 ) | ( n969 & n4691 ) | ( n4690 & n4691 ) ;
  assign n4693 = ( x137 & n3420 ) | ( x137 & n4692 ) | ( n3420 & n4692 ) ;
  assign n4694 = n4693 ^ n1744 ^ n750 ;
  assign n4685 = ( n591 & n2213 ) | ( n591 & n2337 ) | ( n2213 & n2337 ) ;
  assign n4686 = n3502 ^ n1314 ^ n325 ;
  assign n4687 = n4686 ^ n454 ^ 1'b0 ;
  assign n4688 = n4687 ^ n736 ^ 1'b0 ;
  assign n4689 = ( n2564 & n4685 ) | ( n2564 & ~n4688 ) | ( n4685 & ~n4688 ) ;
  assign n4695 = n4694 ^ n4689 ^ x211 ;
  assign n4696 = ( n850 & ~n2743 ) | ( n850 & n3735 ) | ( ~n2743 & n3735 ) ;
  assign n4697 = n4696 ^ n4302 ^ x203 ;
  assign n4698 = n4299 ^ n3924 ^ n2796 ;
  assign n4699 = n4698 ^ n4658 ^ n2038 ;
  assign n4700 = ( n493 & n729 ) | ( n493 & ~n1053 ) | ( n729 & ~n1053 ) ;
  assign n4701 = n1297 ^ n970 ^ n439 ;
  assign n4702 = ( n2705 & n4700 ) | ( n2705 & n4701 ) | ( n4700 & n4701 ) ;
  assign n4703 = ( n1221 & n2844 ) | ( n1221 & ~n4702 ) | ( n2844 & ~n4702 ) ;
  assign n4710 = n3158 ^ n2957 ^ n1312 ;
  assign n4704 = n649 ^ n399 ^ x246 ;
  assign n4705 = x90 ^ x1 ^ 1'b0 ;
  assign n4706 = x3 & n4705 ;
  assign n4707 = ( x179 & ~n939 ) | ( x179 & n4706 ) | ( ~n939 & n4706 ) ;
  assign n4708 = n4707 ^ n3541 ^ n2890 ;
  assign n4709 = ( n2223 & n4704 ) | ( n2223 & n4708 ) | ( n4704 & n4708 ) ;
  assign n4711 = n4710 ^ n4709 ^ x97 ;
  assign n4712 = ( ~n2239 & n2639 ) | ( ~n2239 & n3584 ) | ( n2639 & n3584 ) ;
  assign n4713 = n4712 ^ n3277 ^ x20 ;
  assign n4714 = n3223 ^ n2935 ^ n1945 ;
  assign n4715 = ( n1496 & ~n1757 ) | ( n1496 & n2800 ) | ( ~n1757 & n2800 ) ;
  assign n4716 = x227 & ~n2127 ;
  assign n4717 = n1182 & n4716 ;
  assign n4718 = n4717 ^ n2760 ^ n975 ;
  assign n4719 = n3121 & n4718 ;
  assign n4720 = n4719 ^ n2694 ^ 1'b0 ;
  assign n4721 = ( ~n4714 & n4715 ) | ( ~n4714 & n4720 ) | ( n4715 & n4720 ) ;
  assign n4722 = n2710 ^ n863 ^ 1'b0 ;
  assign n4723 = n4722 ^ n2521 ^ 1'b0 ;
  assign n4735 = ( x104 & ~n1837 ) | ( x104 & n3319 ) | ( ~n1837 & n3319 ) ;
  assign n4724 = n1547 ^ n635 ^ n538 ;
  assign n4725 = ( x170 & n792 ) | ( x170 & ~n949 ) | ( n792 & ~n949 ) ;
  assign n4727 = ( x95 & ~n428 ) | ( x95 & n755 ) | ( ~n428 & n755 ) ;
  assign n4728 = ( x16 & n1590 ) | ( x16 & ~n4727 ) | ( n1590 & ~n4727 ) ;
  assign n4726 = n2410 ^ n2259 ^ 1'b0 ;
  assign n4729 = n4728 ^ n4726 ^ n2041 ;
  assign n4730 = n4725 & n4729 ;
  assign n4731 = n1440 & n4730 ;
  assign n4732 = n3901 ^ n3167 ^ n1955 ;
  assign n4733 = n4732 ^ n3527 ^ n1689 ;
  assign n4734 = ( n4724 & n4731 ) | ( n4724 & ~n4733 ) | ( n4731 & ~n4733 ) ;
  assign n4736 = n4735 ^ n4734 ^ n2641 ;
  assign n4738 = n2564 ^ n1280 ^ n893 ;
  assign n4737 = ( x147 & n3230 ) | ( x147 & n4117 ) | ( n3230 & n4117 ) ;
  assign n4739 = n4738 ^ n4737 ^ n1740 ;
  assign n4740 = n4739 ^ n1981 ^ n544 ;
  assign n4741 = ( n424 & ~n1277 ) | ( n424 & n2564 ) | ( ~n1277 & n2564 ) ;
  assign n4742 = ( n2583 & n4740 ) | ( n2583 & n4741 ) | ( n4740 & n4741 ) ;
  assign n4750 = ( n724 & n2231 ) | ( n724 & ~n3293 ) | ( n2231 & ~n3293 ) ;
  assign n4749 = n3463 ^ n1892 ^ n1420 ;
  assign n4751 = n4750 ^ n4749 ^ n3194 ;
  assign n4747 = n971 ^ x157 ^ 1'b0 ;
  assign n4745 = n3488 ^ x189 ^ x94 ;
  assign n4746 = ( n1285 & n1641 ) | ( n1285 & n4745 ) | ( n1641 & n4745 ) ;
  assign n4743 = n2222 ^ n939 ^ n303 ;
  assign n4744 = n2198 | n4743 ;
  assign n4748 = n4747 ^ n4746 ^ n4744 ;
  assign n4752 = n4751 ^ n4748 ^ n3723 ;
  assign n4753 = n2888 & n4752 ;
  assign n4754 = n4742 & n4753 ;
  assign n4755 = ( x200 & ~x251 ) | ( x200 & n1543 ) | ( ~x251 & n1543 ) ;
  assign n4756 = n4113 ^ n1661 ^ 1'b0 ;
  assign n4757 = n4755 & ~n4756 ;
  assign n4758 = ( n1363 & n3071 ) | ( n1363 & ~n3103 ) | ( n3071 & ~n3103 ) ;
  assign n4759 = n4758 ^ n1536 ^ x108 ;
  assign n4760 = ( n2756 & n4757 ) | ( n2756 & ~n4759 ) | ( n4757 & ~n4759 ) ;
  assign n4761 = ( n1561 & n1950 ) | ( n1561 & ~n3508 ) | ( n1950 & ~n3508 ) ;
  assign n4762 = ( n1456 & n3466 ) | ( n1456 & ~n4761 ) | ( n3466 & ~n4761 ) ;
  assign n4763 = n347 & n3103 ;
  assign n4764 = n579 & n4763 ;
  assign n4765 = n4764 ^ n2893 ^ n1652 ;
  assign n4766 = n4248 & n4765 ;
  assign n4767 = ~n3683 & n4766 ;
  assign n4775 = ( x83 & n2204 ) | ( x83 & ~n4599 ) | ( n2204 & ~n4599 ) ;
  assign n4776 = n4775 ^ n745 ^ x128 ;
  assign n4773 = n1398 & n1509 ;
  assign n4774 = n1673 & n4773 ;
  assign n4770 = ( n481 & n1710 ) | ( n481 & ~n3224 ) | ( n1710 & ~n3224 ) ;
  assign n4771 = n4770 ^ n2690 ^ n2184 ;
  assign n4768 = n2065 ^ n1665 ^ n833 ;
  assign n4769 = ( ~x59 & n3110 ) | ( ~x59 & n4768 ) | ( n3110 & n4768 ) ;
  assign n4772 = n4771 ^ n4769 ^ n3439 ;
  assign n4777 = n4776 ^ n4774 ^ n4772 ;
  assign n4780 = ( n464 & ~n648 ) | ( n464 & n1910 ) | ( ~n648 & n1910 ) ;
  assign n4778 = ( n481 & n1317 ) | ( n481 & ~n1794 ) | ( n1317 & ~n1794 ) ;
  assign n4779 = n4778 ^ n1936 ^ n1840 ;
  assign n4781 = n4780 ^ n4779 ^ n258 ;
  assign n4782 = ~x119 & n407 ;
  assign n4783 = ( ~n699 & n3172 ) | ( ~n699 & n4782 ) | ( n3172 & n4782 ) ;
  assign n4784 = n4783 ^ n2997 ^ 1'b0 ;
  assign n4785 = ( n596 & n1276 ) | ( n596 & ~n4784 ) | ( n1276 & ~n4784 ) ;
  assign n4795 = ( ~n738 & n1219 ) | ( ~n738 & n2795 ) | ( n1219 & n2795 ) ;
  assign n4792 = n1969 ^ n1308 ^ x247 ;
  assign n4793 = ( n384 & n1464 ) | ( n384 & n4792 ) | ( n1464 & n4792 ) ;
  assign n4794 = n4793 ^ n1858 ^ n1670 ;
  assign n4791 = n3634 ^ n3132 ^ n1928 ;
  assign n4796 = n4795 ^ n4794 ^ n4791 ;
  assign n4786 = n4700 ^ n2743 ^ n1545 ;
  assign n4787 = ( n2097 & n2438 ) | ( n2097 & ~n4786 ) | ( n2438 & ~n4786 ) ;
  assign n4788 = ( n671 & ~n3292 ) | ( n671 & n4787 ) | ( ~n3292 & n4787 ) ;
  assign n4789 = n4788 ^ n2768 ^ n1824 ;
  assign n4790 = x121 & n4789 ;
  assign n4797 = n4796 ^ n4790 ^ 1'b0 ;
  assign n4798 = ~n1575 & n4226 ;
  assign n4799 = ( n475 & ~n3785 ) | ( n475 & n4798 ) | ( ~n3785 & n4798 ) ;
  assign n4800 = n2784 ^ n265 ^ 1'b0 ;
  assign n4801 = n535 & ~n4800 ;
  assign n4802 = n4801 ^ n3089 ^ n664 ;
  assign n4803 = n4358 ^ n520 ^ 1'b0 ;
  assign n4804 = ~n4802 & n4803 ;
  assign n4805 = n4804 ^ n2586 ^ n2099 ;
  assign n4806 = n4805 ^ n2510 ^ n378 ;
  assign n4818 = n1151 & n2346 ;
  assign n4819 = ~x167 & n4818 ;
  assign n4816 = n398 & ~n2303 ;
  assign n4815 = n1119 & ~n1172 ;
  assign n4817 = n4816 ^ n4815 ^ 1'b0 ;
  assign n4820 = n4819 ^ n4817 ^ n1199 ;
  assign n4811 = n3467 ^ n1904 ^ n1359 ;
  assign n4808 = n1930 & ~n4293 ;
  assign n4809 = n1745 & n4808 ;
  assign n4807 = n4747 ^ n3792 ^ n1545 ;
  assign n4810 = n4809 ^ n4807 ^ n2362 ;
  assign n4812 = n4811 ^ n4810 ^ n2116 ;
  assign n4813 = x167 & ~n4812 ;
  assign n4814 = ~x240 & n4813 ;
  assign n4821 = n4820 ^ n4814 ^ 1'b0 ;
  assign n4822 = n2714 & ~n4222 ;
  assign n4823 = ~n3007 & n4822 ;
  assign n4824 = n4301 ^ n3613 ^ n2351 ;
  assign n4825 = ( n1646 & ~n4823 ) | ( n1646 & n4824 ) | ( ~n4823 & n4824 ) ;
  assign n4826 = ( ~x10 & n3476 ) | ( ~x10 & n4825 ) | ( n3476 & n4825 ) ;
  assign n4827 = ( n989 & ~n3879 ) | ( n989 & n4826 ) | ( ~n3879 & n4826 ) ;
  assign n4828 = n4027 ^ n3829 ^ n1320 ;
  assign n4829 = ( n650 & n3889 ) | ( n650 & ~n4828 ) | ( n3889 & ~n4828 ) ;
  assign n4830 = n2309 ^ n482 ^ 1'b0 ;
  assign n4831 = ( n297 & n1093 ) | ( n297 & ~n4830 ) | ( n1093 & ~n4830 ) ;
  assign n4832 = ( n399 & n751 ) | ( n399 & ~n1822 ) | ( n751 & ~n1822 ) ;
  assign n4833 = ( n1740 & n4831 ) | ( n1740 & n4832 ) | ( n4831 & n4832 ) ;
  assign n4834 = n1205 ^ n969 ^ n642 ;
  assign n4835 = ( ~n2196 & n2206 ) | ( ~n2196 & n2735 ) | ( n2206 & n2735 ) ;
  assign n4836 = ( ~n3488 & n4834 ) | ( ~n3488 & n4835 ) | ( n4834 & n4835 ) ;
  assign n4837 = ( n1041 & ~n3172 ) | ( n1041 & n4836 ) | ( ~n3172 & n4836 ) ;
  assign n4838 = ~n4833 & n4837 ;
  assign n4839 = n4838 ^ n1101 ^ 1'b0 ;
  assign n4840 = ( ~n2730 & n4829 ) | ( ~n2730 & n4839 ) | ( n4829 & n4839 ) ;
  assign n4841 = n3374 ^ x235 ^ 1'b0 ;
  assign n4842 = ~n301 & n4841 ;
  assign n4843 = ( n3071 & n4606 ) | ( n3071 & n4842 ) | ( n4606 & n4842 ) ;
  assign n4844 = ( n4180 & n4840 ) | ( n4180 & ~n4843 ) | ( n4840 & ~n4843 ) ;
  assign n4845 = ( n1397 & ~n2795 ) | ( n1397 & n3082 ) | ( ~n2795 & n3082 ) ;
  assign n4846 = n3729 ^ n2765 ^ n931 ;
  assign n4847 = n4846 ^ n448 ^ 1'b0 ;
  assign n4848 = n4847 ^ n4430 ^ n2415 ;
  assign n4849 = ( n1846 & n3025 ) | ( n1846 & ~n4848 ) | ( n3025 & ~n4848 ) ;
  assign n4850 = n1869 ^ n1762 ^ n904 ;
  assign n4851 = n4850 ^ n4451 ^ n3367 ;
  assign n4852 = n3541 ^ n1795 ^ n1304 ;
  assign n4853 = n4852 ^ n4802 ^ 1'b0 ;
  assign n4854 = n4851 & n4853 ;
  assign n4868 = ~n971 & n1154 ;
  assign n4869 = n4868 ^ n3381 ^ 1'b0 ;
  assign n4870 = n4869 ^ x31 ^ 1'b0 ;
  assign n4871 = ~n1269 & n4870 ;
  assign n4872 = n4871 ^ n4567 ^ n2146 ;
  assign n4855 = n3901 ^ n2402 ^ x135 ;
  assign n4856 = ( ~n1078 & n2711 ) | ( ~n1078 & n4855 ) | ( n2711 & n4855 ) ;
  assign n4857 = n2444 & n4856 ;
  assign n4858 = n4857 ^ n873 ^ 1'b0 ;
  assign n4859 = ( n4434 & n4727 ) | ( n4434 & n4858 ) | ( n4727 & n4858 ) ;
  assign n4863 = n502 | n610 ;
  assign n4864 = n4863 ^ n4271 ^ x29 ;
  assign n4860 = ( ~x109 & n2936 ) | ( ~x109 & n4580 ) | ( n2936 & n4580 ) ;
  assign n4861 = ( n1002 & n1754 ) | ( n1002 & n3782 ) | ( n1754 & n3782 ) ;
  assign n4862 = ( n2116 & n4860 ) | ( n2116 & ~n4861 ) | ( n4860 & ~n4861 ) ;
  assign n4865 = n4864 ^ n4862 ^ n2340 ;
  assign n4866 = n4859 & ~n4865 ;
  assign n4867 = ~n539 & n4866 ;
  assign n4873 = n4872 ^ n4867 ^ n4449 ;
  assign n4874 = n3103 ^ n1132 ^ n895 ;
  assign n4875 = ( x120 & n1599 ) | ( x120 & n4874 ) | ( n1599 & n4874 ) ;
  assign n4876 = ( n1383 & n2125 ) | ( n1383 & n3719 ) | ( n2125 & n3719 ) ;
  assign n4877 = n1720 ^ n1213 ^ n635 ;
  assign n4878 = ( n4875 & n4876 ) | ( n4875 & ~n4877 ) | ( n4876 & ~n4877 ) ;
  assign n4879 = ( n305 & ~n571 ) | ( n305 & n794 ) | ( ~n571 & n794 ) ;
  assign n4880 = ( x39 & ~n2499 ) | ( x39 & n4879 ) | ( ~n2499 & n4879 ) ;
  assign n4881 = n4880 ^ n2815 ^ 1'b0 ;
  assign n4882 = n4878 & n4881 ;
  assign n4883 = n3118 | n4882 ;
  assign n4884 = ( x60 & n694 ) | ( x60 & ~n2539 ) | ( n694 & ~n2539 ) ;
  assign n4885 = ( n1150 & n1814 ) | ( n1150 & n3560 ) | ( n1814 & n3560 ) ;
  assign n4886 = ( n4712 & n4884 ) | ( n4712 & n4885 ) | ( n4884 & n4885 ) ;
  assign n4887 = n4886 ^ n3320 ^ n1666 ;
  assign n4888 = n4887 ^ n1261 ^ 1'b0 ;
  assign n4890 = n3244 ^ n3108 ^ n1844 ;
  assign n4891 = ( n304 & n2302 ) | ( n304 & ~n4890 ) | ( n2302 & ~n4890 ) ;
  assign n4889 = n1588 ^ n879 ^ n286 ;
  assign n4892 = n4891 ^ n4889 ^ x51 ;
  assign n4893 = n4892 ^ n2062 ^ n990 ;
  assign n4894 = n2152 | n4893 ;
  assign n4895 = n2193 ^ x243 ^ 1'b0 ;
  assign n4896 = ( n617 & ~n4502 ) | ( n617 & n4895 ) | ( ~n4502 & n4895 ) ;
  assign n4897 = n937 ^ x239 ^ x183 ;
  assign n4898 = n1543 & ~n4897 ;
  assign n4899 = n2759 & n4898 ;
  assign n4900 = n3892 | n4899 ;
  assign n4901 = ( n1982 & n4896 ) | ( n1982 & ~n4900 ) | ( n4896 & ~n4900 ) ;
  assign n4907 = n3151 ^ n1260 ^ n368 ;
  assign n4908 = n4907 ^ n4794 ^ n1983 ;
  assign n4904 = ( n1437 & ~n2677 ) | ( n1437 & n2877 ) | ( ~n2677 & n2877 ) ;
  assign n4902 = n925 ^ n905 ^ n784 ;
  assign n4903 = ( ~n1898 & n4876 ) | ( ~n1898 & n4902 ) | ( n4876 & n4902 ) ;
  assign n4905 = n4904 ^ n4903 ^ n4385 ;
  assign n4906 = n706 | n4905 ;
  assign n4909 = n4908 ^ n4906 ^ 1'b0 ;
  assign n4910 = ( ~n421 & n2914 ) | ( ~n421 & n4909 ) | ( n2914 & n4909 ) ;
  assign n4911 = ( n940 & n2879 ) | ( n940 & ~n4565 ) | ( n2879 & ~n4565 ) ;
  assign n4912 = ( n1181 & n4910 ) | ( n1181 & n4911 ) | ( n4910 & n4911 ) ;
  assign n4913 = ~n413 & n3061 ;
  assign n4914 = n3791 ^ n682 ^ n674 ;
  assign n4915 = n4417 ^ n2669 ^ x193 ;
  assign n4916 = n2532 & n4915 ;
  assign n4917 = n4350 ^ n3789 ^ n1409 ;
  assign n4918 = n4917 ^ n2277 ^ n925 ;
  assign n4919 = ( ~n1289 & n4916 ) | ( ~n1289 & n4918 ) | ( n4916 & n4918 ) ;
  assign n4920 = n4919 ^ n416 ^ 1'b0 ;
  assign n4921 = ( ~n4913 & n4914 ) | ( ~n4913 & n4920 ) | ( n4914 & n4920 ) ;
  assign n4924 = ( x61 & n703 ) | ( x61 & ~n1180 ) | ( n703 & ~n1180 ) ;
  assign n4925 = n4924 ^ n4578 ^ n294 ;
  assign n4926 = n4925 ^ n4307 ^ n3656 ;
  assign n4922 = n3117 ^ n1435 ^ n617 ;
  assign n4923 = ( ~n579 & n719 ) | ( ~n579 & n4922 ) | ( n719 & n4922 ) ;
  assign n4927 = n4926 ^ n4923 ^ x13 ;
  assign n4935 = ( ~x16 & n1003 ) | ( ~x16 & n2555 ) | ( n1003 & n2555 ) ;
  assign n4936 = n4935 ^ n2868 ^ n365 ;
  assign n4937 = n4936 ^ n2323 ^ n1352 ;
  assign n4932 = ( n843 & ~n893 ) | ( n843 & n1582 ) | ( ~n893 & n1582 ) ;
  assign n4928 = n397 ^ x94 ^ 1'b0 ;
  assign n4929 = ( n572 & ~n4566 ) | ( n572 & n4928 ) | ( ~n4566 & n4928 ) ;
  assign n4930 = ( n1096 & ~n1489 ) | ( n1096 & n4929 ) | ( ~n1489 & n4929 ) ;
  assign n4931 = n4930 ^ n2045 ^ x113 ;
  assign n4933 = n4932 ^ n4931 ^ n2615 ;
  assign n4934 = n4933 ^ n1048 ^ n1013 ;
  assign n4938 = n4937 ^ n4934 ^ n3855 ;
  assign n4940 = ( n442 & ~n889 ) | ( n442 & n4678 ) | ( ~n889 & n4678 ) ;
  assign n4939 = n2827 ^ n1533 ^ x179 ;
  assign n4941 = n4940 ^ n4939 ^ n1979 ;
  assign n4942 = n1448 & ~n4941 ;
  assign n4956 = n3496 ^ n2328 ^ n2233 ;
  assign n4955 = ( ~n830 & n1552 ) | ( ~n830 & n4018 ) | ( n1552 & n4018 ) ;
  assign n4944 = n1129 ^ n991 ^ n378 ;
  assign n4943 = n1552 ^ n933 ^ n693 ;
  assign n4945 = n4944 ^ n4943 ^ n656 ;
  assign n4946 = n4945 ^ n4643 ^ n2363 ;
  assign n4948 = n3541 ^ n1532 ^ n777 ;
  assign n4947 = n2018 ^ n1187 ^ x40 ;
  assign n4949 = n4948 ^ n4947 ^ n4147 ;
  assign n4950 = ( n569 & n1734 ) | ( n569 & ~n3749 ) | ( n1734 & ~n3749 ) ;
  assign n4951 = n1843 | n4950 ;
  assign n4952 = n4949 & ~n4951 ;
  assign n4953 = n4952 ^ n2969 ^ 1'b0 ;
  assign n4954 = ( n1921 & n4946 ) | ( n1921 & n4953 ) | ( n4946 & n4953 ) ;
  assign n4957 = n4956 ^ n4955 ^ n4954 ;
  assign n4958 = ( ~n1452 & n1710 ) | ( ~n1452 & n3950 ) | ( n1710 & n3950 ) ;
  assign n4959 = n3815 ^ n2159 ^ x196 ;
  assign n4960 = n3432 & n4959 ;
  assign n4961 = n4960 ^ n2945 ^ 1'b0 ;
  assign n4962 = n4961 ^ n414 ^ 1'b0 ;
  assign n4963 = ( n2376 & n4958 ) | ( n2376 & n4962 ) | ( n4958 & n4962 ) ;
  assign n4964 = n4835 ^ n2300 ^ n2154 ;
  assign n4965 = n3284 ^ n2835 ^ n2485 ;
  assign n4966 = n3883 | n4965 ;
  assign n4967 = n4966 ^ n4702 ^ 1'b0 ;
  assign n4968 = ( n1153 & n4964 ) | ( n1153 & ~n4967 ) | ( n4964 & ~n4967 ) ;
  assign n4970 = ( ~n416 & n2257 ) | ( ~n416 & n3089 ) | ( n2257 & n3089 ) ;
  assign n4971 = n4970 ^ n993 ^ n971 ;
  assign n4972 = n4971 ^ n268 ^ 1'b0 ;
  assign n4973 = n1506 & ~n4972 ;
  assign n4969 = ( x135 & n1967 ) | ( x135 & n2089 ) | ( n1967 & n2089 ) ;
  assign n4974 = n4973 ^ n4969 ^ n2190 ;
  assign n4975 = n4974 ^ n2644 ^ n1542 ;
  assign n4992 = n3259 ^ n2033 ^ x221 ;
  assign n4993 = n2621 ^ n1591 ^ n1500 ;
  assign n4994 = ~n4992 & n4993 ;
  assign n4988 = ( ~n295 & n1108 ) | ( ~n295 & n3007 ) | ( n1108 & n3007 ) ;
  assign n4989 = n4988 ^ n2238 ^ n1306 ;
  assign n4990 = n4989 ^ n3225 ^ n2197 ;
  assign n4987 = n2731 ^ n2157 ^ n1943 ;
  assign n4991 = n4990 ^ n4987 ^ 1'b0 ;
  assign n4995 = n4994 ^ n4991 ^ n3043 ;
  assign n4976 = ~x239 & n1288 ;
  assign n4977 = ( n256 & n1071 ) | ( n256 & n2233 ) | ( n1071 & n2233 ) ;
  assign n4978 = ( ~n437 & n4545 ) | ( ~n437 & n4977 ) | ( n4545 & n4977 ) ;
  assign n4979 = n4176 ^ n3558 ^ n1922 ;
  assign n4980 = n4979 ^ n2269 ^ n1864 ;
  assign n4981 = n4980 ^ n2093 ^ n538 ;
  assign n4982 = n1057 & n1862 ;
  assign n4983 = n4982 ^ n2875 ^ 1'b0 ;
  assign n4984 = n4983 ^ n2980 ^ n1662 ;
  assign n4985 = ( n4978 & n4981 ) | ( n4978 & ~n4984 ) | ( n4981 & ~n4984 ) ;
  assign n4986 = ( n2009 & n4976 ) | ( n2009 & n4985 ) | ( n4976 & n4985 ) ;
  assign n4996 = n4995 ^ n4986 ^ n3415 ;
  assign n4997 = n859 ^ n391 ^ n332 ;
  assign n4998 = ( ~x80 & x116 ) | ( ~x80 & n1086 ) | ( x116 & n1086 ) ;
  assign n4999 = ( ~x244 & n3856 ) | ( ~x244 & n4040 ) | ( n3856 & n4040 ) ;
  assign n5000 = ( n4997 & ~n4998 ) | ( n4997 & n4999 ) | ( ~n4998 & n4999 ) ;
  assign n5001 = ( n1358 & n2284 ) | ( n1358 & ~n5000 ) | ( n2284 & ~n5000 ) ;
  assign n5002 = n3384 ^ n2248 ^ 1'b0 ;
  assign n5003 = n5002 ^ n1787 ^ 1'b0 ;
  assign n5004 = n4971 & n5003 ;
  assign n5009 = n1326 ^ n368 ^ n294 ;
  assign n5005 = x247 ^ x213 ^ x1 ;
  assign n5006 = n1902 ^ n1104 ^ x110 ;
  assign n5007 = n5006 ^ n3069 ^ x38 ;
  assign n5008 = ( n3255 & n5005 ) | ( n3255 & n5007 ) | ( n5005 & n5007 ) ;
  assign n5010 = n5009 ^ n5008 ^ n428 ;
  assign n5011 = n5010 ^ n2394 ^ n2044 ;
  assign n5012 = n5004 & n5011 ;
  assign n5013 = n1213 ^ n914 ^ n693 ;
  assign n5014 = n5013 ^ n2603 ^ n2218 ;
  assign n5015 = n5014 ^ n4769 ^ n1194 ;
  assign n5033 = ( n1086 & n2642 ) | ( n1086 & ~n2656 ) | ( n2642 & ~n2656 ) ;
  assign n5034 = n3320 ^ n1467 ^ 1'b0 ;
  assign n5035 = ~n5033 & n5034 ;
  assign n5036 = ( n2031 & ~n2229 ) | ( n2031 & n5035 ) | ( ~n2229 & n5035 ) ;
  assign n5026 = n2705 ^ n1204 ^ n813 ;
  assign n5027 = n4560 ^ n2268 ^ n2169 ;
  assign n5028 = n5027 ^ n955 ^ n467 ;
  assign n5029 = n5028 ^ n2411 ^ n2351 ;
  assign n5030 = n5029 ^ n4663 ^ x31 ;
  assign n5031 = n5030 ^ n2176 ^ 1'b0 ;
  assign n5032 = n5026 & n5031 ;
  assign n5023 = n1653 ^ n1450 ^ n396 ;
  assign n5022 = ( n431 & n1684 ) | ( n431 & n2463 ) | ( n1684 & n2463 ) ;
  assign n5024 = n5023 ^ n5022 ^ n2110 ;
  assign n5019 = ( x109 & n801 ) | ( x109 & ~n4582 ) | ( n801 & ~n4582 ) ;
  assign n5016 = n1370 ^ n487 ^ 1'b0 ;
  assign n5017 = x12 & n5016 ;
  assign n5018 = n2658 & n5017 ;
  assign n5020 = n5019 ^ n5018 ^ 1'b0 ;
  assign n5021 = n5020 ^ n1930 ^ n1250 ;
  assign n5025 = n5024 ^ n5021 ^ n1204 ;
  assign n5037 = n5036 ^ n5032 ^ n5025 ;
  assign n5038 = n1304 ^ n995 ^ 1'b0 ;
  assign n5039 = ( x0 & ~n1114 ) | ( x0 & n5038 ) | ( ~n1114 & n5038 ) ;
  assign n5040 = n3819 ^ n2328 ^ n2241 ;
  assign n5041 = ( ~n4180 & n5039 ) | ( ~n4180 & n5040 ) | ( n5039 & n5040 ) ;
  assign n5042 = ( ~x99 & n2481 ) | ( ~x99 & n5041 ) | ( n2481 & n5041 ) ;
  assign n5061 = n4436 ^ n2011 ^ x192 ;
  assign n5062 = n1345 & n5061 ;
  assign n5063 = n2081 & n5062 ;
  assign n5057 = n1647 ^ n1572 ^ n828 ;
  assign n5058 = ( ~n2314 & n3116 ) | ( ~n2314 & n5057 ) | ( n3116 & n5057 ) ;
  assign n5043 = n1320 & ~n4786 ;
  assign n5044 = n5043 ^ x201 ^ 1'b0 ;
  assign n5045 = ( x222 & ~n1850 ) | ( x222 & n2505 ) | ( ~n1850 & n2505 ) ;
  assign n5046 = n793 | n5040 ;
  assign n5047 = n1440 & ~n5046 ;
  assign n5048 = n5047 ^ n2440 ^ n578 ;
  assign n5049 = n5045 | n5048 ;
  assign n5050 = n5044 & ~n5049 ;
  assign n5051 = ( n326 & ~n446 ) | ( n326 & n812 ) | ( ~n446 & n812 ) ;
  assign n5052 = n325 & ~n5051 ;
  assign n5053 = ~n533 & n5052 ;
  assign n5054 = n2899 & ~n5053 ;
  assign n5055 = n5054 ^ n1601 ^ 1'b0 ;
  assign n5056 = ( n2891 & ~n5050 ) | ( n2891 & n5055 ) | ( ~n5050 & n5055 ) ;
  assign n5059 = n5058 ^ n5056 ^ 1'b0 ;
  assign n5060 = n801 | n5059 ;
  assign n5064 = n5063 ^ n5060 ^ n651 ;
  assign n5065 = ( n894 & n967 ) | ( n894 & ~n4400 ) | ( n967 & ~n4400 ) ;
  assign n5066 = n5065 ^ n2567 ^ n950 ;
  assign n5067 = n5066 ^ n1836 ^ 1'b0 ;
  assign n5068 = ( n581 & n5064 ) | ( n581 & ~n5067 ) | ( n5064 & ~n5067 ) ;
  assign n5075 = n773 ^ x192 ^ 1'b0 ;
  assign n5072 = n2360 ^ n752 ^ n384 ;
  assign n5073 = ( n2427 & ~n2818 ) | ( n2427 & n5072 ) | ( ~n2818 & n5072 ) ;
  assign n5074 = n5073 ^ n2562 ^ x206 ;
  assign n5069 = n2701 ^ n2383 ^ n1911 ;
  assign n5070 = n5069 ^ n737 ^ x243 ;
  assign n5071 = ( x72 & ~n4304 ) | ( x72 & n5070 ) | ( ~n4304 & n5070 ) ;
  assign n5076 = n5075 ^ n5074 ^ n5071 ;
  assign n5077 = n5076 ^ n5069 ^ n2101 ;
  assign n5078 = n3146 ^ n1523 ^ n431 ;
  assign n5079 = n3783 & ~n5078 ;
  assign n5080 = n2999 ^ n587 ^ 1'b0 ;
  assign n5081 = n1647 & ~n5080 ;
  assign n5082 = n3598 ^ n2152 ^ n530 ;
  assign n5083 = n5082 ^ n1682 ^ n1420 ;
  assign n5084 = n698 ^ n663 ^ 1'b0 ;
  assign n5085 = n5084 ^ n1514 ^ x169 ;
  assign n5086 = ( n4244 & n4949 ) | ( n4244 & n5085 ) | ( n4949 & n5085 ) ;
  assign n5087 = ( n1292 & n5083 ) | ( n1292 & n5086 ) | ( n5083 & n5086 ) ;
  assign n5088 = n5087 ^ n4619 ^ n1410 ;
  assign n5089 = ( x83 & ~n1016 ) | ( x83 & n3433 ) | ( ~n1016 & n3433 ) ;
  assign n5096 = n1795 ^ x243 ^ x116 ;
  assign n5093 = ( n943 & n2287 ) | ( n943 & ~n2381 ) | ( n2287 & ~n2381 ) ;
  assign n5094 = n5093 ^ n3248 ^ x72 ;
  assign n5090 = n3541 ^ n2389 ^ n350 ;
  assign n5091 = n5090 ^ n4750 ^ n4545 ;
  assign n5092 = n4595 & ~n5091 ;
  assign n5095 = n5094 ^ n5092 ^ 1'b0 ;
  assign n5097 = n5096 ^ n5095 ^ n4445 ;
  assign n5098 = n5097 ^ n2507 ^ n1602 ;
  assign n5099 = n5089 & ~n5098 ;
  assign n5110 = n1328 ^ n1123 ^ n262 ;
  assign n5100 = x67 & n1810 ;
  assign n5101 = ~x236 & n5100 ;
  assign n5102 = n5101 ^ n3734 ^ 1'b0 ;
  assign n5103 = n346 | n5102 ;
  assign n5104 = n2416 ^ n1311 ^ x214 ;
  assign n5105 = ( ~n2373 & n5103 ) | ( ~n2373 & n5104 ) | ( n5103 & n5104 ) ;
  assign n5106 = ( x211 & n2483 ) | ( x211 & n3677 ) | ( n2483 & n3677 ) ;
  assign n5107 = ( n847 & ~n1086 ) | ( n847 & n5106 ) | ( ~n1086 & n5106 ) ;
  assign n5108 = n5107 ^ n4825 ^ 1'b0 ;
  assign n5109 = ( n4163 & n5105 ) | ( n4163 & ~n5108 ) | ( n5105 & ~n5108 ) ;
  assign n5111 = n5110 ^ n5109 ^ n3899 ;
  assign n5118 = n4129 ^ n2686 ^ 1'b0 ;
  assign n5115 = ( ~n1435 & n2210 ) | ( ~n1435 & n2492 ) | ( n2210 & n2492 ) ;
  assign n5112 = n1018 & ~n1919 ;
  assign n5113 = ~n5028 & n5112 ;
  assign n5114 = n539 & ~n5113 ;
  assign n5116 = n5115 ^ n5114 ^ 1'b0 ;
  assign n5117 = ( n431 & ~n1740 ) | ( n431 & n5116 ) | ( ~n1740 & n5116 ) ;
  assign n5119 = n5118 ^ n5117 ^ 1'b0 ;
  assign n5120 = x0 & n5119 ;
  assign n5121 = n1223 ^ n1098 ^ n997 ;
  assign n5122 = n5121 ^ n1404 ^ n469 ;
  assign n5123 = n2600 ^ n1590 ^ 1'b0 ;
  assign n5124 = n5123 ^ n3620 ^ n669 ;
  assign n5125 = ( ~n1937 & n5122 ) | ( ~n1937 & n5124 ) | ( n5122 & n5124 ) ;
  assign n5126 = ( n1842 & ~n3071 ) | ( n1842 & n4022 ) | ( ~n3071 & n4022 ) ;
  assign n5127 = n4090 ^ n2058 ^ 1'b0 ;
  assign n5128 = n5126 & ~n5127 ;
  assign n5129 = n5128 ^ n4441 ^ n3486 ;
  assign n5130 = n3503 ^ n1167 ^ x118 ;
  assign n5131 = ( n308 & ~n815 ) | ( n308 & n5130 ) | ( ~n815 & n5130 ) ;
  assign n5132 = n4834 & n5131 ;
  assign n5133 = ( ~n1952 & n4509 ) | ( ~n1952 & n5132 ) | ( n4509 & n5132 ) ;
  assign n5134 = n298 | n867 ;
  assign n5135 = ( n1981 & n3451 ) | ( n1981 & ~n4956 ) | ( n3451 & ~n4956 ) ;
  assign n5136 = ( ~n804 & n5134 ) | ( ~n804 & n5135 ) | ( n5134 & n5135 ) ;
  assign n5137 = n2559 | n5136 ;
  assign n5138 = n5137 ^ n2933 ^ 1'b0 ;
  assign n5148 = ( n794 & ~n1471 ) | ( n794 & n3108 ) | ( ~n1471 & n3108 ) ;
  assign n5149 = n5148 ^ n4928 ^ n1491 ;
  assign n5143 = ( n1304 & n2506 ) | ( n1304 & ~n2827 ) | ( n2506 & ~n2827 ) ;
  assign n5144 = n2989 | n5143 ;
  assign n5145 = n3746 & ~n5144 ;
  assign n5146 = ( n929 & ~n4050 ) | ( n929 & n5145 ) | ( ~n4050 & n5145 ) ;
  assign n5147 = n5146 ^ n3635 ^ n3210 ;
  assign n5139 = n2084 & ~n3317 ;
  assign n5140 = n5139 ^ n1682 ^ 1'b0 ;
  assign n5141 = ~n814 & n5140 ;
  assign n5142 = ( n2100 & n4423 ) | ( n2100 & ~n5141 ) | ( n4423 & ~n5141 ) ;
  assign n5150 = n5149 ^ n5147 ^ n5142 ;
  assign n5151 = n4380 ^ n3878 ^ n3268 ;
  assign n5152 = ( n3685 & ~n4657 ) | ( n3685 & n5151 ) | ( ~n4657 & n5151 ) ;
  assign n5153 = n1761 & ~n5152 ;
  assign n5154 = n5150 & n5153 ;
  assign n5155 = ( ~n355 & n2377 ) | ( ~n355 & n2738 ) | ( n2377 & n2738 ) ;
  assign n5156 = n5155 ^ n621 ^ x212 ;
  assign n5157 = n5156 ^ n2899 ^ n1169 ;
  assign n5161 = n5038 ^ n2733 ^ n758 ;
  assign n5162 = n1339 & n2206 ;
  assign n5163 = ~n5161 & n5162 ;
  assign n5164 = n5163 ^ n3889 ^ x241 ;
  assign n5158 = n751 & n1751 ;
  assign n5159 = n5158 ^ n4141 ^ 1'b0 ;
  assign n5160 = n5159 ^ n4533 ^ n3957 ;
  assign n5165 = n5164 ^ n5160 ^ n2785 ;
  assign n5166 = n5165 ^ n540 ^ n349 ;
  assign n5167 = n4916 ^ n1420 ^ n602 ;
  assign n5168 = n5101 ^ x11 ^ 1'b0 ;
  assign n5169 = n5168 ^ n2028 ^ 1'b0 ;
  assign n5170 = ( ~n2360 & n5167 ) | ( ~n2360 & n5169 ) | ( n5167 & n5169 ) ;
  assign n5172 = n2286 ^ n934 ^ x220 ;
  assign n5171 = ( n352 & n4737 ) | ( n352 & n4835 ) | ( n4737 & n4835 ) ;
  assign n5173 = n5172 ^ n5171 ^ n2851 ;
  assign n5174 = ( x171 & n1039 ) | ( x171 & ~n1533 ) | ( n1039 & ~n1533 ) ;
  assign n5178 = ( n1261 & n3445 ) | ( n1261 & n3691 ) | ( n3445 & n3691 ) ;
  assign n5181 = n1160 | n4133 ;
  assign n5182 = n5181 ^ n3374 ^ n3151 ;
  assign n5180 = ( ~n1167 & n1442 ) | ( ~n1167 & n1535 ) | ( n1442 & n1535 ) ;
  assign n5183 = n5182 ^ n5180 ^ n1506 ;
  assign n5179 = ( n1303 & ~n1846 ) | ( n1303 & n3613 ) | ( ~n1846 & n3613 ) ;
  assign n5184 = n5183 ^ n5179 ^ n685 ;
  assign n5185 = ( n2279 & n5178 ) | ( n2279 & n5184 ) | ( n5178 & n5184 ) ;
  assign n5176 = n399 ^ x169 ^ 1'b0 ;
  assign n5177 = ( ~n2488 & n3406 ) | ( ~n2488 & n5176 ) | ( n3406 & n5176 ) ;
  assign n5175 = ( ~n2051 & n2125 ) | ( ~n2051 & n3387 ) | ( n2125 & n3387 ) ;
  assign n5186 = n5185 ^ n5177 ^ n5175 ;
  assign n5192 = n3296 ^ n2240 ^ n1413 ;
  assign n5187 = ( x137 & n3627 ) | ( x137 & n4593 ) | ( n3627 & n4593 ) ;
  assign n5188 = ( n769 & n927 ) | ( n769 & ~n5187 ) | ( n927 & ~n5187 ) ;
  assign n5189 = n5188 ^ n3355 ^ n1730 ;
  assign n5190 = n4836 ^ n4371 ^ 1'b0 ;
  assign n5191 = n5189 & n5190 ;
  assign n5193 = n5192 ^ n5191 ^ n2507 ;
  assign n5196 = n5145 ^ n1663 ^ x89 ;
  assign n5197 = ( x38 & n3284 ) | ( x38 & ~n5196 ) | ( n3284 & ~n5196 ) ;
  assign n5194 = ( n2524 & n2571 ) | ( n2524 & ~n3019 ) | ( n2571 & ~n3019 ) ;
  assign n5195 = n5194 ^ x124 ^ x108 ;
  assign n5198 = n5197 ^ n5195 ^ n3709 ;
  assign n5199 = n4297 ^ n2273 ^ 1'b0 ;
  assign n5201 = n617 & n1426 ;
  assign n5202 = ~n854 & n1362 ;
  assign n5203 = n5201 & n5202 ;
  assign n5204 = ( n395 & n571 ) | ( n395 & n5203 ) | ( n571 & n5203 ) ;
  assign n5200 = ~n3600 & n5073 ;
  assign n5205 = n5204 ^ n5200 ^ 1'b0 ;
  assign n5206 = n5199 | n5205 ;
  assign n5207 = n5206 ^ n4627 ^ n2220 ;
  assign n5208 = x70 & n5179 ;
  assign n5209 = n3658 ^ n2825 ^ n1224 ;
  assign n5210 = ( ~x5 & n1521 ) | ( ~x5 & n5209 ) | ( n1521 & n5209 ) ;
  assign n5217 = n1257 ^ n921 ^ 1'b0 ;
  assign n5218 = n610 & n5217 ;
  assign n5216 = ( n331 & n367 ) | ( n331 & ~n3643 ) | ( n367 & ~n3643 ) ;
  assign n5219 = n5218 ^ n5216 ^ n2462 ;
  assign n5211 = n3183 ^ n897 ^ 1'b0 ;
  assign n5212 = n3508 & n5211 ;
  assign n5213 = ( n1260 & n1997 ) | ( n1260 & ~n2172 ) | ( n1997 & ~n2172 ) ;
  assign n5214 = ( ~x233 & n5212 ) | ( ~x233 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5215 = n955 & n5214 ;
  assign n5220 = n5219 ^ n5215 ^ n2362 ;
  assign n5223 = n3559 ^ n1892 ^ n473 ;
  assign n5221 = ( n1274 & n1605 ) | ( n1274 & ~n4706 ) | ( n1605 & ~n4706 ) ;
  assign n5222 = ( n3095 & n4528 ) | ( n3095 & n5221 ) | ( n4528 & n5221 ) ;
  assign n5224 = n5223 ^ n5222 ^ n3022 ;
  assign n5227 = n1279 | n1830 ;
  assign n5228 = n1222 & ~n5227 ;
  assign n5225 = n2766 ^ n273 ^ x239 ;
  assign n5226 = ( n4271 & n4704 ) | ( n4271 & ~n5225 ) | ( n4704 & ~n5225 ) ;
  assign n5229 = n5228 ^ n5226 ^ n2657 ;
  assign n5230 = ( x174 & n5224 ) | ( x174 & n5229 ) | ( n5224 & n5229 ) ;
  assign n5231 = ( n5210 & ~n5220 ) | ( n5210 & n5230 ) | ( ~n5220 & n5230 ) ;
  assign n5232 = n2769 ^ n1127 ^ n760 ;
  assign n5233 = n5232 ^ n3263 ^ n1910 ;
  assign n5234 = ( n1835 & n2133 ) | ( n1835 & n2332 ) | ( n2133 & n2332 ) ;
  assign n5235 = n1372 ^ x226 ^ x54 ;
  assign n5236 = x121 & ~n3070 ;
  assign n5237 = n2972 & n5236 ;
  assign n5238 = n5237 ^ n1512 ^ 1'b0 ;
  assign n5239 = ( n4287 & ~n5235 ) | ( n4287 & n5238 ) | ( ~n5235 & n5238 ) ;
  assign n5240 = ( n955 & n1659 ) | ( n955 & n5239 ) | ( n1659 & n5239 ) ;
  assign n5241 = x45 & ~n5240 ;
  assign n5242 = n5234 & n5241 ;
  assign n5243 = ( n4038 & n5233 ) | ( n4038 & n5242 ) | ( n5233 & n5242 ) ;
  assign n5244 = ( n523 & n761 ) | ( n523 & ~n1188 ) | ( n761 & ~n1188 ) ;
  assign n5245 = n5244 ^ n1775 ^ x190 ;
  assign n5246 = ~n567 & n4480 ;
  assign n5247 = ~n4244 & n5246 ;
  assign n5248 = ( ~n1487 & n5245 ) | ( ~n1487 & n5247 ) | ( n5245 & n5247 ) ;
  assign n5249 = n4725 ^ n3338 ^ n565 ;
  assign n5250 = n1042 | n2356 ;
  assign n5251 = n5250 ^ n759 ^ 1'b0 ;
  assign n5252 = ( n1112 & ~n1121 ) | ( n1112 & n2703 ) | ( ~n1121 & n2703 ) ;
  assign n5253 = ( x7 & ~n5251 ) | ( x7 & n5252 ) | ( ~n5251 & n5252 ) ;
  assign n5254 = n5253 ^ n3050 ^ 1'b0 ;
  assign n5255 = n3177 & ~n5254 ;
  assign n5256 = ( ~n5248 & n5249 ) | ( ~n5248 & n5255 ) | ( n5249 & n5255 ) ;
  assign n5257 = n277 & n2860 ;
  assign n5258 = n5257 ^ n2286 ^ 1'b0 ;
  assign n5259 = n3941 & n5258 ;
  assign n5260 = n5259 ^ n5186 ^ n1794 ;
  assign n5261 = ( n1426 & n2566 ) | ( n1426 & ~n3366 ) | ( n2566 & ~n3366 ) ;
  assign n5269 = n4433 ^ n3302 ^ 1'b0 ;
  assign n5270 = n5269 ^ n4752 ^ x163 ;
  assign n5262 = n321 | n5188 ;
  assign n5263 = n5262 ^ n2351 ^ n2152 ;
  assign n5264 = ( n980 & n4750 ) | ( n980 & n4795 ) | ( n4750 & n4795 ) ;
  assign n5265 = n4907 ^ n1489 ^ n1332 ;
  assign n5266 = n3256 | n5265 ;
  assign n5267 = n5264 & ~n5266 ;
  assign n5268 = ~n5263 & n5267 ;
  assign n5271 = n5270 ^ n5268 ^ n2105 ;
  assign n5272 = n1836 ^ n1459 ^ x57 ;
  assign n5273 = ( n2041 & n5038 ) | ( n2041 & ~n5272 ) | ( n5038 & ~n5272 ) ;
  assign n5274 = n2013 ^ n545 ^ n469 ;
  assign n5275 = ( n912 & n2711 ) | ( n912 & ~n5274 ) | ( n2711 & ~n5274 ) ;
  assign n5277 = ( n546 & n2336 ) | ( n546 & ~n2552 ) | ( n2336 & ~n2552 ) ;
  assign n5278 = ( n1476 & n1534 ) | ( n1476 & ~n2879 ) | ( n1534 & ~n2879 ) ;
  assign n5279 = ( ~n3710 & n5277 ) | ( ~n3710 & n5278 ) | ( n5277 & n5278 ) ;
  assign n5276 = n3870 ^ n3269 ^ n1104 ;
  assign n5280 = n5279 ^ n5276 ^ 1'b0 ;
  assign n5281 = ( n1415 & ~n5275 ) | ( n1415 & n5280 ) | ( ~n5275 & n5280 ) ;
  assign n5282 = n3764 ^ n978 ^ 1'b0 ;
  assign n5283 = n3757 ^ n3384 ^ n2608 ;
  assign n5284 = n5283 ^ n4269 ^ n459 ;
  assign n5287 = n1394 ^ x245 ^ x48 ;
  assign n5288 = ( ~x83 & n693 ) | ( ~x83 & n5287 ) | ( n693 & n5287 ) ;
  assign n5286 = n440 ^ x183 ^ 1'b0 ;
  assign n5289 = n5288 ^ n5286 ^ n311 ;
  assign n5285 = x47 & ~n340 ;
  assign n5290 = n5289 ^ n5285 ^ n846 ;
  assign n5291 = ( n949 & n2976 ) | ( n949 & ~n5290 ) | ( n2976 & ~n5290 ) ;
  assign n5292 = ( n3117 & n5069 ) | ( n3117 & n5291 ) | ( n5069 & n5291 ) ;
  assign n5293 = n2165 ^ n727 ^ 1'b0 ;
  assign n5294 = n1275 | n5293 ;
  assign n5295 = ( n5284 & n5292 ) | ( n5284 & ~n5294 ) | ( n5292 & ~n5294 ) ;
  assign n5296 = ( n2640 & ~n3034 ) | ( n2640 & n4286 ) | ( ~n3034 & n4286 ) ;
  assign n5297 = n5296 ^ n1682 ^ 1'b0 ;
  assign n5313 = n2862 & n3822 ;
  assign n5314 = ~n2118 & n5313 ;
  assign n5315 = ( n1835 & ~n3646 ) | ( n1835 & n5314 ) | ( ~n3646 & n5314 ) ;
  assign n5301 = n2958 ^ n1816 ^ n1653 ;
  assign n5300 = ( n651 & n2629 ) | ( n651 & n5019 ) | ( n2629 & n5019 ) ;
  assign n5302 = n5301 ^ n5300 ^ n1078 ;
  assign n5298 = ( n558 & n604 ) | ( n558 & ~n4917 ) | ( n604 & ~n4917 ) ;
  assign n5299 = n5298 ^ n1205 ^ x107 ;
  assign n5303 = n5302 ^ n5299 ^ n5143 ;
  assign n5306 = n4755 ^ n727 ^ x108 ;
  assign n5304 = ( n1285 & n2784 ) | ( n1285 & ~n3056 ) | ( n2784 & ~n3056 ) ;
  assign n5305 = ( n2757 & n4048 ) | ( n2757 & ~n5304 ) | ( n4048 & ~n5304 ) ;
  assign n5307 = n5306 ^ n5305 ^ n1307 ;
  assign n5308 = ( n4111 & n5303 ) | ( n4111 & ~n5307 ) | ( n5303 & ~n5307 ) ;
  assign n5309 = ( n289 & n1180 ) | ( n289 & ~n1474 ) | ( n1180 & ~n1474 ) ;
  assign n5310 = ~n4105 & n5309 ;
  assign n5311 = n5308 | n5310 ;
  assign n5312 = n5311 ^ n2362 ^ 1'b0 ;
  assign n5316 = n5315 ^ n5312 ^ n691 ;
  assign n5317 = ( n2291 & n3466 ) | ( n2291 & ~n5316 ) | ( n3466 & ~n5316 ) ;
  assign n5318 = ( n5166 & ~n5297 ) | ( n5166 & n5317 ) | ( ~n5297 & n5317 ) ;
  assign n5319 = n3639 ^ n2563 ^ n947 ;
  assign n5320 = n4222 ^ n1917 ^ 1'b0 ;
  assign n5321 = x109 & ~n5320 ;
  assign n5322 = n5321 ^ n4210 ^ n284 ;
  assign n5323 = ( n360 & ~n3177 ) | ( n360 & n5322 ) | ( ~n3177 & n5322 ) ;
  assign n5324 = n5323 ^ n1910 ^ n644 ;
  assign n5325 = ( ~n1014 & n5319 ) | ( ~n1014 & n5324 ) | ( n5319 & n5324 ) ;
  assign n5326 = ( ~n1269 & n2098 ) | ( ~n1269 & n5304 ) | ( n2098 & n5304 ) ;
  assign n5327 = ( n4472 & n4630 ) | ( n4472 & n5326 ) | ( n4630 & n5326 ) ;
  assign n5328 = n5327 ^ n5050 ^ 1'b0 ;
  assign n5334 = n4856 ^ n2565 ^ n933 ;
  assign n5336 = ( n968 & ~n1639 ) | ( n968 & n3387 ) | ( ~n1639 & n3387 ) ;
  assign n5335 = ~n435 & n4492 ;
  assign n5337 = n5336 ^ n5335 ^ 1'b0 ;
  assign n5338 = ~n2066 & n5337 ;
  assign n5339 = n2157 ^ n1511 ^ n310 ;
  assign n5340 = ( n950 & n965 ) | ( n950 & n5339 ) | ( n965 & n5339 ) ;
  assign n5341 = n1595 ^ n828 ^ n532 ;
  assign n5342 = n5341 ^ n2184 ^ 1'b0 ;
  assign n5343 = ~n5340 & n5342 ;
  assign n5344 = ( ~n518 & n728 ) | ( ~n518 & n3260 ) | ( n728 & n3260 ) ;
  assign n5345 = n5344 ^ n4947 ^ n4594 ;
  assign n5346 = ( ~n5338 & n5343 ) | ( ~n5338 & n5345 ) | ( n5343 & n5345 ) ;
  assign n5347 = ( ~n2253 & n5334 ) | ( ~n2253 & n5346 ) | ( n5334 & n5346 ) ;
  assign n5329 = n1531 ^ n591 ^ n400 ;
  assign n5330 = ( n1477 & n3142 ) | ( n1477 & n5329 ) | ( n3142 & n5329 ) ;
  assign n5331 = n5330 ^ x129 ^ x61 ;
  assign n5332 = n5331 ^ n4013 ^ n1771 ;
  assign n5333 = n4580 | n5332 ;
  assign n5348 = n5347 ^ n5333 ^ 1'b0 ;
  assign n5351 = ( n1566 & n2401 ) | ( n1566 & n2962 ) | ( n2401 & n2962 ) ;
  assign n5352 = ( n1161 & n3302 ) | ( n1161 & n5351 ) | ( n3302 & n5351 ) ;
  assign n5349 = n2687 | n4691 ;
  assign n5350 = n5349 ^ x164 ^ 1'b0 ;
  assign n5353 = n5352 ^ n5350 ^ n2220 ;
  assign n5354 = n3811 ^ n3271 ^ n545 ;
  assign n5358 = ( ~n1693 & n1858 ) | ( ~n1693 & n5022 ) | ( n1858 & n5022 ) ;
  assign n5359 = ( ~n2993 & n4727 ) | ( ~n2993 & n5358 ) | ( n4727 & n5358 ) ;
  assign n5355 = ( n2807 & n3197 ) | ( n2807 & n4820 ) | ( n3197 & n4820 ) ;
  assign n5356 = ( n4104 & ~n4544 ) | ( n4104 & n5355 ) | ( ~n4544 & n5355 ) ;
  assign n5357 = ~n1266 & n5356 ;
  assign n5360 = n5359 ^ n5357 ^ 1'b0 ;
  assign n5361 = n5315 ^ n3378 ^ n1355 ;
  assign n5362 = n2329 & ~n3270 ;
  assign n5363 = n5361 & n5362 ;
  assign n5364 = ( x5 & ~n5302 ) | ( x5 & n5345 ) | ( ~n5302 & n5345 ) ;
  assign n5365 = ( x97 & n3648 ) | ( x97 & n3740 ) | ( n3648 & n3740 ) ;
  assign n5366 = ( n990 & ~n3650 ) | ( n990 & n3776 ) | ( ~n3650 & n3776 ) ;
  assign n5367 = n5366 ^ n4064 ^ n1596 ;
  assign n5368 = ( n1817 & n1953 ) | ( n1817 & n5367 ) | ( n1953 & n5367 ) ;
  assign n5369 = n5368 ^ n2993 ^ n2127 ;
  assign n5370 = ( ~n2381 & n3541 ) | ( ~n2381 & n5369 ) | ( n3541 & n5369 ) ;
  assign n5371 = n1335 & ~n5370 ;
  assign n5372 = n3191 & n5371 ;
  assign n5373 = n5372 ^ n4380 ^ n620 ;
  assign n5383 = ( n761 & ~n1425 ) | ( n761 & n1785 ) | ( ~n1425 & n1785 ) ;
  assign n5381 = n4019 ^ n428 ^ 1'b0 ;
  assign n5382 = n1935 & ~n5381 ;
  assign n5384 = n5383 ^ n5382 ^ 1'b0 ;
  assign n5376 = n1344 ^ x59 ^ 1'b0 ;
  assign n5377 = ( n1783 & n3201 ) | ( n1783 & ~n5376 ) | ( n3201 & ~n5376 ) ;
  assign n5378 = ( n2481 & n3639 ) | ( n2481 & ~n5377 ) | ( n3639 & ~n5377 ) ;
  assign n5375 = n2399 ^ n1800 ^ n395 ;
  assign n5374 = n1012 & ~n2249 ;
  assign n5379 = n5378 ^ n5375 ^ n5374 ;
  assign n5380 = n4424 | n5379 ;
  assign n5385 = n5384 ^ n5380 ^ 1'b0 ;
  assign n5393 = x80 & n4944 ;
  assign n5394 = n5393 ^ n2224 ^ n1558 ;
  assign n5389 = n2314 ^ n1422 ^ 1'b0 ;
  assign n5390 = n3743 & n5389 ;
  assign n5391 = n5390 ^ n3594 ^ x18 ;
  assign n5386 = ( n676 & ~n717 ) | ( n676 & n4582 ) | ( ~n717 & n4582 ) ;
  assign n5387 = n5386 ^ n3319 ^ x127 ;
  assign n5388 = n5387 ^ n4239 ^ n4231 ;
  assign n5392 = n5391 ^ n5388 ^ n1338 ;
  assign n5395 = n5394 ^ n5392 ^ n4752 ;
  assign n5396 = n4727 ^ n3842 ^ n2355 ;
  assign n5397 = n5396 ^ n4079 ^ n3222 ;
  assign n5398 = n5397 ^ n4831 ^ 1'b0 ;
  assign n5399 = n535 & ~n5398 ;
  assign n5400 = ( n651 & n5395 ) | ( n651 & n5399 ) | ( n5395 & n5399 ) ;
  assign n5401 = ( n1278 & n1684 ) | ( n1278 & ~n3052 ) | ( n1684 & ~n3052 ) ;
  assign n5402 = ( n1589 & ~n2370 ) | ( n1589 & n5401 ) | ( ~n2370 & n5401 ) ;
  assign n5403 = ( n650 & n1026 ) | ( n650 & ~n4079 ) | ( n1026 & ~n4079 ) ;
  assign n5404 = n5403 ^ n4465 ^ 1'b0 ;
  assign n5405 = n3292 ^ n1471 ^ x175 ;
  assign n5406 = n5405 ^ n4854 ^ x156 ;
  assign n5407 = n4988 ^ n1700 ^ n609 ;
  assign n5408 = n4688 ^ n3880 ^ 1'b0 ;
  assign n5409 = ( ~n938 & n5407 ) | ( ~n938 & n5408 ) | ( n5407 & n5408 ) ;
  assign n5410 = n3376 & ~n3709 ;
  assign n5411 = n3735 & n5410 ;
  assign n5412 = ( n1921 & ~n4789 ) | ( n1921 & n5411 ) | ( ~n4789 & n5411 ) ;
  assign n5413 = n2514 ^ x239 ^ 1'b0 ;
  assign n5414 = n5413 ^ n2813 ^ n406 ;
  assign n5415 = x77 & n923 ;
  assign n5416 = n3003 & n5415 ;
  assign n5417 = n5416 ^ n5070 ^ n2102 ;
  assign n5418 = ( ~n1054 & n5414 ) | ( ~n1054 & n5417 ) | ( n5414 & n5417 ) ;
  assign n5422 = ( ~n3777 & n5358 ) | ( ~n3777 & n5368 ) | ( n5358 & n5368 ) ;
  assign n5419 = ( n275 & ~n1902 ) | ( n275 & n3742 ) | ( ~n1902 & n3742 ) ;
  assign n5420 = ~n1107 & n5419 ;
  assign n5421 = n5283 & n5420 ;
  assign n5423 = n5422 ^ n5421 ^ n4344 ;
  assign n5424 = ( n951 & n1686 ) | ( n951 & ~n3183 ) | ( n1686 & ~n3183 ) ;
  assign n5425 = n5424 ^ n4492 ^ n2122 ;
  assign n5426 = n3533 ^ n457 ^ 1'b0 ;
  assign n5427 = n4371 & n5426 ;
  assign n5431 = n1640 | n4690 ;
  assign n5432 = n4598 | n5431 ;
  assign n5428 = ( n1664 & n2453 ) | ( n1664 & ~n5083 ) | ( n2453 & ~n5083 ) ;
  assign n5429 = ( ~n2638 & n3266 ) | ( ~n2638 & n5428 ) | ( n3266 & n5428 ) ;
  assign n5430 = ~n1910 & n5429 ;
  assign n5433 = n5432 ^ n5430 ^ 1'b0 ;
  assign n5434 = n5427 | n5433 ;
  assign n5435 = n5434 ^ n4831 ^ n3040 ;
  assign n5437 = n2158 ^ x240 ^ 1'b0 ;
  assign n5438 = n5437 ^ n3864 ^ n3753 ;
  assign n5436 = n589 | n964 ;
  assign n5439 = n5438 ^ n5436 ^ 1'b0 ;
  assign n5440 = n3264 & n5439 ;
  assign n5441 = n5435 & n5440 ;
  assign n5445 = n1368 ^ n296 ^ x238 ;
  assign n5446 = n2317 | n5445 ;
  assign n5447 = n5446 ^ x50 ^ 1'b0 ;
  assign n5448 = ( ~n3305 & n4882 ) | ( ~n3305 & n5447 ) | ( n4882 & n5447 ) ;
  assign n5449 = ( n980 & n1107 ) | ( n980 & n3303 ) | ( n1107 & n3303 ) ;
  assign n5450 = ( n783 & n5448 ) | ( n783 & n5449 ) | ( n5448 & n5449 ) ;
  assign n5442 = ( n1146 & n1511 ) | ( n1146 & ~n1690 ) | ( n1511 & ~n1690 ) ;
  assign n5443 = n1751 & ~n5442 ;
  assign n5444 = n5443 ^ n5161 ^ n3189 ;
  assign n5451 = n5450 ^ n5444 ^ 1'b0 ;
  assign n5452 = n1579 ^ n1540 ^ n1187 ;
  assign n5453 = n5452 ^ n4862 ^ n3238 ;
  assign n5455 = ( n777 & ~n3509 ) | ( n777 & n3815 ) | ( ~n3509 & n3815 ) ;
  assign n5456 = n5455 ^ n2443 ^ n383 ;
  assign n5454 = n4326 & n4909 ;
  assign n5457 = n5456 ^ n5454 ^ 1'b0 ;
  assign n5458 = n5453 | n5457 ;
  assign n5463 = n3236 ^ n2546 ^ n1130 ;
  assign n5464 = n1903 & ~n5463 ;
  assign n5461 = ( n1816 & n1866 ) | ( n1816 & ~n3250 ) | ( n1866 & ~n3250 ) ;
  assign n5462 = ( n418 & ~n1090 ) | ( n418 & n5461 ) | ( ~n1090 & n5461 ) ;
  assign n5459 = n1693 ^ n1348 ^ 1'b0 ;
  assign n5460 = n5459 ^ n1318 ^ n305 ;
  assign n5465 = n5464 ^ n5462 ^ n5460 ;
  assign n5469 = n4598 ^ n3785 ^ 1'b0 ;
  assign n5470 = n1000 | n5469 ;
  assign n5471 = n5470 ^ n5163 ^ n2059 ;
  assign n5466 = ~n1272 & n5002 ;
  assign n5467 = n1330 & n5466 ;
  assign n5468 = ~n4343 & n5467 ;
  assign n5472 = n5471 ^ n5468 ^ n2884 ;
  assign n5473 = n5289 ^ n4726 ^ x18 ;
  assign n5474 = n1361 ^ n1359 ^ n1285 ;
  assign n5475 = ( n1949 & n5339 ) | ( n1949 & n5474 ) | ( n5339 & n5474 ) ;
  assign n5476 = ( n2645 & n4704 ) | ( n2645 & n5475 ) | ( n4704 & n5475 ) ;
  assign n5478 = n3151 & ~n3172 ;
  assign n5479 = n5478 ^ n2951 ^ 1'b0 ;
  assign n5480 = ( n869 & ~n3856 ) | ( n869 & n5479 ) | ( ~n3856 & n5479 ) ;
  assign n5481 = ( n293 & n1651 ) | ( n293 & n5480 ) | ( n1651 & n5480 ) ;
  assign n5482 = n3734 & ~n5481 ;
  assign n5483 = ~x149 & n5482 ;
  assign n5477 = n957 | n3396 ;
  assign n5484 = n5483 ^ n5477 ^ 1'b0 ;
  assign n5485 = n959 & ~n5484 ;
  assign n5486 = x51 & n956 ;
  assign n5487 = ~n5485 & n5486 ;
  assign n5488 = x252 & n4198 ;
  assign n5489 = ~n940 & n5488 ;
  assign n5492 = ( n470 & n973 ) | ( n470 & ~n1101 ) | ( n973 & ~n1101 ) ;
  assign n5493 = n5492 ^ n4232 ^ n1022 ;
  assign n5490 = ( n872 & n3384 ) | ( n872 & n3872 ) | ( n3384 & n3872 ) ;
  assign n5491 = n5490 ^ n3871 ^ n3138 ;
  assign n5494 = n5493 ^ n5491 ^ n1970 ;
  assign n5495 = n558 ^ x173 ^ 1'b0 ;
  assign n5496 = ( x232 & ~n5494 ) | ( x232 & n5495 ) | ( ~n5494 & n5495 ) ;
  assign n5505 = ( n1198 & ~n2519 ) | ( n1198 & n2969 ) | ( ~n2519 & n2969 ) ;
  assign n5498 = ( x63 & n1065 ) | ( x63 & n2736 ) | ( n1065 & n2736 ) ;
  assign n5497 = n1062 | n3372 ;
  assign n5499 = n5498 ^ n5497 ^ 1'b0 ;
  assign n5501 = ~n840 & n1151 ;
  assign n5502 = n5501 ^ n666 ^ x194 ;
  assign n5500 = ( n3382 & n3446 ) | ( n3382 & n4977 ) | ( n3446 & n4977 ) ;
  assign n5503 = n5502 ^ n5500 ^ n1718 ;
  assign n5504 = ( n2290 & n5499 ) | ( n2290 & ~n5503 ) | ( n5499 & ~n5503 ) ;
  assign n5506 = n5505 ^ n5504 ^ 1'b0 ;
  assign n5507 = n5496 & ~n5506 ;
  assign n5508 = ~n3189 & n5507 ;
  assign n5509 = n5489 & n5508 ;
  assign n5510 = ( x66 & ~n1977 ) | ( x66 & n3776 ) | ( ~n1977 & n3776 ) ;
  assign n5511 = ( n1790 & n3140 ) | ( n1790 & ~n5510 ) | ( n3140 & ~n5510 ) ;
  assign n5512 = n5511 ^ n881 ^ n561 ;
  assign n5513 = ( n3632 & n3810 ) | ( n3632 & n5512 ) | ( n3810 & n5512 ) ;
  assign n5515 = n1783 ^ n713 ^ n613 ;
  assign n5514 = ( n1194 & n1624 ) | ( n1194 & ~n3822 ) | ( n1624 & ~n3822 ) ;
  assign n5516 = n5515 ^ n5514 ^ n657 ;
  assign n5521 = n2282 ^ n626 ^ x161 ;
  assign n5518 = ( n826 & n1263 ) | ( n826 & ~n2850 ) | ( n1263 & ~n2850 ) ;
  assign n5517 = n356 & n5006 ;
  assign n5519 = n5518 ^ n5517 ^ 1'b0 ;
  assign n5520 = ( n364 & ~n2771 ) | ( n364 & n5519 ) | ( ~n2771 & n5519 ) ;
  assign n5522 = n5521 ^ n5520 ^ n676 ;
  assign n5523 = n5522 ^ n4308 ^ n263 ;
  assign n5524 = n1184 | n3279 ;
  assign n5529 = n1506 ^ x72 ^ 1'b0 ;
  assign n5530 = n462 & n5529 ;
  assign n5531 = ~n1024 & n2690 ;
  assign n5532 = n541 & n5531 ;
  assign n5533 = ( n1714 & n2304 ) | ( n1714 & ~n5532 ) | ( n2304 & ~n5532 ) ;
  assign n5534 = ( n872 & ~n5530 ) | ( n872 & n5533 ) | ( ~n5530 & n5533 ) ;
  assign n5525 = n5298 ^ n1615 ^ 1'b0 ;
  assign n5526 = n4402 ^ n2899 ^ 1'b0 ;
  assign n5527 = ~n2654 & n5526 ;
  assign n5528 = ~n5525 & n5527 ;
  assign n5535 = n5534 ^ n5528 ^ n1195 ;
  assign n5536 = n3139 & ~n3727 ;
  assign n5537 = n3477 & ~n5536 ;
  assign n5538 = ~n5535 & n5537 ;
  assign n5540 = ( ~n1527 & n4158 ) | ( ~n1527 & n4297 ) | ( n4158 & n4297 ) ;
  assign n5539 = ( n1297 & ~n1850 ) | ( n1297 & n1965 ) | ( ~n1850 & n1965 ) ;
  assign n5541 = n5540 ^ n5539 ^ 1'b0 ;
  assign n5548 = ( ~x0 & x138 ) | ( ~x0 & n4359 ) | ( x138 & n4359 ) ;
  assign n5542 = n1006 ^ n996 ^ 1'b0 ;
  assign n5543 = n1661 & n5542 ;
  assign n5544 = n5543 ^ n465 ^ 1'b0 ;
  assign n5545 = n5544 ^ n5527 ^ n1761 ;
  assign n5546 = n5545 ^ n1796 ^ n276 ;
  assign n5547 = n5546 ^ n4442 ^ n2829 ;
  assign n5549 = n5548 ^ n5547 ^ n3580 ;
  assign n5550 = n4387 ^ n2498 ^ n1459 ;
  assign n5551 = n2744 & n4585 ;
  assign n5552 = n5551 ^ n2164 ^ 1'b0 ;
  assign n5553 = n1003 & ~n2978 ;
  assign n5554 = ( n399 & ~n1579 ) | ( n399 & n4391 ) | ( ~n1579 & n4391 ) ;
  assign n5555 = ( ~n2195 & n5553 ) | ( ~n2195 & n5554 ) | ( n5553 & n5554 ) ;
  assign n5556 = ( x0 & n5552 ) | ( x0 & ~n5555 ) | ( n5552 & ~n5555 ) ;
  assign n5557 = ( ~n1295 & n5550 ) | ( ~n1295 & n5556 ) | ( n5550 & n5556 ) ;
  assign n5573 = n4792 ^ n3579 ^ n2311 ;
  assign n5574 = ( n3023 & n4370 ) | ( n3023 & n5573 ) | ( n4370 & n5573 ) ;
  assign n5564 = n3858 ^ n957 ^ x31 ;
  assign n5565 = n5564 ^ n4584 ^ n2069 ;
  assign n5563 = n1583 ^ n322 ^ 1'b0 ;
  assign n5566 = n5565 ^ n5563 ^ n3134 ;
  assign n5567 = ( n1247 & n4104 ) | ( n1247 & ~n5566 ) | ( n4104 & ~n5566 ) ;
  assign n5568 = ( n641 & n847 ) | ( n641 & n1034 ) | ( n847 & n1034 ) ;
  assign n5569 = n3956 & n5568 ;
  assign n5570 = n2608 & n5569 ;
  assign n5571 = ( ~n646 & n3910 ) | ( ~n646 & n5570 ) | ( n3910 & n5570 ) ;
  assign n5572 = ( n5176 & n5567 ) | ( n5176 & n5571 ) | ( n5567 & n5571 ) ;
  assign n5559 = n3240 ^ n3076 ^ n1236 ;
  assign n5558 = ~n1282 & n2067 ;
  assign n5560 = n5559 ^ n5558 ^ 1'b0 ;
  assign n5561 = n5560 ^ n4622 ^ n945 ;
  assign n5562 = n5561 ^ n5178 ^ n596 ;
  assign n5575 = n5574 ^ n5572 ^ n5562 ;
  assign n5576 = ( n1722 & ~n2173 ) | ( n1722 & n3201 ) | ( ~n2173 & n3201 ) ;
  assign n5577 = ( n619 & n1565 ) | ( n619 & n3205 ) | ( n1565 & n3205 ) ;
  assign n5584 = n1946 ^ n1927 ^ n640 ;
  assign n5581 = n1368 ^ n910 ^ n558 ;
  assign n5582 = n2020 & ~n5581 ;
  assign n5583 = n5582 ^ n2141 ^ 1'b0 ;
  assign n5585 = n5584 ^ n5583 ^ n2260 ;
  assign n5579 = n561 & ~n2661 ;
  assign n5580 = n5579 ^ n1265 ^ 1'b0 ;
  assign n5586 = n5585 ^ n5580 ^ n2309 ;
  assign n5578 = n2629 ^ n1873 ^ n739 ;
  assign n5587 = n5586 ^ n5578 ^ x83 ;
  assign n5588 = ( n3528 & ~n5577 ) | ( n3528 & n5587 ) | ( ~n5577 & n5587 ) ;
  assign n5589 = n5588 ^ n4050 ^ 1'b0 ;
  assign n5590 = n5576 & ~n5589 ;
  assign n5592 = n885 | n3885 ;
  assign n5591 = ( ~n475 & n664 ) | ( ~n475 & n1038 ) | ( n664 & n1038 ) ;
  assign n5593 = n5592 ^ n5591 ^ n4656 ;
  assign n5594 = ( ~n1929 & n1975 ) | ( ~n1929 & n5593 ) | ( n1975 & n5593 ) ;
  assign n5595 = n5594 ^ n504 ^ x0 ;
  assign n5596 = ( n1716 & n2217 ) | ( n1716 & n5595 ) | ( n2217 & n5595 ) ;
  assign n5599 = n5253 ^ n4463 ^ n3350 ;
  assign n5602 = n3716 ^ n711 ^ 1'b0 ;
  assign n5603 = n2171 & ~n5602 ;
  assign n5600 = n4053 ^ n2336 ^ n511 ;
  assign n5601 = ( n584 & n3535 ) | ( n584 & n5600 ) | ( n3535 & n5600 ) ;
  assign n5604 = n5603 ^ n5601 ^ 1'b0 ;
  assign n5605 = n5599 | n5604 ;
  assign n5597 = ( n552 & ~n1940 ) | ( n552 & n2257 ) | ( ~n1940 & n2257 ) ;
  assign n5598 = n5597 ^ n4891 ^ n2930 ;
  assign n5606 = n5605 ^ n5598 ^ n3669 ;
  assign n5621 = ~n2141 & n3027 ;
  assign n5620 = n2564 & n3373 ;
  assign n5622 = n5621 ^ n5620 ^ 1'b0 ;
  assign n5607 = n4205 ^ n2557 ^ n1373 ;
  assign n5608 = n5607 ^ n4693 ^ n2578 ;
  assign n5609 = n4126 ^ n2058 ^ n1384 ;
  assign n5610 = x217 & ~n701 ;
  assign n5611 = n5610 ^ n2872 ^ 1'b0 ;
  assign n5612 = ( n2337 & n5609 ) | ( n2337 & ~n5611 ) | ( n5609 & ~n5611 ) ;
  assign n5613 = ~n5063 & n5612 ;
  assign n5614 = n5613 ^ n2901 ^ 1'b0 ;
  assign n5615 = ( n1076 & n1377 ) | ( n1076 & n4904 ) | ( n1377 & n4904 ) ;
  assign n5616 = ~n4656 & n4860 ;
  assign n5617 = n5615 & ~n5616 ;
  assign n5618 = n5614 & n5617 ;
  assign n5619 = ( ~n4069 & n5608 ) | ( ~n4069 & n5618 ) | ( n5608 & n5618 ) ;
  assign n5623 = n5622 ^ n5619 ^ n4022 ;
  assign n5624 = ( n1419 & ~n3651 ) | ( n1419 & n5382 ) | ( ~n3651 & n5382 ) ;
  assign n5625 = ( n2133 & n2890 ) | ( n2133 & ~n2952 ) | ( n2890 & ~n2952 ) ;
  assign n5626 = ( ~n1274 & n4884 ) | ( ~n1274 & n5332 ) | ( n4884 & n5332 ) ;
  assign n5627 = ( n5624 & n5625 ) | ( n5624 & n5626 ) | ( n5625 & n5626 ) ;
  assign n5628 = n4177 ^ n2205 ^ n319 ;
  assign n5629 = ( n693 & n3984 ) | ( n693 & ~n5628 ) | ( n3984 & ~n5628 ) ;
  assign n5630 = n5629 ^ n3222 ^ n2721 ;
  assign n5631 = n3858 | n5630 ;
  assign n5632 = n5631 ^ n5599 ^ n857 ;
  assign n5633 = ( n3087 & n5194 ) | ( n3087 & ~n5601 ) | ( n5194 & ~n5601 ) ;
  assign n5634 = n3695 ^ n3012 ^ n2445 ;
  assign n5635 = n5634 ^ n4191 ^ x60 ;
  assign n5636 = ( x211 & n1727 ) | ( x211 & n3082 ) | ( n1727 & n3082 ) ;
  assign n5637 = n1845 & n5636 ;
  assign n5638 = ~n5635 & n5637 ;
  assign n5639 = ~n5498 & n5638 ;
  assign n5640 = ( ~n4318 & n5633 ) | ( ~n4318 & n5639 ) | ( n5633 & n5639 ) ;
  assign n5641 = ( ~n3174 & n3200 ) | ( ~n3174 & n5171 ) | ( n3200 & n5171 ) ;
  assign n5642 = ( n1452 & n1589 ) | ( n1452 & ~n2110 ) | ( n1589 & ~n2110 ) ;
  assign n5643 = ( n2609 & n3071 ) | ( n2609 & n5642 ) | ( n3071 & n5642 ) ;
  assign n5656 = n2521 ^ n1033 ^ n1001 ;
  assign n5657 = n5656 ^ n2655 ^ n741 ;
  assign n5658 = n5657 ^ n4123 ^ n3711 ;
  assign n5659 = ~n2914 & n5658 ;
  assign n5654 = n315 & ~n5226 ;
  assign n5655 = n5654 ^ n1754 ^ x71 ;
  assign n5644 = n4352 ^ n3575 ^ n2888 ;
  assign n5645 = n5644 ^ n2672 ^ n288 ;
  assign n5646 = ( n1265 & n3807 ) | ( n1265 & ~n5645 ) | ( n3807 & ~n5645 ) ;
  assign n5647 = ( n1289 & ~n1456 ) | ( n1289 & n5646 ) | ( ~n1456 & n5646 ) ;
  assign n5648 = n3649 ^ n1843 ^ n1515 ;
  assign n5649 = ( x202 & ~n710 ) | ( x202 & n3877 ) | ( ~n710 & n3877 ) ;
  assign n5650 = ( n1759 & ~n5648 ) | ( n1759 & n5649 ) | ( ~n5648 & n5649 ) ;
  assign n5651 = ( n4701 & n5647 ) | ( n4701 & n5650 ) | ( n5647 & n5650 ) ;
  assign n5652 = ( ~n1547 & n5276 ) | ( ~n1547 & n5651 ) | ( n5276 & n5651 ) ;
  assign n5653 = n4298 | n5652 ;
  assign n5660 = n5659 ^ n5655 ^ n5653 ;
  assign n5661 = n2621 ^ n925 ^ n595 ;
  assign n5662 = ( ~n676 & n1262 ) | ( ~n676 & n5661 ) | ( n1262 & n5661 ) ;
  assign n5663 = n5662 ^ n4918 ^ n2782 ;
  assign n5664 = n655 | n1275 ;
  assign n5665 = n4357 | n5664 ;
  assign n5666 = ( x94 & n2511 ) | ( x94 & n3666 ) | ( n2511 & n3666 ) ;
  assign n5667 = ( n2220 & n3012 ) | ( n2220 & n5666 ) | ( n3012 & n5666 ) ;
  assign n5668 = ( n4090 & ~n5665 ) | ( n4090 & n5667 ) | ( ~n5665 & n5667 ) ;
  assign n5669 = ( n3058 & n5663 ) | ( n3058 & ~n5668 ) | ( n5663 & ~n5668 ) ;
  assign n5670 = ( ~n647 & n3007 ) | ( ~n647 & n4039 ) | ( n3007 & n4039 ) ;
  assign n5671 = n5670 ^ n1819 ^ 1'b0 ;
  assign n5672 = n256 & ~n5671 ;
  assign n5673 = n5672 ^ n3855 ^ 1'b0 ;
  assign n5674 = n2296 ^ n932 ^ x104 ;
  assign n5675 = n1696 ^ n1026 ^ x116 ;
  assign n5676 = ~n1757 & n5675 ;
  assign n5677 = n5676 ^ n3025 ^ 1'b0 ;
  assign n5678 = ~n5674 & n5677 ;
  assign n5679 = n5678 ^ n3711 ^ n345 ;
  assign n5680 = ( n1790 & ~n2741 ) | ( n1790 & n4391 ) | ( ~n2741 & n4391 ) ;
  assign n5681 = n5149 ^ n3286 ^ 1'b0 ;
  assign n5682 = n5681 ^ n4134 ^ n2430 ;
  assign n5683 = n5682 ^ n4350 ^ n940 ;
  assign n5684 = ( n3283 & ~n5680 ) | ( n3283 & n5683 ) | ( ~n5680 & n5683 ) ;
  assign n5685 = n5278 ^ n3980 ^ n3570 ;
  assign n5686 = ( x4 & n5684 ) | ( x4 & ~n5685 ) | ( n5684 & ~n5685 ) ;
  assign n5695 = n4856 ^ n2543 ^ n1612 ;
  assign n5687 = n3518 ^ n2273 ^ n907 ;
  assign n5689 = n1660 ^ n546 ^ n334 ;
  assign n5690 = n5689 ^ n2184 ^ n439 ;
  assign n5688 = ( ~x8 & x78 ) | ( ~x8 & n3951 ) | ( x78 & n3951 ) ;
  assign n5691 = n5690 ^ n5688 ^ n2145 ;
  assign n5692 = n1388 | n2799 ;
  assign n5693 = n5691 & ~n5692 ;
  assign n5694 = n5687 & ~n5693 ;
  assign n5696 = n5695 ^ n5694 ^ n3379 ;
  assign n5697 = ~n1469 & n4470 ;
  assign n5698 = ~n5696 & n5697 ;
  assign n5699 = x220 & n898 ;
  assign n5700 = ( x68 & n1095 ) | ( x68 & ~n5699 ) | ( n1095 & ~n5699 ) ;
  assign n5701 = ( n2587 & ~n4326 ) | ( n2587 & n4929 ) | ( ~n4326 & n4929 ) ;
  assign n5704 = n2510 ^ n1497 ^ n1427 ;
  assign n5705 = ( ~n1204 & n2424 ) | ( ~n1204 & n4364 ) | ( n2424 & n4364 ) ;
  assign n5706 = ( n1819 & n2011 ) | ( n1819 & n4198 ) | ( n2011 & n4198 ) ;
  assign n5707 = ( n5693 & n5705 ) | ( n5693 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = n5707 ^ n2378 ^ 1'b0 ;
  assign n5709 = n3079 | n5708 ;
  assign n5710 = ( n5178 & n5704 ) | ( n5178 & ~n5709 ) | ( n5704 & ~n5709 ) ;
  assign n5711 = n2319 ^ x130 ^ 1'b0 ;
  assign n5712 = ~n668 & n5711 ;
  assign n5713 = n5712 ^ n3711 ^ 1'b0 ;
  assign n5714 = ( ~n805 & n5710 ) | ( ~n805 & n5713 ) | ( n5710 & n5713 ) ;
  assign n5702 = n5078 ^ n1691 ^ n339 ;
  assign n5703 = n5702 ^ n2929 ^ 1'b0 ;
  assign n5715 = n5714 ^ n5703 ^ n1580 ;
  assign n5716 = ( n5700 & n5701 ) | ( n5700 & ~n5715 ) | ( n5701 & ~n5715 ) ;
  assign n5717 = n5716 ^ n5470 ^ n4254 ;
  assign n5718 = n3984 ^ n1555 ^ n860 ;
  assign n5719 = n1223 & n1509 ;
  assign n5720 = n796 ^ x2 ^ 1'b0 ;
  assign n5721 = n2598 & ~n5720 ;
  assign n5722 = ( ~x7 & n622 ) | ( ~x7 & n5721 ) | ( n622 & n5721 ) ;
  assign n5723 = ( ~n5718 & n5719 ) | ( ~n5718 & n5722 ) | ( n5719 & n5722 ) ;
  assign n5724 = n1536 ^ n1434 ^ 1'b0 ;
  assign n5725 = n579 & ~n5724 ;
  assign n5726 = ( n752 & n5053 ) | ( n752 & ~n5725 ) | ( n5053 & ~n5725 ) ;
  assign n5727 = n2067 & n5726 ;
  assign n5728 = n667 | n5727 ;
  assign n5729 = ~n5723 & n5728 ;
  assign n5730 = n3502 ^ n1117 ^ x194 ;
  assign n5731 = ( n4589 & ~n5688 ) | ( n4589 & n5730 ) | ( ~n5688 & n5730 ) ;
  assign n5732 = n5731 ^ n2916 ^ n1332 ;
  assign n5733 = n3789 ^ n2567 ^ 1'b0 ;
  assign n5734 = n1644 ^ n285 ^ 1'b0 ;
  assign n5735 = n5238 ^ n1628 ^ n568 ;
  assign n5736 = ( n3262 & n5091 ) | ( n3262 & ~n5735 ) | ( n5091 & ~n5735 ) ;
  assign n5737 = ( n3843 & n5734 ) | ( n3843 & n5736 ) | ( n5734 & n5736 ) ;
  assign n5738 = ( x45 & ~n4394 ) | ( x45 & n4745 ) | ( ~n4394 & n4745 ) ;
  assign n5739 = ( n571 & n873 ) | ( n571 & ~n893 ) | ( n873 & ~n893 ) ;
  assign n5740 = ( n2336 & n5738 ) | ( n2336 & n5739 ) | ( n5738 & n5739 ) ;
  assign n5741 = n2450 ^ n1539 ^ n469 ;
  assign n5742 = n5741 ^ n4544 ^ n1778 ;
  assign n5743 = ( n1770 & n2202 ) | ( n1770 & n5742 ) | ( n2202 & n5742 ) ;
  assign n5744 = n1056 ^ n992 ^ 1'b0 ;
  assign n5745 = ~n4320 & n5744 ;
  assign n5746 = ( n1779 & n1959 ) | ( n1779 & ~n5745 ) | ( n1959 & ~n5745 ) ;
  assign n5747 = n5746 ^ x33 ^ 1'b0 ;
  assign n5748 = ~n4581 & n5747 ;
  assign n5749 = ( n1392 & ~n4275 ) | ( n1392 & n5748 ) | ( ~n4275 & n5748 ) ;
  assign n5750 = ( ~n3590 & n5743 ) | ( ~n3590 & n5749 ) | ( n5743 & n5749 ) ;
  assign n5751 = n1694 ^ n1473 ^ x92 ;
  assign n5752 = ( n3700 & n4095 ) | ( n3700 & n5751 ) | ( n4095 & n5751 ) ;
  assign n5753 = ( ~n485 & n647 ) | ( ~n485 & n5752 ) | ( n647 & n5752 ) ;
  assign n5754 = n371 | n3304 ;
  assign n5755 = n1498 & ~n3893 ;
  assign n5756 = ( n505 & n583 ) | ( n505 & n5755 ) | ( n583 & n5755 ) ;
  assign n5757 = n5756 ^ n1109 ^ n682 ;
  assign n5758 = ( x234 & n3319 ) | ( x234 & n4105 ) | ( n3319 & n4105 ) ;
  assign n5759 = n5758 ^ n4018 ^ 1'b0 ;
  assign n5760 = ( n398 & n3404 ) | ( n398 & ~n5759 ) | ( n3404 & ~n5759 ) ;
  assign n5761 = ( n5754 & n5757 ) | ( n5754 & n5760 ) | ( n5757 & n5760 ) ;
  assign n5762 = ( n3412 & ~n3441 ) | ( n3412 & n5543 ) | ( ~n3441 & n5543 ) ;
  assign n5763 = ( n5753 & n5761 ) | ( n5753 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5764 = ( n5740 & ~n5750 ) | ( n5740 & n5763 ) | ( ~n5750 & n5763 ) ;
  assign n5765 = ( n5733 & ~n5737 ) | ( n5733 & n5764 ) | ( ~n5737 & n5764 ) ;
  assign n5767 = ( x233 & n900 ) | ( x233 & ~n1656 ) | ( n900 & ~n1656 ) ;
  assign n5766 = n5700 ^ n2412 ^ n1392 ;
  assign n5768 = n5767 ^ n5766 ^ n2483 ;
  assign n5769 = n2031 ^ n1276 ^ 1'b0 ;
  assign n5770 = ( n4042 & ~n5768 ) | ( n4042 & n5769 ) | ( ~n5768 & n5769 ) ;
  assign n5777 = n1934 ^ n1670 ^ 1'b0 ;
  assign n5775 = ( n419 & ~n2580 ) | ( n419 & n2765 ) | ( ~n2580 & n2765 ) ;
  assign n5776 = n258 & n5775 ;
  assign n5778 = n5777 ^ n5776 ^ n2555 ;
  assign n5779 = n5778 ^ n5287 ^ n597 ;
  assign n5771 = n2589 & ~n3628 ;
  assign n5772 = n4338 & n5771 ;
  assign n5773 = n4988 | n5772 ;
  assign n5774 = n2838 & ~n5773 ;
  assign n5780 = n5779 ^ n5774 ^ 1'b0 ;
  assign n5781 = ( n1492 & n5770 ) | ( n1492 & n5780 ) | ( n5770 & n5780 ) ;
  assign n5782 = ( ~x15 & n1450 ) | ( ~x15 & n2396 ) | ( n1450 & n2396 ) ;
  assign n5783 = n5782 ^ n5379 ^ n734 ;
  assign n5784 = ( n1030 & n5699 ) | ( n1030 & ~n5783 ) | ( n5699 & ~n5783 ) ;
  assign n5785 = ( n3194 & ~n4331 ) | ( n3194 & n5784 ) | ( ~n4331 & n5784 ) ;
  assign n5786 = ( ~n3651 & n4207 ) | ( ~n3651 & n5204 ) | ( n4207 & n5204 ) ;
  assign n5787 = ( n3789 & n5109 ) | ( n3789 & ~n5786 ) | ( n5109 & ~n5786 ) ;
  assign n5788 = n5787 ^ n2033 ^ n538 ;
  assign n5792 = ( n1437 & n1912 ) | ( n1437 & n4391 ) | ( n1912 & n4391 ) ;
  assign n5789 = ~n854 & n5699 ;
  assign n5790 = n5789 ^ n1308 ^ 1'b0 ;
  assign n5791 = n5790 ^ n4728 ^ n2239 ;
  assign n5793 = n5792 ^ n5791 ^ 1'b0 ;
  assign n5795 = ( n3081 & n4196 ) | ( n3081 & n5748 ) | ( n4196 & n5748 ) ;
  assign n5796 = n2152 & ~n5795 ;
  assign n5798 = ( n1182 & n1655 ) | ( n1182 & n1711 ) | ( n1655 & n1711 ) ;
  assign n5799 = n2260 | n5798 ;
  assign n5797 = n1708 & ~n2160 ;
  assign n5800 = n5799 ^ n5797 ^ 1'b0 ;
  assign n5801 = n5800 ^ n1899 ^ n720 ;
  assign n5802 = ( ~n4655 & n5796 ) | ( ~n4655 & n5801 ) | ( n5796 & n5801 ) ;
  assign n5794 = ( ~x16 & n2825 ) | ( ~x16 & n4593 ) | ( n2825 & n4593 ) ;
  assign n5803 = n5802 ^ n5794 ^ n3740 ;
  assign n5804 = ( n264 & n2200 ) | ( n264 & ~n4415 ) | ( n2200 & ~n4415 ) ;
  assign n5805 = ( n1350 & ~n2246 ) | ( n1350 & n5804 ) | ( ~n2246 & n5804 ) ;
  assign n5806 = ( n4196 & n5803 ) | ( n4196 & n5805 ) | ( n5803 & n5805 ) ;
  assign n5807 = ( n257 & n1368 ) | ( n257 & n3284 ) | ( n1368 & n3284 ) ;
  assign n5808 = ( n2116 & ~n2879 ) | ( n2116 & n5807 ) | ( ~n2879 & n5807 ) ;
  assign n5809 = n4070 ^ n2480 ^ n999 ;
  assign n5810 = n3290 | n5809 ;
  assign n5811 = n423 & ~n5810 ;
  assign n5812 = n5808 & ~n5811 ;
  assign n5813 = n5812 ^ n985 ^ 1'b0 ;
  assign n5814 = n3863 ^ n1866 ^ 1'b0 ;
  assign n5815 = ( n438 & ~n5813 ) | ( n438 & n5814 ) | ( ~n5813 & n5814 ) ;
  assign n5816 = n2635 ^ n2613 ^ n494 ;
  assign n5817 = ( n4717 & ~n4795 ) | ( n4717 & n5816 ) | ( ~n4795 & n5816 ) ;
  assign n5818 = ( n956 & ~n4038 ) | ( n956 & n5817 ) | ( ~n4038 & n5817 ) ;
  assign n5819 = ( ~n3854 & n4880 ) | ( ~n3854 & n5818 ) | ( n4880 & n5818 ) ;
  assign n5820 = n5279 & n5819 ;
  assign n5821 = ( n2664 & n3698 ) | ( n2664 & ~n3815 ) | ( n3698 & ~n3815 ) ;
  assign n5822 = ( n726 & ~n1580 ) | ( n726 & n2776 ) | ( ~n1580 & n2776 ) ;
  assign n5823 = ( n999 & ~n5821 ) | ( n999 & n5822 ) | ( ~n5821 & n5822 ) ;
  assign n5824 = x228 & ~n5823 ;
  assign n5825 = n561 & ~n3479 ;
  assign n5826 = n5825 ^ n273 ^ 1'b0 ;
  assign n5827 = ( n5388 & ~n5824 ) | ( n5388 & n5826 ) | ( ~n5824 & n5826 ) ;
  assign n5843 = n1802 ^ n661 ^ x94 ;
  assign n5842 = ( n1372 & n4668 ) | ( n1372 & ~n5780 ) | ( n4668 & ~n5780 ) ;
  assign n5829 = n1405 ^ n287 ^ x159 ;
  assign n5830 = n5829 ^ n2586 ^ 1'b0 ;
  assign n5831 = n1380 & n5830 ;
  assign n5828 = n4336 ^ n1735 ^ n753 ;
  assign n5832 = n5831 ^ n5828 ^ n4168 ;
  assign n5833 = ( n1705 & ~n2146 ) | ( n1705 & n2698 ) | ( ~n2146 & n2698 ) ;
  assign n5834 = n1379 | n2821 ;
  assign n5835 = ( ~n1130 & n1655 ) | ( ~n1130 & n5834 ) | ( n1655 & n5834 ) ;
  assign n5836 = n5835 ^ n2366 ^ x237 ;
  assign n5837 = n4905 ^ n4542 ^ n1006 ;
  assign n5838 = ( n3458 & n5836 ) | ( n3458 & ~n5837 ) | ( n5836 & ~n5837 ) ;
  assign n5839 = ~n2100 & n5838 ;
  assign n5840 = n5833 & n5839 ;
  assign n5841 = n5832 & ~n5840 ;
  assign n5844 = n5843 ^ n5842 ^ n5841 ;
  assign n5853 = n2219 & ~n4370 ;
  assign n5849 = ( n1078 & n1816 ) | ( n1078 & n3470 ) | ( n1816 & n3470 ) ;
  assign n5850 = ( n1029 & n1048 ) | ( n1029 & ~n5849 ) | ( n1048 & ~n5849 ) ;
  assign n5846 = n788 ^ n565 ^ 1'b0 ;
  assign n5847 = n847 & ~n5846 ;
  assign n5845 = ( n682 & ~n2915 ) | ( n682 & n3095 ) | ( ~n2915 & n3095 ) ;
  assign n5848 = n5847 ^ n5845 ^ n2220 ;
  assign n5851 = n5850 ^ n5848 ^ n2743 ;
  assign n5852 = ~n5596 & n5851 ;
  assign n5854 = n5853 ^ n5852 ^ n5837 ;
  assign n5855 = n949 | n990 ;
  assign n5856 = ( ~n2062 & n2602 ) | ( ~n2062 & n5855 ) | ( n2602 & n5855 ) ;
  assign n5857 = ( x77 & n1158 ) | ( x77 & n5856 ) | ( n1158 & n5856 ) ;
  assign n5858 = ( n452 & ~n2829 ) | ( n452 & n5857 ) | ( ~n2829 & n5857 ) ;
  assign n5859 = n5858 ^ n5750 ^ n4254 ;
  assign n5868 = n3797 ^ n2067 ^ 1'b0 ;
  assign n5869 = ~n1868 & n5868 ;
  assign n5870 = ~n2403 & n5461 ;
  assign n5871 = ( ~n433 & n5869 ) | ( ~n433 & n5870 ) | ( n5869 & n5870 ) ;
  assign n5863 = n3008 ^ n2586 ^ n805 ;
  assign n5864 = ( ~n728 & n1530 ) | ( ~n728 & n5863 ) | ( n1530 & n5863 ) ;
  assign n5865 = n5864 ^ n3706 ^ n2286 ;
  assign n5861 = n1836 ^ n597 ^ 1'b0 ;
  assign n5862 = n5577 & n5861 ;
  assign n5860 = ( n1367 & n1944 ) | ( n1367 & n5624 ) | ( n1944 & n5624 ) ;
  assign n5866 = n5865 ^ n5862 ^ n5860 ;
  assign n5867 = n5866 ^ n4051 ^ n3735 ;
  assign n5872 = n5871 ^ n5867 ^ n2043 ;
  assign n5873 = ( n1244 & ~n5859 ) | ( n1244 & n5872 ) | ( ~n5859 & n5872 ) ;
  assign n5874 = ( n681 & n828 ) | ( n681 & ~n2430 ) | ( n828 & ~n2430 ) ;
  assign n5875 = ( n1464 & ~n1538 ) | ( n1464 & n5492 ) | ( ~n1538 & n5492 ) ;
  assign n5876 = n5767 ^ n4935 ^ n1954 ;
  assign n5877 = ( x41 & n962 ) | ( x41 & n5876 ) | ( n962 & n5876 ) ;
  assign n5878 = ( n5874 & ~n5875 ) | ( n5874 & n5877 ) | ( ~n5875 & n5877 ) ;
  assign n5879 = n5878 ^ n5743 ^ n342 ;
  assign n5880 = ( n1471 & n1745 ) | ( n1471 & n1817 ) | ( n1745 & n1817 ) ;
  assign n5881 = n5880 ^ n955 ^ n763 ;
  assign n5882 = ( n1463 & n1667 ) | ( n1463 & ~n2366 ) | ( n1667 & ~n2366 ) ;
  assign n5883 = n5882 ^ n932 ^ n491 ;
  assign n5884 = ( n1009 & n1522 ) | ( n1009 & ~n2739 ) | ( n1522 & ~n2739 ) ;
  assign n5885 = n5883 & n5884 ;
  assign n5889 = n1106 & ~n1252 ;
  assign n5890 = ( n1339 & n4874 ) | ( n1339 & ~n5889 ) | ( n4874 & ~n5889 ) ;
  assign n5888 = ( x71 & n1711 ) | ( x71 & ~n4706 ) | ( n1711 & ~n4706 ) ;
  assign n5891 = n5890 ^ n5888 ^ n921 ;
  assign n5892 = ( ~n2291 & n2391 ) | ( ~n2291 & n5891 ) | ( n2391 & n5891 ) ;
  assign n5886 = ( n552 & n2804 ) | ( n552 & ~n5263 ) | ( n2804 & ~n5263 ) ;
  assign n5887 = n815 | n5886 ;
  assign n5893 = n5892 ^ n5887 ^ n768 ;
  assign n5894 = ( n5881 & n5885 ) | ( n5881 & ~n5893 ) | ( n5885 & ~n5893 ) ;
  assign n5895 = n2744 ^ n2256 ^ 1'b0 ;
  assign n5896 = n5581 ^ n5152 ^ n1786 ;
  assign n5897 = n4998 | n5896 ;
  assign n5898 = ( n2324 & n5895 ) | ( n2324 & ~n5897 ) | ( n5895 & ~n5897 ) ;
  assign n5899 = n5339 ^ n3572 ^ n2185 ;
  assign n5900 = ( n671 & n1488 ) | ( n671 & n2459 ) | ( n1488 & n2459 ) ;
  assign n5901 = n888 & n5123 ;
  assign n5902 = ( n5705 & n5900 ) | ( n5705 & n5901 ) | ( n5900 & n5901 ) ;
  assign n5903 = ~n5899 & n5902 ;
  assign n5904 = n5666 ^ n1887 ^ 1'b0 ;
  assign n5905 = n4135 ^ n3131 ^ n886 ;
  assign n5906 = n5905 ^ n5535 ^ n1351 ;
  assign n5907 = n3423 ^ n1611 ^ 1'b0 ;
  assign n5908 = n5907 ^ n1732 ^ 1'b0 ;
  assign n5909 = ( n2440 & n3346 ) | ( n2440 & n5908 ) | ( n3346 & n5908 ) ;
  assign n5913 = n2389 ^ n1983 ^ n321 ;
  assign n5914 = n5913 ^ n1866 ^ 1'b0 ;
  assign n5915 = ( n428 & n3901 ) | ( n428 & ~n5914 ) | ( n3901 & ~n5914 ) ;
  assign n5920 = ( ~x217 & n882 ) | ( ~x217 & n2212 ) | ( n882 & n2212 ) ;
  assign n5921 = n5920 ^ n2478 ^ n1497 ;
  assign n5919 = n5455 ^ n1062 ^ n876 ;
  assign n5916 = ( x1 & ~n1693 ) | ( x1 & n3286 ) | ( ~n1693 & n3286 ) ;
  assign n5917 = n2956 ^ n2164 ^ n647 ;
  assign n5918 = ( ~n1356 & n5916 ) | ( ~n1356 & n5917 ) | ( n5916 & n5917 ) ;
  assign n5922 = n5921 ^ n5919 ^ n5918 ;
  assign n5923 = ( n2978 & n5915 ) | ( n2978 & ~n5922 ) | ( n5915 & ~n5922 ) ;
  assign n5910 = ( ~n578 & n1702 ) | ( ~n578 & n2780 ) | ( n1702 & n2780 ) ;
  assign n5911 = ( n858 & n3785 ) | ( n858 & ~n3907 ) | ( n3785 & ~n3907 ) ;
  assign n5912 = ( n702 & n5910 ) | ( n702 & ~n5911 ) | ( n5910 & ~n5911 ) ;
  assign n5924 = n5923 ^ n5912 ^ x122 ;
  assign n5925 = n5277 ^ n1374 ^ n733 ;
  assign n5926 = n2552 | n5925 ;
  assign n5927 = ( n3417 & n4848 ) | ( n3417 & n5926 ) | ( n4848 & n5926 ) ;
  assign n5928 = n5927 ^ n4042 ^ n2942 ;
  assign n5935 = n2850 ^ n1575 ^ n1000 ;
  assign n5929 = n2523 | n3511 ;
  assign n5930 = n5929 ^ n3893 ^ n3192 ;
  assign n5931 = n3040 ^ n885 ^ x113 ;
  assign n5932 = n5931 ^ n3184 ^ 1'b0 ;
  assign n5933 = n5930 & n5932 ;
  assign n5934 = ~n4481 & n5933 ;
  assign n5936 = n5935 ^ n5934 ^ n5060 ;
  assign n5941 = n4375 ^ n2760 ^ n852 ;
  assign n5942 = ( x39 & n5481 ) | ( x39 & n5941 ) | ( n5481 & n5941 ) ;
  assign n5937 = ~n1778 & n4904 ;
  assign n5938 = n5937 ^ n491 ^ 1'b0 ;
  assign n5939 = n3475 & ~n3859 ;
  assign n5940 = n5938 & n5939 ;
  assign n5943 = n5942 ^ n5940 ^ n770 ;
  assign n5944 = n804 & n2044 ;
  assign n5945 = n4749 & n5944 ;
  assign n5946 = n5945 ^ n1772 ^ 1'b0 ;
  assign n5947 = n5946 ^ n2835 ^ n2302 ;
  assign n5948 = n2921 ^ n1165 ^ 1'b0 ;
  assign n5949 = n5948 ^ n4897 ^ n453 ;
  assign n5950 = ( n898 & n5947 ) | ( n898 & n5949 ) | ( n5947 & n5949 ) ;
  assign n5973 = n2306 ^ n2020 ^ n1303 ;
  assign n5951 = n3759 ^ n3116 ^ 1'b0 ;
  assign n5969 = n1531 & n1541 ;
  assign n5961 = ( ~n520 & n2679 ) | ( ~n520 & n5013 ) | ( n2679 & n5013 ) ;
  assign n5962 = ( n1848 & n5889 ) | ( n1848 & n5961 ) | ( n5889 & n5961 ) ;
  assign n5963 = n317 & n2597 ;
  assign n5964 = n5963 ^ x87 ^ 1'b0 ;
  assign n5965 = n5964 ^ n3310 ^ n904 ;
  assign n5966 = ( n1555 & n5962 ) | ( n1555 & ~n5965 ) | ( n5962 & ~n5965 ) ;
  assign n5967 = n5966 ^ n2494 ^ 1'b0 ;
  assign n5968 = n2690 & n5967 ;
  assign n5970 = n5969 ^ n5968 ^ n1984 ;
  assign n5953 = n995 ^ x47 ^ 1'b0 ;
  assign n5955 = n1311 ^ n1142 ^ n649 ;
  assign n5954 = n5741 ^ n3766 ^ n888 ;
  assign n5956 = n5955 ^ n5954 ^ n5030 ;
  assign n5957 = ( n341 & n5953 ) | ( n341 & n5956 ) | ( n5953 & n5956 ) ;
  assign n5952 = n3267 | n4423 ;
  assign n5958 = n5957 ^ n5952 ^ 1'b0 ;
  assign n5959 = n5958 ^ n3700 ^ n2377 ;
  assign n5960 = n5959 ^ n4810 ^ n2470 ;
  assign n5971 = n5970 ^ n5960 ^ n968 ;
  assign n5972 = ( n3407 & ~n5951 ) | ( n3407 & n5971 ) | ( ~n5951 & n5971 ) ;
  assign n5974 = n5973 ^ n5972 ^ x0 ;
  assign n5975 = n5974 ^ n2704 ^ 1'b0 ;
  assign n5976 = n4031 ^ n2705 ^ n851 ;
  assign n5977 = ( ~n2220 & n2940 ) | ( ~n2220 & n5976 ) | ( n2940 & n5976 ) ;
  assign n5985 = n3723 ^ n2831 ^ n602 ;
  assign n5978 = n5289 ^ x159 ^ 1'b0 ;
  assign n5979 = n500 & ~n5978 ;
  assign n5980 = n5979 ^ n5560 ^ n1143 ;
  assign n5981 = ( ~n1341 & n3457 ) | ( ~n1341 & n4835 ) | ( n3457 & n4835 ) ;
  assign n5982 = n1899 & n5981 ;
  assign n5983 = ~n1565 & n5982 ;
  assign n5984 = ( x138 & n5980 ) | ( x138 & ~n5983 ) | ( n5980 & ~n5983 ) ;
  assign n5986 = n5985 ^ n5984 ^ n342 ;
  assign n5987 = n5179 ^ n2844 ^ x233 ;
  assign n5988 = n5987 ^ n3345 ^ n1532 ;
  assign n5989 = n4377 ^ n3872 ^ n1210 ;
  assign n5990 = n5989 ^ n2634 ^ n605 ;
  assign n5991 = ( n1522 & n3991 ) | ( n1522 & n5990 ) | ( n3991 & n5990 ) ;
  assign n5992 = ~n298 & n2344 ;
  assign n5993 = n5992 ^ n4347 ^ 1'b0 ;
  assign n5994 = ( n658 & n3323 ) | ( n658 & ~n5993 ) | ( n3323 & ~n5993 ) ;
  assign n5997 = ( n475 & n1088 ) | ( n475 & n2166 ) | ( n1088 & n2166 ) ;
  assign n5996 = n1220 | n2611 ;
  assign n5998 = n5997 ^ n5996 ^ n5805 ;
  assign n5995 = n4718 ^ n3950 ^ n1239 ;
  assign n5999 = n5998 ^ n5995 ^ 1'b0 ;
  assign n6000 = n5994 | n5999 ;
  assign n6001 = ( n282 & ~n524 ) | ( n282 & n2452 ) | ( ~n524 & n2452 ) ;
  assign n6002 = ( n668 & ~n2388 ) | ( n668 & n6001 ) | ( ~n2388 & n6001 ) ;
  assign n6003 = n6002 ^ n2936 ^ n2922 ;
  assign n6004 = ( n1899 & n4563 ) | ( n1899 & n6003 ) | ( n4563 & n6003 ) ;
  assign n6005 = n6004 ^ n5973 ^ x243 ;
  assign n6007 = n2767 ^ n2192 ^ 1'b0 ;
  assign n6008 = ( ~n349 & n2457 ) | ( ~n349 & n6007 ) | ( n2457 & n6007 ) ;
  assign n6009 = n4214 ^ n2654 ^ n2158 ;
  assign n6010 = n6009 ^ n3195 ^ n899 ;
  assign n6011 = n6010 ^ n2049 ^ n804 ;
  assign n6012 = n6008 & n6011 ;
  assign n6013 = n6012 ^ n3449 ^ 1'b0 ;
  assign n6006 = n880 & n4342 ;
  assign n6014 = n6013 ^ n6006 ^ 1'b0 ;
  assign n6015 = ( n2440 & n3440 ) | ( n2440 & n6014 ) | ( n3440 & n6014 ) ;
  assign n6026 = ~n1655 & n2316 ;
  assign n6027 = n6026 ^ n3625 ^ 1'b0 ;
  assign n6024 = n1722 & n3417 ;
  assign n6025 = n6024 ^ n5675 ^ 1'b0 ;
  assign n6028 = n6027 ^ n6025 ^ n5665 ;
  assign n6029 = n1562 ^ n1229 ^ 1'b0 ;
  assign n6030 = ( ~n2575 & n6028 ) | ( ~n2575 & n6029 ) | ( n6028 & n6029 ) ;
  assign n6018 = n1803 ^ n1677 ^ n843 ;
  assign n6019 = n2204 ^ n1579 ^ n1154 ;
  assign n6020 = ( n965 & n6018 ) | ( n965 & n6019 ) | ( n6018 & n6019 ) ;
  assign n6021 = n6020 ^ n4415 ^ n1415 ;
  assign n6022 = n6021 ^ n1976 ^ n1968 ;
  assign n6016 = ( n1750 & n2488 ) | ( n1750 & ~n4184 ) | ( n2488 & ~n4184 ) ;
  assign n6017 = ( x74 & n1151 ) | ( x74 & n6016 ) | ( n1151 & n6016 ) ;
  assign n6023 = n6022 ^ n6017 ^ n2849 ;
  assign n6031 = n6030 ^ n6023 ^ n4544 ;
  assign n6038 = n4340 ^ n3464 ^ n972 ;
  assign n6039 = n1556 ^ n1418 ^ n1001 ;
  assign n6040 = n2326 & ~n6039 ;
  assign n6041 = ( x47 & n421 ) | ( x47 & n6040 ) | ( n421 & n6040 ) ;
  assign n6042 = ( n1770 & n6038 ) | ( n1770 & ~n6041 ) | ( n6038 & ~n6041 ) ;
  assign n6043 = n4441 & ~n6042 ;
  assign n6044 = n2795 & n6043 ;
  assign n6032 = n1256 & ~n1739 ;
  assign n6033 = ~n2774 & n6032 ;
  assign n6034 = n6033 ^ n1499 ^ x18 ;
  assign n6035 = n6034 ^ n5397 ^ n1112 ;
  assign n6036 = n3968 ^ n2115 ^ 1'b0 ;
  assign n6037 = n6035 & n6036 ;
  assign n6045 = n6044 ^ n6037 ^ 1'b0 ;
  assign n6046 = n2329 ^ n1416 ^ 1'b0 ;
  assign n6047 = ( n1704 & n4448 ) | ( n1704 & ~n6046 ) | ( n4448 & ~n6046 ) ;
  assign n6049 = n2356 ^ n1233 ^ n1139 ;
  assign n6050 = n6049 ^ n2375 ^ n2155 ;
  assign n6048 = n3390 ^ n1851 ^ n848 ;
  assign n6051 = n6050 ^ n6048 ^ n4636 ;
  assign n6052 = n925 & n6051 ;
  assign n6055 = n2758 ^ n1362 ^ x195 ;
  assign n6054 = n3739 & n4528 ;
  assign n6056 = n6055 ^ n6054 ^ 1'b0 ;
  assign n6053 = ( ~n758 & n1213 ) | ( ~n758 & n1460 ) | ( n1213 & n1460 ) ;
  assign n6057 = n6056 ^ n6053 ^ n386 ;
  assign n6058 = ( ~x118 & n6052 ) | ( ~x118 & n6057 ) | ( n6052 & n6057 ) ;
  assign n6059 = x42 & ~n831 ;
  assign n6060 = ~n3043 & n6059 ;
  assign n6064 = n5786 ^ n4370 ^ x226 ;
  assign n6061 = n5481 ^ n1107 ^ 1'b0 ;
  assign n6062 = n6061 ^ n5278 ^ 1'b0 ;
  assign n6063 = n6062 ^ n5220 ^ 1'b0 ;
  assign n6065 = n6064 ^ n6063 ^ n5935 ;
  assign n6068 = n2342 ^ n427 ^ x106 ;
  assign n6066 = n3116 ^ n1500 ^ n981 ;
  assign n6067 = ( n1494 & n4305 ) | ( n1494 & ~n6066 ) | ( n4305 & ~n6066 ) ;
  assign n6069 = n6068 ^ n6067 ^ n4978 ;
  assign n6070 = ( n1631 & ~n4404 ) | ( n1631 & n5387 ) | ( ~n4404 & n5387 ) ;
  assign n6071 = n6070 ^ n1870 ^ n1292 ;
  assign n6072 = ( ~x85 & n2497 ) | ( ~x85 & n6071 ) | ( n2497 & n6071 ) ;
  assign n6073 = n6072 ^ n2722 ^ n1509 ;
  assign n6091 = n2878 ^ x223 ^ x166 ;
  assign n6092 = ( n4303 & n4473 ) | ( n4303 & n6091 ) | ( n4473 & n6091 ) ;
  assign n6093 = ( ~x178 & n1984 ) | ( ~x178 & n6092 ) | ( n1984 & n6092 ) ;
  assign n6094 = n6093 ^ n4069 ^ n3897 ;
  assign n6095 = n6094 ^ n2881 ^ n2373 ;
  assign n6089 = n3320 ^ n1664 ^ n524 ;
  assign n6090 = n6089 ^ n5216 ^ n2163 ;
  assign n6087 = ( ~n1737 & n2309 ) | ( ~n1737 & n3820 ) | ( n2309 & n3820 ) ;
  assign n6088 = n6087 ^ n2956 ^ n682 ;
  assign n6096 = n6095 ^ n6090 ^ n6088 ;
  assign n6097 = ( n3994 & ~n5312 ) | ( n3994 & n6096 ) | ( ~n5312 & n6096 ) ;
  assign n6082 = ( n2793 & n4464 ) | ( n2793 & ~n4746 ) | ( n4464 & ~n4746 ) ;
  assign n6083 = n929 | n2330 ;
  assign n6084 = n6082 | n6083 ;
  assign n6085 = n6084 ^ n5141 ^ n4917 ;
  assign n6076 = ( n846 & n2253 ) | ( n846 & n2390 ) | ( n2253 & n2390 ) ;
  assign n6075 = ( n856 & n2131 ) | ( n856 & ~n2240 ) | ( n2131 & ~n2240 ) ;
  assign n6077 = n6076 ^ n6075 ^ n3168 ;
  assign n6078 = n5809 ^ n4830 ^ n580 ;
  assign n6079 = ( x113 & ~n5818 ) | ( x113 & n6078 ) | ( ~n5818 & n6078 ) ;
  assign n6080 = n6079 ^ n4474 ^ n3873 ;
  assign n6081 = ( n3811 & n6077 ) | ( n3811 & n6080 ) | ( n6077 & n6080 ) ;
  assign n6074 = ( ~n365 & n2172 ) | ( ~n365 & n3391 ) | ( n2172 & n3391 ) ;
  assign n6086 = n6085 ^ n6081 ^ n6074 ;
  assign n6098 = n6097 ^ n6086 ^ n2370 ;
  assign n6099 = n2022 | n3835 ;
  assign n6100 = ( n327 & n1855 ) | ( n327 & n2235 ) | ( n1855 & n2235 ) ;
  assign n6101 = n6100 ^ n5674 ^ n3788 ;
  assign n6102 = n6099 | n6101 ;
  assign n6107 = x93 & ~n2248 ;
  assign n6108 = n6107 ^ n726 ^ 1'b0 ;
  assign n6103 = n1567 & n5515 ;
  assign n6104 = ( n349 & ~n801 ) | ( n349 & n2122 ) | ( ~n801 & n2122 ) ;
  assign n6105 = ( n2493 & ~n6103 ) | ( n2493 & n6104 ) | ( ~n6103 & n6104 ) ;
  assign n6106 = n6105 ^ n3963 ^ n721 ;
  assign n6109 = n6108 ^ n6106 ^ n4063 ;
  assign n6115 = n4943 ^ n1836 ^ 1'b0 ;
  assign n6116 = ( x131 & n909 ) | ( x131 & ~n6115 ) | ( n909 & ~n6115 ) ;
  assign n6111 = n2937 & ~n3815 ;
  assign n6112 = ~n325 & n6111 ;
  assign n6110 = n5688 ^ n2382 ^ n493 ;
  assign n6113 = n6112 ^ n6110 ^ 1'b0 ;
  assign n6114 = n6113 ^ n2999 ^ n2774 ;
  assign n6117 = n6116 ^ n6114 ^ n3493 ;
  assign n6118 = ( n311 & n2068 ) | ( n311 & ~n3963 ) | ( n2068 & ~n3963 ) ;
  assign n6119 = n3547 ^ n3013 ^ n1350 ;
  assign n6120 = n6119 ^ n2749 ^ 1'b0 ;
  assign n6121 = ( n1892 & n5327 ) | ( n1892 & n6120 ) | ( n5327 & n6120 ) ;
  assign n6122 = n2759 ^ n2731 ^ x30 ;
  assign n6123 = ( n521 & ~n4638 ) | ( n521 & n6122 ) | ( ~n4638 & n6122 ) ;
  assign n6124 = n6123 ^ n1563 ^ n1534 ;
  assign n6125 = n3382 & n3809 ;
  assign n6126 = n6125 ^ n5051 ^ 1'b0 ;
  assign n6127 = n1613 | n6126 ;
  assign n6128 = ( ~n6121 & n6124 ) | ( ~n6121 & n6127 ) | ( n6124 & n6127 ) ;
  assign n6129 = ( ~n2857 & n4129 ) | ( ~n2857 & n6128 ) | ( n4129 & n6128 ) ;
  assign n6130 = ( ~n6117 & n6118 ) | ( ~n6117 & n6129 ) | ( n6118 & n6129 ) ;
  assign n6131 = ( n1281 & n1511 ) | ( n1281 & n2308 ) | ( n1511 & n2308 ) ;
  assign n6132 = n1337 & n6131 ;
  assign n6133 = n326 & n2098 ;
  assign n6134 = n2883 & ~n6133 ;
  assign n6135 = n4109 & n6134 ;
  assign n6137 = ( n710 & n1294 ) | ( n710 & n5340 ) | ( n1294 & n5340 ) ;
  assign n6136 = n5283 ^ n4468 ^ x226 ;
  assign n6138 = n6137 ^ n6136 ^ n296 ;
  assign n6139 = n6138 ^ n3977 ^ n2850 ;
  assign n6140 = ( n6132 & n6135 ) | ( n6132 & ~n6139 ) | ( n6135 & ~n6139 ) ;
  assign n6147 = n2783 ^ n1387 ^ x145 ;
  assign n6148 = n6147 ^ n2944 ^ n1688 ;
  assign n6149 = ( n259 & n2052 ) | ( n259 & ~n3000 ) | ( n2052 & ~n3000 ) ;
  assign n6150 = ( n2139 & n6148 ) | ( n2139 & ~n6149 ) | ( n6148 & ~n6149 ) ;
  assign n6143 = n3865 ^ n2914 ^ x46 ;
  assign n6141 = ( n511 & n1469 ) | ( n511 & ~n6123 ) | ( n1469 & ~n6123 ) ;
  assign n6142 = ( n1004 & n1423 ) | ( n1004 & ~n6141 ) | ( n1423 & ~n6141 ) ;
  assign n6144 = n6143 ^ n6142 ^ 1'b0 ;
  assign n6145 = n6144 ^ n5536 ^ n1981 ;
  assign n6146 = n1358 & n6145 ;
  assign n6151 = n6150 ^ n6146 ^ 1'b0 ;
  assign n6155 = n4588 ^ n3614 ^ n2166 ;
  assign n6156 = n6155 ^ n3843 ^ n2102 ;
  assign n6152 = n3246 ^ n349 ^ x121 ;
  assign n6153 = n6152 ^ n1994 ^ 1'b0 ;
  assign n6154 = n3042 | n6153 ;
  assign n6157 = n6156 ^ n6154 ^ x103 ;
  assign n6179 = x28 & n1897 ;
  assign n6180 = n2577 & n6179 ;
  assign n6177 = n5180 ^ n2892 ^ x160 ;
  assign n6172 = n2722 ^ x254 ^ x214 ;
  assign n6173 = ( n1335 & n2316 ) | ( n1335 & ~n6172 ) | ( n2316 & ~n6172 ) ;
  assign n6174 = ( n354 & ~n1057 ) | ( n354 & n6173 ) | ( ~n1057 & n6173 ) ;
  assign n6175 = ( ~n2494 & n5237 ) | ( ~n2494 & n6174 ) | ( n5237 & n6174 ) ;
  assign n6176 = ( ~n4357 & n4398 ) | ( ~n4357 & n6175 ) | ( n4398 & n6175 ) ;
  assign n6168 = n587 | n3322 ;
  assign n6169 = n6168 ^ n5832 ^ n654 ;
  assign n6170 = n6169 ^ n2717 ^ n1924 ;
  assign n6171 = n6170 ^ n1042 ^ n724 ;
  assign n6178 = n6177 ^ n6176 ^ n6171 ;
  assign n6158 = n1095 ^ n690 ^ n378 ;
  assign n6159 = n6158 ^ n936 ^ 1'b0 ;
  assign n6160 = ~n1804 & n6159 ;
  assign n6164 = n3067 ^ n2511 ^ n856 ;
  assign n6165 = ( n4692 & n4948 ) | ( n4692 & n6164 ) | ( n4948 & n6164 ) ;
  assign n6161 = ( x119 & n2473 ) | ( x119 & n4452 ) | ( n2473 & n4452 ) ;
  assign n6162 = n6161 ^ n5748 ^ n1362 ;
  assign n6163 = n3600 | n6162 ;
  assign n6166 = n6165 ^ n6163 ^ 1'b0 ;
  assign n6167 = ( ~x41 & n6160 ) | ( ~x41 & n6166 ) | ( n6160 & n6166 ) ;
  assign n6181 = n6180 ^ n6178 ^ n6167 ;
  assign n6182 = ( n4109 & ~n4217 ) | ( n4109 & n4885 ) | ( ~n4217 & n4885 ) ;
  assign n6183 = n2438 ^ n1828 ^ n1474 ;
  assign n6184 = n3552 | n6183 ;
  assign n6185 = n2372 | n6184 ;
  assign n6186 = n6185 ^ n3143 ^ 1'b0 ;
  assign n6187 = n1670 ^ x210 ^ 1'b0 ;
  assign n6188 = ( ~n6164 & n6186 ) | ( ~n6164 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6189 = n3095 ^ n1664 ^ n1014 ;
  assign n6190 = n491 ^ x244 ^ 1'b0 ;
  assign n6191 = ~n1817 & n6190 ;
  assign n6192 = n6191 ^ n3864 ^ n2173 ;
  assign n6193 = n1813 | n6192 ;
  assign n6194 = ( n1166 & n6189 ) | ( n1166 & ~n6193 ) | ( n6189 & ~n6193 ) ;
  assign n6195 = n6194 ^ n6170 ^ n905 ;
  assign n6196 = x36 ^ x13 ^ 1'b0 ;
  assign n6197 = n284 & n6196 ;
  assign n6198 = n6197 ^ n3968 ^ n374 ;
  assign n6199 = n6198 ^ n4211 ^ n1326 ;
  assign n6200 = n1471 ^ n1430 ^ n1343 ;
  assign n6201 = ( x66 & ~n834 ) | ( x66 & n936 ) | ( ~n834 & n936 ) ;
  assign n6202 = ( ~n2365 & n6200 ) | ( ~n2365 & n6201 ) | ( n6200 & n6201 ) ;
  assign n6203 = ~x111 & n491 ;
  assign n6204 = n903 & ~n1587 ;
  assign n6205 = n6203 & n6204 ;
  assign n6206 = ( n1329 & n3782 ) | ( n1329 & n6205 ) | ( n3782 & n6205 ) ;
  assign n6207 = ( n880 & n6202 ) | ( n880 & n6206 ) | ( n6202 & n6206 ) ;
  assign n6208 = n6207 ^ n3316 ^ n1710 ;
  assign n6209 = ( ~n4523 & n6199 ) | ( ~n4523 & n6208 ) | ( n6199 & n6208 ) ;
  assign n6210 = n1018 & n3589 ;
  assign n6211 = ~x20 & n6210 ;
  assign n6214 = n4079 ^ n522 ^ x11 ;
  assign n6212 = n321 & n2016 ;
  assign n6213 = n6212 ^ n3734 ^ 1'b0 ;
  assign n6215 = n6214 ^ n6213 ^ n3706 ;
  assign n6216 = n4466 ^ n4287 ^ n2328 ;
  assign n6217 = ( x242 & ~n885 ) | ( x242 & n1134 ) | ( ~n885 & n1134 ) ;
  assign n6218 = n6217 ^ n5255 ^ n2006 ;
  assign n6219 = ( ~n1877 & n3616 ) | ( ~n1877 & n6218 ) | ( n3616 & n6218 ) ;
  assign n6220 = ( n6215 & n6216 ) | ( n6215 & n6219 ) | ( n6216 & n6219 ) ;
  assign n6221 = ( n387 & ~n1983 ) | ( n387 & n2456 ) | ( ~n1983 & n2456 ) ;
  assign n6222 = n6221 ^ n1887 ^ x80 ;
  assign n6223 = n719 | n6222 ;
  assign n6224 = n5543 ^ n2859 ^ n2640 ;
  assign n6225 = ( n434 & ~n6223 ) | ( n434 & n6224 ) | ( ~n6223 & n6224 ) ;
  assign n6226 = n3124 ^ n1248 ^ n887 ;
  assign n6227 = ( ~n1827 & n1997 ) | ( ~n1827 & n2350 ) | ( n1997 & n2350 ) ;
  assign n6228 = ( n887 & n6226 ) | ( n887 & n6227 ) | ( n6226 & n6227 ) ;
  assign n6229 = ( x79 & n4679 ) | ( x79 & n6228 ) | ( n4679 & n6228 ) ;
  assign n6232 = n4145 ^ n1561 ^ n283 ;
  assign n6233 = ( ~x251 & n2922 ) | ( ~x251 & n4048 ) | ( n2922 & n4048 ) ;
  assign n6234 = ( ~x170 & n6232 ) | ( ~x170 & n6233 ) | ( n6232 & n6233 ) ;
  assign n6230 = ( n440 & n2510 ) | ( n440 & ~n2614 ) | ( n2510 & ~n2614 ) ;
  assign n6231 = ( n2878 & ~n4168 ) | ( n2878 & n6230 ) | ( ~n4168 & n6230 ) ;
  assign n6235 = n6234 ^ n6231 ^ n4076 ;
  assign n6241 = n1775 ^ n646 ^ n535 ;
  assign n6237 = n1803 ^ n801 ^ x211 ;
  assign n6236 = n388 & ~n1024 ;
  assign n6238 = n6237 ^ n6236 ^ 1'b0 ;
  assign n6239 = n6238 ^ n3300 ^ 1'b0 ;
  assign n6240 = ( ~n1233 & n1771 ) | ( ~n1233 & n6239 ) | ( n1771 & n6239 ) ;
  assign n6242 = n6241 ^ n6240 ^ n800 ;
  assign n6243 = ( n6229 & ~n6235 ) | ( n6229 & n6242 ) | ( ~n6235 & n6242 ) ;
  assign n6244 = n5662 ^ n4167 ^ n3245 ;
  assign n6245 = n6244 ^ n4864 ^ n4443 ;
  assign n6246 = ~n1686 & n6245 ;
  assign n6247 = n6246 ^ n5815 ^ 1'b0 ;
  assign n6248 = n2374 | n2736 ;
  assign n6249 = ( n538 & ~n1792 ) | ( n538 & n3593 ) | ( ~n1792 & n3593 ) ;
  assign n6253 = ( n838 & n2538 ) | ( n838 & ~n3552 ) | ( n2538 & ~n3552 ) ;
  assign n6254 = ( n1214 & n1395 ) | ( n1214 & ~n6253 ) | ( n1395 & ~n6253 ) ;
  assign n6255 = n3222 ^ n1318 ^ n910 ;
  assign n6256 = ( n5498 & ~n6254 ) | ( n5498 & n6255 ) | ( ~n6254 & n6255 ) ;
  assign n6257 = n6256 ^ n3724 ^ n2072 ;
  assign n6250 = n5040 ^ n2804 ^ n1443 ;
  assign n6251 = ( x128 & n523 ) | ( x128 & ~n4347 ) | ( n523 & ~n4347 ) ;
  assign n6252 = ( n5966 & ~n6250 ) | ( n5966 & n6251 ) | ( ~n6250 & n6251 ) ;
  assign n6258 = n6257 ^ n6252 ^ 1'b0 ;
  assign n6262 = ( x54 & n361 ) | ( x54 & n4487 ) | ( n361 & n4487 ) ;
  assign n6259 = n6254 ^ n2519 ^ 1'b0 ;
  assign n6260 = ( n849 & n1595 ) | ( n849 & n6259 ) | ( n1595 & n6259 ) ;
  assign n6261 = ( n2375 & n2521 ) | ( n2375 & ~n6260 ) | ( n2521 & ~n6260 ) ;
  assign n6263 = n6262 ^ n6261 ^ n1680 ;
  assign n6264 = n2783 ^ n1240 ^ n435 ;
  assign n6265 = ~n1654 & n6264 ;
  assign n6266 = n6263 & n6265 ;
  assign n6267 = ( ~n1601 & n2006 ) | ( ~n1601 & n6266 ) | ( n2006 & n6266 ) ;
  assign n6268 = n5500 ^ n2508 ^ 1'b0 ;
  assign n6269 = n5689 | n6268 ;
  assign n6270 = ~n6106 & n6269 ;
  assign n6271 = ( n3251 & n6267 ) | ( n3251 & ~n6270 ) | ( n6267 & ~n6270 ) ;
  assign n6272 = n2670 & ~n3887 ;
  assign n6273 = ( n3658 & ~n5388 ) | ( n3658 & n6272 ) | ( ~n5388 & n6272 ) ;
  assign n6276 = ( ~n343 & n741 ) | ( ~n343 & n3256 ) | ( n741 & n3256 ) ;
  assign n6277 = n6276 ^ n2974 ^ n2674 ;
  assign n6278 = ~n2245 & n3181 ;
  assign n6279 = n6278 ^ n1823 ^ 1'b0 ;
  assign n6280 = n5691 | n6279 ;
  assign n6281 = n6277 & ~n6280 ;
  assign n6274 = n4264 ^ n1688 ^ 1'b0 ;
  assign n6275 = ~n869 & n6274 ;
  assign n6282 = n6281 ^ n6275 ^ n5156 ;
  assign n6286 = ( ~n610 & n767 ) | ( ~n610 & n777 ) | ( n767 & n777 ) ;
  assign n6287 = ( ~n1426 & n5849 ) | ( ~n1426 & n6286 ) | ( n5849 & n6286 ) ;
  assign n6288 = ( x111 & ~n2451 ) | ( x111 & n6287 ) | ( ~n2451 & n6287 ) ;
  assign n6289 = n6288 ^ n5322 ^ n1452 ;
  assign n6284 = n5017 ^ n3859 ^ n2832 ;
  assign n6283 = ( n3848 & n4910 ) | ( n3848 & ~n6033 ) | ( n4910 & ~n6033 ) ;
  assign n6285 = n6284 ^ n6283 ^ n419 ;
  assign n6290 = n6289 ^ n6285 ^ n1673 ;
  assign n6294 = ( n663 & ~n684 ) | ( n663 & n2878 ) | ( ~n684 & n2878 ) ;
  assign n6295 = n5751 ^ n4832 ^ 1'b0 ;
  assign n6296 = n6294 & ~n6295 ;
  assign n6291 = ( ~n334 & n3856 ) | ( ~n334 & n4322 ) | ( n3856 & n4322 ) ;
  assign n6292 = n4029 ^ n1285 ^ n759 ;
  assign n6293 = ( n4218 & ~n6291 ) | ( n4218 & n6292 ) | ( ~n6291 & n6292 ) ;
  assign n6297 = n6296 ^ n6293 ^ 1'b0 ;
  assign n6298 = n4156 ^ n1473 ^ n315 ;
  assign n6299 = n6298 ^ n2596 ^ n1959 ;
  assign n6300 = n6299 ^ n1454 ^ n659 ;
  assign n6301 = n6300 ^ n1598 ^ n1217 ;
  assign n6302 = ( x92 & n367 ) | ( x92 & ~n4936 ) | ( n367 & ~n4936 ) ;
  assign n6303 = n4293 ^ n3329 ^ n1634 ;
  assign n6304 = ( n6301 & n6302 ) | ( n6301 & n6303 ) | ( n6302 & n6303 ) ;
  assign n6306 = n5143 ^ n519 ^ 1'b0 ;
  assign n6307 = n636 & n6306 ;
  assign n6308 = n5185 ^ n1658 ^ 1'b0 ;
  assign n6309 = ( n6200 & ~n6307 ) | ( n6200 & n6308 ) | ( ~n6307 & n6308 ) ;
  assign n6305 = n947 & n4535 ;
  assign n6310 = n6309 ^ n6305 ^ 1'b0 ;
  assign n6316 = ( ~n468 & n2098 ) | ( ~n468 & n6133 ) | ( n2098 & n6133 ) ;
  assign n6312 = x231 ^ x183 ^ 1'b0 ;
  assign n6313 = ( x47 & n2879 ) | ( x47 & n6312 ) | ( n2879 & n6312 ) ;
  assign n6314 = n602 & ~n2229 ;
  assign n6315 = ~n6313 & n6314 ;
  assign n6311 = n5984 ^ n3720 ^ n3505 ;
  assign n6317 = n6316 ^ n6315 ^ n6311 ;
  assign n6318 = n1803 ^ n872 ^ n870 ;
  assign n6319 = n2699 ^ n645 ^ n283 ;
  assign n6320 = ( ~n992 & n1949 ) | ( ~n992 & n4915 ) | ( n1949 & n4915 ) ;
  assign n6321 = n6320 ^ n3716 ^ n2376 ;
  assign n6322 = ( n6318 & ~n6319 ) | ( n6318 & n6321 ) | ( ~n6319 & n6321 ) ;
  assign n6323 = n4444 ^ n687 ^ 1'b0 ;
  assign n6324 = ( n2870 & n3840 ) | ( n2870 & n6323 ) | ( n3840 & n6323 ) ;
  assign n6325 = ~x4 & n6324 ;
  assign n6326 = n3171 ^ n3070 ^ n2975 ;
  assign n6327 = n1034 ^ n1022 ^ n522 ;
  assign n6328 = n2171 ^ n487 ^ n468 ;
  assign n6329 = ~n3819 & n6328 ;
  assign n6330 = n6327 & n6329 ;
  assign n6331 = n6326 | n6330 ;
  assign n6332 = n6325 & ~n6331 ;
  assign n6333 = n6332 ^ n1573 ^ n1145 ;
  assign n6334 = ( n1267 & n1533 ) | ( n1267 & n2658 ) | ( n1533 & n2658 ) ;
  assign n6335 = ( ~n317 & n914 ) | ( ~n317 & n1013 ) | ( n914 & n1013 ) ;
  assign n6336 = ~n2290 & n6335 ;
  assign n6337 = n6336 ^ n5438 ^ n4431 ;
  assign n6338 = ( n2445 & n6334 ) | ( n2445 & ~n6337 ) | ( n6334 & ~n6337 ) ;
  assign n6340 = n5587 ^ n5075 ^ n3185 ;
  assign n6339 = n3840 ^ n2011 ^ 1'b0 ;
  assign n6341 = n6340 ^ n6339 ^ n5460 ;
  assign n6342 = n6338 & n6341 ;
  assign n6347 = n2350 ^ n2153 ^ n1566 ;
  assign n6345 = ( n802 & n847 ) | ( n802 & n1318 ) | ( n847 & n1318 ) ;
  assign n6343 = n4708 ^ n1941 ^ 1'b0 ;
  assign n6344 = ~n2087 & n6343 ;
  assign n6346 = n6345 ^ n6344 ^ n4281 ;
  assign n6348 = n6347 ^ n6346 ^ 1'b0 ;
  assign n6349 = ~n4557 & n6348 ;
  assign n6350 = ( n2251 & n2972 ) | ( n2251 & ~n5624 ) | ( n2972 & ~n5624 ) ;
  assign n6351 = n6350 ^ n4282 ^ n1484 ;
  assign n6352 = ( n2212 & n2403 ) | ( n2212 & n3131 ) | ( n2403 & n3131 ) ;
  assign n6353 = n4816 ^ n4071 ^ n1195 ;
  assign n6354 = ( ~n3395 & n6352 ) | ( ~n3395 & n6353 ) | ( n6352 & n6353 ) ;
  assign n6355 = n430 & ~n6354 ;
  assign n6359 = n5455 ^ n763 ^ 1'b0 ;
  assign n6360 = n2324 ^ n2169 ^ n1199 ;
  assign n6361 = n6360 ^ n3058 ^ 1'b0 ;
  assign n6362 = n6361 ^ n5705 ^ n337 ;
  assign n6363 = n6362 ^ n5235 ^ n2777 ;
  assign n6364 = n6359 | n6363 ;
  assign n6365 = n713 & ~n6364 ;
  assign n6366 = ( n627 & n5899 ) | ( n627 & ~n6365 ) | ( n5899 & ~n6365 ) ;
  assign n6356 = n2850 ^ n671 ^ 1'b0 ;
  assign n6357 = n6356 ^ n1601 ^ n1401 ;
  assign n6358 = ~n2395 & n6357 ;
  assign n6367 = n6366 ^ n6358 ^ 1'b0 ;
  assign n6368 = n6367 ^ n4373 ^ n3581 ;
  assign n6369 = n1067 ^ n565 ^ n337 ;
  assign n6370 = n6369 ^ n3100 ^ n2365 ;
  assign n6371 = n6040 ^ n5690 ^ n4180 ;
  assign n6372 = n6371 ^ n5630 ^ n2513 ;
  assign n6375 = n848 ^ n772 ^ x173 ;
  assign n6373 = ( ~n648 & n1472 ) | ( ~n648 & n2967 ) | ( n1472 & n2967 ) ;
  assign n6374 = ( ~n3307 & n3823 ) | ( ~n3307 & n6373 ) | ( n3823 & n6373 ) ;
  assign n6376 = n6375 ^ n6374 ^ 1'b0 ;
  assign n6380 = ~n921 & n1553 ;
  assign n6381 = ~n4236 & n6380 ;
  assign n6377 = n2790 ^ n927 ^ x41 ;
  assign n6378 = n6377 ^ n1579 ^ n1282 ;
  assign n6379 = n6378 ^ n5856 ^ n3944 ;
  assign n6382 = n6381 ^ n6379 ^ n2291 ;
  assign n6383 = n1423 ^ n1265 ^ n552 ;
  assign n6384 = n1607 & n3343 ;
  assign n6385 = n6384 ^ n2866 ^ n1729 ;
  assign n6386 = ( n619 & ~n6264 ) | ( n619 & n6385 ) | ( ~n6264 & n6385 ) ;
  assign n6387 = ( ~n1355 & n6383 ) | ( ~n1355 & n6386 ) | ( n6383 & n6386 ) ;
  assign n6388 = n6387 ^ n1201 ^ n611 ;
  assign n6389 = n3805 ^ n3075 ^ 1'b0 ;
  assign n6390 = ( ~n1664 & n1705 ) | ( ~n1664 & n6389 ) | ( n1705 & n6389 ) ;
  assign n6401 = n2044 ^ n1236 ^ n1169 ;
  assign n6399 = n4426 ^ n1874 ^ n1015 ;
  assign n6400 = n6399 ^ n3195 ^ x70 ;
  assign n6395 = n3252 ^ n1601 ^ n792 ;
  assign n6396 = n4064 ^ n3367 ^ n1290 ;
  assign n6397 = n6396 ^ n5247 ^ n4828 ;
  assign n6398 = n6395 & ~n6397 ;
  assign n6402 = n6401 ^ n6400 ^ n6398 ;
  assign n6391 = n663 & n5578 ;
  assign n6392 = n6391 ^ n4217 ^ n1172 ;
  assign n6393 = ~n6116 & n6392 ;
  assign n6394 = ~n619 & n6393 ;
  assign n6403 = n6402 ^ n6394 ^ n5856 ;
  assign n6408 = n1585 | n5727 ;
  assign n6409 = n6408 ^ n4224 ^ n2054 ;
  assign n6406 = n5177 ^ n3508 ^ n391 ;
  assign n6404 = n2680 | n5335 ;
  assign n6405 = n4396 | n6404 ;
  assign n6407 = n6406 ^ n6405 ^ n1517 ;
  assign n6410 = n6409 ^ n6407 ^ n1702 ;
  assign n6411 = n6410 ^ n4833 ^ 1'b0 ;
  assign n6412 = n1489 & ~n2068 ;
  assign n6413 = n3217 & n6412 ;
  assign n6414 = ( n3338 & ~n5245 ) | ( n3338 & n5530 ) | ( ~n5245 & n5530 ) ;
  assign n6415 = ( x207 & n323 ) | ( x207 & n349 ) | ( n323 & n349 ) ;
  assign n6416 = ( n1924 & n2689 ) | ( n1924 & n3139 ) | ( n2689 & n3139 ) ;
  assign n6417 = ( n3348 & ~n6415 ) | ( n3348 & n6416 ) | ( ~n6415 & n6416 ) ;
  assign n6418 = ( ~n1089 & n1489 ) | ( ~n1089 & n6417 ) | ( n1489 & n6417 ) ;
  assign n6419 = ( n6413 & n6414 ) | ( n6413 & ~n6418 ) | ( n6414 & ~n6418 ) ;
  assign n6420 = ( n2263 & n3294 ) | ( n2263 & n4275 ) | ( n3294 & n4275 ) ;
  assign n6421 = n6420 ^ n4644 ^ n1570 ;
  assign n6422 = n445 | n2803 ;
  assign n6423 = ( n5096 & n6421 ) | ( n5096 & ~n6422 ) | ( n6421 & ~n6422 ) ;
  assign n6424 = n6423 ^ n4281 ^ n2015 ;
  assign n6428 = n5351 ^ n1127 ^ n485 ;
  assign n6425 = ( ~n789 & n1688 ) | ( ~n789 & n1926 ) | ( n1688 & n1926 ) ;
  assign n6426 = ( n2280 & n3220 ) | ( n2280 & ~n6425 ) | ( n3220 & ~n6425 ) ;
  assign n6427 = n6426 ^ n1958 ^ 1'b0 ;
  assign n6429 = n6428 ^ n6427 ^ 1'b0 ;
  assign n6430 = x214 & n6429 ;
  assign n6431 = ( n4944 & ~n6424 ) | ( n4944 & n6430 ) | ( ~n6424 & n6430 ) ;
  assign n6432 = ( x131 & ~n1060 ) | ( x131 & n2147 ) | ( ~n1060 & n2147 ) ;
  assign n6433 = n1074 ^ n1063 ^ n668 ;
  assign n6434 = n6432 | n6433 ;
  assign n6435 = n1145 | n6434 ;
  assign n6436 = n1603 & n6435 ;
  assign n6437 = ( x5 & n4816 ) | ( x5 & n6436 ) | ( n4816 & n6436 ) ;
  assign n6438 = n1099 & ~n2226 ;
  assign n6439 = ~n941 & n6438 ;
  assign n6440 = n878 | n2070 ;
  assign n6441 = ( n1443 & ~n6439 ) | ( n1443 & n6440 ) | ( ~n6439 & n6440 ) ;
  assign n6442 = n3184 ^ n1172 ^ 1'b0 ;
  assign n6443 = ( x158 & n3843 ) | ( x158 & ~n4582 ) | ( n3843 & ~n4582 ) ;
  assign n6444 = n6443 ^ n2739 ^ n2502 ;
  assign n6445 = n4656 ^ n331 ^ 1'b0 ;
  assign n6446 = n5216 | n6445 ;
  assign n6447 = n2698 & ~n5690 ;
  assign n6448 = ( n1949 & n6446 ) | ( n1949 & n6447 ) | ( n6446 & n6447 ) ;
  assign n6449 = ~n365 & n521 ;
  assign n6450 = n3479 & n6449 ;
  assign n6454 = n2978 ^ n2515 ^ x175 ;
  assign n6453 = ( n1591 & n3569 ) | ( n1591 & ~n5642 ) | ( n3569 & ~n5642 ) ;
  assign n6451 = n2737 ^ n2485 ^ n1573 ;
  assign n6452 = ( n1793 & n4112 ) | ( n1793 & n6451 ) | ( n4112 & n6451 ) ;
  assign n6455 = n6454 ^ n6453 ^ n6452 ;
  assign n6456 = ( ~n1928 & n6450 ) | ( ~n1928 & n6455 ) | ( n6450 & n6455 ) ;
  assign n6457 = ( n1680 & ~n4250 ) | ( n1680 & n5511 ) | ( ~n4250 & n5511 ) ;
  assign n6458 = ( x170 & n838 ) | ( x170 & ~n6457 ) | ( n838 & ~n6457 ) ;
  assign n6459 = n6458 ^ n2534 ^ n2306 ;
  assign n6460 = x108 & n4191 ;
  assign n6461 = n6460 ^ n1200 ^ 1'b0 ;
  assign n6462 = n6461 ^ n3750 ^ n1188 ;
  assign n6463 = ( n2051 & ~n2151 ) | ( n2051 & n5661 ) | ( ~n2151 & n5661 ) ;
  assign n6464 = ( n3252 & ~n6462 ) | ( n3252 & n6463 ) | ( ~n6462 & n6463 ) ;
  assign n6465 = n4013 ^ n3139 ^ n3119 ;
  assign n6466 = n6465 ^ n3547 ^ n1452 ;
  assign n6467 = ( n786 & n1405 ) | ( n786 & n5699 ) | ( n1405 & n5699 ) ;
  assign n6468 = n6467 ^ n2658 ^ n1829 ;
  assign n6469 = ( n751 & n4073 ) | ( n751 & ~n6468 ) | ( n4073 & ~n6468 ) ;
  assign n6470 = ( x94 & n356 ) | ( x94 & ~n6469 ) | ( n356 & ~n6469 ) ;
  assign n6471 = ( n3998 & n5426 ) | ( n3998 & n5435 ) | ( n5426 & n5435 ) ;
  assign n6477 = n3140 ^ n490 ^ 1'b0 ;
  assign n6472 = n4902 ^ n1822 ^ n1044 ;
  assign n6473 = ~n842 & n2822 ;
  assign n6474 = n3462 & n6473 ;
  assign n6475 = n6472 & n6474 ;
  assign n6476 = ( n321 & ~n810 ) | ( n321 & n6475 ) | ( ~n810 & n6475 ) ;
  assign n6478 = n6477 ^ n6476 ^ n4978 ;
  assign n6500 = n3960 ^ n3259 ^ 1'b0 ;
  assign n6501 = n1588 & n6500 ;
  assign n6502 = n6501 ^ n5252 ^ n2334 ;
  assign n6485 = n4842 ^ n4439 ^ n4376 ;
  assign n6486 = ( ~n826 & n1821 ) | ( ~n826 & n6485 ) | ( n1821 & n6485 ) ;
  assign n6487 = n3117 ^ n1852 ^ n1818 ;
  assign n6488 = n6487 ^ n2914 ^ n1123 ;
  assign n6489 = ( n3004 & n6486 ) | ( n3004 & n6488 ) | ( n6486 & n6488 ) ;
  assign n6494 = ( ~x46 & n561 ) | ( ~x46 & n1967 ) | ( n561 & n1967 ) ;
  assign n6495 = n6494 ^ n828 ^ 1'b0 ;
  assign n6496 = n2333 | n6495 ;
  assign n6497 = n6496 ^ n5247 ^ n3564 ;
  assign n6491 = n1536 ^ n700 ^ n629 ;
  assign n6492 = ( x151 & n556 ) | ( x151 & ~n6491 ) | ( n556 & ~n6491 ) ;
  assign n6490 = n3810 ^ n1153 ^ n816 ;
  assign n6493 = n6492 ^ n6490 ^ n2235 ;
  assign n6498 = n6497 ^ n6493 ^ n1233 ;
  assign n6499 = ( n2015 & ~n6489 ) | ( n2015 & n6498 ) | ( ~n6489 & n6498 ) ;
  assign n6482 = ( n560 & ~n1489 ) | ( n560 & n2088 ) | ( ~n1489 & n2088 ) ;
  assign n6479 = ( n2023 & n3734 ) | ( n2023 & ~n3783 ) | ( n3734 & ~n3783 ) ;
  assign n6480 = n2875 ^ n1789 ^ n1309 ;
  assign n6481 = ( ~n3016 & n6479 ) | ( ~n3016 & n6480 ) | ( n6479 & n6480 ) ;
  assign n6483 = n6482 ^ n6481 ^ n539 ;
  assign n6484 = n6483 ^ n3749 ^ n2475 ;
  assign n6503 = n6502 ^ n6499 ^ n6484 ;
  assign n6504 = ( n1344 & ~n6299 ) | ( n1344 & n6503 ) | ( ~n6299 & n6503 ) ;
  assign n6505 = ( n3934 & n6478 ) | ( n3934 & ~n6504 ) | ( n6478 & ~n6504 ) ;
  assign n6506 = n3278 ^ n3103 ^ n2131 ;
  assign n6507 = ( ~n3348 & n4810 ) | ( ~n3348 & n6506 ) | ( n4810 & n6506 ) ;
  assign n6509 = n2080 ^ x4 ^ 1'b0 ;
  assign n6508 = n5393 ^ n4875 ^ n947 ;
  assign n6510 = n6509 ^ n6508 ^ n2035 ;
  assign n6511 = n4586 & ~n6510 ;
  assign n6520 = ( n465 & ~n2324 ) | ( n465 & n3974 ) | ( ~n2324 & n3974 ) ;
  assign n6521 = n6520 ^ n6133 ^ n286 ;
  assign n6516 = ( ~x192 & n1342 ) | ( ~x192 & n4522 ) | ( n1342 & n4522 ) ;
  assign n6517 = ( n1436 & n2788 ) | ( n1436 & ~n6516 ) | ( n2788 & ~n6516 ) ;
  assign n6518 = n1081 & ~n4925 ;
  assign n6519 = ~n6517 & n6518 ;
  assign n6512 = ( n1986 & n2330 ) | ( n1986 & ~n4625 ) | ( n2330 & ~n4625 ) ;
  assign n6513 = n6512 ^ n4639 ^ n4464 ;
  assign n6514 = ( ~n675 & n2098 ) | ( ~n675 & n6513 ) | ( n2098 & n6513 ) ;
  assign n6515 = n643 & n6514 ;
  assign n6522 = n6521 ^ n6519 ^ n6515 ;
  assign n6526 = n4259 ^ n1533 ^ n1044 ;
  assign n6523 = ( n2521 & ~n4000 ) | ( n2521 & n4418 ) | ( ~n4000 & n4418 ) ;
  assign n6524 = n6523 ^ n3479 ^ n851 ;
  assign n6525 = n460 & n6524 ;
  assign n6527 = n6526 ^ n6525 ^ n4137 ;
  assign n6532 = n1718 ^ n1567 ^ n1186 ;
  assign n6533 = n983 | n2761 ;
  assign n6534 = n6532 & ~n6533 ;
  assign n6531 = n6198 ^ n3262 ^ n340 ;
  assign n6535 = n6534 ^ n6531 ^ n6413 ;
  assign n6528 = n4594 ^ n2643 ^ n1528 ;
  assign n6529 = n6528 ^ n6477 ^ n1081 ;
  assign n6530 = n6529 ^ n5457 ^ n5156 ;
  assign n6536 = n6535 ^ n6530 ^ n1494 ;
  assign n6537 = n4197 ^ n2637 ^ n1521 ;
  assign n6538 = n3716 ^ n2936 ^ n1977 ;
  assign n6539 = ( n1048 & n6537 ) | ( n1048 & n6538 ) | ( n6537 & n6538 ) ;
  assign n6540 = ( ~n1104 & n1298 ) | ( ~n1104 & n3220 ) | ( n1298 & n3220 ) ;
  assign n6541 = n3522 | n6540 ;
  assign n6553 = ( n1537 & ~n2420 ) | ( n1537 & n4582 ) | ( ~n2420 & n4582 ) ;
  assign n6556 = n3064 & n5662 ;
  assign n6557 = n6556 ^ n4077 ^ 1'b0 ;
  assign n6554 = n2425 ^ n2312 ^ n1016 ;
  assign n6555 = n6554 ^ n2253 ^ n1252 ;
  assign n6558 = n6557 ^ n6555 ^ n791 ;
  assign n6559 = ( n5306 & n6553 ) | ( n5306 & ~n6558 ) | ( n6553 & ~n6558 ) ;
  assign n6550 = n2510 ^ n1259 ^ n1224 ;
  assign n6551 = n6550 ^ n4862 ^ n4812 ;
  assign n6552 = n6551 ^ n3203 ^ n280 ;
  assign n6547 = n6260 ^ n3522 ^ 1'b0 ;
  assign n6548 = ~n2842 & n6547 ;
  assign n6542 = n1800 | n2195 ;
  assign n6543 = n6542 ^ n933 ^ 1'b0 ;
  assign n6544 = ( n2268 & n2952 ) | ( n2268 & n6543 ) | ( n2952 & n6543 ) ;
  assign n6545 = ( n4010 & n4308 ) | ( n4010 & n6544 ) | ( n4308 & n6544 ) ;
  assign n6546 = ( n3350 & ~n6147 ) | ( n3350 & n6545 ) | ( ~n6147 & n6545 ) ;
  assign n6549 = n6548 ^ n6546 ^ n2948 ;
  assign n6560 = n6559 ^ n6552 ^ n6549 ;
  assign n6561 = ( n3356 & n6541 ) | ( n3356 & ~n6560 ) | ( n6541 & ~n6560 ) ;
  assign n6562 = n6561 ^ n1661 ^ 1'b0 ;
  assign n6563 = ~n6539 & n6562 ;
  assign n6564 = n2056 ^ n1764 ^ n1673 ;
  assign n6565 = n1781 ^ x241 ^ x2 ;
  assign n6566 = n6565 ^ n6545 ^ 1'b0 ;
  assign n6567 = n6228 & n6566 ;
  assign n6568 = n6406 & n6567 ;
  assign n6569 = n6568 ^ n4366 ^ 1'b0 ;
  assign n6573 = n4126 ^ n2639 ^ x129 ;
  assign n6574 = n349 & ~n6573 ;
  assign n6570 = ( ~n515 & n1613 ) | ( ~n515 & n4816 ) | ( n1613 & n4816 ) ;
  assign n6571 = n6570 ^ n5681 ^ 1'b0 ;
  assign n6572 = n1217 & n6571 ;
  assign n6575 = n6574 ^ n6572 ^ 1'b0 ;
  assign n6576 = n4728 ^ n2098 ^ n953 ;
  assign n6577 = x90 & n6576 ;
  assign n6578 = ( n3655 & ~n4118 ) | ( n3655 & n6577 ) | ( ~n4118 & n6577 ) ;
  assign n6579 = n5309 ^ n4830 ^ n4405 ;
  assign n6585 = ( n1607 & n1992 ) | ( n1607 & ~n2704 ) | ( n1992 & ~n2704 ) ;
  assign n6580 = n4820 ^ n3436 ^ 1'b0 ;
  assign n6581 = ( ~n1195 & n1718 ) | ( ~n1195 & n1998 ) | ( n1718 & n1998 ) ;
  assign n6582 = ~n5265 & n6581 ;
  assign n6583 = ~n3085 & n6582 ;
  assign n6584 = ( n3129 & n6580 ) | ( n3129 & n6583 ) | ( n6580 & n6583 ) ;
  assign n6586 = n6585 ^ n6584 ^ n2526 ;
  assign n6587 = n2239 | n5528 ;
  assign n6588 = ( n6579 & n6586 ) | ( n6579 & ~n6587 ) | ( n6586 & ~n6587 ) ;
  assign n6589 = ( x67 & n2892 ) | ( x67 & ~n4150 ) | ( n2892 & ~n4150 ) ;
  assign n6590 = n1137 ^ n945 ^ 1'b0 ;
  assign n6591 = n6589 & ~n6590 ;
  assign n6592 = ( n3431 & n4556 ) | ( n3431 & n6591 ) | ( n4556 & n6591 ) ;
  assign n6593 = n6592 ^ n935 ^ 1'b0 ;
  assign n6608 = n1348 ^ n1268 ^ n1025 ;
  assign n6609 = n4598 ^ n2105 ^ n1678 ;
  assign n6610 = ( n1061 & ~n6608 ) | ( n1061 & n6609 ) | ( ~n6608 & n6609 ) ;
  assign n6606 = ( n617 & n743 ) | ( n617 & n2775 ) | ( n743 & n2775 ) ;
  assign n6605 = ( x154 & n3353 ) | ( x154 & ~n4575 ) | ( n3353 & ~n4575 ) ;
  assign n6594 = n4460 ^ n1459 ^ n1269 ;
  assign n6595 = n1360 & ~n6594 ;
  assign n6596 = ( x38 & n705 ) | ( x38 & n1618 ) | ( n705 & n1618 ) ;
  assign n6598 = n3537 ^ n1760 ^ n1677 ;
  assign n6597 = n1204 | n1827 ;
  assign n6599 = n6598 ^ n6597 ^ 1'b0 ;
  assign n6600 = n6599 ^ n3220 ^ n2634 ;
  assign n6601 = n6596 & n6600 ;
  assign n6602 = ( x51 & n6595 ) | ( x51 & n6601 ) | ( n6595 & n6601 ) ;
  assign n6603 = x29 & ~n6602 ;
  assign n6604 = n6603 ^ n4119 ^ 1'b0 ;
  assign n6607 = n6606 ^ n6605 ^ n6604 ;
  assign n6611 = n6610 ^ n6607 ^ n2287 ;
  assign n6612 = n684 | n5929 ;
  assign n6613 = n6612 ^ n720 ^ 1'b0 ;
  assign n6614 = n6613 ^ n3489 ^ 1'b0 ;
  assign n6617 = n5020 ^ n3728 ^ n1697 ;
  assign n6618 = n6617 ^ n4002 ^ n1198 ;
  assign n6615 = n2791 & ~n4233 ;
  assign n6616 = n6615 ^ n2955 ^ n2539 ;
  assign n6619 = n6618 ^ n6616 ^ 1'b0 ;
  assign n6620 = n6614 & ~n6619 ;
  assign n6624 = n289 & n2201 ;
  assign n6625 = ~n532 & n6624 ;
  assign n6626 = n6625 ^ n2987 ^ n256 ;
  assign n6627 = ( x71 & n1922 ) | ( x71 & ~n6626 ) | ( n1922 & ~n6626 ) ;
  assign n6628 = n6627 ^ n3009 ^ n1024 ;
  assign n6621 = n2967 ^ n2162 ^ 1'b0 ;
  assign n6622 = ( n1426 & n3468 ) | ( n1426 & n6621 ) | ( n3468 & n6621 ) ;
  assign n6623 = ( n3555 & n4192 ) | ( n3555 & n6622 ) | ( n4192 & n6622 ) ;
  assign n6629 = n6628 ^ n6623 ^ n3772 ;
  assign n6631 = ( n1925 & n2935 ) | ( n1925 & n3057 ) | ( n2935 & n3057 ) ;
  assign n6632 = ~n2611 & n6631 ;
  assign n6633 = n6632 ^ n1011 ^ 1'b0 ;
  assign n6634 = n3194 | n6633 ;
  assign n6630 = n6498 ^ n3007 ^ 1'b0 ;
  assign n6635 = n6634 ^ n6630 ^ n3025 ;
  assign n6636 = n6635 ^ n298 ^ 1'b0 ;
  assign n6637 = n6636 ^ n3240 ^ 1'b0 ;
  assign n6647 = n2993 ^ n1088 ^ 1'b0 ;
  assign n6648 = n1894 & n6647 ;
  assign n6645 = ( n1522 & n3276 ) | ( n1522 & ~n4496 ) | ( n3276 & ~n4496 ) ;
  assign n6646 = ( x1 & ~n3076 ) | ( x1 & n6645 ) | ( ~n3076 & n6645 ) ;
  assign n6638 = ( n3022 & n4178 ) | ( n3022 & n5419 ) | ( n4178 & n5419 ) ;
  assign n6639 = ( n1371 & n2103 ) | ( n1371 & ~n6638 ) | ( n2103 & ~n6638 ) ;
  assign n6640 = ( ~n399 & n2394 ) | ( ~n399 & n4070 ) | ( n2394 & n4070 ) ;
  assign n6641 = n6640 ^ n4271 ^ n2649 ;
  assign n6642 = ~n3902 & n6105 ;
  assign n6643 = ~n6641 & n6642 ;
  assign n6644 = ( n350 & ~n6639 ) | ( n350 & n6643 ) | ( ~n6639 & n6643 ) ;
  assign n6649 = n6648 ^ n6646 ^ n6644 ;
  assign n6655 = ( n1363 & ~n2450 ) | ( n1363 & n4463 ) | ( ~n2450 & n4463 ) ;
  assign n6650 = n1905 & n2809 ;
  assign n6651 = n6650 ^ n4540 ^ 1'b0 ;
  assign n6652 = n4128 & ~n6651 ;
  assign n6653 = n6652 ^ n1152 ^ n321 ;
  assign n6654 = n6653 ^ n4189 ^ n1443 ;
  assign n6656 = n6655 ^ n6654 ^ n1124 ;
  assign n6657 = ( n2902 & n4709 ) | ( n2902 & n6656 ) | ( n4709 & n6656 ) ;
  assign n6659 = ( n870 & ~n4459 ) | ( n870 & n5700 ) | ( ~n4459 & n5700 ) ;
  assign n6660 = ( n1881 & ~n5796 ) | ( n1881 & n6659 ) | ( ~n5796 & n6659 ) ;
  assign n6658 = n1961 | n3897 ;
  assign n6661 = n6660 ^ n6658 ^ 1'b0 ;
  assign n6675 = n4031 ^ n1255 ^ n648 ;
  assign n6676 = n6675 ^ n6147 ^ n2049 ;
  assign n6663 = n5691 ^ n5527 ^ n3523 ;
  assign n6664 = n4196 ^ n2605 ^ n2363 ;
  assign n6665 = n5447 ^ n2284 ^ n302 ;
  assign n6666 = n4347 ^ n3211 ^ 1'b0 ;
  assign n6667 = n6665 & ~n6666 ;
  assign n6668 = n705 ^ x129 ^ x36 ;
  assign n6669 = n6668 ^ n6214 ^ n2599 ;
  assign n6670 = n3899 & n6669 ;
  assign n6671 = n6670 ^ n5105 ^ 1'b0 ;
  assign n6672 = ( n6664 & n6667 ) | ( n6664 & ~n6671 ) | ( n6667 & ~n6671 ) ;
  assign n6673 = n6663 | n6672 ;
  assign n6674 = n6673 ^ n454 ^ 1'b0 ;
  assign n6662 = n4436 ^ n4069 ^ 1'b0 ;
  assign n6677 = n6676 ^ n6674 ^ n6662 ;
  assign n6678 = ( ~n868 & n938 ) | ( ~n868 & n4910 ) | ( n938 & n4910 ) ;
  assign n6680 = n852 ^ n578 ^ x192 ;
  assign n6679 = n4128 ^ n2711 ^ n1621 ;
  assign n6681 = n6680 ^ n6679 ^ n3600 ;
  assign n6682 = n6678 | n6681 ;
  assign n6699 = ( n824 & n1511 ) | ( n824 & n3630 ) | ( n1511 & n3630 ) ;
  assign n6683 = ( x149 & ~n826 ) | ( x149 & n3048 ) | ( ~n826 & n3048 ) ;
  assign n6684 = ~n312 & n6683 ;
  assign n6685 = ( ~x123 & n1382 ) | ( ~x123 & n1659 ) | ( n1382 & n1659 ) ;
  assign n6686 = n6685 ^ n1352 ^ x225 ;
  assign n6690 = ( n711 & n808 ) | ( n711 & n3393 ) | ( n808 & n3393 ) ;
  assign n6691 = n871 ^ x142 ^ 1'b0 ;
  assign n6692 = n6690 & ~n6691 ;
  assign n6693 = n6692 ^ n2844 ^ 1'b0 ;
  assign n6688 = n3180 ^ n2360 ^ n1164 ;
  assign n6689 = n2962 & n6688 ;
  assign n6694 = n6693 ^ n6689 ^ n2023 ;
  assign n6695 = ( ~n1041 & n5163 ) | ( ~n1041 & n6694 ) | ( n5163 & n6694 ) ;
  assign n6687 = ~n1766 & n4301 ;
  assign n6696 = n6695 ^ n6687 ^ 1'b0 ;
  assign n6697 = ( ~n820 & n6686 ) | ( ~n820 & n6696 ) | ( n6686 & n6696 ) ;
  assign n6698 = ( n991 & ~n6684 ) | ( n991 & n6697 ) | ( ~n6684 & n6697 ) ;
  assign n6700 = n6699 ^ n6698 ^ n5326 ;
  assign n6702 = n1671 ^ n1008 ^ n884 ;
  assign n6701 = n2853 ^ n1084 ^ n933 ;
  assign n6703 = n6702 ^ n6701 ^ n436 ;
  assign n6712 = ~n782 & n4184 ;
  assign n6713 = n6712 ^ n1797 ^ 1'b0 ;
  assign n6714 = n6713 ^ n4345 ^ n1316 ;
  assign n6707 = ( n339 & n1232 ) | ( n339 & ~n4522 ) | ( n1232 & ~n4522 ) ;
  assign n6704 = n1555 ^ n785 ^ n297 ;
  assign n6705 = ( ~n417 & n1898 ) | ( ~n417 & n6704 ) | ( n1898 & n6704 ) ;
  assign n6706 = n6705 ^ n6147 ^ n358 ;
  assign n6708 = n6707 ^ n6706 ^ n1539 ;
  assign n6709 = n6708 ^ n2569 ^ n1922 ;
  assign n6710 = n6709 ^ n3410 ^ n2955 ;
  assign n6711 = ( ~n2441 & n5017 ) | ( ~n2441 & n6710 ) | ( n5017 & n6710 ) ;
  assign n6715 = n6714 ^ n6711 ^ n3720 ;
  assign n6716 = n5731 ^ n4715 ^ x158 ;
  assign n6717 = ( ~n5583 & n5650 ) | ( ~n5583 & n6716 ) | ( n5650 & n6716 ) ;
  assign n6718 = n4056 & n6717 ;
  assign n6719 = n1928 | n6718 ;
  assign n6720 = n6715 | n6719 ;
  assign n6721 = ( x198 & ~x217 ) | ( x198 & n1758 ) | ( ~x217 & n1758 ) ;
  assign n6722 = ( n365 & n3687 ) | ( n365 & ~n4560 ) | ( n3687 & ~n4560 ) ;
  assign n6723 = ( n5784 & n6721 ) | ( n5784 & ~n6722 ) | ( n6721 & ~n6722 ) ;
  assign n6732 = n4364 ^ n3942 ^ n3056 ;
  assign n6733 = ( n1914 & n2832 ) | ( n1914 & n6732 ) | ( n2832 & n6732 ) ;
  assign n6724 = n4399 ^ n3796 ^ n516 ;
  assign n6725 = ( n4507 & ~n6313 ) | ( n4507 & n6724 ) | ( ~n6313 & n6724 ) ;
  assign n6726 = n2332 ^ n1668 ^ n318 ;
  assign n6727 = ( n374 & n1819 ) | ( n374 & ~n6420 ) | ( n1819 & ~n6420 ) ;
  assign n6728 = n4336 ^ n2535 ^ n2100 ;
  assign n6729 = ( n2537 & n6727 ) | ( n2537 & ~n6728 ) | ( n6727 & ~n6728 ) ;
  assign n6730 = n6726 & ~n6729 ;
  assign n6731 = ~n6725 & n6730 ;
  assign n6734 = n6733 ^ n6731 ^ 1'b0 ;
  assign n6736 = ( n484 & ~n1982 ) | ( n484 & n4834 ) | ( ~n1982 & n4834 ) ;
  assign n6737 = n4144 ^ n1329 ^ 1'b0 ;
  assign n6738 = ( ~n4520 & n6736 ) | ( ~n4520 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6735 = n4265 ^ n3706 ^ n1527 ;
  assign n6739 = n6738 ^ n6735 ^ n2770 ;
  assign n6746 = n4913 ^ n2567 ^ n830 ;
  assign n6747 = n6746 ^ n805 ^ x35 ;
  assign n6748 = n6747 ^ n6075 ^ n2609 ;
  assign n6745 = n657 & ~n2377 ;
  assign n6742 = n6177 ^ n3627 ^ n2847 ;
  assign n6743 = ( ~n1706 & n4465 ) | ( ~n1706 & n6742 ) | ( n4465 & n6742 ) ;
  assign n6740 = n5113 ^ n3567 ^ 1'b0 ;
  assign n6741 = n6740 ^ n6344 ^ n1895 ;
  assign n6744 = n6743 ^ n6741 ^ 1'b0 ;
  assign n6749 = n6748 ^ n6745 ^ n6744 ;
  assign n6750 = ~n2585 & n6194 ;
  assign n6751 = ~n3212 & n6750 ;
  assign n6752 = n6553 ^ n2865 ^ x242 ;
  assign n6753 = n6752 ^ n4495 ^ n1229 ;
  assign n6754 = n6753 ^ n2911 ^ n435 ;
  assign n6755 = ( n2068 & ~n6751 ) | ( n2068 & n6754 ) | ( ~n6751 & n6754 ) ;
  assign n6756 = n6112 ^ x17 ^ 1'b0 ;
  assign n6757 = n4401 ^ n1398 ^ n1162 ;
  assign n6758 = n3706 | n4054 ;
  assign n6759 = n6758 ^ n4749 ^ 1'b0 ;
  assign n6761 = ( n292 & n3363 ) | ( n292 & n6638 ) | ( n3363 & n6638 ) ;
  assign n6760 = n3406 ^ n2158 ^ n641 ;
  assign n6762 = n6761 ^ n6760 ^ n2086 ;
  assign n6763 = n3429 ^ n1539 ^ x160 ;
  assign n6764 = n6763 ^ n3772 ^ 1'b0 ;
  assign n6765 = n6762 & n6764 ;
  assign n6773 = ~n473 & n3240 ;
  assign n6774 = ~n451 & n6773 ;
  assign n6775 = ( n1702 & n2831 ) | ( n1702 & n2892 ) | ( n2831 & n2892 ) ;
  assign n6776 = ( n6486 & n6774 ) | ( n6486 & n6775 ) | ( n6774 & n6775 ) ;
  assign n6769 = n3460 ^ n3457 ^ n395 ;
  assign n6770 = n3841 | n6769 ;
  assign n6766 = n3292 ^ n1109 ^ n968 ;
  assign n6767 = ( n762 & ~n2527 ) | ( n762 & n6766 ) | ( ~n2527 & n6766 ) ;
  assign n6768 = n6767 ^ n4057 ^ n601 ;
  assign n6771 = n6770 ^ n6768 ^ 1'b0 ;
  assign n6772 = n4389 | n6771 ;
  assign n6777 = n6776 ^ n6772 ^ n309 ;
  assign n6778 = ( ~n6759 & n6765 ) | ( ~n6759 & n6777 ) | ( n6765 & n6777 ) ;
  assign n6779 = n1036 ^ n489 ^ 1'b0 ;
  assign n6780 = n581 & n6779 ;
  assign n6781 = n1632 | n3115 ;
  assign n6782 = n6780 | n6781 ;
  assign n6783 = ( n721 & ~n6027 ) | ( n721 & n6782 ) | ( ~n6027 & n6782 ) ;
  assign n6784 = n6783 ^ n1292 ^ 1'b0 ;
  assign n6785 = ( n1061 & ~n6778 ) | ( n1061 & n6784 ) | ( ~n6778 & n6784 ) ;
  assign n6786 = n2982 ^ n1060 ^ n839 ;
  assign n6787 = n6786 ^ n6084 ^ n3489 ;
  assign n6788 = ( ~n927 & n1537 ) | ( ~n927 & n3445 ) | ( n1537 & n3445 ) ;
  assign n6790 = n885 ^ n436 ^ n407 ;
  assign n6791 = n6790 ^ n2085 ^ n1324 ;
  assign n6792 = ( ~n1653 & n6017 ) | ( ~n1653 & n6791 ) | ( n6017 & n6791 ) ;
  assign n6789 = ( n451 & n3102 ) | ( n451 & n6473 ) | ( n3102 & n6473 ) ;
  assign n6793 = n6792 ^ n6789 ^ n6581 ;
  assign n6794 = n6788 & ~n6793 ;
  assign n6795 = n6787 & n6794 ;
  assign n6796 = n5966 ^ n4037 ^ 1'b0 ;
  assign n6798 = n1777 ^ n1540 ^ x233 ;
  assign n6799 = n6798 ^ n2611 ^ n1758 ;
  assign n6797 = x100 & ~n5294 ;
  assign n6800 = n6799 ^ n6797 ^ 1'b0 ;
  assign n6804 = ( n365 & ~n563 ) | ( n365 & n1281 ) | ( ~n563 & n1281 ) ;
  assign n6805 = n6804 ^ n5533 ^ n4070 ;
  assign n6801 = ( n1060 & n2602 ) | ( n1060 & ~n3874 ) | ( n2602 & ~n3874 ) ;
  assign n6802 = n6801 ^ n3407 ^ n1394 ;
  assign n6803 = ( n2003 & n5808 ) | ( n2003 & ~n6802 ) | ( n5808 & ~n6802 ) ;
  assign n6806 = n6805 ^ n6803 ^ n2797 ;
  assign n6807 = ( n5089 & n5918 ) | ( n5089 & n6806 ) | ( n5918 & n6806 ) ;
  assign n6808 = n2838 ^ n1050 ^ n1039 ;
  assign n6809 = ( n6425 & n6807 ) | ( n6425 & ~n6808 ) | ( n6807 & ~n6808 ) ;
  assign n6810 = ( n1534 & n3072 ) | ( n1534 & ~n4602 ) | ( n3072 & ~n4602 ) ;
  assign n6811 = ( ~n1695 & n2875 ) | ( ~n1695 & n3130 ) | ( n2875 & n3130 ) ;
  assign n6812 = n5296 & n6811 ;
  assign n6813 = n4007 ^ n2269 ^ 1'b0 ;
  assign n6814 = ~n1036 & n6813 ;
  assign n6815 = ( ~x210 & n445 ) | ( ~x210 & n3743 ) | ( n445 & n3743 ) ;
  assign n6816 = ( n569 & n967 ) | ( n569 & ~n6369 ) | ( n967 & ~n6369 ) ;
  assign n6817 = n3115 | n6816 ;
  assign n6818 = n6817 ^ n3735 ^ 1'b0 ;
  assign n6819 = ( ~n2070 & n2138 ) | ( ~n2070 & n6818 ) | ( n2138 & n6818 ) ;
  assign n6820 = ~n642 & n6819 ;
  assign n6821 = n3997 & n6820 ;
  assign n6822 = ( n367 & ~n6815 ) | ( n367 & n6821 ) | ( ~n6815 & n6821 ) ;
  assign n6823 = ( n6639 & n6814 ) | ( n6639 & n6822 ) | ( n6814 & n6822 ) ;
  assign n6841 = n6401 ^ n2260 ^ n1836 ;
  assign n6840 = ( ~n331 & n1117 ) | ( ~n331 & n4427 ) | ( n1117 & n4427 ) ;
  assign n6838 = n1662 ^ n1431 ^ n456 ;
  assign n6839 = n6838 ^ n5232 ^ n2214 ;
  assign n6842 = n6841 ^ n6840 ^ n6839 ;
  assign n6843 = n6842 ^ n3741 ^ n1559 ;
  assign n6834 = n2975 ^ n1777 ^ n654 ;
  assign n6835 = n6834 ^ n2573 ^ n1650 ;
  assign n6833 = n6028 ^ n1436 ^ 1'b0 ;
  assign n6836 = n6835 ^ n6833 ^ n5382 ;
  assign n6831 = ( n568 & n4564 ) | ( n568 & n5019 ) | ( n4564 & n5019 ) ;
  assign n6832 = ~n1924 & n6831 ;
  assign n6837 = n6836 ^ n6832 ^ n5005 ;
  assign n6824 = ~n1292 & n2682 ;
  assign n6825 = ( n987 & ~n3893 ) | ( n987 & n6824 ) | ( ~n3893 & n6824 ) ;
  assign n6826 = n2701 ^ n1596 ^ n1059 ;
  assign n6827 = ( n814 & ~n1195 ) | ( n814 & n5689 ) | ( ~n1195 & n5689 ) ;
  assign n6828 = ( n762 & n1013 ) | ( n762 & n6827 ) | ( n1013 & n6827 ) ;
  assign n6829 = ( n3990 & n6826 ) | ( n3990 & ~n6828 ) | ( n6826 & ~n6828 ) ;
  assign n6830 = ( n2380 & n6825 ) | ( n2380 & ~n6829 ) | ( n6825 & ~n6829 ) ;
  assign n6844 = n6843 ^ n6837 ^ n6830 ;
  assign n6848 = n2751 ^ n2209 ^ n971 ;
  assign n6847 = n4698 ^ n3859 ^ n1344 ;
  assign n6845 = n1362 ^ n1344 ^ n1239 ;
  assign n6846 = ( ~n940 & n2639 ) | ( ~n940 & n6845 ) | ( n2639 & n6845 ) ;
  assign n6849 = n6848 ^ n6847 ^ n6846 ;
  assign n6850 = n6849 ^ n6068 ^ x223 ;
  assign n6852 = ( n1762 & ~n3809 ) | ( n1762 & n4232 ) | ( ~n3809 & n4232 ) ;
  assign n6851 = n3296 ^ n1704 ^ n401 ;
  assign n6853 = n6852 ^ n6851 ^ 1'b0 ;
  assign n6854 = ( x190 & n5107 ) | ( x190 & ~n6853 ) | ( n5107 & ~n6853 ) ;
  assign n6855 = ( n3894 & ~n6699 ) | ( n3894 & n6854 ) | ( ~n6699 & n6854 ) ;
  assign n6856 = ~n546 & n4792 ;
  assign n6857 = n6856 ^ n2599 ^ 1'b0 ;
  assign n6858 = ( n1357 & n2977 ) | ( n1357 & ~n3541 ) | ( n2977 & ~n3541 ) ;
  assign n6859 = ( n2557 & n2732 ) | ( n2557 & n6858 ) | ( n2732 & n6858 ) ;
  assign n6860 = ( n3711 & ~n6857 ) | ( n3711 & n6859 ) | ( ~n6857 & n6859 ) ;
  assign n6869 = n3585 & ~n5558 ;
  assign n6870 = n6141 & n6869 ;
  assign n6864 = ( n1592 & n2949 ) | ( n1592 & ~n6432 ) | ( n2949 & ~n6432 ) ;
  assign n6865 = ( n900 & ~n1794 ) | ( n900 & n1931 ) | ( ~n1794 & n1931 ) ;
  assign n6866 = ( n1413 & n1927 ) | ( n1413 & ~n6865 ) | ( n1927 & ~n6865 ) ;
  assign n6867 = n6866 ^ n277 ^ x132 ;
  assign n6868 = ~n6864 & n6867 ;
  assign n6861 = n3493 ^ x41 ^ 1'b0 ;
  assign n6862 = ~n5010 & n6861 ;
  assign n6863 = n6862 ^ n3256 ^ 1'b0 ;
  assign n6871 = n6870 ^ n6868 ^ n6863 ;
  assign n6872 = n6871 ^ n4654 ^ n3926 ;
  assign n6873 = ( n535 & ~n1864 ) | ( n535 & n3296 ) | ( ~n1864 & n3296 ) ;
  assign n6874 = ( n542 & n2509 ) | ( n542 & ~n5544 ) | ( n2509 & ~n5544 ) ;
  assign n6875 = n3600 ^ n1490 ^ n1117 ;
  assign n6876 = ( n4275 & n6269 ) | ( n4275 & ~n6875 ) | ( n6269 & ~n6875 ) ;
  assign n6877 = ( n3771 & n6874 ) | ( n3771 & n6876 ) | ( n6874 & n6876 ) ;
  assign n6878 = ( n577 & n6873 ) | ( n577 & ~n6877 ) | ( n6873 & ~n6877 ) ;
  assign n6879 = ( n6148 & ~n6715 ) | ( n6148 & n6878 ) | ( ~n6715 & n6878 ) ;
  assign n6880 = n825 ^ x66 ^ 1'b0 ;
  assign n6881 = ( n1348 & n2819 ) | ( n1348 & ~n6880 ) | ( n2819 & ~n6880 ) ;
  assign n6882 = ( n1200 & n4345 ) | ( n1200 & ~n6881 ) | ( n4345 & ~n6881 ) ;
  assign n6884 = n6585 ^ n4801 ^ 1'b0 ;
  assign n6883 = ( n3066 & n3114 ) | ( n3066 & n4890 ) | ( n3114 & n4890 ) ;
  assign n6885 = n6884 ^ n6883 ^ n6598 ;
  assign n6886 = n5351 | n6885 ;
  assign n6887 = n6886 ^ n2226 ^ n959 ;
  assign n6888 = ( n1074 & n4485 ) | ( n1074 & n6882 ) | ( n4485 & n6882 ) ;
  assign n6892 = ( n1816 & ~n2156 ) | ( n1816 & n2307 ) | ( ~n2156 & n2307 ) ;
  assign n6889 = n6301 ^ n3506 ^ n2097 ;
  assign n6890 = n3945 ^ n2236 ^ 1'b0 ;
  assign n6891 = ( n6320 & ~n6889 ) | ( n6320 & n6890 ) | ( ~n6889 & n6890 ) ;
  assign n6893 = n6892 ^ n6891 ^ n2444 ;
  assign n6894 = ( ~x4 & n3052 ) | ( ~x4 & n3950 ) | ( n3052 & n3950 ) ;
  assign n6895 = n6053 & n6894 ;
  assign n6896 = ( n4872 & ~n6496 ) | ( n4872 & n6895 ) | ( ~n6496 & n6895 ) ;
  assign n6902 = ( n762 & n857 ) | ( n762 & ~n5285 ) | ( n857 & ~n5285 ) ;
  assign n6903 = ( ~n1149 & n3591 ) | ( ~n1149 & n6902 ) | ( n3591 & n6902 ) ;
  assign n6897 = x78 & ~n1893 ;
  assign n6898 = n6897 ^ n1845 ^ x177 ;
  assign n6899 = n6898 ^ n3452 ^ 1'b0 ;
  assign n6900 = n4167 & ~n6899 ;
  assign n6901 = n6900 ^ n5433 ^ n3173 ;
  assign n6904 = n6903 ^ n6901 ^ n3685 ;
  assign n6905 = ( n1265 & n1393 ) | ( n1265 & ~n6206 ) | ( n1393 & ~n6206 ) ;
  assign n6906 = ( n705 & n4219 ) | ( n705 & ~n5009 ) | ( n4219 & ~n5009 ) ;
  assign n6907 = n6906 ^ n3016 ^ n676 ;
  assign n6908 = n4341 ^ n2433 ^ n1437 ;
  assign n6909 = n3443 | n4693 ;
  assign n6910 = n6908 | n6909 ;
  assign n6911 = ( n1454 & n3303 ) | ( n1454 & ~n4514 ) | ( n3303 & ~n4514 ) ;
  assign n6912 = ( n6907 & ~n6910 ) | ( n6907 & n6911 ) | ( ~n6910 & n6911 ) ;
  assign n6913 = ( n3410 & ~n6905 ) | ( n3410 & n6912 ) | ( ~n6905 & n6912 ) ;
  assign n6914 = ( ~n949 & n2879 ) | ( ~n949 & n3558 ) | ( n2879 & n3558 ) ;
  assign n6915 = n4956 ^ n1931 ^ n1279 ;
  assign n6916 = n6915 ^ n514 ^ 1'b0 ;
  assign n6917 = n266 & ~n6916 ;
  assign n6918 = n4123 ^ n3112 ^ n1150 ;
  assign n6919 = n6918 ^ n1829 ^ n711 ;
  assign n6920 = n3131 ^ n1097 ^ 1'b0 ;
  assign n6921 = n680 | n6920 ;
  assign n6922 = n6921 ^ n1153 ^ 1'b0 ;
  assign n6923 = ( n2133 & n3088 ) | ( n2133 & ~n6922 ) | ( n3088 & ~n6922 ) ;
  assign n6924 = ( n6917 & ~n6919 ) | ( n6917 & n6923 ) | ( ~n6919 & n6923 ) ;
  assign n6925 = ( n5818 & n6914 ) | ( n5818 & ~n6924 ) | ( n6914 & ~n6924 ) ;
  assign n6926 = n6925 ^ n6543 ^ 1'b0 ;
  assign n6927 = ( n5138 & n6913 ) | ( n5138 & ~n6926 ) | ( n6913 & ~n6926 ) ;
  assign n6933 = n1410 ^ n686 ^ 1'b0 ;
  assign n6934 = ( n2279 & n3921 ) | ( n2279 & ~n6933 ) | ( n3921 & ~n6933 ) ;
  assign n6935 = n6934 ^ n5796 ^ n4547 ;
  assign n6931 = ( ~n2180 & n4042 ) | ( ~n2180 & n5735 ) | ( n4042 & n5735 ) ;
  assign n6930 = n3406 ^ n1510 ^ n1315 ;
  assign n6928 = ( n715 & n2310 ) | ( n715 & ~n3757 ) | ( n2310 & ~n3757 ) ;
  assign n6929 = ( ~n1618 & n3796 ) | ( ~n1618 & n6928 ) | ( n3796 & n6928 ) ;
  assign n6932 = n6931 ^ n6930 ^ n6929 ;
  assign n6936 = n6935 ^ n6932 ^ 1'b0 ;
  assign n6937 = n762 & n6936 ;
  assign n6938 = n6780 ^ n6020 ^ n1073 ;
  assign n6939 = ( ~n2485 & n3092 ) | ( ~n2485 & n6938 ) | ( n3092 & n6938 ) ;
  assign n6940 = ( n2349 & n5383 ) | ( n2349 & ~n5510 ) | ( n5383 & ~n5510 ) ;
  assign n6941 = n6940 ^ n6801 ^ n2844 ;
  assign n6942 = ( ~n2542 & n6939 ) | ( ~n2542 & n6941 ) | ( n6939 & n6941 ) ;
  assign n6943 = ( ~n3670 & n4518 ) | ( ~n3670 & n6942 ) | ( n4518 & n6942 ) ;
  assign n6944 = n4663 ^ n577 ^ 1'b0 ;
  assign n6945 = n1602 | n6944 ;
  assign n6946 = ~n4990 & n5403 ;
  assign n6947 = n2867 & n6946 ;
  assign n6948 = ( n5387 & n6945 ) | ( n5387 & ~n6947 ) | ( n6945 & ~n6947 ) ;
  assign n6949 = n6884 ^ n2529 ^ n1605 ;
  assign n6950 = ( n1717 & ~n1910 ) | ( n1717 & n1954 ) | ( ~n1910 & n1954 ) ;
  assign n6951 = ( x34 & n1853 ) | ( x34 & ~n6774 ) | ( n1853 & ~n6774 ) ;
  assign n6952 = n6951 ^ n5265 ^ n1299 ;
  assign n6953 = n6952 ^ n1556 ^ 1'b0 ;
  assign n6954 = n6950 & ~n6953 ;
  assign n6957 = n5563 ^ n2568 ^ n1535 ;
  assign n6958 = n2715 ^ n2656 ^ n2246 ;
  assign n6959 = ( n402 & ~n6957 ) | ( n402 & n6958 ) | ( ~n6957 & n6958 ) ;
  assign n6960 = n6959 ^ n6320 ^ n1052 ;
  assign n6955 = ( n427 & ~n4879 ) | ( n427 & n6663 ) | ( ~n4879 & n6663 ) ;
  assign n6956 = n6955 ^ n5828 ^ n4109 ;
  assign n6961 = n6960 ^ n6956 ^ n1049 ;
  assign n6962 = n2679 ^ n842 ^ n756 ;
  assign n6963 = ( n1594 & n5131 ) | ( n1594 & n6066 ) | ( n5131 & n6066 ) ;
  assign n6964 = ( n1118 & n6962 ) | ( n1118 & n6963 ) | ( n6962 & n6963 ) ;
  assign n6965 = n3886 & ~n4076 ;
  assign n6966 = n4469 & n6965 ;
  assign n6967 = n701 ^ n532 ^ n520 ;
  assign n6968 = ~n929 & n6967 ;
  assign n6969 = n6966 & n6968 ;
  assign n6970 = n6969 ^ n4947 ^ n4047 ;
  assign n6976 = ( n1338 & n1734 ) | ( n1338 & ~n3809 ) | ( n1734 & ~n3809 ) ;
  assign n6977 = ( n787 & n6858 ) | ( n787 & n6976 ) | ( n6858 & n6976 ) ;
  assign n6975 = n3549 | n4521 ;
  assign n6971 = n6690 ^ n5131 ^ n4336 ;
  assign n6972 = n6971 ^ n3457 ^ n2915 ;
  assign n6973 = n6625 ^ n2195 ^ 1'b0 ;
  assign n6974 = ( n5282 & n6972 ) | ( n5282 & ~n6973 ) | ( n6972 & ~n6973 ) ;
  assign n6978 = n6977 ^ n6975 ^ n6974 ;
  assign n6979 = n1393 ^ n449 ^ 1'b0 ;
  assign n6980 = n6979 ^ n1262 ^ n686 ;
  assign n6981 = x218 & ~n1224 ;
  assign n6982 = n6981 ^ n1310 ^ n1072 ;
  assign n6983 = ( n727 & n6980 ) | ( n727 & ~n6982 ) | ( n6980 & ~n6982 ) ;
  assign n6985 = ( n2597 & n3232 ) | ( n2597 & ~n6501 ) | ( n3232 & ~n6501 ) ;
  assign n6986 = n6985 ^ n6082 ^ n741 ;
  assign n6984 = n6950 ^ n4182 ^ n949 ;
  assign n6987 = n6986 ^ n6984 ^ x171 ;
  assign n6988 = n3894 ^ n1957 ^ n1574 ;
  assign n6989 = n6988 ^ n4203 ^ n836 ;
  assign n6990 = n6989 ^ n5299 ^ n3484 ;
  assign n6995 = n3533 ^ n850 ^ n484 ;
  assign n6994 = n1924 ^ n1739 ^ n522 ;
  assign n6991 = x240 & ~n1662 ;
  assign n6992 = n2063 ^ n1242 ^ 1'b0 ;
  assign n6993 = ~n6991 & n6992 ;
  assign n6996 = n6995 ^ n6994 ^ n6993 ;
  assign n6997 = n6996 ^ n6684 ^ n2831 ;
  assign n6998 = ~n4403 & n6997 ;
  assign n7003 = n1663 & n2649 ;
  assign n6999 = n3559 ^ n2431 ^ n2218 ;
  assign n7000 = ( n1581 & ~n3711 ) | ( n1581 & n6999 ) | ( ~n3711 & n6999 ) ;
  assign n7001 = ( n2584 & n2870 ) | ( n2584 & n7000 ) | ( n2870 & n7000 ) ;
  assign n7002 = n1368 & ~n7001 ;
  assign n7004 = n7003 ^ n7002 ^ n3415 ;
  assign n7005 = n488 & n7004 ;
  assign n7006 = n5257 ^ n4535 ^ 1'b0 ;
  assign n7011 = ( ~n1414 & n2980 ) | ( ~n1414 & n4690 ) | ( n2980 & n4690 ) ;
  assign n7012 = n7011 ^ n436 ^ x203 ;
  assign n7009 = ( ~n3064 & n5047 ) | ( ~n3064 & n6289 ) | ( n5047 & n6289 ) ;
  assign n7007 = ( x151 & n878 ) | ( x151 & n5027 ) | ( n878 & n5027 ) ;
  assign n7008 = n4961 & ~n7007 ;
  assign n7010 = n7009 ^ n7008 ^ 1'b0 ;
  assign n7013 = n7012 ^ n7010 ^ n1825 ;
  assign n7014 = ( ~n1148 & n4370 ) | ( ~n1148 & n4472 ) | ( n4370 & n4472 ) ;
  assign n7016 = n6261 ^ n2124 ^ x99 ;
  assign n7015 = n3393 ^ n1430 ^ n1192 ;
  assign n7017 = n7016 ^ n7015 ^ 1'b0 ;
  assign n7018 = ~n7014 & n7017 ;
  assign n7028 = ( n823 & n2141 ) | ( n823 & ~n2439 ) | ( n2141 & ~n2439 ) ;
  assign n7029 = ( ~n1506 & n2986 ) | ( ~n1506 & n7028 ) | ( n2986 & n7028 ) ;
  assign n7019 = n2667 & n2866 ;
  assign n7022 = ( ~n2336 & n4245 ) | ( ~n2336 & n5426 ) | ( n4245 & n5426 ) ;
  assign n7023 = n2320 & n7022 ;
  assign n7024 = n4149 & n7023 ;
  assign n7020 = n5474 ^ n5143 ^ n866 ;
  assign n7021 = n7020 ^ n4228 ^ n3680 ;
  assign n7025 = n7024 ^ n7021 ^ n6257 ;
  assign n7026 = n7019 & n7025 ;
  assign n7027 = n5756 & n7026 ;
  assign n7030 = n7029 ^ n7027 ^ 1'b0 ;
  assign n7031 = n4780 ^ n1172 ^ n896 ;
  assign n7032 = n7031 ^ n2370 ^ n2110 ;
  assign n7033 = ( ~x55 & n2749 ) | ( ~x55 & n7032 ) | ( n2749 & n7032 ) ;
  assign n7034 = n7033 ^ n1953 ^ n1345 ;
  assign n7035 = n2292 ^ n490 ^ 1'b0 ;
  assign n7036 = ( n639 & n739 ) | ( n639 & n7035 ) | ( n739 & n7035 ) ;
  assign n7037 = ( n1471 & n4039 ) | ( n1471 & ~n6921 ) | ( n4039 & ~n6921 ) ;
  assign n7038 = ( n1093 & n1907 ) | ( n1093 & ~n7037 ) | ( n1907 & ~n7037 ) ;
  assign n7039 = ( n1737 & n4191 ) | ( n1737 & ~n7038 ) | ( n4191 & ~n7038 ) ;
  assign n7040 = ( n5301 & ~n6878 ) | ( n5301 & n7039 ) | ( ~n6878 & n7039 ) ;
  assign n7041 = n2067 & n7040 ;
  assign n7042 = ~n6058 & n7041 ;
  assign n7043 = n1922 ^ n1641 ^ x30 ;
  assign n7044 = n7043 ^ n3031 ^ x209 ;
  assign n7045 = n6553 ^ n4241 ^ n1476 ;
  assign n7046 = n5790 ^ n4745 ^ n4424 ;
  assign n7047 = n7046 ^ n6627 ^ n753 ;
  assign n7048 = n7047 ^ n4233 ^ n756 ;
  assign n7049 = ( n309 & n2918 ) | ( n309 & ~n7048 ) | ( n2918 & ~n7048 ) ;
  assign n7050 = ( n7044 & n7045 ) | ( n7044 & n7049 ) | ( n7045 & n7049 ) ;
  assign n7051 = n5741 ^ n3565 ^ n2675 ;
  assign n7052 = n7051 ^ n3215 ^ 1'b0 ;
  assign n7053 = ( n1358 & ~n1442 ) | ( n1358 & n7052 ) | ( ~n1442 & n7052 ) ;
  assign n7054 = ( ~n794 & n1757 ) | ( ~n794 & n2150 ) | ( n1757 & n2150 ) ;
  assign n7055 = ( n1109 & n1927 ) | ( n1109 & n7054 ) | ( n1927 & n7054 ) ;
  assign n7056 = n7055 ^ n2945 ^ 1'b0 ;
  assign n7057 = n2275 | n7056 ;
  assign n7058 = n7057 ^ n4031 ^ n1132 ;
  assign n7064 = n2251 ^ x235 ^ x141 ;
  assign n7065 = n4271 ^ n2898 ^ 1'b0 ;
  assign n7066 = n1551 & ~n7065 ;
  assign n7067 = ( n1540 & n7064 ) | ( n1540 & n7066 ) | ( n7064 & n7066 ) ;
  assign n7059 = ( n300 & ~n1418 ) | ( n300 & n3490 ) | ( ~n1418 & n3490 ) ;
  assign n7060 = n2721 ^ n1544 ^ n998 ;
  assign n7061 = n7060 ^ n5703 ^ n2242 ;
  assign n7062 = ( n2607 & ~n2858 ) | ( n2607 & n7061 ) | ( ~n2858 & n7061 ) ;
  assign n7063 = ( x91 & n7059 ) | ( x91 & ~n7062 ) | ( n7059 & ~n7062 ) ;
  assign n7068 = n7067 ^ n7063 ^ 1'b0 ;
  assign n7071 = ( n625 & ~n2112 ) | ( n625 & n4643 ) | ( ~n2112 & n4643 ) ;
  assign n7072 = n1394 | n1981 ;
  assign n7073 = ( n4422 & n7071 ) | ( n4422 & ~n7072 ) | ( n7071 & ~n7072 ) ;
  assign n7069 = ~n2546 & n3322 ;
  assign n7070 = n7069 ^ n6544 ^ 1'b0 ;
  assign n7074 = n7073 ^ n7070 ^ 1'b0 ;
  assign n7075 = n1288 & ~n7074 ;
  assign n7076 = n1238 ^ n862 ^ n641 ;
  assign n7077 = ( ~n1531 & n4134 ) | ( ~n1531 & n7076 ) | ( n4134 & n7076 ) ;
  assign n7078 = ( ~n1887 & n4377 ) | ( ~n1887 & n4593 ) | ( n4377 & n4593 ) ;
  assign n7079 = ~n2994 & n7078 ;
  assign n7080 = n5674 & n7079 ;
  assign n7081 = ( n759 & n7077 ) | ( n759 & n7080 ) | ( n7077 & n7080 ) ;
  assign n7082 = n2108 ^ n1707 ^ n1509 ;
  assign n7083 = n7082 ^ n4776 ^ x242 ;
  assign n7084 = n7083 ^ n6504 ^ n3484 ;
  assign n7085 = n4726 ^ n904 ^ n842 ;
  assign n7086 = n3384 ^ x39 ^ 1'b0 ;
  assign n7097 = n6908 ^ n1647 ^ x159 ;
  assign n7087 = ( ~n1496 & n4129 ) | ( ~n1496 & n5979 ) | ( n4129 & n5979 ) ;
  assign n7093 = n1678 ^ n1469 ^ 1'b0 ;
  assign n7094 = n2039 | n7093 ;
  assign n7089 = n5687 ^ n2633 ^ n2265 ;
  assign n7088 = ( n974 & n1481 ) | ( n974 & n1674 ) | ( n1481 & n1674 ) ;
  assign n7090 = n7089 ^ n7088 ^ n2101 ;
  assign n7091 = n7090 ^ n5962 ^ 1'b0 ;
  assign n7092 = ~n1476 & n7091 ;
  assign n7095 = n7094 ^ n7092 ^ 1'b0 ;
  assign n7096 = ( n4970 & n7087 ) | ( n4970 & ~n7095 ) | ( n7087 & ~n7095 ) ;
  assign n7098 = n7097 ^ n7096 ^ n3286 ;
  assign n7099 = ( n7085 & n7086 ) | ( n7085 & ~n7098 ) | ( n7086 & ~n7098 ) ;
  assign n7100 = ( ~n1497 & n4472 ) | ( ~n1497 & n5091 ) | ( n4472 & n5091 ) ;
  assign n7101 = n7100 ^ n6508 ^ n5378 ;
  assign n7102 = ( n656 & ~n2722 ) | ( n656 & n4064 ) | ( ~n2722 & n4064 ) ;
  assign n7103 = ( ~n2911 & n3210 ) | ( ~n2911 & n3390 ) | ( n3210 & n3390 ) ;
  assign n7104 = n6458 & ~n7103 ;
  assign n7105 = ~n7102 & n7104 ;
  assign n7106 = ( n6648 & ~n7101 ) | ( n6648 & n7105 ) | ( ~n7101 & n7105 ) ;
  assign n7107 = n3191 ^ n1840 ^ n1115 ;
  assign n7108 = n7107 ^ n6367 ^ n2096 ;
  assign n7109 = n6788 & ~n7108 ;
  assign n7131 = ~n2172 & n2569 ;
  assign n7132 = ~n2268 & n7131 ;
  assign n7133 = n631 | n7132 ;
  assign n7134 = n7133 ^ n3236 ^ 1'b0 ;
  assign n7135 = ( n1410 & n1797 ) | ( n1410 & ~n7134 ) | ( n1797 & ~n7134 ) ;
  assign n7128 = n3125 ^ n1099 ^ n796 ;
  assign n7127 = ~n2819 & n4586 ;
  assign n7129 = n7128 ^ n7127 ^ n407 ;
  assign n7130 = n7129 ^ n3217 ^ x162 ;
  assign n7123 = ( ~n957 & n1391 ) | ( ~n957 & n1556 ) | ( n1391 & n1556 ) ;
  assign n7124 = n7123 ^ n3317 ^ n431 ;
  assign n7120 = ( n359 & ~n2049 ) | ( n359 & n7020 ) | ( ~n2049 & n7020 ) ;
  assign n7121 = n3709 ^ n1779 ^ 1'b0 ;
  assign n7122 = n7120 | n7121 ;
  assign n7125 = n7124 ^ n7122 ^ n1131 ;
  assign n7110 = ( ~n1814 & n2038 ) | ( ~n1814 & n2858 ) | ( n2038 & n2858 ) ;
  assign n7111 = ( n907 & n4467 ) | ( n907 & n7110 ) | ( n4467 & n7110 ) ;
  assign n7112 = ( n2744 & n3224 ) | ( n2744 & n3400 ) | ( n3224 & n3400 ) ;
  assign n7113 = n7112 ^ n1620 ^ n854 ;
  assign n7114 = n1869 ^ n1756 ^ 1'b0 ;
  assign n7115 = n7114 ^ n1658 ^ n1534 ;
  assign n7116 = ~n5490 & n7115 ;
  assign n7117 = ~n7113 & n7116 ;
  assign n7118 = ( n2031 & n7111 ) | ( n2031 & ~n7117 ) | ( n7111 & ~n7117 ) ;
  assign n7119 = n7118 ^ n5799 ^ n3908 ;
  assign n7126 = n7125 ^ n7119 ^ n748 ;
  assign n7136 = n7135 ^ n7130 ^ n7126 ;
  assign n7137 = ( n675 & ~n826 ) | ( n675 & n1278 ) | ( ~n826 & n1278 ) ;
  assign n7138 = n7137 ^ n2185 ^ n550 ;
  assign n7139 = n7138 ^ n5277 ^ n5009 ;
  assign n7140 = ( x18 & ~n2696 ) | ( x18 & n3153 ) | ( ~n2696 & n3153 ) ;
  assign n7141 = n7140 ^ n1460 ^ 1'b0 ;
  assign n7142 = n711 & ~n7141 ;
  assign n7143 = ( n1361 & n7139 ) | ( n1361 & ~n7142 ) | ( n7139 & ~n7142 ) ;
  assign n7144 = ( n4260 & ~n5261 ) | ( n4260 & n7143 ) | ( ~n5261 & n7143 ) ;
  assign n7147 = n2571 ^ n1697 ^ n1272 ;
  assign n7145 = ( n702 & ~n1336 ) | ( n702 & n4428 ) | ( ~n1336 & n4428 ) ;
  assign n7146 = n7145 ^ n5212 ^ n3755 ;
  assign n7148 = n7147 ^ n7146 ^ x48 ;
  assign n7149 = n7148 ^ n1919 ^ n1425 ;
  assign n7150 = n2970 & n5443 ;
  assign n7151 = n7149 | n7150 ;
  assign n7152 = n5090 & ~n7151 ;
  assign n7155 = n4971 ^ n290 ^ 1'b0 ;
  assign n7153 = n3069 ^ n2396 ^ n1983 ;
  assign n7154 = ( n3400 & n4627 ) | ( n3400 & n7153 ) | ( n4627 & n7153 ) ;
  assign n7156 = n7155 ^ n7154 ^ n2698 ;
  assign n7157 = n7156 ^ n580 ^ 1'b0 ;
  assign n7158 = n7157 ^ n5908 ^ n4001 ;
  assign n7159 = n3522 ^ n2523 ^ n356 ;
  assign n7160 = ( n4496 & ~n6150 ) | ( n4496 & n7159 ) | ( ~n6150 & n7159 ) ;
  assign n7161 = n7160 ^ n5413 ^ n1109 ;
  assign n7171 = n4663 ^ n3139 ^ 1'b0 ;
  assign n7162 = n1681 ^ n1235 ^ 1'b0 ;
  assign n7163 = n2742 ^ n288 ^ x120 ;
  assign n7164 = n7163 ^ n5267 ^ x220 ;
  assign n7165 = n6627 ^ n5459 ^ n2234 ;
  assign n7166 = n5700 ^ n2140 ^ n1394 ;
  assign n7167 = n7166 ^ n4899 ^ n3153 ;
  assign n7168 = ( n2286 & n7165 ) | ( n2286 & ~n7167 ) | ( n7165 & ~n7167 ) ;
  assign n7169 = n2985 & ~n7168 ;
  assign n7170 = ( n7162 & n7164 ) | ( n7162 & ~n7169 ) | ( n7164 & ~n7169 ) ;
  assign n7172 = n7171 ^ n7170 ^ n3389 ;
  assign n7175 = ( ~n935 & n1569 ) | ( ~n935 & n5009 ) | ( n1569 & n5009 ) ;
  assign n7173 = n1009 | n1151 ;
  assign n7174 = n685 & n7173 ;
  assign n7176 = n7175 ^ n7174 ^ 1'b0 ;
  assign n7177 = n7176 ^ n3980 ^ n1926 ;
  assign n7188 = n4141 ^ n1790 ^ n1308 ;
  assign n7187 = n4980 ^ n2859 ^ n2316 ;
  assign n7181 = n1956 ^ n1119 ^ 1'b0 ;
  assign n7183 = ( ~n1586 & n4691 ) | ( ~n1586 & n5007 ) | ( n4691 & n5007 ) ;
  assign n7182 = n2000 ^ n1016 ^ n897 ;
  assign n7184 = n7183 ^ n7182 ^ n585 ;
  assign n7185 = ( n3150 & ~n7181 ) | ( n3150 & n7184 ) | ( ~n7181 & n7184 ) ;
  assign n7186 = ( n3601 & n4734 ) | ( n3601 & ~n7185 ) | ( n4734 & ~n7185 ) ;
  assign n7189 = n7188 ^ n7187 ^ n7186 ;
  assign n7178 = n5525 ^ n1917 ^ n326 ;
  assign n7179 = n7178 ^ n5580 ^ n5527 ;
  assign n7180 = ( n1232 & n2056 ) | ( n1232 & n7179 ) | ( n2056 & n7179 ) ;
  assign n7190 = n7189 ^ n7180 ^ n1965 ;
  assign n7191 = ( ~n1738 & n7177 ) | ( ~n1738 & n7190 ) | ( n7177 & n7190 ) ;
  assign n7192 = ( ~n3500 & n3816 ) | ( ~n3500 & n6142 ) | ( n3816 & n6142 ) ;
  assign n7193 = n7192 ^ n1661 ^ n1631 ;
  assign n7194 = n7193 ^ n6276 ^ n3690 ;
  assign n7195 = ( n1416 & ~n1596 ) | ( n1416 & n1869 ) | ( ~n1596 & n1869 ) ;
  assign n7196 = n6279 ^ n4080 ^ n2767 ;
  assign n7197 = ( n2385 & n7195 ) | ( n2385 & n7196 ) | ( n7195 & n7196 ) ;
  assign n7198 = n4579 ^ n523 ^ 1'b0 ;
  assign n7201 = n3123 ^ n1880 ^ n536 ;
  assign n7202 = n7201 ^ n3083 ^ n1075 ;
  assign n7199 = n1478 ^ n1063 ^ n563 ;
  assign n7200 = ( n1939 & n5722 ) | ( n1939 & ~n7199 ) | ( n5722 & ~n7199 ) ;
  assign n7203 = n7202 ^ n7200 ^ n3462 ;
  assign n7204 = n7203 ^ n4447 ^ n1375 ;
  assign n7208 = ( n2463 & ~n2910 ) | ( n2463 & n6791 ) | ( ~n2910 & n6791 ) ;
  assign n7205 = ( ~n614 & n720 ) | ( ~n614 & n3345 ) | ( n720 & n3345 ) ;
  assign n7206 = n7205 ^ n3216 ^ n3198 ;
  assign n7207 = ( n4420 & ~n5976 ) | ( n4420 & n7206 ) | ( ~n5976 & n7206 ) ;
  assign n7209 = n7208 ^ n7207 ^ n5759 ;
  assign n7213 = x104 & ~n1962 ;
  assign n7214 = n7213 ^ n1244 ^ 1'b0 ;
  assign n7210 = n5101 ^ n4172 ^ 1'b0 ;
  assign n7211 = ~n7103 & n7210 ;
  assign n7212 = ( x172 & n3756 ) | ( x172 & ~n7211 ) | ( n3756 & ~n7211 ) ;
  assign n7215 = n7214 ^ n7212 ^ n1762 ;
  assign n7225 = n5223 ^ n4917 ^ n1011 ;
  assign n7226 = ~n1910 & n7225 ;
  assign n7227 = n7226 ^ n2536 ^ 1'b0 ;
  assign n7223 = n6811 ^ n2817 ^ 1'b0 ;
  assign n7224 = ( n1301 & n6450 ) | ( n1301 & ~n7223 ) | ( n6450 & ~n7223 ) ;
  assign n7216 = n4492 ^ n3283 ^ n1282 ;
  assign n7217 = n4387 ^ n1948 ^ x192 ;
  assign n7218 = n7217 ^ n4087 ^ n842 ;
  assign n7219 = ( n2593 & n3457 ) | ( n2593 & ~n7218 ) | ( n3457 & ~n7218 ) ;
  assign n7220 = n4241 & n7219 ;
  assign n7221 = n7216 & n7220 ;
  assign n7222 = n7221 ^ n4391 ^ 1'b0 ;
  assign n7228 = n7227 ^ n7224 ^ n7222 ;
  assign n7229 = ( n541 & n7215 ) | ( n541 & n7228 ) | ( n7215 & n7228 ) ;
  assign n7230 = x78 & n7229 ;
  assign n7231 = n7230 ^ n6841 ^ 1'b0 ;
  assign n7237 = n2869 ^ n2506 ^ 1'b0 ;
  assign n7238 = n7237 ^ n6921 ^ n3259 ;
  assign n7239 = ( n516 & ~n970 ) | ( n516 & n7238 ) | ( ~n970 & n7238 ) ;
  assign n7240 = n7239 ^ n1628 ^ n287 ;
  assign n7235 = n6087 ^ n2402 ^ 1'b0 ;
  assign n7236 = n2437 & n7235 ;
  assign n7233 = n6426 ^ n6161 ^ n1949 ;
  assign n7234 = ( n1590 & n4049 ) | ( n1590 & n7233 ) | ( n4049 & n7233 ) ;
  assign n7241 = n7240 ^ n7236 ^ n7234 ;
  assign n7232 = n5271 & n6853 ;
  assign n7242 = n7241 ^ n7232 ^ 1'b0 ;
  assign n7243 = ( ~x69 & n490 ) | ( ~x69 & n2591 ) | ( n490 & n2591 ) ;
  assign n7244 = ( n3348 & n3480 ) | ( n3348 & n6488 ) | ( n3480 & n6488 ) ;
  assign n7245 = ( n6421 & ~n7243 ) | ( n6421 & n7244 ) | ( ~n7243 & n7244 ) ;
  assign n7246 = n7245 ^ n6789 ^ n859 ;
  assign n7247 = n747 ^ n436 ^ n351 ;
  assign n7248 = n7247 ^ n959 ^ n358 ;
  assign n7249 = n5115 ^ n2618 ^ n1308 ;
  assign n7250 = ( ~n1381 & n3534 ) | ( ~n1381 & n7249 ) | ( n3534 & n7249 ) ;
  assign n7251 = ( n1023 & n2140 ) | ( n1023 & ~n3023 ) | ( n2140 & ~n3023 ) ;
  assign n7252 = ~n7216 & n7251 ;
  assign n7253 = n7252 ^ n6770 ^ n2500 ;
  assign n7254 = ( ~n7248 & n7250 ) | ( ~n7248 & n7253 ) | ( n7250 & n7253 ) ;
  assign n7255 = ( n1994 & n4204 ) | ( n1994 & n7254 ) | ( n4204 & n7254 ) ;
  assign n7256 = ( n3469 & ~n7246 ) | ( n3469 & n7255 ) | ( ~n7246 & n7255 ) ;
  assign n7257 = n6844 ^ n3043 ^ n887 ;
  assign n7258 = n1526 ^ n489 ^ 1'b0 ;
  assign n7259 = n7258 ^ n6103 ^ n1931 ;
  assign n7260 = n5836 ^ n2344 ^ 1'b0 ;
  assign n7261 = ( ~n4477 & n7259 ) | ( ~n4477 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7262 = n3503 ^ n1361 ^ n401 ;
  assign n7263 = ~n4816 & n7262 ;
  assign n7264 = ~n1758 & n7263 ;
  assign n7265 = n5701 ^ n4390 ^ n1637 ;
  assign n7266 = n7265 ^ n5966 ^ n2721 ;
  assign n7267 = ( n2871 & n7264 ) | ( n2871 & ~n7266 ) | ( n7264 & ~n7266 ) ;
  assign n7268 = ( n1926 & n7261 ) | ( n1926 & ~n7267 ) | ( n7261 & ~n7267 ) ;
  assign n7269 = n4469 ^ n3706 ^ 1'b0 ;
  assign n7270 = n4235 & n7269 ;
  assign n7271 = n565 & n7270 ;
  assign n7272 = ~n3963 & n7271 ;
  assign n7273 = ( n792 & n6216 ) | ( n792 & n7272 ) | ( n6216 & n7272 ) ;
  assign n7274 = n1392 | n1530 ;
  assign n7275 = ( n969 & n2069 ) | ( n969 & n3059 ) | ( n2069 & n3059 ) ;
  assign n7278 = n3194 ^ n1786 ^ n788 ;
  assign n7279 = ( n3432 & n4012 ) | ( n3432 & ~n7278 ) | ( n4012 & ~n7278 ) ;
  assign n7280 = n940 ^ x65 ^ 1'b0 ;
  assign n7281 = ~n7279 & n7280 ;
  assign n7276 = n4298 ^ n3498 ^ n3247 ;
  assign n7277 = ( x182 & n3083 ) | ( x182 & n7276 ) | ( n3083 & n7276 ) ;
  assign n7282 = n7281 ^ n7277 ^ n5088 ;
  assign n7289 = n2043 ^ n938 ^ 1'b0 ;
  assign n7288 = n6938 ^ n4098 ^ n1231 ;
  assign n7290 = n7289 ^ n7288 ^ 1'b0 ;
  assign n7286 = ( ~n2555 & n3005 ) | ( ~n2555 & n5644 ) | ( n3005 & n5644 ) ;
  assign n7283 = n2151 ^ n2044 ^ n957 ;
  assign n7284 = n4024 ^ n902 ^ n297 ;
  assign n7285 = ~n7283 & n7284 ;
  assign n7287 = n7286 ^ n7285 ^ 1'b0 ;
  assign n7291 = n7290 ^ n7287 ^ 1'b0 ;
  assign n7292 = n3124 & n7291 ;
  assign n7293 = n1829 ^ n1746 ^ n560 ;
  assign n7294 = n7293 ^ n5143 ^ 1'b0 ;
  assign n7295 = ( n753 & n2511 ) | ( n753 & ~n7294 ) | ( n2511 & ~n7294 ) ;
  assign n7296 = ( n3367 & ~n5044 ) | ( n3367 & n6396 ) | ( ~n5044 & n6396 ) ;
  assign n7297 = ( ~n285 & n3234 ) | ( ~n285 & n7296 ) | ( n3234 & n7296 ) ;
  assign n7298 = ( n1596 & ~n7295 ) | ( n1596 & n7297 ) | ( ~n7295 & n7297 ) ;
  assign n7299 = ( n999 & n7236 ) | ( n999 & n7298 ) | ( n7236 & n7298 ) ;
  assign n7300 = n7299 ^ n5292 ^ 1'b0 ;
  assign n7301 = n7292 & ~n7300 ;
  assign n7302 = n5351 ^ n4315 ^ n1014 ;
  assign n7303 = n7302 ^ n2539 ^ n2527 ;
  assign n7304 = ( n980 & n1608 ) | ( n980 & ~n3901 ) | ( n1608 & ~n3901 ) ;
  assign n7305 = n7304 ^ n308 ^ 1'b0 ;
  assign n7306 = n1195 | n7305 ;
  assign n7307 = n7306 ^ n3988 ^ n449 ;
  assign n7308 = ( n3065 & n3818 ) | ( n3065 & n6010 ) | ( n3818 & n6010 ) ;
  assign n7309 = n7308 ^ n3279 ^ 1'b0 ;
  assign n7310 = ~n7307 & n7309 ;
  assign n7313 = n2681 ^ n2102 ^ n858 ;
  assign n7311 = x253 & ~n1633 ;
  assign n7312 = n7311 ^ n3746 ^ 1'b0 ;
  assign n7314 = n7313 ^ n7312 ^ 1'b0 ;
  assign n7315 = n7314 ^ n4224 ^ 1'b0 ;
  assign n7316 = n1895 & ~n5889 ;
  assign n7318 = n2340 ^ n720 ^ 1'b0 ;
  assign n7319 = n2529 & ~n7318 ;
  assign n7317 = n315 | n1725 ;
  assign n7320 = n7319 ^ n7317 ^ 1'b0 ;
  assign n7321 = n7320 ^ n3904 ^ n2611 ;
  assign n7322 = ( x0 & n4243 ) | ( x0 & ~n7321 ) | ( n4243 & ~n7321 ) ;
  assign n7323 = n7316 & ~n7322 ;
  assign n7324 = n1527 ^ n534 ^ n463 ;
  assign n7325 = n7324 ^ n4877 ^ n4801 ;
  assign n7326 = n7325 ^ n4618 ^ 1'b0 ;
  assign n7346 = n4196 ^ n2679 ^ n1562 ;
  assign n7347 = n7346 ^ n4823 ^ 1'b0 ;
  assign n7348 = n2828 & ~n7347 ;
  assign n7343 = n3210 ^ n2344 ^ n1507 ;
  assign n7344 = ( n702 & n1162 ) | ( n702 & n2052 ) | ( n1162 & n2052 ) ;
  assign n7345 = ( n1337 & ~n7343 ) | ( n1337 & n7344 ) | ( ~n7343 & n7344 ) ;
  assign n7327 = n4169 ^ n2614 ^ 1'b0 ;
  assign n7328 = n7211 & n7327 ;
  assign n7329 = ( ~n3204 & n4604 ) | ( ~n3204 & n7328 ) | ( n4604 & n7328 ) ;
  assign n7330 = ( n815 & n2708 ) | ( n815 & n5918 ) | ( n2708 & n5918 ) ;
  assign n7331 = n7330 ^ x105 ^ 1'b0 ;
  assign n7332 = n7329 | n7331 ;
  assign n7338 = ~x78 & n1130 ;
  assign n7335 = ( n700 & n3316 ) | ( n700 & ~n6803 ) | ( n3316 & ~n6803 ) ;
  assign n7336 = n7319 & ~n7335 ;
  assign n7337 = n7336 ^ n5595 ^ 1'b0 ;
  assign n7333 = n4508 ^ n4156 ^ n1171 ;
  assign n7334 = ( n3115 & n5212 ) | ( n3115 & n7333 ) | ( n5212 & n7333 ) ;
  assign n7339 = n7338 ^ n7337 ^ n7334 ;
  assign n7340 = ~n7332 & n7339 ;
  assign n7341 = n7340 ^ n6185 ^ 1'b0 ;
  assign n7342 = n7341 ^ n2835 ^ n1737 ;
  assign n7349 = n7348 ^ n7345 ^ n7342 ;
  assign n7350 = n3212 ^ n1677 ^ n1014 ;
  assign n7351 = ( n2154 & ~n6550 ) | ( n2154 & n7350 ) | ( ~n6550 & n7350 ) ;
  assign n7352 = n5900 ^ n5240 ^ n781 ;
  assign n7353 = n2475 & ~n7352 ;
  assign n7354 = ( ~n743 & n1257 ) | ( ~n743 & n2489 ) | ( n1257 & n2489 ) ;
  assign n7355 = ( n3135 & n3753 ) | ( n3135 & n7354 ) | ( n3753 & n7354 ) ;
  assign n7356 = n7355 ^ n2433 ^ 1'b0 ;
  assign n7357 = n7353 | n7356 ;
  assign n7358 = ( n1189 & ~n1802 ) | ( n1189 & n4785 ) | ( ~n1802 & n4785 ) ;
  assign n7359 = n7358 ^ x240 ^ x54 ;
  assign n7360 = ( n7351 & n7357 ) | ( n7351 & n7359 ) | ( n7357 & n7359 ) ;
  assign n7361 = n1098 ^ n426 ^ 1'b0 ;
  assign n7362 = n7361 ^ n7221 ^ n2528 ;
  assign n7363 = n3932 & ~n7362 ;
  assign n7365 = n5257 ^ n1869 ^ 1'b0 ;
  assign n7366 = n7365 ^ n5309 ^ 1'b0 ;
  assign n7367 = n847 & n7366 ;
  assign n7368 = ( n438 & n4750 ) | ( n438 & ~n7367 ) | ( n4750 & ~n7367 ) ;
  assign n7369 = n7368 ^ n3735 ^ n2224 ;
  assign n7364 = ~n3339 & n4939 ;
  assign n7370 = n7369 ^ n7364 ^ 1'b0 ;
  assign n7371 = n7370 ^ n6218 ^ n1836 ;
  assign n7372 = n5182 ^ n1517 ^ n1228 ;
  assign n7373 = ( n360 & ~n989 ) | ( n360 & n6917 ) | ( ~n989 & n6917 ) ;
  assign n7374 = ( ~n4696 & n7372 ) | ( ~n4696 & n7373 ) | ( n7372 & n7373 ) ;
  assign n7375 = n5384 ^ n1909 ^ n281 ;
  assign n7380 = ( ~n1023 & n2263 ) | ( ~n1023 & n2776 ) | ( n2263 & n2776 ) ;
  assign n7381 = ( n337 & n2291 ) | ( n337 & ~n4309 ) | ( n2291 & ~n4309 ) ;
  assign n7382 = n7380 | n7381 ;
  assign n7383 = n7382 ^ n711 ^ 1'b0 ;
  assign n7378 = ( ~n507 & n2673 ) | ( ~n507 & n5126 ) | ( n2673 & n5126 ) ;
  assign n7376 = ~n5994 & n6574 ;
  assign n7377 = n7376 ^ n3223 ^ 1'b0 ;
  assign n7379 = n7378 ^ n7377 ^ n1165 ;
  assign n7384 = n7383 ^ n7379 ^ n6863 ;
  assign n7385 = ( n850 & ~n3003 ) | ( n850 & n3859 ) | ( ~n3003 & n3859 ) ;
  assign n7386 = n5105 | n7385 ;
  assign n7387 = n2551 | n7386 ;
  assign n7388 = n7387 ^ n3332 ^ n484 ;
  assign n7389 = ( n3304 & n4319 ) | ( n3304 & n4919 ) | ( n4319 & n4919 ) ;
  assign n7390 = n7389 ^ n5521 ^ 1'b0 ;
  assign n7391 = n7390 ^ n5292 ^ 1'b0 ;
  assign n7392 = ~n7388 & n7391 ;
  assign n7393 = n7392 ^ n4331 ^ n1262 ;
  assign n7394 = ( n2486 & n7384 ) | ( n2486 & n7393 ) | ( n7384 & n7393 ) ;
  assign n7395 = ( ~n3268 & n4729 ) | ( ~n3268 & n5753 ) | ( n4729 & n5753 ) ;
  assign n7399 = n1827 ^ n1342 ^ n351 ;
  assign n7400 = n7399 ^ n2278 ^ n2021 ;
  assign n7396 = n1421 ^ n809 ^ 1'b0 ;
  assign n7397 = n7396 ^ n2080 ^ n525 ;
  assign n7398 = n7397 ^ n1232 ^ n598 ;
  assign n7401 = n7400 ^ n7398 ^ n7114 ;
  assign n7402 = ( ~n4224 & n7395 ) | ( ~n4224 & n7401 ) | ( n7395 & n7401 ) ;
  assign n7403 = n5788 ^ n1946 ^ 1'b0 ;
  assign n7404 = ( n2769 & ~n3303 ) | ( n2769 & n3555 ) | ( ~n3303 & n3555 ) ;
  assign n7405 = n3962 ^ n3210 ^ n1917 ;
  assign n7406 = ~n341 & n7205 ;
  assign n7407 = n7406 ^ n2088 ^ 1'b0 ;
  assign n7408 = ( n7153 & n7405 ) | ( n7153 & ~n7407 ) | ( n7405 & ~n7407 ) ;
  assign n7409 = n1196 & n7343 ;
  assign n7410 = n7408 & ~n7409 ;
  assign n7411 = ~n7404 & n7410 ;
  assign n7412 = n3659 ^ n812 ^ x133 ;
  assign n7413 = x68 & ~n7412 ;
  assign n7414 = n7413 ^ n1218 ^ 1'b0 ;
  assign n7415 = ( n281 & n1784 ) | ( n281 & n7414 ) | ( n1784 & n7414 ) ;
  assign n7416 = n785 | n3650 ;
  assign n7417 = ( n1623 & n3653 ) | ( n1623 & n7416 ) | ( n3653 & n7416 ) ;
  assign n7418 = ( n671 & n5194 ) | ( n671 & ~n6851 ) | ( n5194 & ~n6851 ) ;
  assign n7419 = ( n3857 & n7417 ) | ( n3857 & ~n7418 ) | ( n7417 & ~n7418 ) ;
  assign n7420 = ( n1684 & n2139 ) | ( n1684 & n7419 ) | ( n2139 & n7419 ) ;
  assign n7425 = ( ~n1932 & n2019 ) | ( ~n1932 & n6136 ) | ( n2019 & n6136 ) ;
  assign n7426 = n7425 ^ n7066 ^ n5278 ;
  assign n7421 = n1915 ^ n362 ^ 1'b0 ;
  assign n7422 = n1418 & ~n7421 ;
  assign n7423 = ( n597 & ~n2910 ) | ( n597 & n4978 ) | ( ~n2910 & n4978 ) ;
  assign n7424 = ( n1058 & n7422 ) | ( n1058 & n7423 ) | ( n7422 & n7423 ) ;
  assign n7427 = n7426 ^ n7424 ^ n7167 ;
  assign n7429 = x168 & n3199 ;
  assign n7430 = n7429 ^ n4415 ^ 1'b0 ;
  assign n7428 = ( n2006 & n2686 ) | ( n2006 & n2807 ) | ( n2686 & n2807 ) ;
  assign n7431 = n7430 ^ n7428 ^ n4481 ;
  assign n7432 = n3287 ^ n2957 ^ n1819 ;
  assign n7433 = n7432 ^ n5690 ^ n3204 ;
  assign n7434 = n3218 ^ n3130 ^ n2219 ;
  assign n7435 = ( n2436 & n3091 ) | ( n2436 & n7434 ) | ( n3091 & n7434 ) ;
  assign n7436 = ( n2597 & n6446 ) | ( n2597 & n7435 ) | ( n6446 & n7435 ) ;
  assign n7437 = x176 & ~n7436 ;
  assign n7438 = ~n4398 & n7437 ;
  assign n7439 = n7433 & ~n7438 ;
  assign n7440 = n3866 & n6087 ;
  assign n7441 = n7440 ^ n3253 ^ 1'b0 ;
  assign n7442 = ~n658 & n3471 ;
  assign n7443 = ( n4509 & n7441 ) | ( n4509 & n7442 ) | ( n7441 & n7442 ) ;
  assign n7444 = ( n1098 & n3829 ) | ( n1098 & n6197 ) | ( n3829 & n6197 ) ;
  assign n7445 = ~n1784 & n7444 ;
  assign n7446 = ~n7443 & n7445 ;
  assign n7447 = n6328 ^ n5428 ^ n796 ;
  assign n7448 = ( x251 & n1121 ) | ( x251 & n3082 ) | ( n1121 & n3082 ) ;
  assign n7457 = ( x27 & ~n479 ) | ( x27 & n2251 ) | ( ~n479 & n2251 ) ;
  assign n7449 = ( n1161 & ~n1888 ) | ( n1161 & n2834 ) | ( ~n1888 & n2834 ) ;
  assign n7451 = n5624 ^ n815 ^ 1'b0 ;
  assign n7452 = n7451 ^ n6664 ^ 1'b0 ;
  assign n7453 = ( n3679 & ~n5795 ) | ( n3679 & n7452 ) | ( ~n5795 & n7452 ) ;
  assign n7450 = ~n1308 & n2887 ;
  assign n7454 = n7453 ^ n7450 ^ 1'b0 ;
  assign n7455 = ( n3500 & ~n5437 ) | ( n3500 & n6993 ) | ( ~n5437 & n6993 ) ;
  assign n7456 = ( n7449 & n7454 ) | ( n7449 & ~n7455 ) | ( n7454 & ~n7455 ) ;
  assign n7458 = n7457 ^ n7456 ^ 1'b0 ;
  assign n7459 = n7448 | n7458 ;
  assign n7460 = ( n4814 & n7447 ) | ( n4814 & n7459 ) | ( n7447 & n7459 ) ;
  assign n7461 = ( n1407 & ~n6283 ) | ( n1407 & n7092 ) | ( ~n6283 & n7092 ) ;
  assign n7475 = n4049 ^ n2621 ^ n1221 ;
  assign n7476 = ( ~n2271 & n5413 ) | ( ~n2271 & n7475 ) | ( n5413 & n7475 ) ;
  assign n7474 = n1373 | n5414 ;
  assign n7477 = n7476 ^ n7474 ^ 1'b0 ;
  assign n7471 = ( n2267 & ~n2855 ) | ( n2267 & n3742 ) | ( ~n2855 & n3742 ) ;
  assign n7472 = n1015 ^ n398 ^ x231 ;
  assign n7473 = ( ~n4040 & n7471 ) | ( ~n4040 & n7472 ) | ( n7471 & n7472 ) ;
  assign n7478 = n7477 ^ n7473 ^ n7196 ;
  assign n7464 = ( ~n2376 & n4032 ) | ( ~n2376 & n5634 ) | ( n4032 & n5634 ) ;
  assign n7462 = n6492 ^ n2356 ^ n659 ;
  assign n7463 = ( n6454 & n7202 ) | ( n6454 & n7462 ) | ( n7202 & n7462 ) ;
  assign n7465 = n7464 ^ n7463 ^ n4662 ;
  assign n7466 = ( n575 & ~n2302 ) | ( n575 & n6008 ) | ( ~n2302 & n6008 ) ;
  assign n7467 = ( n2044 & n5987 ) | ( n2044 & ~n6206 ) | ( n5987 & ~n6206 ) ;
  assign n7468 = n7467 ^ n3103 ^ n2454 ;
  assign n7469 = ( n1368 & ~n7466 ) | ( n1368 & n7468 ) | ( ~n7466 & n7468 ) ;
  assign n7470 = ( ~n3920 & n7465 ) | ( ~n3920 & n7469 ) | ( n7465 & n7469 ) ;
  assign n7479 = n7478 ^ n7470 ^ n1383 ;
  assign n7491 = n4712 ^ n3720 ^ 1'b0 ;
  assign n7492 = n1233 & ~n7491 ;
  assign n7480 = n5309 ^ n2112 ^ n1490 ;
  assign n7481 = ( n1435 & n4201 ) | ( n1435 & ~n7480 ) | ( n4201 & ~n7480 ) ;
  assign n7482 = n7481 ^ n3699 ^ 1'b0 ;
  assign n7487 = ( ~n2781 & n5084 ) | ( ~n2781 & n5895 ) | ( n5084 & n5895 ) ;
  assign n7483 = n4347 ^ n2021 ^ n1689 ;
  assign n7484 = ( n575 & n1106 ) | ( n575 & ~n4385 ) | ( n1106 & ~n4385 ) ;
  assign n7485 = n7483 & ~n7484 ;
  assign n7486 = n5597 & n7485 ;
  assign n7488 = n7487 ^ n7486 ^ n1805 ;
  assign n7489 = n7482 & n7488 ;
  assign n7490 = n7489 ^ n3458 ^ n2067 ;
  assign n7493 = n7492 ^ n7490 ^ n6002 ;
  assign n7494 = ( n3612 & n3780 ) | ( n3612 & n7128 ) | ( n3780 & n7128 ) ;
  assign n7495 = n7494 ^ n2548 ^ n1695 ;
  assign n7496 = n7495 ^ n3580 ^ n1504 ;
  assign n7497 = n1862 ^ n938 ^ n638 ;
  assign n7498 = n7497 ^ n2872 ^ 1'b0 ;
  assign n7499 = n738 & ~n7498 ;
  assign n7500 = n6327 ^ n1682 ^ n518 ;
  assign n7501 = n7499 & n7500 ;
  assign n7502 = ( n449 & ~n7496 ) | ( n449 & n7501 ) | ( ~n7496 & n7501 ) ;
  assign n7503 = ( n2881 & n5826 ) | ( n2881 & n7502 ) | ( n5826 & n7502 ) ;
  assign n7504 = n5161 ^ n1468 ^ 1'b0 ;
  assign n7505 = n4240 & ~n7504 ;
  assign n7506 = n7505 ^ n4748 ^ n926 ;
  assign n7507 = x131 | n7506 ;
  assign n7508 = ( n310 & n4144 ) | ( n310 & ~n7507 ) | ( n4144 & ~n7507 ) ;
  assign n7509 = ( n1102 & n1469 ) | ( n1102 & ~n4700 ) | ( n1469 & ~n4700 ) ;
  assign n7510 = ( n508 & n3726 ) | ( n508 & ~n7509 ) | ( n3726 & ~n7509 ) ;
  assign n7532 = ( n673 & ~n1652 ) | ( n673 & n6567 ) | ( ~n1652 & n6567 ) ;
  assign n7526 = n6783 ^ n3533 ^ x210 ;
  assign n7527 = ( ~n1499 & n3134 ) | ( ~n1499 & n7526 ) | ( n3134 & n7526 ) ;
  assign n7524 = n6194 ^ n5171 ^ n2963 ;
  assign n7525 = n7524 ^ n5752 ^ n294 ;
  assign n7528 = n7527 ^ n7525 ^ n1917 ;
  assign n7529 = ( n584 & ~n4182 ) | ( n584 & n4707 ) | ( ~n4182 & n4707 ) ;
  assign n7530 = n3457 & n7529 ;
  assign n7531 = n7528 & n7530 ;
  assign n7512 = n3082 | n3756 ;
  assign n7513 = n7512 ^ n2450 ^ 1'b0 ;
  assign n7511 = ( ~n1983 & n2737 ) | ( ~n1983 & n3914 ) | ( n2737 & n3914 ) ;
  assign n7514 = n7513 ^ n7511 ^ n2364 ;
  assign n7515 = ( n2012 & n2268 ) | ( n2012 & n2706 ) | ( n2268 & n2706 ) ;
  assign n7516 = n5069 ^ n4746 ^ n2487 ;
  assign n7517 = n7516 ^ n5968 ^ n1781 ;
  assign n7518 = ( ~n4899 & n7515 ) | ( ~n4899 & n7517 ) | ( n7515 & n7517 ) ;
  assign n7519 = ( n1535 & ~n7514 ) | ( n1535 & n7518 ) | ( ~n7514 & n7518 ) ;
  assign n7520 = n7519 ^ n5880 ^ x29 ;
  assign n7521 = n2526 ^ n413 ^ 1'b0 ;
  assign n7522 = n296 & ~n7521 ;
  assign n7523 = ( n5915 & n7520 ) | ( n5915 & n7522 ) | ( n7520 & n7522 ) ;
  assign n7533 = n7532 ^ n7531 ^ n7523 ;
  assign n7534 = ( n2098 & n7510 ) | ( n2098 & ~n7533 ) | ( n7510 & ~n7533 ) ;
  assign n7535 = ( ~n3210 & n7508 ) | ( ~n3210 & n7534 ) | ( n7508 & n7534 ) ;
  assign n7536 = ( n2697 & ~n2780 ) | ( n2697 & n4669 ) | ( ~n2780 & n4669 ) ;
  assign n7537 = n3866 ^ n3412 ^ 1'b0 ;
  assign n7538 = n7537 ^ n5607 ^ 1'b0 ;
  assign n7539 = ( ~n3848 & n7536 ) | ( ~n3848 & n7538 ) | ( n7536 & n7538 ) ;
  assign n7540 = n2762 ^ n1877 ^ x237 ;
  assign n7541 = ( n1974 & n3566 ) | ( n1974 & n5270 ) | ( n3566 & n5270 ) ;
  assign n7542 = n7541 ^ n3924 ^ n3623 ;
  assign n7543 = ( n2537 & n7540 ) | ( n2537 & ~n7542 ) | ( n7540 & ~n7542 ) ;
  assign n7544 = ( ~n5772 & n7539 ) | ( ~n5772 & n7543 ) | ( n7539 & n7543 ) ;
  assign n7545 = ( n578 & ~n5675 ) | ( n578 & n5860 ) | ( ~n5675 & n5860 ) ;
  assign n7546 = n7545 ^ n4740 ^ 1'b0 ;
  assign n7547 = n309 & n2684 ;
  assign n7552 = ( ~n1165 & n1399 ) | ( ~n1165 & n7399 ) | ( n1399 & n7399 ) ;
  assign n7550 = n1551 & n2774 ;
  assign n7551 = ~n4583 & n7550 ;
  assign n7553 = n7552 ^ n7551 ^ n449 ;
  assign n7554 = ( n2405 & n7032 ) | ( n2405 & ~n7553 ) | ( n7032 & ~n7553 ) ;
  assign n7555 = n7554 ^ n5145 ^ 1'b0 ;
  assign n7556 = n1392 & n7555 ;
  assign n7548 = ( x225 & n1088 ) | ( x225 & n1864 ) | ( n1088 & n1864 ) ;
  assign n7549 = n7548 ^ n4016 ^ 1'b0 ;
  assign n7557 = n7556 ^ n7549 ^ n5394 ;
  assign n7558 = n5931 ^ n5823 ^ n3373 ;
  assign n7559 = ( ~n3585 & n5395 ) | ( ~n3585 & n7558 ) | ( n5395 & n7558 ) ;
  assign n7560 = ( n4227 & ~n7557 ) | ( n4227 & n7559 ) | ( ~n7557 & n7559 ) ;
  assign n7561 = n7560 ^ n5347 ^ 1'b0 ;
  assign n7562 = n2410 & ~n7561 ;
  assign n7563 = n7208 ^ n6496 ^ n2428 ;
  assign n7564 = n7563 ^ n3768 ^ n2966 ;
  assign n7566 = ( ~n1283 & n1571 ) | ( ~n1283 & n3541 ) | ( n1571 & n3541 ) ;
  assign n7567 = ( n2228 & n2865 ) | ( n2228 & ~n7566 ) | ( n2865 & ~n7566 ) ;
  assign n7568 = n7567 ^ n5184 ^ n2225 ;
  assign n7565 = n5145 ^ n4485 ^ 1'b0 ;
  assign n7569 = n7568 ^ n7565 ^ n6814 ;
  assign n7570 = n7186 ^ n1261 ^ 1'b0 ;
  assign n7571 = x212 & n7570 ;
  assign n7574 = n6940 ^ n4331 ^ n4277 ;
  assign n7575 = ~n5667 & n7574 ;
  assign n7576 = n7575 ^ n382 ^ 1'b0 ;
  assign n7572 = ~n6255 & n6291 ;
  assign n7573 = ( n732 & ~n4651 ) | ( n732 & n7572 ) | ( ~n4651 & n7572 ) ;
  assign n7577 = n7576 ^ n7573 ^ n3895 ;
  assign n7578 = ( ~n6913 & n7118 ) | ( ~n6913 & n7577 ) | ( n7118 & n7577 ) ;
  assign n7579 = ( n2993 & n4436 ) | ( n2993 & n5759 ) | ( n4436 & n5759 ) ;
  assign n7580 = n6665 ^ n4536 ^ 1'b0 ;
  assign n7581 = n3842 & ~n7580 ;
  assign n7582 = ( ~n2126 & n3532 ) | ( ~n2126 & n7581 ) | ( n3532 & n7581 ) ;
  assign n7583 = n7579 & ~n7582 ;
  assign n7591 = n5009 ^ n4855 ^ n1173 ;
  assign n7592 = n3307 ^ n1039 ^ n496 ;
  assign n7593 = ( ~n278 & n7591 ) | ( ~n278 & n7592 ) | ( n7591 & n7592 ) ;
  assign n7594 = n2996 | n7593 ;
  assign n7595 = n5567 | n7594 ;
  assign n7588 = n2905 ^ n1317 ^ n1026 ;
  assign n7587 = ( ~n2038 & n3975 ) | ( ~n2038 & n4054 ) | ( n3975 & n4054 ) ;
  assign n7589 = n7588 ^ n7587 ^ 1'b0 ;
  assign n7590 = n675 & ~n7589 ;
  assign n7584 = n2112 ^ n1321 ^ x49 ;
  assign n7585 = n7584 ^ n1338 ^ x53 ;
  assign n7586 = n7585 ^ n7584 ^ n2046 ;
  assign n7596 = n7595 ^ n7590 ^ n7586 ;
  assign n7598 = n6027 ^ n938 ^ n537 ;
  assign n7597 = ( ~n480 & n1003 ) | ( ~n480 & n1580 ) | ( n1003 & n1580 ) ;
  assign n7599 = n7598 ^ n7597 ^ n4627 ;
  assign n7600 = ( n399 & n5834 ) | ( n399 & ~n7599 ) | ( n5834 & ~n7599 ) ;
  assign n7601 = ( n7583 & n7596 ) | ( n7583 & ~n7600 ) | ( n7596 & ~n7600 ) ;
  assign n7602 = n1561 ^ n1261 ^ x202 ;
  assign n7603 = ( ~n2202 & n6834 ) | ( ~n2202 & n7602 ) | ( n6834 & n7602 ) ;
  assign n7604 = ( ~n1016 & n2168 ) | ( ~n1016 & n4286 ) | ( n2168 & n4286 ) ;
  assign n7605 = n7604 ^ n5209 ^ n896 ;
  assign n7606 = ( x46 & ~n7603 ) | ( x46 & n7605 ) | ( ~n7603 & n7605 ) ;
  assign n7607 = n1858 ^ n640 ^ x197 ;
  assign n7608 = n2833 ^ n2718 ^ 1'b0 ;
  assign n7609 = ( n609 & ~n1510 ) | ( n609 & n7608 ) | ( ~n1510 & n7608 ) ;
  assign n7610 = ( n3889 & ~n7607 ) | ( n3889 & n7609 ) | ( ~n7607 & n7609 ) ;
  assign n7611 = n1469 | n7610 ;
  assign n7612 = ( n1302 & n7606 ) | ( n1302 & ~n7611 ) | ( n7606 & ~n7611 ) ;
  assign n7613 = ( ~n3591 & n4220 ) | ( ~n3591 & n7612 ) | ( n4220 & n7612 ) ;
  assign n7614 = ( n2470 & n2571 ) | ( n2470 & n4864 ) | ( n2571 & n4864 ) ;
  assign n7615 = ( n1456 & ~n3837 ) | ( n1456 & n5247 ) | ( ~n3837 & n5247 ) ;
  assign n7616 = n7615 ^ n5184 ^ 1'b0 ;
  assign n7617 = n7616 ^ n5403 ^ n396 ;
  assign n7625 = n7163 ^ n2163 ^ n1500 ;
  assign n7626 = n7625 ^ n7045 ^ n1577 ;
  assign n7619 = n4528 ^ n2068 ^ n1894 ;
  assign n7620 = n7619 ^ n2761 ^ 1'b0 ;
  assign n7621 = n2372 & ~n7620 ;
  assign n7618 = n4945 ^ n1309 ^ n1215 ;
  assign n7622 = n7621 ^ n7618 ^ 1'b0 ;
  assign n7623 = ( n1178 & ~n3284 ) | ( n1178 & n7622 ) | ( ~n3284 & n7622 ) ;
  assign n7624 = ( ~n1817 & n7481 ) | ( ~n1817 & n7623 ) | ( n7481 & n7623 ) ;
  assign n7627 = n7626 ^ n7624 ^ n2436 ;
  assign n7628 = n7627 ^ n7308 ^ n6321 ;
  assign n7629 = ( n3100 & n3355 ) | ( n3100 & ~n7513 ) | ( n3355 & ~n7513 ) ;
  assign n7632 = n536 | n1278 ;
  assign n7633 = n6217 | n7632 ;
  assign n7634 = ( n784 & ~n2962 ) | ( n784 & n7633 ) | ( ~n2962 & n7633 ) ;
  assign n7635 = n7634 ^ n4312 ^ n3034 ;
  assign n7630 = n4779 & ~n5961 ;
  assign n7631 = n3863 & n7630 ;
  assign n7636 = n7635 ^ n7631 ^ n342 ;
  assign n7637 = ( ~n3221 & n4314 ) | ( ~n3221 & n6918 ) | ( n4314 & n6918 ) ;
  assign n7638 = n7637 ^ n6279 ^ n3265 ;
  assign n7650 = ( n656 & n4037 ) | ( n656 & n7066 ) | ( n4037 & n7066 ) ;
  assign n7642 = n4564 ^ n2717 ^ 1'b0 ;
  assign n7643 = n3643 ^ n389 ^ n305 ;
  assign n7644 = ( n2197 & n3491 ) | ( n2197 & n4746 ) | ( n3491 & n4746 ) ;
  assign n7645 = n7644 ^ n6841 ^ n1196 ;
  assign n7646 = ( n504 & n3653 ) | ( n504 & ~n7645 ) | ( n3653 & ~n7645 ) ;
  assign n7647 = ( n2681 & n7643 ) | ( n2681 & n7646 ) | ( n7643 & n7646 ) ;
  assign n7648 = ( ~n2223 & n7642 ) | ( ~n2223 & n7647 ) | ( n7642 & n7647 ) ;
  assign n7639 = n5491 ^ n513 ^ 1'b0 ;
  assign n7640 = ~n5882 & n7639 ;
  assign n7641 = n7640 ^ n4807 ^ n1142 ;
  assign n7649 = n7648 ^ n7641 ^ n6240 ;
  assign n7651 = n7650 ^ n7649 ^ n496 ;
  assign n7652 = ( n298 & n2159 ) | ( n298 & n3623 ) | ( n2159 & n3623 ) ;
  assign n7653 = n2956 ^ n2488 ^ n639 ;
  assign n7654 = ( n1310 & n4575 ) | ( n1310 & n5921 ) | ( n4575 & n5921 ) ;
  assign n7655 = n3972 & ~n5964 ;
  assign n7656 = ( n4083 & n7654 ) | ( n4083 & ~n7655 ) | ( n7654 & ~n7655 ) ;
  assign n7657 = ( n6681 & ~n7653 ) | ( n6681 & n7656 ) | ( ~n7653 & n7656 ) ;
  assign n7658 = n7652 & n7657 ;
  assign n7659 = ( n1406 & ~n4050 ) | ( n1406 & n7658 ) | ( ~n4050 & n7658 ) ;
  assign n7661 = n5177 ^ n3006 ^ n1907 ;
  assign n7660 = n6049 ^ n3565 ^ n678 ;
  assign n7662 = n7661 ^ n7660 ^ n614 ;
  assign n7668 = n6192 ^ n5751 ^ n1090 ;
  assign n7669 = ( n4290 & n6041 ) | ( n4290 & n7668 ) | ( n6041 & n7668 ) ;
  assign n7664 = n2866 ^ n742 ^ 1'b0 ;
  assign n7665 = n2966 & n7664 ;
  assign n7666 = ( n556 & n984 ) | ( n556 & ~n6216 ) | ( n984 & ~n6216 ) ;
  assign n7667 = ( n6751 & n7665 ) | ( n6751 & ~n7666 ) | ( n7665 & ~n7666 ) ;
  assign n7663 = n6096 ^ n3585 ^ n1538 ;
  assign n7670 = n7669 ^ n7667 ^ n7663 ;
  assign n7671 = n4403 ^ n3052 ^ n2658 ;
  assign n7672 = ( n856 & ~n1938 ) | ( n856 & n7607 ) | ( ~n1938 & n7607 ) ;
  assign n7673 = n7672 ^ n7452 ^ n5093 ;
  assign n7674 = ( n1809 & ~n7671 ) | ( n1809 & n7673 ) | ( ~n7671 & n7673 ) ;
  assign n7675 = ( n295 & n1282 ) | ( n295 & ~n1595 ) | ( n1282 & ~n1595 ) ;
  assign n7676 = n7675 ^ n1548 ^ 1'b0 ;
  assign n7677 = ~n7674 & n7676 ;
  assign n7678 = n5642 ^ n2745 ^ n569 ;
  assign n7679 = n3307 ^ x67 ^ 1'b0 ;
  assign n7680 = n2257 & n7679 ;
  assign n7681 = ( ~n1343 & n5458 ) | ( ~n1343 & n7680 ) | ( n5458 & n7680 ) ;
  assign n7682 = n5473 | n6934 ;
  assign n7683 = ( n1084 & n3466 ) | ( n1084 & n7682 ) | ( n3466 & n7682 ) ;
  assign n7684 = n5824 ^ n3336 ^ n1542 ;
  assign n7690 = ( ~n1052 & n2452 ) | ( ~n1052 & n2774 ) | ( n2452 & n2774 ) ;
  assign n7691 = n7690 ^ n3658 ^ n1683 ;
  assign n7692 = ( x45 & n2987 ) | ( x45 & ~n7691 ) | ( n2987 & ~n7691 ) ;
  assign n7685 = n2196 ^ n759 ^ x250 ;
  assign n7686 = ( n4616 & ~n6852 ) | ( n4616 & n7685 ) | ( ~n6852 & n7685 ) ;
  assign n7687 = n5777 ^ n3040 ^ 1'b0 ;
  assign n7688 = n7686 | n7687 ;
  assign n7689 = n7688 ^ n5359 ^ x202 ;
  assign n7693 = n7692 ^ n7689 ^ 1'b0 ;
  assign n7694 = n3177 & n7693 ;
  assign n7695 = n7694 ^ n3543 ^ 1'b0 ;
  assign n7696 = ~n7684 & n7695 ;
  assign n7697 = n7696 ^ n7196 ^ 1'b0 ;
  assign n7700 = ( n534 & ~n2809 ) | ( n534 & n6345 ) | ( ~n2809 & n6345 ) ;
  assign n7701 = n2093 ^ n1892 ^ 1'b0 ;
  assign n7702 = ~n1397 & n7701 ;
  assign n7703 = n7702 ^ n4041 ^ n2549 ;
  assign n7704 = ( n5701 & ~n7700 ) | ( n5701 & n7703 ) | ( ~n7700 & n7703 ) ;
  assign n7705 = n1619 & ~n3513 ;
  assign n7706 = ~n7704 & n7705 ;
  assign n7707 = n5298 ^ n2221 ^ n2173 ;
  assign n7708 = n7706 | n7707 ;
  assign n7698 = ( ~n2977 & n3511 ) | ( ~n2977 & n4549 ) | ( n3511 & n4549 ) ;
  assign n7699 = ( n2359 & n7284 ) | ( n2359 & n7698 ) | ( n7284 & n7698 ) ;
  assign n7709 = n7708 ^ n7699 ^ n376 ;
  assign n7713 = n646 | n2373 ;
  assign n7714 = n696 & ~n7713 ;
  assign n7715 = ( x103 & n2863 ) | ( x103 & n7714 ) | ( n2863 & n7714 ) ;
  assign n7710 = n3199 ^ n319 ^ n261 ;
  assign n7711 = n2874 ^ n2420 ^ n1231 ;
  assign n7712 = ( ~n3731 & n7710 ) | ( ~n3731 & n7711 ) | ( n7710 & n7711 ) ;
  assign n7716 = n7715 ^ n7712 ^ 1'b0 ;
  assign n7717 = n5691 | n7716 ;
  assign n7718 = n7717 ^ n3066 ^ n740 ;
  assign n7721 = ( ~x48 & x58 ) | ( ~x48 & n1079 ) | ( x58 & n1079 ) ;
  assign n7722 = ~n5104 & n7721 ;
  assign n7723 = n3944 & n7722 ;
  assign n7719 = ( n3303 & ~n4955 ) | ( n3303 & n5548 ) | ( ~n4955 & n5548 ) ;
  assign n7720 = ( ~n937 & n7475 ) | ( ~n937 & n7719 ) | ( n7475 & n7719 ) ;
  assign n7724 = n7723 ^ n7720 ^ n2004 ;
  assign n7725 = ( n1683 & n2365 ) | ( n1683 & ~n5502 ) | ( n2365 & ~n5502 ) ;
  assign n7726 = ~n1479 & n7725 ;
  assign n7727 = n4770 & n7726 ;
  assign n7728 = ( n538 & n3971 ) | ( n538 & n4326 ) | ( n3971 & n4326 ) ;
  assign n7729 = ( n2541 & n6363 ) | ( n2541 & ~n7728 ) | ( n6363 & ~n7728 ) ;
  assign n7730 = ( n4677 & n7727 ) | ( n4677 & n7729 ) | ( n7727 & n7729 ) ;
  assign n7741 = n4134 ^ n2509 ^ n1201 ;
  assign n7737 = ( n830 & ~n2969 ) | ( n830 & n3272 ) | ( ~n2969 & n3272 ) ;
  assign n7738 = n7737 ^ n5746 ^ n3696 ;
  assign n7734 = ( ~x180 & n1740 ) | ( ~x180 & n6727 ) | ( n1740 & n6727 ) ;
  assign n7735 = ( x29 & x188 ) | ( x29 & n7734 ) | ( x188 & n7734 ) ;
  assign n7736 = n7735 ^ n2271 ^ 1'b0 ;
  assign n7739 = n7738 ^ n7736 ^ n659 ;
  assign n7740 = n7739 ^ n6417 ^ n5622 ;
  assign n7731 = n5069 ^ n3460 ^ n378 ;
  assign n7732 = ( n3870 & n5896 ) | ( n3870 & n7731 ) | ( n5896 & n7731 ) ;
  assign n7733 = n7732 ^ n7644 ^ n5942 ;
  assign n7742 = n7741 ^ n7740 ^ n7733 ;
  assign n7743 = n3539 ^ n3188 ^ n1436 ;
  assign n7744 = n7743 ^ n2484 ^ n1976 ;
  assign n7745 = ( n4352 & n5121 ) | ( n4352 & n7499 ) | ( n5121 & n7499 ) ;
  assign n7746 = n4453 ^ n4043 ^ n310 ;
  assign n7747 = n7154 ^ n5321 ^ n2571 ;
  assign n7748 = n6250 ^ n4345 ^ 1'b0 ;
  assign n7749 = ( ~n7746 & n7747 ) | ( ~n7746 & n7748 ) | ( n7747 & n7748 ) ;
  assign n7750 = n7490 ^ n6589 ^ 1'b0 ;
  assign n7751 = ( ~n7745 & n7749 ) | ( ~n7745 & n7750 ) | ( n7749 & n7750 ) ;
  assign n7755 = n3054 ^ n1103 ^ x171 ;
  assign n7756 = n7755 ^ n5286 ^ n3347 ;
  assign n7757 = ( n2015 & ~n7293 ) | ( n2015 & n7756 ) | ( ~n7293 & n7756 ) ;
  assign n7758 = n7757 ^ n3233 ^ 1'b0 ;
  assign n7759 = n2061 & n7758 ;
  assign n7760 = n7759 ^ n6665 ^ n283 ;
  assign n7752 = ( n312 & n1112 ) | ( n312 & ~n2105 ) | ( n1112 & ~n2105 ) ;
  assign n7753 = ( n514 & n1886 ) | ( n514 & n7752 ) | ( n1886 & n7752 ) ;
  assign n7754 = ( n5439 & n5701 ) | ( n5439 & n7753 ) | ( n5701 & n7753 ) ;
  assign n7761 = n7760 ^ n7754 ^ n3810 ;
  assign n7762 = n5159 | n6320 ;
  assign n7763 = n3283 | n7762 ;
  assign n7765 = n704 & n3553 ;
  assign n7766 = n7765 ^ n7163 ^ 1'b0 ;
  assign n7764 = n4012 ^ n383 ^ x108 ;
  assign n7767 = n7766 ^ n7764 ^ n3977 ;
  assign n7768 = ~n3130 & n7767 ;
  assign n7769 = n7275 ^ n1605 ^ 1'b0 ;
  assign n7770 = n5163 ^ n891 ^ n607 ;
  assign n7771 = n3843 ^ n3781 ^ n2715 ;
  assign n7772 = n7771 ^ n3244 ^ n2647 ;
  assign n7773 = n7772 ^ n4514 ^ 1'b0 ;
  assign n7774 = ~n6824 & n7773 ;
  assign n7775 = ( n6068 & ~n7770 ) | ( n6068 & n7774 ) | ( ~n7770 & n7774 ) ;
  assign n7776 = n5194 ^ n2875 ^ n2640 ;
  assign n7777 = n555 ^ x167 ^ 1'b0 ;
  assign n7778 = n7776 | n7777 ;
  assign n7784 = n3639 ^ n751 ^ n320 ;
  assign n7785 = ( n2695 & n5980 ) | ( n2695 & ~n6197 ) | ( n5980 & ~n6197 ) ;
  assign n7786 = ( ~n2456 & n7784 ) | ( ~n2456 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7787 = n7786 ^ n1024 ^ 1'b0 ;
  assign n7779 = ( ~n690 & n1122 ) | ( ~n690 & n2621 ) | ( n1122 & n2621 ) ;
  assign n7780 = n5938 ^ n1430 ^ 1'b0 ;
  assign n7781 = n7780 ^ x49 ^ 1'b0 ;
  assign n7782 = n7779 & n7781 ;
  assign n7783 = n7782 ^ n6373 ^ x61 ;
  assign n7788 = n7787 ^ n7783 ^ n345 ;
  assign n7789 = ( n323 & n2393 ) | ( n323 & ~n2838 ) | ( n2393 & ~n2838 ) ;
  assign n7790 = n5501 ^ n2141 ^ x200 ;
  assign n7791 = n7790 ^ n3443 ^ 1'b0 ;
  assign n7792 = ( n3183 & n7789 ) | ( n3183 & n7791 ) | ( n7789 & n7791 ) ;
  assign n7793 = n4922 ^ n1059 ^ n542 ;
  assign n7800 = ( n262 & ~n294 ) | ( n262 & n2099 ) | ( ~n294 & n2099 ) ;
  assign n7801 = n7800 ^ n2097 ^ 1'b0 ;
  assign n7802 = n317 & ~n7801 ;
  assign n7794 = ( ~n1159 & n1279 ) | ( ~n1159 & n1990 ) | ( n1279 & n1990 ) ;
  assign n7795 = ( n2514 & ~n5368 ) | ( n2514 & n7794 ) | ( ~n5368 & n7794 ) ;
  assign n7796 = n6934 ^ n1837 ^ 1'b0 ;
  assign n7797 = ~n7795 & n7796 ;
  assign n7798 = n329 & n7797 ;
  assign n7799 = n7798 ^ n1415 ^ 1'b0 ;
  assign n7803 = n7802 ^ n7799 ^ n1689 ;
  assign n7804 = n6705 ^ n827 ^ n493 ;
  assign n7805 = ( n5169 & ~n6592 ) | ( n5169 & n7804 ) | ( ~n6592 & n7804 ) ;
  assign n7806 = ( n323 & n2982 ) | ( n323 & n6827 ) | ( n2982 & n6827 ) ;
  assign n7807 = n7806 ^ n5319 ^ n829 ;
  assign n7808 = ( n2701 & n3526 ) | ( n2701 & n5869 ) | ( n3526 & n5869 ) ;
  assign n7809 = ( ~n4320 & n4823 ) | ( ~n4320 & n5401 ) | ( n4823 & n5401 ) ;
  assign n7811 = ( x112 & ~x210 ) | ( x112 & n534 ) | ( ~x210 & n534 ) ;
  assign n7810 = n2476 ^ n1770 ^ n406 ;
  assign n7812 = n7811 ^ n7810 ^ n3650 ;
  assign n7813 = ( ~n7808 & n7809 ) | ( ~n7808 & n7812 ) | ( n7809 & n7812 ) ;
  assign n7814 = ( ~n3811 & n6257 ) | ( ~n3811 & n7813 ) | ( n6257 & n7813 ) ;
  assign n7815 = n6143 ^ n1411 ^ n490 ;
  assign n7816 = ( n1540 & n4502 ) | ( n1540 & n7494 ) | ( n4502 & n7494 ) ;
  assign n7817 = n7816 ^ n1563 ^ n1278 ;
  assign n7818 = n7817 ^ n2166 ^ 1'b0 ;
  assign n7819 = ( ~n297 & n7815 ) | ( ~n297 & n7818 ) | ( n7815 & n7818 ) ;
  assign n7820 = ( n7807 & n7814 ) | ( n7807 & ~n7819 ) | ( n7814 & ~n7819 ) ;
  assign n7821 = n7388 ^ n6137 ^ n1349 ;
  assign n7824 = n2462 ^ n1081 ^ 1'b0 ;
  assign n7822 = ( n1784 & ~n4439 ) | ( n1784 & n7735 ) | ( ~n4439 & n7735 ) ;
  assign n7823 = ( n946 & ~n4981 ) | ( n946 & n7822 ) | ( ~n4981 & n7822 ) ;
  assign n7825 = n7824 ^ n7823 ^ n7286 ;
  assign n7826 = n7483 & ~n7825 ;
  assign n7827 = ~n1220 & n7826 ;
  assign n7828 = n4744 ^ n2540 ^ n817 ;
  assign n7829 = n1071 | n7828 ;
  assign n7830 = n7829 ^ n6798 ^ n4144 ;
  assign n7831 = n7830 ^ n7760 ^ n3296 ;
  assign n7832 = n351 & ~n1573 ;
  assign n7833 = n7832 ^ n1840 ^ n1061 ;
  assign n7834 = ( ~n3779 & n4133 ) | ( ~n3779 & n7833 ) | ( n4133 & n7833 ) ;
  assign n7837 = n3594 ^ n3530 ^ n2119 ;
  assign n7838 = ( ~n736 & n5110 ) | ( ~n736 & n7837 ) | ( n5110 & n7837 ) ;
  assign n7839 = n7838 ^ n6654 ^ n1789 ;
  assign n7835 = n5642 ^ n4459 ^ n2527 ;
  assign n7836 = n1298 | n7835 ;
  assign n7840 = n7839 ^ n7836 ^ 1'b0 ;
  assign n7850 = n6792 ^ n6610 ^ n1199 ;
  assign n7848 = ( n1042 & n1360 ) | ( n1042 & ~n4620 ) | ( n1360 & ~n4620 ) ;
  assign n7847 = ( n5288 & n6594 ) | ( n5288 & n7475 ) | ( n6594 & n7475 ) ;
  assign n7846 = n4412 ^ n3956 ^ 1'b0 ;
  assign n7849 = n7848 ^ n7847 ^ n7846 ;
  assign n7841 = ( n1950 & ~n3110 ) | ( n1950 & n6485 ) | ( ~n3110 & n6485 ) ;
  assign n7842 = n7841 ^ n2984 ^ n2687 ;
  assign n7843 = n1458 ^ n684 ^ 1'b0 ;
  assign n7844 = n7196 | n7843 ;
  assign n7845 = ( ~n4324 & n7842 ) | ( ~n4324 & n7844 ) | ( n7842 & n7844 ) ;
  assign n7851 = n7850 ^ n7849 ^ n7845 ;
  assign n7855 = n5033 ^ n4732 ^ x20 ;
  assign n7852 = n4000 ^ n1864 ^ 1'b0 ;
  assign n7853 = n6683 & ~n7852 ;
  assign n7854 = n7853 ^ n6867 ^ n2441 ;
  assign n7856 = n7855 ^ n7854 ^ n6804 ;
  assign n7857 = ( n956 & n3332 ) | ( n956 & ~n3791 ) | ( n3332 & ~n3791 ) ;
  assign n7858 = ( x112 & n1233 ) | ( x112 & ~n7857 ) | ( n1233 & ~n7857 ) ;
  assign n7859 = ( n303 & ~n1263 ) | ( n303 & n6840 ) | ( ~n1263 & n6840 ) ;
  assign n7860 = n7859 ^ n7237 ^ n2443 ;
  assign n7861 = n7860 ^ n5218 ^ n3216 ;
  assign n7862 = ( n4417 & ~n7858 ) | ( n4417 & n7861 ) | ( ~n7858 & n7861 ) ;
  assign n7863 = n3815 ^ n2662 ^ n638 ;
  assign n7864 = n7863 ^ n3154 ^ n1570 ;
  assign n7865 = n4123 ^ n2224 ^ n1294 ;
  assign n7866 = n5177 ^ n2715 ^ n678 ;
  assign n7867 = ( n3215 & n7865 ) | ( n3215 & ~n7866 ) | ( n7865 & ~n7866 ) ;
  assign n7868 = ( ~n4320 & n7864 ) | ( ~n4320 & n7867 ) | ( n7864 & n7867 ) ;
  assign n7869 = n6391 ^ n4748 ^ n1479 ;
  assign n7870 = ~n6832 & n7869 ;
  assign n7871 = n7870 ^ n6993 ^ n1006 ;
  assign n7872 = n7611 ^ n5030 ^ n3062 ;
  assign n7873 = ( n465 & n7205 ) | ( n465 & n7872 ) | ( n7205 & n7872 ) ;
  assign n7874 = n1534 & ~n7873 ;
  assign n7875 = n5543 ^ n1093 ^ n386 ;
  assign n7876 = ( ~n6293 & n6351 ) | ( ~n6293 & n7875 ) | ( n6351 & n7875 ) ;
  assign n7880 = n1157 ^ n1042 ^ n1001 ;
  assign n7877 = ( n367 & n1281 ) | ( n367 & n2234 ) | ( n1281 & n2234 ) ;
  assign n7878 = n7877 ^ n357 ^ 1'b0 ;
  assign n7879 = n6792 & ~n7878 ;
  assign n7881 = n7880 ^ n7879 ^ n5029 ;
  assign n7898 = n323 ^ n269 ^ 1'b0 ;
  assign n7897 = ( n1651 & ~n2884 ) | ( n1651 & n5808 ) | ( ~n2884 & n5808 ) ;
  assign n7899 = n7898 ^ n7897 ^ n1598 ;
  assign n7895 = n5007 ^ n823 ^ 1'b0 ;
  assign n7892 = n6999 ^ n2287 ^ 1'b0 ;
  assign n7891 = n6695 | n7680 ;
  assign n7893 = n7892 ^ n7891 ^ n2716 ;
  assign n7885 = n410 | n2655 ;
  assign n7886 = n7885 ^ n4316 ^ 1'b0 ;
  assign n7887 = n7886 ^ n6598 ^ n2070 ;
  assign n7888 = n1976 ^ n1762 ^ n1272 ;
  assign n7889 = n4701 ^ n3216 ^ n1191 ;
  assign n7890 = ( n7887 & n7888 ) | ( n7887 & ~n7889 ) | ( n7888 & ~n7889 ) ;
  assign n7884 = n2470 | n7650 ;
  assign n7894 = n7893 ^ n7890 ^ n7884 ;
  assign n7896 = n7895 ^ n7894 ^ n5854 ;
  assign n7882 = n2614 ^ n1547 ^ 1'b0 ;
  assign n7883 = n7882 ^ n6982 ^ 1'b0 ;
  assign n7900 = n7899 ^ n7896 ^ n7883 ;
  assign n7901 = n6103 ^ n4263 ^ n702 ;
  assign n7902 = ( n3622 & n7401 ) | ( n3622 & ~n7901 ) | ( n7401 & ~n7901 ) ;
  assign n7903 = n3171 ^ n1716 ^ n1335 ;
  assign n7904 = n7903 ^ n6545 ^ n5780 ;
  assign n7908 = n1562 ^ n1080 ^ n874 ;
  assign n7905 = ( n1874 & n4606 ) | ( n1874 & n4775 ) | ( n4606 & n4775 ) ;
  assign n7906 = n4196 | n7905 ;
  assign n7907 = ( n3451 & n4776 ) | ( n3451 & n7906 ) | ( n4776 & n7906 ) ;
  assign n7909 = n7908 ^ n7907 ^ n7457 ;
  assign n7910 = ( n1810 & n4422 ) | ( n1810 & n6494 ) | ( n4422 & n6494 ) ;
  assign n7911 = ( x180 & n3764 ) | ( x180 & n7910 ) | ( n3764 & n7910 ) ;
  assign n7912 = ( n964 & ~n2875 ) | ( n964 & n7911 ) | ( ~n2875 & n7911 ) ;
  assign n7913 = n2369 | n7912 ;
  assign n7914 = n1206 & ~n7913 ;
  assign n7915 = ( ~n7423 & n7909 ) | ( ~n7423 & n7914 ) | ( n7909 & n7914 ) ;
  assign n7918 = n4222 ^ n736 ^ n496 ;
  assign n7917 = n3834 & ~n6935 ;
  assign n7919 = n7918 ^ n7917 ^ 1'b0 ;
  assign n7916 = ( n621 & n1497 ) | ( n621 & ~n2037 ) | ( n1497 & ~n2037 ) ;
  assign n7920 = n7919 ^ n7916 ^ n1505 ;
  assign n7925 = ( x94 & n938 ) | ( x94 & ~n1473 ) | ( n938 & ~n1473 ) ;
  assign n7921 = n4685 ^ n1587 ^ x64 ;
  assign n7922 = ( n2666 & n5944 ) | ( n2666 & ~n7921 ) | ( n5944 & ~n7921 ) ;
  assign n7923 = ( ~x21 & n1742 ) | ( ~x21 & n7922 ) | ( n1742 & n7922 ) ;
  assign n7924 = n7923 ^ n2780 ^ n1343 ;
  assign n7926 = n7925 ^ n7924 ^ n773 ;
  assign n7927 = ( n646 & ~n2337 ) | ( n646 & n7926 ) | ( ~n2337 & n7926 ) ;
  assign n7928 = ( n3929 & n6166 ) | ( n3929 & n7927 ) | ( n6166 & n7927 ) ;
  assign n7930 = n2195 ^ n1511 ^ n694 ;
  assign n7929 = n3501 ^ n2938 ^ n1048 ;
  assign n7931 = n7930 ^ n7929 ^ n3731 ;
  assign n7932 = ( ~x26 & n1468 ) | ( ~x26 & n3950 ) | ( n1468 & n3950 ) ;
  assign n7933 = ( n1069 & ~n4322 ) | ( n1069 & n7932 ) | ( ~n4322 & n7932 ) ;
  assign n7934 = n7933 ^ n2464 ^ x25 ;
  assign n7935 = n7931 & ~n7934 ;
  assign n7936 = n7935 ^ n7283 ^ 1'b0 ;
  assign n7937 = n7936 ^ n2287 ^ n1239 ;
  assign n7938 = n7618 ^ n7595 ^ 1'b0 ;
  assign n7939 = ( x250 & n3427 ) | ( x250 & ~n7553 ) | ( n3427 & ~n7553 ) ;
  assign n7940 = n7939 ^ n4487 ^ n744 ;
  assign n7941 = ( n1927 & n1991 ) | ( n1927 & n7940 ) | ( n1991 & n7940 ) ;
  assign n7942 = ( ~n7683 & n7938 ) | ( ~n7683 & n7941 ) | ( n7938 & n7941 ) ;
  assign n7943 = n4638 ^ n3512 ^ n487 ;
  assign n7944 = ( n789 & ~n1663 ) | ( n789 & n6425 ) | ( ~n1663 & n6425 ) ;
  assign n7945 = n7944 ^ n6945 ^ 1'b0 ;
  assign n7946 = ( ~n5310 & n7943 ) | ( ~n5310 & n7945 ) | ( n7943 & n7945 ) ;
  assign n7947 = n5915 ^ n4969 ^ n2570 ;
  assign n7948 = n4915 ^ n2207 ^ n830 ;
  assign n7949 = ( n6090 & ~n7947 ) | ( n6090 & n7948 ) | ( ~n7947 & n7948 ) ;
  assign n7958 = ( n558 & ~n5094 ) | ( n558 & n7120 ) | ( ~n5094 & n7120 ) ;
  assign n7955 = n5759 ^ n4638 ^ n1345 ;
  assign n7956 = ( n626 & ~n5351 ) | ( n626 & n7955 ) | ( ~n5351 & n7955 ) ;
  assign n7957 = ( n998 & n2679 ) | ( n998 & ~n7956 ) | ( n2679 & ~n7956 ) ;
  assign n7959 = n7958 ^ n7957 ^ n1862 ;
  assign n7952 = n4201 ^ n591 ^ n486 ;
  assign n7953 = ( ~n1210 & n3566 ) | ( ~n1210 & n7952 ) | ( n3566 & n7952 ) ;
  assign n7950 = n804 & ~n6132 ;
  assign n7951 = n7950 ^ n1527 ^ 1'b0 ;
  assign n7954 = n7953 ^ n7951 ^ n2675 ;
  assign n7960 = n7959 ^ n7954 ^ n1898 ;
  assign n7961 = ~n1233 & n1976 ;
  assign n7962 = ( ~n3797 & n6979 ) | ( ~n3797 & n7790 ) | ( n6979 & n7790 ) ;
  assign n7963 = n2327 ^ n1152 ^ x78 ;
  assign n7964 = n7963 ^ n2758 ^ n1778 ;
  assign n7965 = n7964 ^ n6328 ^ n6148 ;
  assign n7966 = ( ~n1108 & n7962 ) | ( ~n1108 & n7965 ) | ( n7962 & n7965 ) ;
  assign n7972 = n4439 ^ n828 ^ x153 ;
  assign n7971 = n1309 ^ n1210 ^ 1'b0 ;
  assign n7973 = n7972 ^ n7971 ^ n4427 ;
  assign n7974 = n5597 & n7973 ;
  assign n7967 = n1701 ^ n1576 ^ n945 ;
  assign n7968 = ( n722 & n5860 ) | ( n722 & n7967 ) | ( n5860 & n7967 ) ;
  assign n7969 = n6170 ^ n3334 ^ n1596 ;
  assign n7970 = ~n7968 & n7969 ;
  assign n7975 = n7974 ^ n7970 ^ 1'b0 ;
  assign n7976 = n1784 | n5383 ;
  assign n7977 = n7976 ^ n4782 ^ 1'b0 ;
  assign n7978 = ( n806 & n2241 ) | ( n806 & n2572 ) | ( n2241 & n2572 ) ;
  assign n7980 = ( x10 & ~x156 ) | ( x10 & n2067 ) | ( ~x156 & n2067 ) ;
  assign n7979 = ~n3762 & n4460 ;
  assign n7981 = n7980 ^ n7979 ^ n1777 ;
  assign n7982 = ( n7977 & ~n7978 ) | ( n7977 & n7981 ) | ( ~n7978 & n7981 ) ;
  assign n7983 = n7982 ^ n3135 ^ 1'b0 ;
  assign n7984 = n4206 & n7983 ;
  assign n7985 = n6441 ^ n6189 ^ 1'b0 ;
  assign n7986 = n6663 | n7985 ;
  assign n7994 = n3363 ^ n973 ^ n461 ;
  assign n7995 = n6996 & ~n7994 ;
  assign n7991 = ( n1471 & n1664 ) | ( n1471 & n4331 ) | ( n1664 & n4331 ) ;
  assign n7992 = n7991 ^ n3560 ^ x215 ;
  assign n7987 = n6237 ^ n666 ^ x44 ;
  assign n7988 = n7987 ^ n2001 ^ n1215 ;
  assign n7989 = n7988 ^ n5457 ^ n4506 ;
  assign n7990 = n7989 ^ n5253 ^ n1902 ;
  assign n7993 = n7992 ^ n7990 ^ n4504 ;
  assign n7996 = n7995 ^ n7993 ^ n4169 ;
  assign n7998 = n3723 | n5500 ;
  assign n7999 = ( ~n3701 & n7857 ) | ( ~n3701 & n7998 ) | ( n7857 & n7998 ) ;
  assign n7997 = n7378 ^ n6802 ^ n1518 ;
  assign n8000 = n7999 ^ n7997 ^ n1296 ;
  assign n8001 = ( n1774 & ~n5985 ) | ( n1774 & n8000 ) | ( ~n5985 & n8000 ) ;
  assign n8002 = n6884 ^ n5660 ^ n1749 ;
  assign n8013 = n3705 ^ n747 ^ x73 ;
  assign n8014 = ( ~n2013 & n7064 ) | ( ~n2013 & n8013 ) | ( n7064 & n8013 ) ;
  assign n8003 = ( n2905 & n3406 ) | ( n2905 & ~n3889 ) | ( n3406 & ~n3889 ) ;
  assign n8004 = ( ~n1926 & n3954 ) | ( ~n1926 & n8003 ) | ( n3954 & n8003 ) ;
  assign n8005 = n2108 ^ n622 ^ n609 ;
  assign n8006 = n8005 ^ n7933 ^ n4171 ;
  assign n8007 = ( n1134 & n3067 ) | ( n1134 & n8006 ) | ( n3067 & n8006 ) ;
  assign n8008 = ( n264 & n404 ) | ( n264 & n8007 ) | ( n404 & n8007 ) ;
  assign n8009 = ( x150 & n781 ) | ( x150 & n8008 ) | ( n781 & n8008 ) ;
  assign n8010 = n8009 ^ n6095 ^ x131 ;
  assign n8011 = ( ~n4134 & n4308 ) | ( ~n4134 & n5306 ) | ( n4308 & n5306 ) ;
  assign n8012 = ( ~n8004 & n8010 ) | ( ~n8004 & n8011 ) | ( n8010 & n8011 ) ;
  assign n8015 = n8014 ^ n8012 ^ n6516 ;
  assign n8016 = ( n334 & n2125 ) | ( n334 & n4093 ) | ( n2125 & n4093 ) ;
  assign n8017 = n8016 ^ n5855 ^ n882 ;
  assign n8018 = n8017 ^ n7215 ^ n6119 ;
  assign n8019 = n6051 | n8018 ;
  assign n8020 = n2263 & n2724 ;
  assign n8021 = n3922 ^ n759 ^ 1'b0 ;
  assign n8022 = x160 & n8021 ;
  assign n8023 = ( n3098 & n3449 ) | ( n3098 & ~n8022 ) | ( n3449 & ~n8022 ) ;
  assign n8024 = n6501 ^ n5699 ^ 1'b0 ;
  assign n8025 = n6174 ^ n6049 ^ n5397 ;
  assign n8026 = ( x244 & n2814 ) | ( x244 & n8025 ) | ( n2814 & n8025 ) ;
  assign n8027 = ( n7354 & n8024 ) | ( n7354 & ~n8026 ) | ( n8024 & ~n8026 ) ;
  assign n8028 = ~n473 & n5424 ;
  assign n8029 = ( ~n1445 & n1725 ) | ( ~n1445 & n7991 ) | ( n1725 & n7991 ) ;
  assign n8030 = n3019 ^ n532 ^ x205 ;
  assign n8031 = n5238 ^ n4094 ^ x199 ;
  assign n8032 = n8031 ^ x251 ^ 1'b0 ;
  assign n8033 = n8032 ^ n2877 ^ n288 ;
  assign n8034 = ( n7500 & n8030 ) | ( n7500 & n8033 ) | ( n8030 & n8033 ) ;
  assign n8035 = n4627 ^ n2757 ^ x149 ;
  assign n8036 = n8035 ^ n2861 ^ n1701 ;
  assign n8037 = n4625 ^ n3688 ^ n3643 ;
  assign n8038 = ~n2238 & n8037 ;
  assign n8039 = ~n8036 & n8038 ;
  assign n8040 = ( n1362 & ~n1622 ) | ( n1362 & n2110 ) | ( ~n1622 & n2110 ) ;
  assign n8041 = n8040 ^ n6840 ^ n5405 ;
  assign n8042 = ( n1470 & n5742 ) | ( n1470 & ~n8041 ) | ( n5742 & ~n8041 ) ;
  assign n8043 = n8042 ^ n5011 ^ n4993 ;
  assign n8044 = ( n2586 & ~n3893 ) | ( n2586 & n4988 ) | ( ~n3893 & n4988 ) ;
  assign n8046 = ~n6091 & n6191 ;
  assign n8047 = n8046 ^ n2493 ^ 1'b0 ;
  assign n8045 = n2074 ^ n1647 ^ x131 ;
  assign n8048 = n8047 ^ n8045 ^ n6020 ;
  assign n8049 = ( n5790 & ~n8044 ) | ( n5790 & n8048 ) | ( ~n8044 & n8048 ) ;
  assign n8050 = ( ~n3666 & n4682 ) | ( ~n3666 & n6048 ) | ( n4682 & n6048 ) ;
  assign n8051 = n4024 & n8050 ;
  assign n8052 = n8051 ^ n6120 ^ 1'b0 ;
  assign n8053 = x114 & ~n2510 ;
  assign n8054 = n8053 ^ n4712 ^ n1418 ;
  assign n8060 = n4248 ^ n3691 ^ n2640 ;
  assign n8055 = n1033 | n7714 ;
  assign n8056 = ( ~n1695 & n7449 ) | ( ~n1695 & n8055 ) | ( n7449 & n8055 ) ;
  assign n8057 = n8056 ^ n2978 ^ x25 ;
  assign n8058 = n8057 ^ n5585 ^ n1859 ;
  assign n8059 = n8058 ^ n5418 ^ n3183 ;
  assign n8061 = n8060 ^ n8059 ^ 1'b0 ;
  assign n8062 = n8054 | n8061 ;
  assign n8063 = n1816 ^ n969 ^ 1'b0 ;
  assign n8064 = ~n1406 & n8063 ;
  assign n8065 = n3126 ^ n3115 ^ n1404 ;
  assign n8066 = n3486 ^ n2015 ^ n512 ;
  assign n8067 = ( n2940 & ~n3891 ) | ( n2940 & n7147 ) | ( ~n3891 & n7147 ) ;
  assign n8068 = ( ~n8065 & n8066 ) | ( ~n8065 & n8067 ) | ( n8066 & n8067 ) ;
  assign n8069 = ( n4445 & n8064 ) | ( n4445 & ~n8068 ) | ( n8064 & ~n8068 ) ;
  assign n8070 = n6864 ^ n5644 ^ n1191 ;
  assign n8071 = ( x30 & n3365 ) | ( x30 & n3464 ) | ( n3365 & n3464 ) ;
  assign n8072 = n8071 ^ n7553 ^ 1'b0 ;
  assign n8073 = ( n2054 & n8070 ) | ( n2054 & n8072 ) | ( n8070 & n8072 ) ;
  assign n8074 = n8073 ^ n991 ^ x79 ;
  assign n8075 = n8074 ^ n4717 ^ n2022 ;
  assign n8076 = ~n1373 & n2844 ;
  assign n8077 = ~n1153 & n6752 ;
  assign n8078 = n1088 & n8077 ;
  assign n8079 = n1919 | n2914 ;
  assign n8080 = ( n2860 & ~n8078 ) | ( n2860 & n8079 ) | ( ~n8078 & n8079 ) ;
  assign n8081 = n8080 ^ n7367 ^ n6021 ;
  assign n8082 = ( n2783 & n6465 ) | ( n2783 & n8081 ) | ( n6465 & n8081 ) ;
  assign n8083 = ( x33 & n664 ) | ( x33 & n1374 ) | ( n664 & n1374 ) ;
  assign n8084 = n7745 ^ n5330 ^ n687 ;
  assign n8089 = ~n2611 & n2860 ;
  assign n8090 = n8089 ^ n6609 ^ 1'b0 ;
  assign n8085 = ( ~n1238 & n1499 ) | ( ~n1238 & n2997 ) | ( n1499 & n2997 ) ;
  assign n8086 = n815 & n1981 ;
  assign n8087 = n8086 ^ n3031 ^ 1'b0 ;
  assign n8088 = ( n4509 & n8085 ) | ( n4509 & n8087 ) | ( n8085 & n8087 ) ;
  assign n8091 = n8090 ^ n8088 ^ 1'b0 ;
  assign n8092 = n1976 & n8091 ;
  assign n8093 = n8092 ^ n6951 ^ n4580 ;
  assign n8094 = ( n8083 & ~n8084 ) | ( n8083 & n8093 ) | ( ~n8084 & n8093 ) ;
  assign n8112 = n1430 ^ n1319 ^ n536 ;
  assign n8113 = n8112 ^ n4746 ^ n666 ;
  assign n8109 = n6727 ^ n4807 ^ n2058 ;
  assign n8110 = n1365 | n8109 ;
  assign n8111 = n8110 ^ n1098 ^ 1'b0 ;
  assign n8095 = ( n5145 & ~n5240 ) | ( n5145 & n5369 ) | ( ~n5240 & n5369 ) ;
  assign n8096 = n8095 ^ n6360 ^ n2244 ;
  assign n8104 = ( n699 & ~n2718 ) | ( n699 & n7211 ) | ( ~n2718 & n7211 ) ;
  assign n8101 = n4638 ^ n4295 ^ n3911 ;
  assign n8102 = ( ~n971 & n2689 ) | ( ~n971 & n5396 ) | ( n2689 & n5396 ) ;
  assign n8103 = ( n532 & n8101 ) | ( n532 & ~n8102 ) | ( n8101 & ~n8102 ) ;
  assign n8105 = n8104 ^ n8103 ^ n2601 ;
  assign n8106 = ( ~n2619 & n6473 ) | ( ~n2619 & n8105 ) | ( n6473 & n8105 ) ;
  assign n8097 = n5674 ^ n1159 ^ n702 ;
  assign n8098 = ( n3448 & n4746 ) | ( n3448 & n8097 ) | ( n4746 & n8097 ) ;
  assign n8099 = ( n403 & n1724 ) | ( n403 & n2865 ) | ( n1724 & n2865 ) ;
  assign n8100 = n8098 | n8099 ;
  assign n8107 = n8106 ^ n8100 ^ 1'b0 ;
  assign n8108 = ( n7825 & ~n8096 ) | ( n7825 & n8107 ) | ( ~n8096 & n8107 ) ;
  assign n8114 = n8113 ^ n8111 ^ n8108 ;
  assign n8116 = ( ~x96 & n286 ) | ( ~x96 & n2059 ) | ( n286 & n2059 ) ;
  assign n8117 = ( n1229 & n5662 ) | ( n1229 & n8116 ) | ( n5662 & n8116 ) ;
  assign n8118 = n8117 ^ n4748 ^ n2076 ;
  assign n8119 = n8118 ^ n5958 ^ n450 ;
  assign n8115 = n2499 ^ n1739 ^ n1289 ;
  assign n8120 = n8119 ^ n8115 ^ n6286 ;
  assign n8123 = n3347 ^ n2253 ^ x86 ;
  assign n8121 = n6079 ^ n5222 ^ n903 ;
  assign n8122 = ( n1076 & ~n6406 ) | ( n1076 & n8121 ) | ( ~n6406 & n8121 ) ;
  assign n8124 = n8123 ^ n8122 ^ n831 ;
  assign n8125 = n5204 ^ n4899 ^ 1'b0 ;
  assign n8126 = n8125 ^ n5587 ^ 1'b0 ;
  assign n8127 = n8126 ^ n6728 ^ n4002 ;
  assign n8128 = n8127 ^ n5966 ^ n858 ;
  assign n8129 = ( ~n2505 & n3272 ) | ( ~n2505 & n3907 ) | ( n3272 & n3907 ) ;
  assign n8130 = n8129 ^ n819 ^ n718 ;
  assign n8131 = n8130 ^ n1801 ^ n1310 ;
  assign n8132 = n8131 ^ n5280 ^ n1599 ;
  assign n8134 = ( n2920 & n3974 ) | ( n2920 & ~n4112 ) | ( n3974 & ~n4112 ) ;
  assign n8135 = ~n1761 & n3458 ;
  assign n8136 = ~n8134 & n8135 ;
  assign n8137 = n3473 & ~n8136 ;
  assign n8138 = n8137 ^ n2611 ^ 1'b0 ;
  assign n8133 = ( ~n703 & n2006 ) | ( ~n703 & n6301 ) | ( n2006 & n6301 ) ;
  assign n8139 = n8138 ^ n8133 ^ n3238 ;
  assign n8140 = ( n2368 & n2422 ) | ( n2368 & n2677 ) | ( n2422 & n2677 ) ;
  assign n8141 = ( n623 & n1283 ) | ( n623 & ~n6100 ) | ( n1283 & ~n6100 ) ;
  assign n8142 = n8141 ^ n7780 ^ n1671 ;
  assign n8143 = ( n2823 & ~n8140 ) | ( n2823 & n8142 ) | ( ~n8140 & n8142 ) ;
  assign n8144 = ( n1443 & ~n4427 ) | ( n1443 & n8143 ) | ( ~n4427 & n8143 ) ;
  assign n8145 = n8144 ^ n1291 ^ 1'b0 ;
  assign n8146 = ( n1115 & ~n1848 ) | ( n1115 & n3904 ) | ( ~n1848 & n3904 ) ;
  assign n8147 = ( ~n4034 & n4935 ) | ( ~n4034 & n8146 ) | ( n4935 & n8146 ) ;
  assign n8148 = ( n319 & ~n472 ) | ( n319 & n8147 ) | ( ~n472 & n8147 ) ;
  assign n8149 = ( n1940 & n2837 ) | ( n1940 & n4415 ) | ( n2837 & n4415 ) ;
  assign n8150 = ~n7573 & n7809 ;
  assign n8151 = ( n8044 & n8149 ) | ( n8044 & n8150 ) | ( n8149 & n8150 ) ;
  assign n8152 = n3116 ^ n1912 ^ n904 ;
  assign n8153 = ( ~n272 & n1086 ) | ( ~n272 & n8152 ) | ( n1086 & n8152 ) ;
  assign n8154 = n3078 ^ n3047 ^ 1'b0 ;
  assign n8155 = n8154 ^ n5256 ^ n782 ;
  assign n8156 = ( n3730 & n4487 ) | ( n3730 & n6908 ) | ( n4487 & n6908 ) ;
  assign n8157 = n5969 ^ n4259 ^ n2441 ;
  assign n8158 = ( n5984 & ~n8156 ) | ( n5984 & n8157 ) | ( ~n8156 & n8157 ) ;
  assign n8159 = n5993 ^ n1255 ^ x129 ;
  assign n8160 = ( n3717 & n4828 ) | ( n3717 & ~n8159 ) | ( n4828 & ~n8159 ) ;
  assign n8161 = n8160 ^ n5110 ^ n4277 ;
  assign n8162 = ( n4545 & n6601 ) | ( n4545 & ~n8161 ) | ( n6601 & ~n8161 ) ;
  assign n8163 = ( ~n6720 & n8158 ) | ( ~n6720 & n8162 ) | ( n8158 & n8162 ) ;
  assign n8164 = ( n8153 & n8155 ) | ( n8153 & ~n8163 ) | ( n8155 & ~n8163 ) ;
  assign n8165 = n7906 ^ n1459 ^ n296 ;
  assign n8166 = n8165 ^ n3850 ^ n1440 ;
  assign n8167 = n8166 ^ n3363 ^ n1537 ;
  assign n8168 = ( n6084 & ~n7748 ) | ( n6084 & n8167 ) | ( ~n7748 & n8167 ) ;
  assign n8169 = n8168 ^ n4991 ^ 1'b0 ;
  assign n8174 = ( n2505 & n3446 ) | ( n2505 & ~n6906 ) | ( n3446 & ~n6906 ) ;
  assign n8170 = n7147 ^ n2044 ^ n277 ;
  assign n8171 = ( x191 & n4480 ) | ( x191 & n8170 ) | ( n4480 & n8170 ) ;
  assign n8172 = ( n1469 & n3219 ) | ( n1469 & n8171 ) | ( n3219 & n8171 ) ;
  assign n8173 = ~n7014 & n8172 ;
  assign n8175 = n8174 ^ n8173 ^ 1'b0 ;
  assign n8176 = n4408 ^ n2975 ^ n294 ;
  assign n8181 = ~n601 & n4819 ;
  assign n8177 = n5705 ^ n4722 ^ 1'b0 ;
  assign n8178 = ~n1197 & n8177 ;
  assign n8179 = ( n3131 & n7392 ) | ( n3131 & n8178 ) | ( n7392 & n8178 ) ;
  assign n8180 = n8179 ^ n4609 ^ n1184 ;
  assign n8182 = n8181 ^ n8180 ^ n3764 ;
  assign n8194 = ( ~n679 & n1214 ) | ( ~n679 & n4863 ) | ( n1214 & n4863 ) ;
  assign n8195 = n5727 & n8194 ;
  assign n8187 = n446 | n2100 ;
  assign n8188 = n3218 | n8187 ;
  assign n8189 = n8188 ^ n5019 ^ x69 ;
  assign n8190 = n554 & n8189 ;
  assign n8191 = n8190 ^ n4156 ^ 1'b0 ;
  assign n8186 = ( n299 & ~n1266 ) | ( n299 & n2545 ) | ( ~n1266 & n2545 ) ;
  assign n8192 = n8191 ^ n8186 ^ 1'b0 ;
  assign n8193 = n6427 & n8192 ;
  assign n8196 = n8195 ^ n8193 ^ n6878 ;
  assign n8183 = ( n4261 & ~n6276 ) | ( n4261 & n8017 ) | ( ~n6276 & n8017 ) ;
  assign n8184 = n8183 ^ n2863 ^ n1059 ;
  assign n8185 = ( x170 & n4672 ) | ( x170 & n8184 ) | ( n4672 & n8184 ) ;
  assign n8197 = n8196 ^ n8185 ^ n632 ;
  assign n8199 = ( n387 & ~n1265 ) | ( n387 & n2728 ) | ( ~n1265 & n2728 ) ;
  assign n8198 = ( ~n324 & n471 ) | ( ~n324 & n5804 ) | ( n471 & n5804 ) ;
  assign n8200 = n8199 ^ n8198 ^ n7869 ;
  assign n8203 = n2217 ^ n706 ^ x26 ;
  assign n8204 = n6259 & ~n8203 ;
  assign n8205 = n3767 ^ n2222 ^ x94 ;
  assign n8206 = n8205 ^ n7045 ^ 1'b0 ;
  assign n8207 = n8204 & n8206 ;
  assign n8201 = ( ~n1865 & n2858 ) | ( ~n1865 & n7532 ) | ( n2858 & n7532 ) ;
  assign n8202 = n571 & n8201 ;
  assign n8208 = n8207 ^ n8202 ^ 1'b0 ;
  assign n8209 = n8208 ^ n6838 ^ n1425 ;
  assign n8210 = n8209 ^ n5894 ^ n2891 ;
  assign n8211 = ~n4420 & n8210 ;
  assign n8215 = ( x68 & n989 ) | ( x68 & ~n3080 ) | ( n989 & ~n3080 ) ;
  assign n8216 = n8215 ^ n4025 ^ n867 ;
  assign n8212 = ( n2597 & ~n3201 ) | ( n2597 & n5179 ) | ( ~n3201 & n5179 ) ;
  assign n8213 = n6034 ^ n688 ^ 1'b0 ;
  assign n8214 = n8212 & ~n8213 ;
  assign n8217 = n8216 ^ n8214 ^ n1659 ;
  assign n8218 = n7591 ^ n5899 ^ 1'b0 ;
  assign n8219 = n8217 | n8218 ;
  assign n8231 = ( ~n918 & n979 ) | ( ~n918 & n5247 ) | ( n979 & n5247 ) ;
  assign n8232 = ( n1634 & n7264 ) | ( n1634 & ~n8231 ) | ( n7264 & ~n8231 ) ;
  assign n8233 = n8232 ^ n7811 ^ n827 ;
  assign n8220 = n8188 ^ n6260 ^ n3727 ;
  assign n8225 = ( x46 & n747 ) | ( x46 & ~n3535 ) | ( n747 & ~n3535 ) ;
  assign n8221 = n2874 ^ n769 ^ n620 ;
  assign n8222 = n8221 ^ n4331 ^ n955 ;
  assign n8223 = ( ~n1199 & n3087 ) | ( ~n1199 & n5467 ) | ( n3087 & n5467 ) ;
  assign n8224 = n8222 | n8223 ;
  assign n8226 = n8225 ^ n8224 ^ 1'b0 ;
  assign n8227 = ~n944 & n8226 ;
  assign n8228 = ( n464 & n8220 ) | ( n464 & ~n8227 ) | ( n8220 & ~n8227 ) ;
  assign n8229 = ( ~n2718 & n7169 ) | ( ~n2718 & n8228 ) | ( n7169 & n8228 ) ;
  assign n8230 = ( n2292 & n3272 ) | ( n2292 & n8229 ) | ( n3272 & n8229 ) ;
  assign n8234 = n8233 ^ n8230 ^ n2430 ;
  assign n8235 = n8234 ^ n3115 ^ n2378 ;
  assign n8236 = ( n1717 & ~n3717 ) | ( n1717 & n4772 ) | ( ~n3717 & n4772 ) ;
  assign n8246 = n5521 ^ n5298 ^ n1956 ;
  assign n8247 = n8246 ^ n3650 ^ 1'b0 ;
  assign n8248 = n5558 | n8247 ;
  assign n8249 = n8248 ^ n6827 ^ n1470 ;
  assign n8237 = ( ~n515 & n3232 ) | ( ~n515 & n3317 ) | ( n3232 & n3317 ) ;
  assign n8238 = n8237 ^ n1899 ^ n624 ;
  assign n8239 = ( n1410 & n2677 ) | ( n1410 & ~n2833 ) | ( n2677 & ~n2833 ) ;
  assign n8240 = ( n2585 & n3283 ) | ( n2585 & ~n8239 ) | ( n3283 & ~n8239 ) ;
  assign n8241 = ( n691 & ~n1781 ) | ( n691 & n6171 ) | ( ~n1781 & n6171 ) ;
  assign n8242 = n8240 & n8241 ;
  assign n8243 = ~n607 & n8242 ;
  assign n8244 = n8238 & ~n8243 ;
  assign n8245 = n4567 & n8244 ;
  assign n8250 = n8249 ^ n8245 ^ 1'b0 ;
  assign n8251 = ( n8157 & n8236 ) | ( n8157 & ~n8250 ) | ( n8236 & ~n8250 ) ;
  assign n8252 = x201 & ~n876 ;
  assign n8253 = n8252 ^ n2064 ^ 1'b0 ;
  assign n8254 = n8253 ^ n1404 ^ 1'b0 ;
  assign n8255 = ( n4654 & ~n7094 ) | ( n4654 & n8254 ) | ( ~n7094 & n8254 ) ;
  assign n8259 = n760 ^ x175 ^ 1'b0 ;
  assign n8260 = ( n6399 & ~n7494 ) | ( n6399 & n8259 ) | ( ~n7494 & n8259 ) ;
  assign n8257 = n2979 ^ n2424 ^ 1'b0 ;
  assign n8256 = ( ~x66 & n602 ) | ( ~x66 & n783 ) | ( n602 & n783 ) ;
  assign n8258 = n8257 ^ n8256 ^ n6963 ;
  assign n8261 = n8260 ^ n8258 ^ 1'b0 ;
  assign n8262 = ( n5969 & ~n8255 ) | ( n5969 & n8261 ) | ( ~n8255 & n8261 ) ;
  assign n8263 = ( n2124 & n3675 ) | ( n2124 & ~n8125 ) | ( n3675 & ~n8125 ) ;
  assign n8264 = n8053 ^ n5444 ^ 1'b0 ;
  assign n8265 = n6766 | n8264 ;
  assign n8271 = ( n840 & n2984 ) | ( n840 & n6467 ) | ( n2984 & n6467 ) ;
  assign n8272 = n1503 & n8271 ;
  assign n8273 = ( x100 & n6852 ) | ( x100 & n8272 ) | ( n6852 & n8272 ) ;
  assign n8274 = ( n937 & ~n3011 ) | ( n937 & n8273 ) | ( ~n3011 & n8273 ) ;
  assign n8266 = ~n2521 & n4670 ;
  assign n8267 = n831 & n8266 ;
  assign n8268 = n6318 ^ n2046 ^ x50 ;
  assign n8269 = ( x36 & n968 ) | ( x36 & ~n8268 ) | ( n968 & ~n8268 ) ;
  assign n8270 = ( n3796 & n8267 ) | ( n3796 & n8269 ) | ( n8267 & n8269 ) ;
  assign n8275 = n8274 ^ n8270 ^ 1'b0 ;
  assign n8276 = ~n8265 & n8275 ;
  assign n8282 = n487 & n2471 ;
  assign n8283 = ~n865 & n8282 ;
  assign n8284 = n914 | n4354 ;
  assign n8285 = ( n6433 & n8283 ) | ( n6433 & n8284 ) | ( n8283 & n8284 ) ;
  assign n8286 = n8285 ^ n6933 ^ n6038 ;
  assign n8277 = n2754 ^ n744 ^ n556 ;
  assign n8278 = n8277 ^ n4940 ^ 1'b0 ;
  assign n8279 = n5518 & ~n8278 ;
  assign n8280 = ~n6487 & n8279 ;
  assign n8281 = n5751 & n8280 ;
  assign n8287 = n8286 ^ n8281 ^ n1399 ;
  assign n8288 = ( ~n1370 & n1853 ) | ( ~n1370 & n4886 ) | ( n1853 & n4886 ) ;
  assign n8289 = n2880 ^ n1529 ^ n1297 ;
  assign n8290 = ( x64 & n1327 ) | ( x64 & n8289 ) | ( n1327 & n8289 ) ;
  assign n8291 = n8290 ^ n5131 ^ 1'b0 ;
  assign n8292 = ( n1579 & n2305 ) | ( n1579 & n8291 ) | ( n2305 & n8291 ) ;
  assign n8293 = n4701 ^ n567 ^ n368 ;
  assign n8294 = ( n665 & n3864 ) | ( n665 & ~n8293 ) | ( n3864 & ~n8293 ) ;
  assign n8295 = n3247 & n8294 ;
  assign n8296 = ~n8292 & n8295 ;
  assign n8297 = n3731 ^ n1408 ^ n607 ;
  assign n8298 = n8297 ^ n7312 ^ n2564 ;
  assign n8299 = ( n6240 & n8296 ) | ( n6240 & ~n8298 ) | ( n8296 & ~n8298 ) ;
  assign n8300 = ( n2598 & n5558 ) | ( n2598 & ~n8299 ) | ( n5558 & ~n8299 ) ;
  assign n8301 = ( n2381 & n2664 ) | ( n2381 & n5900 ) | ( n2664 & n5900 ) ;
  assign n8302 = ( n1090 & n1119 ) | ( n1090 & ~n6902 ) | ( n1119 & ~n6902 ) ;
  assign n8303 = ( ~n527 & n1781 ) | ( ~n527 & n8302 ) | ( n1781 & n8302 ) ;
  assign n8304 = n8303 ^ n2204 ^ 1'b0 ;
  assign n8305 = ~n8301 & n8304 ;
  assign n8306 = ( n7744 & n8300 ) | ( n7744 & n8305 ) | ( n8300 & n8305 ) ;
  assign n8307 = n7603 ^ n6205 ^ n791 ;
  assign n8308 = ( n435 & n7602 ) | ( n435 & ~n8307 ) | ( n7602 & ~n8307 ) ;
  assign n8309 = n8308 ^ n8013 ^ x163 ;
  assign n8310 = ( n817 & ~n2874 ) | ( n817 & n8309 ) | ( ~n2874 & n8309 ) ;
  assign n8311 = ( n2065 & n2858 ) | ( n2065 & ~n5543 ) | ( n2858 & ~n5543 ) ;
  assign n8312 = ( n1858 & n2775 ) | ( n1858 & n8311 ) | ( n2775 & n8311 ) ;
  assign n8313 = ( n261 & n4580 ) | ( n261 & ~n8312 ) | ( n4580 & ~n8312 ) ;
  assign n8314 = ( ~n581 & n1118 ) | ( ~n581 & n6156 ) | ( n1118 & n6156 ) ;
  assign n8315 = ( n315 & ~n5558 ) | ( n315 & n8314 ) | ( ~n5558 & n8314 ) ;
  assign n8316 = n8313 | n8315 ;
  assign n8317 = n261 | n8316 ;
  assign n8318 = n8255 ^ n2948 ^ n953 ;
  assign n8319 = ( ~n1399 & n1905 ) | ( ~n1399 & n3635 ) | ( n1905 & n3635 ) ;
  assign n8320 = n7886 ^ n970 ^ 1'b0 ;
  assign n8321 = ( n765 & ~n1219 ) | ( n765 & n8320 ) | ( ~n1219 & n8320 ) ;
  assign n8322 = n8321 ^ n3400 ^ 1'b0 ;
  assign n8323 = x126 & ~n8322 ;
  assign n8324 = ( x81 & n3618 ) | ( x81 & n8323 ) | ( n3618 & n8323 ) ;
  assign n8325 = ( n402 & ~n1636 ) | ( n402 & n3192 ) | ( ~n1636 & n3192 ) ;
  assign n8326 = ( n8319 & ~n8324 ) | ( n8319 & n8325 ) | ( ~n8324 & n8325 ) ;
  assign n8332 = n3004 ^ n1417 ^ 1'b0 ;
  assign n8333 = n1719 | n8332 ;
  assign n8327 = n478 ^ n276 ^ 1'b0 ;
  assign n8328 = n2238 ^ n793 ^ 1'b0 ;
  assign n8329 = n8327 & n8328 ;
  assign n8330 = n8329 ^ n3666 ^ n479 ;
  assign n8331 = ( n6233 & n6481 ) | ( n6233 & n8330 ) | ( n6481 & n8330 ) ;
  assign n8334 = n8333 ^ n8331 ^ n4433 ;
  assign n8335 = n7120 ^ n2229 ^ 1'b0 ;
  assign n8336 = ( n4219 & n5346 ) | ( n4219 & n6827 ) | ( n5346 & n6827 ) ;
  assign n8338 = ( n437 & n6864 ) | ( n437 & n8329 ) | ( n6864 & n8329 ) ;
  assign n8337 = n1741 ^ n1729 ^ n588 ;
  assign n8339 = n8338 ^ n8337 ^ 1'b0 ;
  assign n8340 = ~n5048 & n8339 ;
  assign n8341 = ( n7797 & n8336 ) | ( n7797 & n8340 ) | ( n8336 & n8340 ) ;
  assign n8342 = n8341 ^ n5705 ^ n3370 ;
  assign n8343 = ( ~n2945 & n8335 ) | ( ~n2945 & n8342 ) | ( n8335 & n8342 ) ;
  assign n8344 = ( n1552 & ~n1863 ) | ( n1552 & n2102 ) | ( ~n1863 & n2102 ) ;
  assign n8345 = ( x97 & n2452 ) | ( x97 & n3803 ) | ( n2452 & n3803 ) ;
  assign n8346 = n8345 ^ n1529 ^ n511 ;
  assign n8347 = ( n1351 & ~n5714 ) | ( n1351 & n8346 ) | ( ~n5714 & n8346 ) ;
  assign n8358 = n6921 ^ n2718 ^ n651 ;
  assign n8354 = ( ~n947 & n2952 ) | ( ~n947 & n6356 ) | ( n2952 & n6356 ) ;
  assign n8352 = n4047 & ~n8223 ;
  assign n8353 = ~n615 & n8352 ;
  assign n8355 = n8354 ^ n8353 ^ n7786 ;
  assign n8356 = ( x34 & ~n918 ) | ( x34 & n2356 ) | ( ~n918 & n2356 ) ;
  assign n8357 = ( n880 & ~n8355 ) | ( n880 & n8356 ) | ( ~n8355 & n8356 ) ;
  assign n8349 = ( n2320 & ~n2637 ) | ( n2320 & n5134 ) | ( ~n2637 & n5134 ) ;
  assign n8350 = n8349 ^ n4104 ^ n681 ;
  assign n8348 = ( x74 & x79 ) | ( x74 & n4094 ) | ( x79 & n4094 ) ;
  assign n8351 = n8350 ^ n8348 ^ n7702 ;
  assign n8359 = n8358 ^ n8357 ^ n8351 ;
  assign n8360 = ( n8344 & n8347 ) | ( n8344 & n8359 ) | ( n8347 & n8359 ) ;
  assign n8361 = ( n1114 & ~n1733 ) | ( n1114 & n2234 ) | ( ~n1733 & n2234 ) ;
  assign n8362 = n2744 & n8246 ;
  assign n8363 = n6496 & n8362 ;
  assign n8364 = n1082 ^ n937 ^ 1'b0 ;
  assign n8365 = ( ~n1041 & n8363 ) | ( ~n1041 & n8364 ) | ( n8363 & n8364 ) ;
  assign n8366 = ( ~n1358 & n8361 ) | ( ~n1358 & n8365 ) | ( n8361 & n8365 ) ;
  assign n8367 = ( n404 & n2644 ) | ( n404 & n8366 ) | ( n2644 & n8366 ) ;
  assign n8368 = n6538 & n7425 ;
  assign n8369 = n5044 ^ n2243 ^ n769 ;
  assign n8370 = n8369 ^ n3339 ^ n2254 ;
  assign n8371 = n8370 ^ n3688 ^ n3628 ;
  assign n8372 = x90 & n2011 ;
  assign n8373 = n1976 & ~n8372 ;
  assign n8374 = n4944 & n8373 ;
  assign n8378 = ( n668 & n2222 ) | ( n668 & n3328 ) | ( n2222 & n3328 ) ;
  assign n8379 = n8378 ^ n2591 ^ n2118 ;
  assign n8380 = n8379 ^ n6884 ^ n2113 ;
  assign n8375 = n922 | n3628 ;
  assign n8376 = n2856 | n8375 ;
  assign n8377 = ( n2157 & n4727 ) | ( n2157 & ~n8376 ) | ( n4727 & ~n8376 ) ;
  assign n8381 = n8380 ^ n8377 ^ 1'b0 ;
  assign n8382 = ( n1245 & ~n8374 ) | ( n1245 & n8381 ) | ( ~n8374 & n8381 ) ;
  assign n8383 = n1030 & n1823 ;
  assign n8384 = n8383 ^ n6106 ^ n2060 ;
  assign n8385 = ( n1608 & n4112 ) | ( n1608 & ~n7396 ) | ( n4112 & ~n7396 ) ;
  assign n8386 = ( n2152 & ~n3492 ) | ( n2152 & n4085 ) | ( ~n3492 & n4085 ) ;
  assign n8387 = n8386 ^ n2413 ^ n2073 ;
  assign n8388 = ( n2443 & ~n8385 ) | ( n2443 & n8387 ) | ( ~n8385 & n8387 ) ;
  assign n8402 = ( n698 & n4862 ) | ( n698 & n5985 ) | ( n4862 & n5985 ) ;
  assign n8400 = n5239 ^ n2515 ^ 1'b0 ;
  assign n8401 = n8400 ^ n6838 ^ n3230 ;
  assign n8395 = n7159 ^ x1 ^ 1'b0 ;
  assign n8396 = n3944 & ~n8395 ;
  assign n8397 = n6923 & n8396 ;
  assign n8398 = n8397 ^ n940 ^ 1'b0 ;
  assign n8392 = n8116 ^ n5264 ^ n3061 ;
  assign n8393 = n8392 ^ n1390 ^ n1137 ;
  assign n8389 = n5326 & n6680 ;
  assign n8390 = ~n2892 & n8389 ;
  assign n8391 = n7786 | n8390 ;
  assign n8394 = n8393 ^ n8391 ^ 1'b0 ;
  assign n8399 = n8398 ^ n8394 ^ n2031 ;
  assign n8403 = n8402 ^ n8401 ^ n8399 ;
  assign n8404 = n4706 ^ n2399 ^ n1352 ;
  assign n8405 = ( ~n3811 & n6799 ) | ( ~n3811 & n8404 ) | ( n6799 & n8404 ) ;
  assign n8406 = n1513 ^ n1458 ^ n650 ;
  assign n8407 = ( n1096 & n3739 ) | ( n1096 & n8406 ) | ( n3739 & n8406 ) ;
  assign n8408 = ( x199 & n1264 ) | ( x199 & ~n8407 ) | ( n1264 & ~n8407 ) ;
  assign n8409 = ( n486 & ~n3866 ) | ( n486 & n8408 ) | ( ~n3866 & n8408 ) ;
  assign n8410 = ( n4826 & ~n8405 ) | ( n4826 & n8409 ) | ( ~n8405 & n8409 ) ;
  assign n8411 = n4093 ^ n3404 ^ 1'b0 ;
  assign n8412 = n6865 ^ n4371 ^ n2595 ;
  assign n8413 = ~n7308 & n8412 ;
  assign n8414 = n2033 ^ n1601 ^ n1184 ;
  assign n8415 = n8414 ^ n4476 ^ n1748 ;
  assign n8416 = n7368 | n8415 ;
  assign n8417 = n8416 ^ n3959 ^ 1'b0 ;
  assign n8418 = n8417 ^ n6859 ^ n1402 ;
  assign n8419 = ~n1147 & n8418 ;
  assign n8420 = n8413 & n8419 ;
  assign n8421 = ( n3078 & n6381 ) | ( n3078 & ~n6659 ) | ( n6381 & ~n6659 ) ;
  assign n8422 = ( n1459 & ~n1539 ) | ( n1459 & n8421 ) | ( ~n1539 & n8421 ) ;
  assign n8423 = n8422 ^ n4697 ^ n3008 ;
  assign n8424 = ( n1889 & n4293 ) | ( n1889 & n6581 ) | ( n4293 & n6581 ) ;
  assign n8429 = ( n1280 & n1557 ) | ( n1280 & ~n1762 ) | ( n1557 & ~n1762 ) ;
  assign n8430 = n8429 ^ n4350 ^ n2309 ;
  assign n8431 = ( n1262 & n5414 ) | ( n1262 & ~n8430 ) | ( n5414 & ~n8430 ) ;
  assign n8425 = ( n5369 & ~n5512 ) | ( n5369 & n7988 ) | ( ~n5512 & n7988 ) ;
  assign n8426 = ( ~n3760 & n7588 ) | ( ~n3760 & n8425 ) | ( n7588 & n8425 ) ;
  assign n8427 = n8426 ^ n7428 ^ 1'b0 ;
  assign n8428 = ~n360 & n8427 ;
  assign n8432 = n8431 ^ n8428 ^ n3237 ;
  assign n8433 = n8432 ^ n5835 ^ n5416 ;
  assign n8434 = n6827 ^ n2252 ^ 1'b0 ;
  assign n8435 = n8434 ^ n868 ^ 1'b0 ;
  assign n8436 = ( n8424 & n8433 ) | ( n8424 & ~n8435 ) | ( n8433 & ~n8435 ) ;
  assign n8437 = ( n559 & ~n4646 ) | ( n559 & n5693 ) | ( ~n4646 & n5693 ) ;
  assign n8438 = n1141 | n8437 ;
  assign n8439 = n8438 ^ n7698 ^ n4527 ;
  assign n8440 = n6675 ^ n1304 ^ x232 ;
  assign n8441 = ( n4977 & ~n7484 ) | ( n4977 & n8440 ) | ( ~n7484 & n8440 ) ;
  assign n8442 = n5030 ^ n1524 ^ 1'b0 ;
  assign n8443 = ( n6436 & ~n8441 ) | ( n6436 & n8442 ) | ( ~n8441 & n8442 ) ;
  assign n8447 = ( n1809 & ~n5475 ) | ( n1809 & n6589 ) | ( ~n5475 & n6589 ) ;
  assign n8448 = n8447 ^ n4916 ^ 1'b0 ;
  assign n8449 = x41 & n6825 ;
  assign n8450 = n8449 ^ n1191 ^ 1'b0 ;
  assign n8451 = n8450 ^ n4473 ^ n2586 ;
  assign n8452 = ( n5790 & ~n8448 ) | ( n5790 & n8451 ) | ( ~n8448 & n8451 ) ;
  assign n8444 = ( ~n880 & n3339 ) | ( ~n880 & n4978 ) | ( n3339 & n4978 ) ;
  assign n8445 = n8444 ^ n7998 ^ 1'b0 ;
  assign n8446 = n3898 & n8445 ;
  assign n8453 = n8452 ^ n8446 ^ n7343 ;
  assign n8454 = ( n5226 & ~n7153 ) | ( n5226 & n8414 ) | ( ~n7153 & n8414 ) ;
  assign n8455 = n3382 & n4597 ;
  assign n8456 = n8455 ^ n561 ^ 1'b0 ;
  assign n8457 = ( n1235 & ~n5122 ) | ( n1235 & n8456 ) | ( ~n5122 & n8456 ) ;
  assign n8458 = n2912 & ~n8457 ;
  assign n8459 = n8454 | n8458 ;
  assign n8460 = n1448 | n8459 ;
  assign n8461 = ( n6722 & n8453 ) | ( n6722 & ~n8460 ) | ( n8453 & ~n8460 ) ;
  assign n8468 = n6689 ^ n2576 ^ n813 ;
  assign n8469 = n8468 ^ n4156 ^ n2997 ;
  assign n8467 = n7124 ^ n4036 ^ n3414 ;
  assign n8464 = n2107 ^ n1872 ^ x120 ;
  assign n8463 = ( ~n975 & n5662 ) | ( ~n975 & n7487 ) | ( n5662 & n7487 ) ;
  assign n8465 = n8464 ^ n8463 ^ n8183 ;
  assign n8462 = n1601 & n7278 ;
  assign n8466 = n8465 ^ n8462 ^ 1'b0 ;
  assign n8470 = n8469 ^ n8467 ^ n8466 ;
  assign n8471 = ( n1136 & ~n8361 ) | ( n1136 & n8470 ) | ( ~n8361 & n8470 ) ;
  assign n8473 = n2618 ^ n2611 ^ n1505 ;
  assign n8474 = ( n561 & n1640 ) | ( n561 & n8473 ) | ( n1640 & n8473 ) ;
  assign n8472 = n3228 ^ n2445 ^ n2244 ;
  assign n8475 = n8474 ^ n8472 ^ n3534 ;
  assign n8476 = n8475 ^ n5685 ^ n1114 ;
  assign n8477 = n8476 ^ n8188 ^ n488 ;
  assign n8478 = ( ~n1858 & n6286 ) | ( ~n1858 & n7019 ) | ( n6286 & n7019 ) ;
  assign n8479 = ( n333 & n464 ) | ( n333 & ~n2156 ) | ( n464 & ~n2156 ) ;
  assign n8480 = n8479 ^ n7328 ^ n1135 ;
  assign n8481 = n8480 ^ n1256 ^ 1'b0 ;
  assign n8482 = ~n371 & n8481 ;
  assign n8483 = ( ~n5702 & n8478 ) | ( ~n5702 & n8482 ) | ( n8478 & n8482 ) ;
  assign n8484 = ( n4144 & ~n5474 ) | ( n4144 & n5727 ) | ( ~n5474 & n5727 ) ;
  assign n8485 = n8040 ^ n6679 ^ n2022 ;
  assign n8486 = ( n4557 & n8484 ) | ( n4557 & n8485 ) | ( n8484 & n8485 ) ;
  assign n8487 = ( ~x100 & x252 ) | ( ~x100 & n4879 ) | ( x252 & n4879 ) ;
  assign n8488 = n8487 ^ n3544 ^ n1834 ;
  assign n8489 = n8488 ^ n4814 ^ n2675 ;
  assign n8490 = ( n374 & ~n3476 ) | ( n374 & n8489 ) | ( ~n3476 & n8489 ) ;
  assign n8491 = n8490 ^ n8052 ^ n6596 ;
  assign n8492 = ~n2439 & n5298 ;
  assign n8493 = n8492 ^ n7547 ^ 1'b0 ;
  assign n8494 = ( n345 & ~n1950 ) | ( n345 & n2792 ) | ( ~n1950 & n2792 ) ;
  assign n8495 = ( n1129 & n4105 ) | ( n1129 & ~n6743 ) | ( n4105 & ~n6743 ) ;
  assign n8496 = ( n1432 & n2417 ) | ( n1432 & n2591 ) | ( n2417 & n2591 ) ;
  assign n8497 = n2475 ^ n2080 ^ 1'b0 ;
  assign n8498 = n1688 & ~n8497 ;
  assign n8499 = ( ~x70 & n345 ) | ( ~x70 & n3992 ) | ( n345 & n3992 ) ;
  assign n8500 = n8499 ^ n8225 ^ n6260 ;
  assign n8501 = ( n1770 & n4792 ) | ( n1770 & ~n8500 ) | ( n4792 & ~n8500 ) ;
  assign n8502 = ( n8496 & n8498 ) | ( n8496 & ~n8501 ) | ( n8498 & ~n8501 ) ;
  assign n8503 = n5377 ^ n3225 ^ 1'b0 ;
  assign n8504 = n8502 | n8503 ;
  assign n8505 = ( ~n6334 & n6348 ) | ( ~n6334 & n7685 ) | ( n6348 & n7685 ) ;
  assign n8506 = ( n4301 & n8504 ) | ( n4301 & n8505 ) | ( n8504 & n8505 ) ;
  assign n8507 = ( n8494 & n8495 ) | ( n8494 & ~n8506 ) | ( n8495 & ~n8506 ) ;
  assign n8508 = ( n655 & ~n2521 ) | ( n655 & n5366 ) | ( ~n2521 & n5366 ) ;
  assign n8509 = ( n2401 & n2579 ) | ( n2401 & n2842 ) | ( n2579 & n2842 ) ;
  assign n8510 = n8509 ^ n3604 ^ n3081 ;
  assign n8511 = ( ~n2286 & n8508 ) | ( ~n2286 & n8510 ) | ( n8508 & n8510 ) ;
  assign n8512 = ( ~n674 & n1210 ) | ( ~n674 & n4133 ) | ( n1210 & n4133 ) ;
  assign n8513 = n8512 ^ n5726 ^ n1830 ;
  assign n8515 = n7176 ^ n2607 ^ n1171 ;
  assign n8514 = ( n488 & ~n4411 ) | ( n488 & n7684 ) | ( ~n4411 & n7684 ) ;
  assign n8516 = n8515 ^ n8514 ^ n5150 ;
  assign n8517 = n6044 ^ n2210 ^ x147 ;
  assign n8518 = n6804 ^ n6610 ^ n2935 ;
  assign n8519 = n8518 ^ n7590 ^ 1'b0 ;
  assign n8520 = ~n1487 & n8519 ;
  assign n8527 = ~n1215 & n2495 ;
  assign n8521 = n7551 ^ n7444 ^ n5874 ;
  assign n8522 = n6939 ^ n6493 ^ n5222 ;
  assign n8523 = ( n954 & n1195 ) | ( n954 & ~n1634 ) | ( n1195 & ~n1634 ) ;
  assign n8524 = n8523 ^ n4999 ^ n2310 ;
  assign n8525 = n8524 ^ n3533 ^ 1'b0 ;
  assign n8526 = ( n8521 & ~n8522 ) | ( n8521 & n8525 ) | ( ~n8522 & n8525 ) ;
  assign n8528 = n8527 ^ n8526 ^ n3245 ;
  assign n8529 = n3756 ^ n1233 ^ 1'b0 ;
  assign n8530 = n3584 & ~n8529 ;
  assign n8531 = n8530 ^ n7293 ^ n578 ;
  assign n8532 = n8531 ^ n5741 ^ 1'b0 ;
  assign n8533 = n4140 & ~n8532 ;
  assign n8534 = n3184 ^ n2720 ^ n2689 ;
  assign n8535 = n7176 ^ n3345 ^ n1819 ;
  assign n8536 = ( ~n1569 & n8534 ) | ( ~n1569 & n8535 ) | ( n8534 & n8535 ) ;
  assign n8537 = n2834 ^ n1889 ^ n970 ;
  assign n8538 = n1787 | n8265 ;
  assign n8539 = ( n8536 & ~n8537 ) | ( n8536 & n8538 ) | ( ~n8537 & n8538 ) ;
  assign n8540 = ( n2524 & n8533 ) | ( n2524 & ~n8539 ) | ( n8533 & ~n8539 ) ;
  assign n8545 = ~n7046 & n7163 ;
  assign n8546 = n8545 ^ n3713 ^ 1'b0 ;
  assign n8547 = n6087 ^ n5634 ^ n2249 ;
  assign n8548 = ( ~n3413 & n3723 ) | ( ~n3413 & n8547 ) | ( n3723 & n8547 ) ;
  assign n8549 = ( x202 & n8546 ) | ( x202 & n8548 ) | ( n8546 & n8548 ) ;
  assign n8543 = ( ~n3972 & n5522 ) | ( ~n3972 & n7279 ) | ( n5522 & n7279 ) ;
  assign n8544 = ( ~n1214 & n6042 ) | ( ~n1214 & n8543 ) | ( n6042 & n8543 ) ;
  assign n8541 = n8426 ^ n5987 ^ 1'b0 ;
  assign n8542 = ( n2840 & ~n7293 ) | ( n2840 & n8541 ) | ( ~n7293 & n8541 ) ;
  assign n8550 = n8549 ^ n8544 ^ n8542 ;
  assign n8567 = ( n1958 & n4504 ) | ( n1958 & ~n5164 ) | ( n4504 & ~n5164 ) ;
  assign n8558 = ( x70 & n752 ) | ( x70 & n6203 ) | ( n752 & n6203 ) ;
  assign n8559 = ~n3571 & n8558 ;
  assign n8560 = n6543 & n8559 ;
  assign n8561 = ( n1096 & ~n1501 ) | ( n1096 & n2644 ) | ( ~n1501 & n2644 ) ;
  assign n8562 = n2061 & n8561 ;
  assign n8563 = ~n2711 & n8562 ;
  assign n8564 = n8563 ^ n5584 ^ n3576 ;
  assign n8565 = ( n1364 & n8560 ) | ( n1364 & n8564 ) | ( n8560 & n8564 ) ;
  assign n8566 = ( n931 & ~n4565 ) | ( n931 & n8565 ) | ( ~n4565 & n8565 ) ;
  assign n8555 = n8055 ^ n1887 ^ n502 ;
  assign n8556 = n6034 & ~n8555 ;
  assign n8551 = n1745 | n4890 ;
  assign n8552 = n8551 ^ n2966 ^ 1'b0 ;
  assign n8553 = ( n2998 & ~n3413 ) | ( n2998 & n8552 ) | ( ~n3413 & n8552 ) ;
  assign n8554 = ( ~n4441 & n4653 ) | ( ~n4441 & n8553 ) | ( n4653 & n8553 ) ;
  assign n8557 = n8556 ^ n8554 ^ n710 ;
  assign n8568 = n8567 ^ n8566 ^ n8557 ;
  assign n8569 = n8568 ^ n5146 ^ n3205 ;
  assign n8570 = n6690 & n8569 ;
  assign n8575 = ~n534 & n3504 ;
  assign n8576 = n8575 ^ n3819 ^ 1'b0 ;
  assign n8577 = ( n1673 & ~n4333 ) | ( n1673 & n8576 ) | ( ~n4333 & n8576 ) ;
  assign n8571 = n1630 ^ x223 ^ 1'b0 ;
  assign n8572 = ~n2952 & n8571 ;
  assign n8573 = n8572 ^ n1655 ^ 1'b0 ;
  assign n8574 = ( n2115 & n2837 ) | ( n2115 & ~n8573 ) | ( n2837 & ~n8573 ) ;
  assign n8578 = n8577 ^ n8574 ^ n1979 ;
  assign n8579 = n5098 & n8578 ;
  assign n8580 = n8579 ^ n3998 ^ n3212 ;
  assign n8581 = n3680 ^ n3333 ^ 1'b0 ;
  assign n8582 = ~n3867 & n8581 ;
  assign n8583 = n8582 ^ n4396 ^ x155 ;
  assign n8588 = ( n4549 & ~n5931 ) | ( n4549 & n7625 ) | ( ~n5931 & n7625 ) ;
  assign n8585 = n2543 ^ n2212 ^ x127 ;
  assign n8586 = n8585 ^ n4410 ^ x59 ;
  assign n8587 = ( ~n1296 & n3686 ) | ( ~n1296 & n8586 ) | ( n3686 & n8586 ) ;
  assign n8589 = n8588 ^ n8587 ^ 1'b0 ;
  assign n8584 = n8097 ^ n3838 ^ n3319 ;
  assign n8590 = n8589 ^ n8584 ^ n7042 ;
  assign n8591 = n3995 ^ n3625 ^ n1277 ;
  assign n8592 = ( n916 & n1829 ) | ( n916 & n3013 ) | ( n1829 & n3013 ) ;
  assign n8593 = n8592 ^ n2941 ^ n793 ;
  assign n8594 = ( ~n6672 & n7653 ) | ( ~n6672 & n8593 ) | ( n7653 & n8593 ) ;
  assign n8595 = n8594 ^ n3194 ^ n359 ;
  assign n8603 = n7457 ^ n6312 ^ n3127 ;
  assign n8596 = n7054 ^ n691 ^ n579 ;
  assign n8597 = n8596 ^ n1971 ^ 1'b0 ;
  assign n8600 = n3073 ^ n1472 ^ n1135 ;
  assign n8598 = ( ~n527 & n1502 ) | ( ~n527 & n6699 ) | ( n1502 & n6699 ) ;
  assign n8599 = n2651 | n8598 ;
  assign n8601 = n8600 ^ n8599 ^ 1'b0 ;
  assign n8602 = n8597 & n8601 ;
  assign n8604 = n8603 ^ n8602 ^ 1'b0 ;
  assign n8605 = n1762 ^ n1557 ^ n508 ;
  assign n8606 = x120 & ~n2178 ;
  assign n8607 = n8605 & n8606 ;
  assign n8608 = ( n6430 & ~n8604 ) | ( n6430 & n8607 ) | ( ~n8604 & n8607 ) ;
  assign n8609 = ( n5527 & ~n8595 ) | ( n5527 & n8608 ) | ( ~n8595 & n8608 ) ;
  assign n8610 = n8609 ^ n2658 ^ 1'b0 ;
  assign n8611 = n4211 ^ n1413 ^ n671 ;
  assign n8612 = ( n1439 & n7242 ) | ( n1439 & ~n8611 ) | ( n7242 & ~n8611 ) ;
  assign n8613 = ( n612 & n2358 ) | ( n612 & n3537 ) | ( n2358 & n3537 ) ;
  assign n8614 = n5221 ^ n1980 ^ n784 ;
  assign n8615 = n8614 ^ n8117 ^ n1526 ;
  assign n8616 = n3407 ^ n1350 ^ 1'b0 ;
  assign n8617 = ( n4846 & n8501 ) | ( n4846 & n8616 ) | ( n8501 & n8616 ) ;
  assign n8618 = ( n2034 & n4010 ) | ( n2034 & n6782 ) | ( n4010 & n6782 ) ;
  assign n8619 = n1558 ^ x32 ^ 1'b0 ;
  assign n8620 = ( n5914 & ~n8618 ) | ( n5914 & n8619 ) | ( ~n8618 & n8619 ) ;
  assign n8621 = ( n3212 & n4926 ) | ( n3212 & n8620 ) | ( n4926 & n8620 ) ;
  assign n8622 = n8621 ^ n6479 ^ x16 ;
  assign n8623 = ( ~n8615 & n8617 ) | ( ~n8615 & n8622 ) | ( n8617 & n8622 ) ;
  assign n8624 = ( n8040 & ~n8613 ) | ( n8040 & n8623 ) | ( ~n8613 & n8623 ) ;
  assign n8625 = n4581 ^ n3588 ^ n2127 ;
  assign n8626 = ( n2246 & ~n4134 ) | ( n2246 & n8625 ) | ( ~n4134 & n8625 ) ;
  assign n8637 = ( n554 & n2097 ) | ( n554 & n6215 ) | ( n2097 & n6215 ) ;
  assign n8627 = ( n2842 & ~n3942 ) | ( n2842 & n4309 ) | ( ~n3942 & n4309 ) ;
  assign n8628 = n8627 ^ n5206 ^ n2608 ;
  assign n8629 = ( ~n1266 & n1341 ) | ( ~n1266 & n6287 ) | ( n1341 & n6287 ) ;
  assign n8630 = n8629 ^ n3286 ^ 1'b0 ;
  assign n8631 = ~n4885 & n8630 ;
  assign n8632 = n8631 ^ x133 ^ 1'b0 ;
  assign n8633 = n8632 ^ n4703 ^ n3458 ;
  assign n8634 = n8633 ^ n5328 ^ n2651 ;
  assign n8635 = n8634 ^ n2203 ^ n1963 ;
  assign n8636 = ( n8454 & n8628 ) | ( n8454 & ~n8635 ) | ( n8628 & ~n8635 ) ;
  assign n8638 = n8637 ^ n8636 ^ n457 ;
  assign n8639 = n8308 ^ n6736 ^ n1969 ;
  assign n8640 = n8639 ^ n2689 ^ n1164 ;
  assign n8642 = n5636 & ~n6253 ;
  assign n8641 = n2158 ^ n1781 ^ x209 ;
  assign n8643 = n8642 ^ n8641 ^ 1'b0 ;
  assign n8644 = n8640 | n8643 ;
  assign n8645 = n3259 ^ n2552 ^ 1'b0 ;
  assign n8646 = n8645 ^ n4831 ^ n2893 ;
  assign n8647 = n8646 ^ n8338 ^ n8301 ;
  assign n8648 = n8647 ^ n7188 ^ n5033 ;
  assign n8649 = ( ~n2282 & n5750 ) | ( ~n2282 & n6191 ) | ( n5750 & n6191 ) ;
  assign n8651 = ( n574 & n837 ) | ( n574 & n1475 ) | ( n837 & n1475 ) ;
  assign n8652 = n2261 ^ n813 ^ 1'b0 ;
  assign n8653 = n294 | n8652 ;
  assign n8654 = ( ~n378 & n5876 ) | ( ~n378 & n8653 ) | ( n5876 & n8653 ) ;
  assign n8655 = ( x10 & ~n8651 ) | ( x10 & n8654 ) | ( ~n8651 & n8654 ) ;
  assign n8650 = n2984 & ~n4021 ;
  assign n8656 = n8655 ^ n8650 ^ 1'b0 ;
  assign n8658 = n6259 ^ n1277 ^ n1081 ;
  assign n8657 = n4379 ^ n2325 ^ n1293 ;
  assign n8659 = n8658 ^ n8657 ^ n6683 ;
  assign n8660 = ( x70 & n1463 ) | ( x70 & ~n1928 ) | ( n1463 & ~n1928 ) ;
  assign n8661 = n8660 ^ n4472 ^ x44 ;
  assign n8662 = ~n1589 & n5126 ;
  assign n8663 = ~n1359 & n8662 ;
  assign n8664 = ( n1676 & ~n2877 ) | ( n1676 & n8663 ) | ( ~n2877 & n8663 ) ;
  assign n8665 = n8664 ^ n7422 ^ n3592 ;
  assign n8668 = ( n485 & n1458 ) | ( n485 & ~n6690 ) | ( n1458 & ~n6690 ) ;
  assign n8669 = n8668 ^ n3616 ^ n2310 ;
  assign n8670 = n8669 ^ n6084 ^ n4063 ;
  assign n8666 = ( n2133 & ~n2862 ) | ( n2133 & n6544 ) | ( ~n2862 & n6544 ) ;
  assign n8667 = ( n4591 & n7442 ) | ( n4591 & n8666 ) | ( n7442 & n8666 ) ;
  assign n8671 = n8670 ^ n8667 ^ n5048 ;
  assign n8672 = ( n8661 & n8665 ) | ( n8661 & n8671 ) | ( n8665 & n8671 ) ;
  assign n8690 = n3205 ^ n2387 ^ n2274 ;
  assign n8691 = n8690 ^ n3705 ^ n415 ;
  assign n8675 = n1164 & ~n1796 ;
  assign n8676 = n8675 ^ n2727 ^ 1'b0 ;
  assign n8677 = n8676 ^ n1166 ^ 1'b0 ;
  assign n8678 = n3181 & ~n8677 ;
  assign n8679 = n8678 ^ n1894 ^ n1762 ;
  assign n8673 = ( n302 & ~n4141 ) | ( n302 & n4192 ) | ( ~n4141 & n4192 ) ;
  assign n8674 = ( n4375 & n7591 ) | ( n4375 & n8673 ) | ( n7591 & n8673 ) ;
  assign n8680 = n8679 ^ n8674 ^ n2811 ;
  assign n8683 = ( n2681 & n2723 ) | ( n2681 & ~n5884 ) | ( n2723 & ~n5884 ) ;
  assign n8684 = ~n336 & n8683 ;
  assign n8685 = n8684 ^ n7880 ^ 1'b0 ;
  assign n8681 = n2790 ^ n1423 ^ n881 ;
  assign n8682 = ( n1594 & n6483 ) | ( n1594 & ~n8681 ) | ( n6483 & ~n8681 ) ;
  assign n8686 = n8685 ^ n8682 ^ n5287 ;
  assign n8687 = ( n4043 & ~n5264 ) | ( n4043 & n8686 ) | ( ~n5264 & n8686 ) ;
  assign n8688 = ( n5662 & n8680 ) | ( n5662 & n8687 ) | ( n8680 & n8687 ) ;
  assign n8689 = ( n2957 & n6421 ) | ( n2957 & n8688 ) | ( n6421 & n8688 ) ;
  assign n8692 = n8691 ^ n8689 ^ n7802 ;
  assign n8693 = n6491 ^ n755 ^ 1'b0 ;
  assign n8694 = n5369 ^ n3709 ^ n2267 ;
  assign n8695 = ( n2724 & n3624 ) | ( n2724 & n8694 ) | ( n3624 & n8694 ) ;
  assign n8696 = ( ~n3728 & n6223 ) | ( ~n3728 & n8695 ) | ( n6223 & n8695 ) ;
  assign n8697 = n4467 ^ n1936 ^ n1793 ;
  assign n8698 = ( n1631 & n7756 ) | ( n1631 & ~n8697 ) | ( n7756 & ~n8697 ) ;
  assign n8699 = ( n5811 & n8696 ) | ( n5811 & n8698 ) | ( n8696 & n8698 ) ;
  assign n8700 = ( n2045 & n2234 ) | ( n2045 & ~n8699 ) | ( n2234 & ~n8699 ) ;
  assign n8701 = ( ~n2480 & n8693 ) | ( ~n2480 & n8700 ) | ( n8693 & n8700 ) ;
  assign n8702 = n3779 ^ x70 ^ x17 ;
  assign n8703 = ( ~n1988 & n7343 ) | ( ~n1988 & n8702 ) | ( n7343 & n8702 ) ;
  assign n8704 = ( n6149 & n7529 ) | ( n6149 & ~n8703 ) | ( n7529 & ~n8703 ) ;
  assign n8705 = ( n6132 & n8701 ) | ( n6132 & ~n8704 ) | ( n8701 & ~n8704 ) ;
  assign n8707 = n1573 ^ n628 ^ x175 ;
  assign n8706 = n6980 ^ n6911 ^ n4324 ;
  assign n8708 = n8707 ^ n8706 ^ n2534 ;
  assign n8712 = n8379 ^ n7858 ^ n821 ;
  assign n8709 = n4861 ^ n2510 ^ 1'b0 ;
  assign n8710 = n8709 ^ n2565 ^ n1749 ;
  assign n8711 = n8710 ^ n6220 ^ 1'b0 ;
  assign n8713 = n8712 ^ n8711 ^ n8148 ;
  assign n8714 = n2863 ^ n2611 ^ n1086 ;
  assign n8715 = n539 & n8714 ;
  assign n8716 = ~n8501 & n8715 ;
  assign n8717 = ( n5515 & n6976 ) | ( n5515 & ~n8716 ) | ( n6976 & ~n8716 ) ;
  assign n8721 = ~n3635 & n6770 ;
  assign n8722 = ~n5223 & n8721 ;
  assign n8723 = n6573 | n8722 ;
  assign n8724 = n2538 & ~n8723 ;
  assign n8720 = ( ~x125 & n2856 ) | ( ~x125 & n5794 ) | ( n2856 & n5794 ) ;
  assign n8725 = n8724 ^ n8720 ^ n4080 ;
  assign n8718 = n7224 ^ n2498 ^ 1'b0 ;
  assign n8719 = n3694 | n8718 ;
  assign n8726 = n8725 ^ n8719 ^ 1'b0 ;
  assign n8727 = n5288 ^ n1831 ^ 1'b0 ;
  assign n8728 = ( n1683 & n2160 ) | ( n1683 & ~n2971 ) | ( n2160 & ~n2971 ) ;
  assign n8729 = ( ~n4695 & n8727 ) | ( ~n4695 & n8728 ) | ( n8727 & n8728 ) ;
  assign n8730 = n4345 & ~n7357 ;
  assign n8731 = n8730 ^ n5339 ^ 1'b0 ;
  assign n8732 = n3127 & ~n8731 ;
  assign n8733 = n8499 ^ n3425 ^ n761 ;
  assign n8735 = n3004 ^ n1752 ^ x2 ;
  assign n8736 = n8735 ^ n8286 ^ n3680 ;
  assign n8734 = ( ~n936 & n3652 ) | ( ~n936 & n7790 ) | ( n3652 & n7790 ) ;
  assign n8737 = n8736 ^ n8734 ^ n4306 ;
  assign n8738 = n8737 ^ n8130 ^ n5323 ;
  assign n8739 = ~x188 & n2695 ;
  assign n8741 = n3822 ^ n1515 ^ n745 ;
  assign n8740 = n2941 ^ n2737 ^ n1970 ;
  assign n8742 = n8741 ^ n8740 ^ n322 ;
  assign n8743 = ( ~n872 & n1602 ) | ( ~n872 & n8742 ) | ( n1602 & n8742 ) ;
  assign n8744 = ~n8739 & n8743 ;
  assign n8745 = ( n8733 & ~n8738 ) | ( n8733 & n8744 ) | ( ~n8738 & n8744 ) ;
  assign n8746 = n5183 ^ n3878 ^ 1'b0 ;
  assign n8747 = n2856 & n8746 ;
  assign n8748 = n8747 ^ n5926 ^ n1392 ;
  assign n8751 = n1418 ^ n294 ^ n260 ;
  assign n8749 = n2081 ^ n1818 ^ x237 ;
  assign n8750 = ( n4948 & ~n6487 ) | ( n4948 & n8749 ) | ( ~n6487 & n8749 ) ;
  assign n8752 = n8751 ^ n8750 ^ n1973 ;
  assign n8753 = n1875 & n8752 ;
  assign n8754 = ( ~n5938 & n8748 ) | ( ~n5938 & n8753 ) | ( n8748 & n8753 ) ;
  assign n8758 = ( n1385 & n3183 ) | ( n1385 & n5828 ) | ( n3183 & n5828 ) ;
  assign n8759 = n8345 ^ n7593 ^ 1'b0 ;
  assign n8760 = n5367 & ~n8759 ;
  assign n8761 = n8758 & ~n8760 ;
  assign n8762 = n8761 ^ n2117 ^ x27 ;
  assign n8763 = n2020 | n8762 ;
  assign n8756 = n1440 | n4056 ;
  assign n8757 = ( ~n3997 & n5351 ) | ( ~n3997 & n8756 ) | ( n5351 & n8756 ) ;
  assign n8755 = ( n1696 & ~n5053 ) | ( n1696 & n6259 ) | ( ~n5053 & n6259 ) ;
  assign n8764 = n8763 ^ n8757 ^ n8755 ;
  assign n8765 = n6917 ^ n4048 ^ n1581 ;
  assign n8766 = n6594 ^ n2108 ^ 1'b0 ;
  assign n8767 = ( n1546 & ~n6068 ) | ( n1546 & n8766 ) | ( ~n6068 & n8766 ) ;
  assign n8768 = ( ~n368 & n3250 ) | ( ~n368 & n8253 ) | ( n3250 & n8253 ) ;
  assign n8769 = ( n6788 & ~n8767 ) | ( n6788 & n8768 ) | ( ~n8767 & n8768 ) ;
  assign n8770 = n8769 ^ n6283 ^ 1'b0 ;
  assign n8771 = n8765 & n8770 ;
  assign n8772 = ( n4584 & n4943 ) | ( n4584 & ~n6640 ) | ( n4943 & ~n6640 ) ;
  assign n8773 = n7738 ^ n7546 ^ n7424 ;
  assign n8774 = ( n6050 & n8772 ) | ( n6050 & n8773 ) | ( n8772 & n8773 ) ;
  assign n8775 = ( n1557 & n3306 ) | ( n1557 & n3432 ) | ( n3306 & n3432 ) ;
  assign n8776 = n1898 & ~n8775 ;
  assign n8777 = ( n4151 & n6401 ) | ( n4151 & ~n8776 ) | ( n6401 & ~n8776 ) ;
  assign n8778 = n8777 ^ n8429 ^ n5352 ;
  assign n8779 = n8778 ^ n3317 ^ n2832 ;
  assign n8780 = n3114 & n6272 ;
  assign n8787 = n6496 ^ n3487 ^ n2891 ;
  assign n8785 = n6068 ^ n2311 ^ 1'b0 ;
  assign n8786 = n5525 & ~n8785 ;
  assign n8788 = n8787 ^ n8786 ^ 1'b0 ;
  assign n8782 = ( n1650 & n2452 ) | ( n1650 & n6608 ) | ( n2452 & n6608 ) ;
  assign n8783 = n8782 ^ n1030 ^ n643 ;
  assign n8784 = ( x24 & ~n3385 ) | ( x24 & n8783 ) | ( ~n3385 & n8783 ) ;
  assign n8789 = n8788 ^ n8784 ^ n2556 ;
  assign n8781 = n2234 & n5087 ;
  assign n8790 = n8789 ^ n8781 ^ 1'b0 ;
  assign n8791 = ( n4298 & ~n7120 ) | ( n4298 & n8790 ) | ( ~n7120 & n8790 ) ;
  assign n8795 = n2854 & n2919 ;
  assign n8792 = n2295 & ~n2438 ;
  assign n8793 = n8792 ^ n2517 ^ 1'b0 ;
  assign n8794 = ( x153 & n2521 ) | ( x153 & ~n8793 ) | ( n2521 & ~n8793 ) ;
  assign n8796 = n8795 ^ n8794 ^ n1025 ;
  assign n8797 = n8796 ^ n8225 ^ n2226 ;
  assign n8799 = n1816 ^ n1812 ^ n1396 ;
  assign n8798 = n2267 ^ n1603 ^ x1 ;
  assign n8800 = n8799 ^ n8798 ^ n1343 ;
  assign n8809 = n8358 ^ n7265 ^ n1898 ;
  assign n8810 = n8809 ^ n7995 ^ n7540 ;
  assign n8811 = n8810 ^ n5561 ^ n5505 ;
  assign n8801 = ~n854 & n4961 ;
  assign n8802 = n8801 ^ n522 ^ 1'b0 ;
  assign n8803 = n6497 ^ n1058 ^ n987 ;
  assign n8804 = n8803 ^ n6841 ^ n3910 ;
  assign n8805 = n8804 ^ n3832 ^ n687 ;
  assign n8806 = n7519 | n8805 ;
  assign n8807 = n4355 & ~n8806 ;
  assign n8808 = ( n693 & n8802 ) | ( n693 & n8807 ) | ( n8802 & n8807 ) ;
  assign n8812 = n8811 ^ n8808 ^ n266 ;
  assign n8818 = ( n1220 & n1507 ) | ( n1220 & n6520 ) | ( n1507 & n6520 ) ;
  assign n8819 = ( n3068 & n6035 ) | ( n3068 & n8818 ) | ( n6035 & n8818 ) ;
  assign n8815 = ( n5069 & n6600 ) | ( n5069 & ~n8323 ) | ( n6600 & ~n8323 ) ;
  assign n8813 = n7163 ^ n6222 ^ n1076 ;
  assign n8814 = n6244 | n8813 ;
  assign n8816 = n8815 ^ n8814 ^ 1'b0 ;
  assign n8817 = ( n6648 & n8746 ) | ( n6648 & n8816 ) | ( n8746 & n8816 ) ;
  assign n8820 = n8819 ^ n8817 ^ n2166 ;
  assign n8821 = n8820 ^ n7173 ^ n442 ;
  assign n8826 = ( n2373 & n3353 ) | ( n2373 & ~n5635 ) | ( n3353 & ~n5635 ) ;
  assign n8827 = ( ~x223 & n4680 ) | ( ~x223 & n8826 ) | ( n4680 & n8826 ) ;
  assign n8822 = n4976 ^ n3028 ^ n2679 ;
  assign n8823 = n6938 | n8822 ;
  assign n8824 = n8823 ^ n4213 ^ 1'b0 ;
  assign n8825 = ( ~n2448 & n8078 ) | ( ~n2448 & n8824 ) | ( n8078 & n8824 ) ;
  assign n8828 = n8827 ^ n8825 ^ n6775 ;
  assign n8835 = ( n794 & n1829 ) | ( n794 & ~n4536 ) | ( n1829 & ~n4536 ) ;
  assign n8829 = n7886 ^ n1118 ^ n1097 ;
  assign n8830 = ( n1130 & ~n3830 ) | ( n1130 & n8829 ) | ( ~n3830 & n8829 ) ;
  assign n8831 = ( n1528 & n2121 ) | ( n1528 & n5376 ) | ( n2121 & n5376 ) ;
  assign n8832 = ~n5916 & n7499 ;
  assign n8833 = n8832 ^ n2721 ^ 1'b0 ;
  assign n8834 = ( ~n8830 & n8831 ) | ( ~n8830 & n8833 ) | ( n8831 & n8833 ) ;
  assign n8836 = n8835 ^ n8834 ^ 1'b0 ;
  assign n8837 = n3076 & ~n8836 ;
  assign n8838 = ( n3065 & ~n5136 ) | ( n3065 & n8547 ) | ( ~n5136 & n8547 ) ;
  assign n8839 = ( n1636 & n6198 ) | ( n1636 & n8838 ) | ( n6198 & n8838 ) ;
  assign n8840 = n8839 ^ n7129 ^ n6978 ;
  assign n8862 = ( n2013 & n2398 ) | ( n2013 & ~n5814 ) | ( n2398 & ~n5814 ) ;
  assign n8842 = ( n3132 & n3954 ) | ( n3132 & ~n5775 ) | ( n3954 & ~n5775 ) ;
  assign n8841 = n8066 ^ n7987 ^ n2392 ;
  assign n8843 = n8842 ^ n8841 ^ n5275 ;
  assign n8844 = n7123 ^ n1831 ^ n692 ;
  assign n8845 = n871 ^ n633 ^ 1'b0 ;
  assign n8846 = ~n8844 & n8845 ;
  assign n8847 = n8846 ^ n6994 ^ 1'b0 ;
  assign n8848 = n6996 & n8847 ;
  assign n8857 = n4856 & n6287 ;
  assign n8858 = n8857 ^ n815 ^ n646 ;
  assign n8855 = ( n383 & n1016 ) | ( n383 & n3379 ) | ( n1016 & n3379 ) ;
  assign n8856 = n8855 ^ n3718 ^ n3302 ;
  assign n8859 = n8858 ^ n8856 ^ n1104 ;
  assign n8851 = x132 & n1160 ;
  assign n8852 = n8851 ^ n1191 ^ 1'b0 ;
  assign n8853 = ( n1454 & n2597 ) | ( n1454 & n8852 ) | ( n2597 & n8852 ) ;
  assign n8854 = n8853 ^ n2251 ^ n1787 ;
  assign n8849 = n1746 ^ n940 ^ x109 ;
  assign n8850 = ( n1086 & ~n2246 ) | ( n1086 & n8849 ) | ( ~n2246 & n8849 ) ;
  assign n8860 = n8859 ^ n8854 ^ n8850 ;
  assign n8861 = ( ~n8843 & n8848 ) | ( ~n8843 & n8860 ) | ( n8848 & n8860 ) ;
  assign n8863 = n8862 ^ n8861 ^ n3638 ;
  assign n8873 = n7907 ^ n770 ^ 1'b0 ;
  assign n8870 = n7785 ^ n3578 ^ n1823 ;
  assign n8871 = ( n2085 & n3924 ) | ( n2085 & ~n8870 ) | ( n3924 & ~n8870 ) ;
  assign n8867 = ( n2470 & n3148 ) | ( n2470 & n4403 ) | ( n3148 & n4403 ) ;
  assign n8868 = n4776 ^ n4167 ^ 1'b0 ;
  assign n8869 = ( n947 & ~n8867 ) | ( n947 & n8868 ) | ( ~n8867 & n8868 ) ;
  assign n8872 = n8871 ^ n8869 ^ n8222 ;
  assign n8874 = n8873 ^ n8872 ^ n7929 ;
  assign n8864 = ( n4630 & n5191 ) | ( n4630 & ~n5955 ) | ( n5191 & ~n5955 ) ;
  assign n8865 = n8864 ^ n6089 ^ n2368 ;
  assign n8866 = n4105 & n8865 ;
  assign n8875 = n8874 ^ n8866 ^ 1'b0 ;
  assign n8876 = n3893 ^ n2499 ^ n2153 ;
  assign n8877 = ( n1979 & ~n2485 ) | ( n1979 & n6488 ) | ( ~n2485 & n6488 ) ;
  assign n8878 = ( n5354 & n8876 ) | ( n5354 & ~n8877 ) | ( n8876 & ~n8877 ) ;
  assign n8879 = ( n2739 & ~n3628 ) | ( n2739 & n6957 ) | ( ~n3628 & n6957 ) ;
  assign n8880 = n8879 ^ n2351 ^ 1'b0 ;
  assign n8881 = ( n4147 & n4903 ) | ( n4147 & n8880 ) | ( n4903 & n8880 ) ;
  assign n8882 = ( n5367 & n5755 ) | ( n5367 & n8881 ) | ( n5755 & n8881 ) ;
  assign n8886 = ( x34 & n890 ) | ( x34 & n4302 ) | ( n890 & n4302 ) ;
  assign n8883 = ~n3771 & n5585 ;
  assign n8884 = n8883 ^ n6451 ^ 1'b0 ;
  assign n8885 = n8884 ^ n7908 ^ n5680 ;
  assign n8887 = n8886 ^ n8885 ^ n5755 ;
  assign n8888 = n1416 | n8887 ;
  assign n8889 = n8882 | n8888 ;
  assign n8890 = ( n1122 & n1810 ) | ( n1122 & ~n4198 ) | ( n1810 & ~n4198 ) ;
  assign n8891 = n5777 ^ n3012 ^ n1401 ;
  assign n8892 = ( ~n3265 & n8890 ) | ( ~n3265 & n8891 ) | ( n8890 & n8891 ) ;
  assign n8893 = n8892 ^ n7767 ^ n2268 ;
  assign n8894 = ( n2296 & ~n3956 ) | ( n2296 & n6262 ) | ( ~n3956 & n6262 ) ;
  assign n8895 = n8894 ^ n6381 ^ n1722 ;
  assign n8896 = ( n4172 & n4807 ) | ( n4172 & ~n8895 ) | ( n4807 & ~n8895 ) ;
  assign n8897 = n8896 ^ n2193 ^ n898 ;
  assign n8898 = ( n7546 & n8143 ) | ( n7546 & n8897 ) | ( n8143 & n8897 ) ;
  assign n8902 = n5115 ^ n1988 ^ 1'b0 ;
  assign n8899 = ( n598 & n1556 ) | ( n598 & ~n2980 ) | ( n1556 & ~n2980 ) ;
  assign n8900 = ( n1346 & n2145 ) | ( n1346 & ~n4889 ) | ( n2145 & ~n4889 ) ;
  assign n8901 = ( n1541 & n8899 ) | ( n1541 & n8900 ) | ( n8899 & n8900 ) ;
  assign n8903 = n8902 ^ n8901 ^ n831 ;
  assign n8904 = n5276 ^ n1302 ^ x206 ;
  assign n8905 = ( n6004 & n8903 ) | ( n6004 & n8904 ) | ( n8903 & n8904 ) ;
  assign n8907 = n4158 ^ n847 ^ 1'b0 ;
  assign n8908 = n8907 ^ n4400 ^ n2338 ;
  assign n8906 = n463 & n2695 ;
  assign n8909 = n8908 ^ n8906 ^ 1'b0 ;
  assign n8910 = ( n524 & n980 ) | ( n524 & ~n3211 ) | ( n980 & ~n3211 ) ;
  assign n8911 = n4668 ^ n4070 ^ n1188 ;
  assign n8912 = n8911 ^ n4835 ^ n1008 ;
  assign n8913 = ( n551 & ~n3131 ) | ( n551 & n4168 ) | ( ~n3131 & n4168 ) ;
  assign n8914 = ( n8233 & ~n8912 ) | ( n8233 & n8913 ) | ( ~n8912 & n8913 ) ;
  assign n8915 = ( n3269 & ~n8611 ) | ( n3269 & n8914 ) | ( ~n8611 & n8914 ) ;
  assign n8918 = ( n1308 & ~n1843 ) | ( n1308 & n3770 ) | ( ~n1843 & n3770 ) ;
  assign n8919 = n8918 ^ n5938 ^ n335 ;
  assign n8916 = n5197 ^ n2796 ^ n2282 ;
  assign n8917 = ( ~n2328 & n2642 ) | ( ~n2328 & n8916 ) | ( n2642 & n8916 ) ;
  assign n8920 = n8919 ^ n8917 ^ n1396 ;
  assign n8926 = ~n2128 & n7088 ;
  assign n8927 = n8926 ^ n4100 ^ 1'b0 ;
  assign n8928 = n2431 | n8927 ;
  assign n8929 = ( ~n407 & n2647 ) | ( ~n407 & n8928 ) | ( n2647 & n8928 ) ;
  assign n8924 = n2180 ^ n715 ^ 1'b0 ;
  assign n8925 = ( n362 & n3523 ) | ( n362 & ~n8924 ) | ( n3523 & ~n8924 ) ;
  assign n8930 = n8929 ^ n8925 ^ n851 ;
  assign n8931 = ( x100 & ~n4363 ) | ( x100 & n8930 ) | ( ~n4363 & n8930 ) ;
  assign n8932 = n7149 & ~n8931 ;
  assign n8921 = ( n424 & n970 ) | ( n424 & n4687 ) | ( n970 & n4687 ) ;
  assign n8922 = ( n2536 & n7656 ) | ( n2536 & n8921 ) | ( n7656 & n8921 ) ;
  assign n8923 = n8922 ^ n820 ^ n782 ;
  assign n8933 = n8932 ^ n8923 ^ 1'b0 ;
  assign n8934 = ~n5840 & n8933 ;
  assign n8935 = n4583 ^ n2859 ^ 1'b0 ;
  assign n8939 = n2563 ^ n2319 ^ n1312 ;
  assign n8936 = n7587 ^ n5422 ^ 1'b0 ;
  assign n8937 = ~n2889 & n8936 ;
  assign n8938 = ( n5544 & n8816 ) | ( n5544 & n8937 ) | ( n8816 & n8937 ) ;
  assign n8940 = n8939 ^ n8938 ^ 1'b0 ;
  assign n8941 = ( n2718 & n8935 ) | ( n2718 & ~n8940 ) | ( n8935 & ~n8940 ) ;
  assign n8942 = n8034 ^ n3393 ^ n1222 ;
  assign n8968 = n2534 ^ n2246 ^ n665 ;
  assign n8969 = n8968 ^ n6288 ^ n5329 ;
  assign n8970 = n8969 ^ n6554 ^ n1134 ;
  assign n8967 = n486 & ~n5299 ;
  assign n8971 = n8970 ^ n8967 ^ 1'b0 ;
  assign n8961 = n1949 ^ n1221 ^ 1'b0 ;
  assign n8962 = ~n8560 & n8961 ;
  assign n8963 = x92 & n417 ;
  assign n8964 = ~x197 & n8963 ;
  assign n8965 = n8964 ^ n7483 ^ 1'b0 ;
  assign n8966 = n8962 & ~n8965 ;
  assign n8943 = ( x43 & x199 ) | ( x43 & ~n2935 ) | ( x199 & ~n2935 ) ;
  assign n8944 = n8943 ^ n8429 ^ n1075 ;
  assign n8945 = ( n500 & ~n3803 ) | ( n500 & n8944 ) | ( ~n3803 & n8944 ) ;
  assign n8953 = n3920 ^ n2136 ^ x147 ;
  assign n8954 = n1015 & n7880 ;
  assign n8955 = n8954 ^ n6409 ^ 1'b0 ;
  assign n8956 = n8618 & n8955 ;
  assign n8957 = ~n8953 & n8956 ;
  assign n8958 = n8957 ^ n5870 ^ n4899 ;
  assign n8946 = n2426 ^ n1614 ^ n1232 ;
  assign n8947 = ( n5345 & n6469 ) | ( n5345 & ~n8946 ) | ( n6469 & ~n8946 ) ;
  assign n8948 = ( ~n2386 & n4654 ) | ( ~n2386 & n8947 ) | ( n4654 & n8947 ) ;
  assign n8950 = ( ~n1153 & n1702 ) | ( ~n1153 & n2662 ) | ( n1702 & n2662 ) ;
  assign n8949 = n1315 ^ x199 ^ x163 ;
  assign n8951 = n8950 ^ n8949 ^ n3731 ;
  assign n8952 = n8948 & n8951 ;
  assign n8959 = n8958 ^ n8952 ^ 1'b0 ;
  assign n8960 = ( n4692 & n8945 ) | ( n4692 & n8959 ) | ( n8945 & n8959 ) ;
  assign n8972 = n8971 ^ n8966 ^ n8960 ;
  assign n8973 = n3856 ^ n2652 ^ n1418 ;
  assign n8974 = ( n1243 & n1318 ) | ( n1243 & ~n6131 ) | ( n1318 & ~n6131 ) ;
  assign n8975 = ( n4945 & n5310 ) | ( n4945 & ~n8974 ) | ( n5310 & ~n8974 ) ;
  assign n8976 = ( n8112 & n8973 ) | ( n8112 & n8975 ) | ( n8973 & n8975 ) ;
  assign n8986 = n7434 ^ n4928 ^ n1927 ;
  assign n8984 = ( n1457 & n1895 ) | ( n1457 & ~n3352 ) | ( n1895 & ~n3352 ) ;
  assign n8982 = ( n848 & n4231 ) | ( n848 & n8697 ) | ( n4231 & n8697 ) ;
  assign n8983 = n8982 ^ n7112 ^ n5759 ;
  assign n8985 = n8984 ^ n8983 ^ 1'b0 ;
  assign n8977 = n1436 ^ n565 ^ 1'b0 ;
  assign n8978 = n3372 ^ n2251 ^ n542 ;
  assign n8979 = n8978 ^ n3151 ^ n2000 ;
  assign n8980 = n7142 ^ n6608 ^ 1'b0 ;
  assign n8981 = ( ~n8977 & n8979 ) | ( ~n8977 & n8980 ) | ( n8979 & n8980 ) ;
  assign n8987 = n8986 ^ n8985 ^ n8981 ;
  assign n8988 = n8987 ^ n3245 ^ n2919 ;
  assign n8989 = ( n1078 & n8976 ) | ( n1078 & n8988 ) | ( n8976 & n8988 ) ;
  assign n8996 = ( n358 & n6010 ) | ( n358 & n6851 ) | ( n6010 & n6851 ) ;
  assign n8993 = n7714 ^ n3758 ^ n1225 ;
  assign n8994 = ( n4765 & n6922 ) | ( n4765 & ~n8993 ) | ( n6922 & ~n8993 ) ;
  assign n8995 = n8994 ^ n3477 ^ n715 ;
  assign n8990 = ( n3691 & ~n5304 ) | ( n3691 & n7908 ) | ( ~n5304 & n7908 ) ;
  assign n8991 = ( n2000 & n7132 ) | ( n2000 & n8990 ) | ( n7132 & n8990 ) ;
  assign n8992 = ( n5128 & ~n8489 ) | ( n5128 & n8991 ) | ( ~n8489 & n8991 ) ;
  assign n8997 = n8996 ^ n8995 ^ n8992 ;
  assign n8998 = ( n1028 & n1698 ) | ( n1028 & n8997 ) | ( n1698 & n8997 ) ;
  assign n9002 = ( n288 & n1176 ) | ( n288 & ~n1536 ) | ( n1176 & ~n1536 ) ;
  assign n9003 = n9002 ^ n7128 ^ n5237 ;
  assign n9004 = n9003 ^ n6031 ^ n3958 ;
  assign n8999 = ( n1771 & n4093 ) | ( n1771 & n5650 ) | ( n4093 & n5650 ) ;
  assign n9000 = ( x29 & n4687 ) | ( x29 & n8999 ) | ( n4687 & n8999 ) ;
  assign n9001 = ~n3384 & n9000 ;
  assign n9005 = n9004 ^ n9001 ^ 1'b0 ;
  assign n9006 = n6326 ^ n4856 ^ n4672 ;
  assign n9007 = n6089 ^ n1766 ^ 1'b0 ;
  assign n9008 = n2290 | n9007 ;
  assign n9009 = n9006 & ~n9008 ;
  assign n9010 = n9009 ^ n1768 ^ 1'b0 ;
  assign n9011 = n6530 & n9010 ;
  assign n9012 = ( n7756 & n8765 ) | ( n7756 & n9011 ) | ( n8765 & n9011 ) ;
  assign n9013 = ~n1383 & n9012 ;
  assign n9014 = ( x182 & n2544 ) | ( x182 & n4156 ) | ( n2544 & n4156 ) ;
  assign n9015 = ( n1167 & ~n5084 ) | ( n1167 & n9014 ) | ( ~n5084 & n9014 ) ;
  assign n9016 = ( n1439 & ~n8178 ) | ( n1439 & n9015 ) | ( ~n8178 & n9015 ) ;
  assign n9017 = n9016 ^ n3748 ^ n2731 ;
  assign n9018 = ( n285 & n6975 ) | ( n285 & ~n9017 ) | ( n6975 & ~n9017 ) ;
  assign n9025 = n3552 ^ n1892 ^ n1427 ;
  assign n9026 = ( n3432 & n5938 ) | ( n3432 & n9025 ) | ( n5938 & n9025 ) ;
  assign n9027 = n9026 ^ n6803 ^ n3252 ;
  assign n9028 = ( n498 & ~n6272 ) | ( n498 & n9027 ) | ( ~n6272 & n9027 ) ;
  assign n9022 = ( n448 & ~n621 ) | ( n448 & n1164 ) | ( ~n621 & n1164 ) ;
  assign n9023 = n9022 ^ n2739 ^ n1793 ;
  assign n9021 = n6558 ^ n3688 ^ x107 ;
  assign n9024 = n9023 ^ n9021 ^ n8426 ;
  assign n9019 = n7816 ^ n3239 ^ 1'b0 ;
  assign n9020 = ~n8762 & n9019 ;
  assign n9029 = n9028 ^ n9024 ^ n9020 ;
  assign n9035 = n4097 ^ n1889 ^ n1539 ;
  assign n9036 = ( ~n4647 & n6256 ) | ( ~n4647 & n6534 ) | ( n6256 & n6534 ) ;
  assign n9037 = n9036 ^ n4542 ^ n1250 ;
  assign n9038 = ( n5880 & n9035 ) | ( n5880 & ~n9037 ) | ( n9035 & ~n9037 ) ;
  assign n9033 = n7842 ^ n4318 ^ n915 ;
  assign n9030 = n8181 ^ n6826 ^ n2293 ;
  assign n9031 = n9030 ^ n7548 ^ n669 ;
  assign n9032 = ( n727 & n3274 ) | ( n727 & n9031 ) | ( n3274 & n9031 ) ;
  assign n9034 = n9033 ^ n9032 ^ x81 ;
  assign n9039 = n9038 ^ n9034 ^ 1'b0 ;
  assign n9040 = n5776 ^ n2977 ^ n1941 ;
  assign n9041 = ( ~n2016 & n3622 ) | ( ~n2016 & n4676 ) | ( n3622 & n4676 ) ;
  assign n9042 = n5020 ^ n1819 ^ n622 ;
  assign n9043 = n3405 ^ n2518 ^ 1'b0 ;
  assign n9044 = ~n9042 & n9043 ;
  assign n9045 = ( n9040 & n9041 ) | ( n9040 & ~n9044 ) | ( n9041 & ~n9044 ) ;
  assign n9046 = n4426 | n5146 ;
  assign n9047 = n8437 & ~n9046 ;
  assign n9048 = n2758 ^ n1300 ^ n579 ;
  assign n9049 = n3596 & ~n9048 ;
  assign n9050 = n6286 & n9049 ;
  assign n9055 = n3484 ^ n1435 ^ n1332 ;
  assign n9052 = n3345 ^ n2072 ^ n539 ;
  assign n9053 = ( n3395 & ~n3810 ) | ( n3395 & n9052 ) | ( ~n3810 & n9052 ) ;
  assign n9051 = n6276 ^ n5107 ^ n1921 ;
  assign n9054 = n9053 ^ n9051 ^ n4751 ;
  assign n9056 = n9055 ^ n9054 ^ 1'b0 ;
  assign n9057 = n9050 & n9056 ;
  assign n9058 = ( n4449 & n8150 ) | ( n4449 & ~n9057 ) | ( n8150 & ~n9057 ) ;
  assign n9059 = n2202 ^ n1212 ^ x68 ;
  assign n9060 = ( n2080 & n6320 ) | ( n2080 & n9059 ) | ( n6320 & n9059 ) ;
  assign n9061 = ( ~n3982 & n6686 ) | ( ~n3982 & n6837 ) | ( n6686 & n6837 ) ;
  assign n9062 = ~n9060 & n9061 ;
  assign n9083 = n5334 ^ n4946 ^ n3452 ;
  assign n9084 = n9083 ^ n7112 ^ n5345 ;
  assign n9085 = n3808 ^ n2764 ^ 1'b0 ;
  assign n9086 = n9084 | n9085 ;
  assign n9063 = ( x147 & n821 ) | ( x147 & n2389 ) | ( n821 & n2389 ) ;
  assign n9065 = ( ~n737 & n860 ) | ( ~n737 & n4161 ) | ( n860 & n4161 ) ;
  assign n9064 = n6704 ^ n6645 ^ x66 ;
  assign n9066 = n9065 ^ n9064 ^ n5535 ;
  assign n9067 = n9066 ^ n3213 ^ n1971 ;
  assign n9068 = n2670 & ~n3736 ;
  assign n9069 = ~n7882 & n9068 ;
  assign n9070 = ( n510 & ~n621 ) | ( n510 & n2196 ) | ( ~n621 & n2196 ) ;
  assign n9071 = n9070 ^ n5665 ^ x184 ;
  assign n9072 = n2647 ^ n1036 ^ n680 ;
  assign n9073 = ( n1821 & n5141 ) | ( n1821 & ~n8022 ) | ( n5141 & ~n8022 ) ;
  assign n9074 = ( ~n4502 & n7715 ) | ( ~n4502 & n9073 ) | ( n7715 & n9073 ) ;
  assign n9075 = ~n3277 & n3664 ;
  assign n9076 = ~n527 & n9075 ;
  assign n9077 = ( n1595 & ~n6907 ) | ( n1595 & n9076 ) | ( ~n6907 & n9076 ) ;
  assign n9078 = n9077 ^ n8925 ^ n2837 ;
  assign n9079 = ( n9072 & ~n9074 ) | ( n9072 & n9078 ) | ( ~n9074 & n9078 ) ;
  assign n9080 = ( n9069 & n9071 ) | ( n9069 & n9079 ) | ( n9071 & n9079 ) ;
  assign n9081 = ( n9063 & ~n9067 ) | ( n9063 & n9080 ) | ( ~n9067 & n9080 ) ;
  assign n9082 = n9081 ^ n4045 ^ n2885 ;
  assign n9087 = n9086 ^ n9082 ^ n2679 ;
  assign n9088 = n8485 ^ n6283 ^ n3381 ;
  assign n9089 = ( n604 & n8592 ) | ( n604 & n9088 ) | ( n8592 & n9088 ) ;
  assign n9091 = n6659 ^ n5530 ^ n623 ;
  assign n9090 = ~x75 & n2251 ;
  assign n9092 = n9091 ^ n9090 ^ n6724 ;
  assign n9093 = ( n3608 & ~n9089 ) | ( n3608 & n9092 ) | ( ~n9089 & n9092 ) ;
  assign n9094 = n1621 ^ n1282 ^ x66 ;
  assign n9095 = ( n1784 & n4993 ) | ( n1784 & n9094 ) | ( n4993 & n9094 ) ;
  assign n9096 = ( ~n6202 & n6746 ) | ( ~n6202 & n9095 ) | ( n6746 & n9095 ) ;
  assign n9097 = n7987 ^ n7857 ^ n566 ;
  assign n9098 = n4876 ^ n2631 ^ n391 ;
  assign n9105 = ~n319 & n1991 ;
  assign n9104 = n6173 ^ n3276 ^ n2530 ;
  assign n9099 = n3376 | n5369 ;
  assign n9100 = n6114 ^ n3349 ^ 1'b0 ;
  assign n9101 = ( n4213 & n9099 ) | ( n4213 & n9100 ) | ( n9099 & n9100 ) ;
  assign n9102 = ( n3168 & n6617 ) | ( n3168 & ~n9101 ) | ( n6617 & ~n9101 ) ;
  assign n9103 = ( ~n3240 & n3604 ) | ( ~n3240 & n9102 ) | ( n3604 & n9102 ) ;
  assign n9106 = n9105 ^ n9104 ^ n9103 ;
  assign n9107 = ( n1083 & ~n9098 ) | ( n1083 & n9106 ) | ( ~n9098 & n9106 ) ;
  assign n9108 = ( ~n6001 & n9097 ) | ( ~n6001 & n9107 ) | ( n9097 & n9107 ) ;
  assign n9110 = n2862 ^ n2166 ^ n1924 ;
  assign n9109 = ( ~n627 & n3433 ) | ( ~n627 & n4998 ) | ( n3433 & n4998 ) ;
  assign n9111 = n9110 ^ n9109 ^ n5844 ;
  assign n9112 = ( x88 & n3873 ) | ( x88 & n8378 ) | ( n3873 & n8378 ) ;
  assign n9113 = n9112 ^ n4208 ^ n1609 ;
  assign n9114 = n4965 ^ n4726 ^ n476 ;
  assign n9115 = n495 ^ x253 ^ 1'b0 ;
  assign n9116 = n6733 | n9115 ;
  assign n9117 = n9114 | n9116 ;
  assign n9118 = n470 | n9117 ;
  assign n9119 = n5558 ^ n2954 ^ 1'b0 ;
  assign n9120 = n9119 ^ n5759 ^ n2468 ;
  assign n9121 = ( n2249 & ~n4564 ) | ( n2249 & n7505 ) | ( ~n4564 & n7505 ) ;
  assign n9122 = ( n4612 & ~n5649 ) | ( n4612 & n9121 ) | ( ~n5649 & n9121 ) ;
  assign n9123 = n3899 | n9122 ;
  assign n9124 = ( ~n2911 & n3664 ) | ( ~n2911 & n4383 ) | ( n3664 & n4383 ) ;
  assign n9125 = ( x180 & ~n3400 ) | ( x180 & n8429 ) | ( ~n3400 & n8429 ) ;
  assign n9126 = n9125 ^ n4492 ^ n1031 ;
  assign n9127 = ( n7217 & ~n9124 ) | ( n7217 & n9126 ) | ( ~n9124 & n9126 ) ;
  assign n9128 = ( n397 & n487 ) | ( n397 & n1956 ) | ( n487 & n1956 ) ;
  assign n9129 = ( n1911 & n4585 ) | ( n1911 & n9128 ) | ( n4585 & n9128 ) ;
  assign n9130 = n9129 ^ n7043 ^ n6777 ;
  assign n9131 = ( n4370 & ~n4780 ) | ( n4370 & n9128 ) | ( ~n4780 & n9128 ) ;
  assign n9132 = ( ~n1884 & n2089 ) | ( ~n1884 & n6699 ) | ( n2089 & n6699 ) ;
  assign n9133 = ( n3827 & ~n4258 ) | ( n3827 & n9132 ) | ( ~n4258 & n9132 ) ;
  assign n9134 = n9071 ^ n4462 ^ n3680 ;
  assign n9135 = ( ~n7771 & n9133 ) | ( ~n7771 & n9134 ) | ( n9133 & n9134 ) ;
  assign n9146 = ( n3349 & n4129 ) | ( n3349 & ~n6526 ) | ( n4129 & ~n6526 ) ;
  assign n9147 = n6530 | n9146 ;
  assign n9143 = n6312 ^ n2892 ^ n1756 ;
  assign n9141 = ( n2736 & n3524 ) | ( n2736 & ~n4693 ) | ( n3524 & ~n4693 ) ;
  assign n9142 = n9141 ^ n3105 ^ n2129 ;
  assign n9144 = n9143 ^ n9142 ^ n4778 ;
  assign n9139 = n5124 ^ n3272 ^ n853 ;
  assign n9140 = n9139 ^ n5383 ^ n4029 ;
  assign n9136 = ( n3632 & ~n4113 ) | ( n3632 & n5492 ) | ( ~n4113 & n5492 ) ;
  assign n9137 = n7087 ^ n2054 ^ 1'b0 ;
  assign n9138 = n9136 & n9137 ;
  assign n9145 = n9144 ^ n9140 ^ n9138 ;
  assign n9148 = n9147 ^ n9145 ^ n4698 ;
  assign n9149 = ( n9131 & ~n9135 ) | ( n9131 & n9148 ) | ( ~n9135 & n9148 ) ;
  assign n9150 = ( n421 & ~n996 ) | ( n421 & n4378 ) | ( ~n996 & n4378 ) ;
  assign n9155 = ( n333 & ~n2282 ) | ( n333 & n3719 ) | ( ~n2282 & n3719 ) ;
  assign n9152 = n301 | n5413 ;
  assign n9153 = n1394 & ~n9152 ;
  assign n9151 = n4990 ^ n3688 ^ n2001 ;
  assign n9154 = n9153 ^ n9151 ^ n4416 ;
  assign n9156 = n9155 ^ n9154 ^ n2401 ;
  assign n9157 = n9156 ^ n6516 ^ n5691 ;
  assign n9158 = ~n320 & n1844 ;
  assign n9159 = n9158 ^ n5289 ^ 1'b0 ;
  assign n9160 = ( n3452 & ~n3498 ) | ( n3452 & n9159 ) | ( ~n3498 & n9159 ) ;
  assign n9161 = n9160 ^ n8349 ^ n539 ;
  assign n9164 = n2721 ^ n758 ^ n755 ;
  assign n9163 = n4984 ^ n3426 ^ n2013 ;
  assign n9162 = ( n1147 & n5377 ) | ( n1147 & ~n6237 ) | ( n5377 & ~n6237 ) ;
  assign n9165 = n9164 ^ n9163 ^ n9162 ;
  assign n9166 = n8257 ^ n1541 ^ n1409 ;
  assign n9167 = ( n449 & n4011 ) | ( n449 & ~n5654 ) | ( n4011 & ~n5654 ) ;
  assign n9168 = ( n9165 & n9166 ) | ( n9165 & n9167 ) | ( n9166 & n9167 ) ;
  assign n9169 = n3475 & n6160 ;
  assign n9170 = n9169 ^ n3941 ^ n1172 ;
  assign n9171 = ( n1399 & n3601 ) | ( n1399 & n6115 ) | ( n3601 & n6115 ) ;
  assign n9172 = n8527 ^ n6707 ^ 1'b0 ;
  assign n9173 = ~n2580 & n9172 ;
  assign n9185 = n5954 ^ n5201 ^ n2439 ;
  assign n9184 = n4079 ^ n2474 ^ n598 ;
  assign n9182 = ( ~n1010 & n1687 ) | ( ~n1010 & n5567 ) | ( n1687 & n5567 ) ;
  assign n9181 = ( n3886 & n4698 ) | ( n3886 & n8654 ) | ( n4698 & n8654 ) ;
  assign n9179 = ( ~n1966 & n2750 ) | ( ~n1966 & n4168 ) | ( n2750 & n4168 ) ;
  assign n9174 = ( ~n450 & n1409 ) | ( ~n450 & n3067 ) | ( n1409 & n3067 ) ;
  assign n9175 = n4260 ^ n3856 ^ n3257 ;
  assign n9176 = ( n1519 & ~n9174 ) | ( n1519 & n9175 ) | ( ~n9174 & n9175 ) ;
  assign n9177 = ( n6051 & n7978 ) | ( n6051 & ~n9176 ) | ( n7978 & ~n9176 ) ;
  assign n9178 = ( x160 & ~n2494 ) | ( x160 & n9177 ) | ( ~n2494 & n9177 ) ;
  assign n9180 = n9179 ^ n9178 ^ n417 ;
  assign n9183 = n9182 ^ n9181 ^ n9180 ;
  assign n9186 = n9185 ^ n9184 ^ n9183 ;
  assign n9187 = ( ~n9171 & n9173 ) | ( ~n9171 & n9186 ) | ( n9173 & n9186 ) ;
  assign n9188 = ( ~x251 & n1196 ) | ( ~x251 & n3634 ) | ( n1196 & n3634 ) ;
  assign n9189 = ( n2521 & n3461 ) | ( n2521 & n3567 ) | ( n3461 & n3567 ) ;
  assign n9203 = ( n578 & n1281 ) | ( n578 & ~n5074 ) | ( n1281 & ~n5074 ) ;
  assign n9204 = ( ~n1160 & n3772 ) | ( ~n1160 & n9203 ) | ( n3772 & n9203 ) ;
  assign n9205 = ( n4837 & ~n7066 ) | ( n4837 & n9204 ) | ( ~n7066 & n9204 ) ;
  assign n9202 = n7488 ^ n3059 ^ n809 ;
  assign n9206 = n9205 ^ n9202 ^ n319 ;
  assign n9196 = n5134 ^ n2469 ^ n404 ;
  assign n9197 = n9196 ^ n4419 ^ n2284 ;
  assign n9198 = n9197 ^ n5719 ^ n2125 ;
  assign n9199 = ( n3354 & n7526 ) | ( n3354 & n9198 ) | ( n7526 & n9198 ) ;
  assign n9195 = x72 & ~n6476 ;
  assign n9200 = n9199 ^ n9195 ^ 1'b0 ;
  assign n9192 = ( x180 & ~n1238 ) | ( x180 & n6288 ) | ( ~n1238 & n6288 ) ;
  assign n9190 = ( x87 & x194 ) | ( x87 & n7752 ) | ( x194 & n7752 ) ;
  assign n9191 = n9190 ^ n4526 ^ n3248 ;
  assign n9193 = n9192 ^ n9191 ^ n830 ;
  assign n9194 = n9193 ^ n7573 ^ n2179 ;
  assign n9201 = n9200 ^ n9194 ^ 1'b0 ;
  assign n9207 = n9206 ^ n9201 ^ n293 ;
  assign n9208 = ( n9188 & n9189 ) | ( n9188 & ~n9207 ) | ( n9189 & ~n9207 ) ;
  assign n9209 = n3159 ^ n3013 ^ x12 ;
  assign n9210 = ( n1580 & ~n2704 ) | ( n1580 & n9209 ) | ( ~n2704 & n9209 ) ;
  assign n9211 = ( n467 & ~n1484 ) | ( n467 & n9210 ) | ( ~n1484 & n9210 ) ;
  assign n9212 = ( n2752 & ~n7618 ) | ( n2752 & n9211 ) | ( ~n7618 & n9211 ) ;
  assign n9213 = n9212 ^ n7846 ^ n3668 ;
  assign n9214 = n9213 ^ n2403 ^ 1'b0 ;
  assign n9225 = ( ~n1182 & n2241 ) | ( ~n1182 & n3197 ) | ( n2241 & n3197 ) ;
  assign n9226 = n9225 ^ n2551 ^ n326 ;
  assign n9227 = ( n924 & ~n5047 ) | ( n924 & n9226 ) | ( ~n5047 & n9226 ) ;
  assign n9215 = ( n3883 & n7061 ) | ( n3883 & ~n7748 ) | ( n7061 & ~n7748 ) ;
  assign n9216 = x112 & ~n929 ;
  assign n9217 = ~n1722 & n9216 ;
  assign n9218 = n3164 ^ n2573 ^ x246 ;
  assign n9219 = n5603 ^ n4043 ^ n3692 ;
  assign n9220 = ( ~n5124 & n9218 ) | ( ~n5124 & n9219 ) | ( n9218 & n9219 ) ;
  assign n9221 = n9220 ^ n5285 ^ n3891 ;
  assign n9222 = ( n7622 & n9217 ) | ( n7622 & n9221 ) | ( n9217 & n9221 ) ;
  assign n9223 = ( n1255 & n9215 ) | ( n1255 & ~n9222 ) | ( n9215 & ~n9222 ) ;
  assign n9224 = ( ~n4407 & n6777 ) | ( ~n4407 & n9223 ) | ( n6777 & n9223 ) ;
  assign n9228 = n9227 ^ n9224 ^ n3929 ;
  assign n9229 = n6194 ^ n1962 ^ n1063 ;
  assign n9230 = n9229 ^ n5167 ^ 1'b0 ;
  assign n9231 = n9230 ^ n7158 ^ n2437 ;
  assign n9232 = n2997 ^ n863 ^ n717 ;
  assign n9233 = n8330 ^ n7932 ^ n7073 ;
  assign n9234 = n9233 ^ n5655 ^ n2353 ;
  assign n9235 = n9232 | n9234 ;
  assign n9236 = n9235 ^ n2861 ^ 1'b0 ;
  assign n9237 = ( n4863 & n6564 ) | ( n4863 & ~n9236 ) | ( n6564 & ~n9236 ) ;
  assign n9238 = n8674 ^ n5384 ^ n1622 ;
  assign n9239 = n3266 & n7154 ;
  assign n9240 = n9238 & n9239 ;
  assign n9241 = ~n2596 & n4903 ;
  assign n9242 = n9241 ^ n3415 ^ n1422 ;
  assign n9243 = n8578 & n9242 ;
  assign n9244 = n6932 & n9243 ;
  assign n9245 = n9244 ^ n3585 ^ n3214 ;
  assign n9246 = n9245 ^ n4216 ^ 1'b0 ;
  assign n9249 = ( n830 & n1671 ) | ( n830 & n6747 ) | ( n1671 & n6747 ) ;
  assign n9250 = ( n1731 & n5756 ) | ( n1731 & n6213 ) | ( n5756 & n6213 ) ;
  assign n9251 = n9250 ^ n4079 ^ n3950 ;
  assign n9252 = ( ~n290 & n9249 ) | ( ~n290 & n9251 ) | ( n9249 & n9251 ) ;
  assign n9247 = ~n1613 & n5923 ;
  assign n9248 = ~n3419 & n9247 ;
  assign n9253 = n9252 ^ n9248 ^ n318 ;
  assign n9268 = n8494 ^ n7603 ^ n4395 ;
  assign n9269 = n9268 ^ n8690 ^ x134 ;
  assign n9265 = ( x165 & n1570 ) | ( x165 & ~n2956 ) | ( n1570 & ~n2956 ) ;
  assign n9264 = x179 & n807 ;
  assign n9266 = n9265 ^ n9264 ^ 1'b0 ;
  assign n9256 = x15 & n1426 ;
  assign n9257 = ( n1350 & n1818 ) | ( n1350 & ~n9256 ) | ( n1818 & ~n9256 ) ;
  assign n9254 = ( x116 & n1777 ) | ( x116 & n5498 ) | ( n1777 & n5498 ) ;
  assign n9255 = ~n1262 & n9254 ;
  assign n9258 = n9257 ^ n9255 ^ 1'b0 ;
  assign n9259 = ( n1557 & n3748 ) | ( n1557 & n5701 ) | ( n3748 & n5701 ) ;
  assign n9260 = ( n464 & n5276 ) | ( n464 & n9259 ) | ( n5276 & n9259 ) ;
  assign n9261 = n5071 & n9260 ;
  assign n9262 = n1120 & ~n3713 ;
  assign n9263 = ( n9258 & n9261 ) | ( n9258 & ~n9262 ) | ( n9261 & ~n9262 ) ;
  assign n9267 = n9266 ^ n9263 ^ n7990 ;
  assign n9270 = n9269 ^ n9267 ^ n2627 ;
  assign n9271 = ( ~n1239 & n9253 ) | ( ~n1239 & n9270 ) | ( n9253 & n9270 ) ;
  assign n9272 = ( n365 & ~n3580 ) | ( n365 & n8732 ) | ( ~n3580 & n8732 ) ;
  assign n9273 = ( n2381 & n4647 ) | ( n2381 & ~n5833 ) | ( n4647 & ~n5833 ) ;
  assign n9274 = ( ~n500 & n2811 ) | ( ~n500 & n8775 ) | ( n2811 & n8775 ) ;
  assign n9275 = n6175 ^ n1760 ^ n303 ;
  assign n9276 = ( n8258 & ~n8849 ) | ( n8258 & n9275 ) | ( ~n8849 & n9275 ) ;
  assign n9291 = n2987 ^ n2393 ^ n1598 ;
  assign n9292 = n9291 ^ n7822 ^ 1'b0 ;
  assign n9293 = ~n548 & n9292 ;
  assign n9287 = ( n3103 & ~n3687 ) | ( n3103 & n6019 ) | ( ~n3687 & n6019 ) ;
  assign n9288 = ~n2218 & n9287 ;
  assign n9289 = n9288 ^ n4287 ^ 1'b0 ;
  assign n9277 = ( n711 & n5755 ) | ( n711 & ~n6640 ) | ( n5755 & ~n6640 ) ;
  assign n9278 = n6094 ^ n1021 ^ n751 ;
  assign n9279 = ( ~n823 & n1158 ) | ( ~n823 & n1365 ) | ( n1158 & n1365 ) ;
  assign n9280 = ( n2254 & n6041 ) | ( n2254 & n9279 ) | ( n6041 & n9279 ) ;
  assign n9281 = ( n1796 & ~n8749 ) | ( n1796 & n9280 ) | ( ~n8749 & n9280 ) ;
  assign n9282 = ( n5160 & n9278 ) | ( n5160 & n9281 ) | ( n9278 & n9281 ) ;
  assign n9283 = ( n8826 & ~n9277 ) | ( n8826 & n9282 ) | ( ~n9277 & n9282 ) ;
  assign n9284 = n9283 ^ n1633 ^ 1'b0 ;
  assign n9285 = n758 | n9284 ;
  assign n9286 = n6147 | n9285 ;
  assign n9290 = n9289 ^ n9286 ^ 1'b0 ;
  assign n9294 = n9293 ^ n9290 ^ n6551 ;
  assign n9296 = n4816 ^ n3883 ^ n781 ;
  assign n9295 = n6051 ^ n1426 ^ n1156 ;
  assign n9297 = n9296 ^ n9295 ^ n2690 ;
  assign n9298 = ( x111 & n666 ) | ( x111 & n3448 ) | ( n666 & n3448 ) ;
  assign n9299 = ( ~n2426 & n2633 ) | ( ~n2426 & n9298 ) | ( n2633 & n9298 ) ;
  assign n9300 = n2275 | n4905 ;
  assign n9301 = n9300 ^ n3326 ^ 1'b0 ;
  assign n9302 = n3719 & n6863 ;
  assign n9303 = n9301 & n9302 ;
  assign n9304 = ( ~n7736 & n9299 ) | ( ~n7736 & n9303 ) | ( n9299 & n9303 ) ;
  assign n9306 = n8161 ^ n7258 ^ n6803 ;
  assign n9305 = n1162 & n8508 ;
  assign n9307 = n9306 ^ n9305 ^ 1'b0 ;
  assign n9308 = n889 & n1776 ;
  assign n9309 = ( n3790 & n5511 ) | ( n3790 & n9308 ) | ( n5511 & n9308 ) ;
  assign n9310 = ( n2296 & n4545 ) | ( n2296 & n8546 ) | ( n4545 & n8546 ) ;
  assign n9311 = n7509 | n7532 ;
  assign n9312 = ( n1107 & n9310 ) | ( n1107 & n9311 ) | ( n9310 & n9311 ) ;
  assign n9313 = ( n1064 & n5863 ) | ( n1064 & n9277 ) | ( n5863 & n9277 ) ;
  assign n9314 = n2014 & ~n9038 ;
  assign n9320 = n6855 ^ n6646 ^ n2839 ;
  assign n9315 = ( ~n1221 & n2518 ) | ( ~n1221 & n5559 ) | ( n2518 & n5559 ) ;
  assign n9316 = ( n2159 & ~n4267 ) | ( n2159 & n9315 ) | ( ~n4267 & n9315 ) ;
  assign n9317 = n9316 ^ n7711 ^ n3387 ;
  assign n9318 = n9317 ^ n3854 ^ n2293 ;
  assign n9319 = ( n301 & ~n8505 ) | ( n301 & n9318 ) | ( ~n8505 & n9318 ) ;
  assign n9321 = n9320 ^ n9319 ^ n8495 ;
  assign n9322 = ( n552 & ~n4094 ) | ( n552 & n6011 ) | ( ~n4094 & n6011 ) ;
  assign n9323 = n9322 ^ n8183 ^ n533 ;
  assign n9324 = n1439 & ~n8011 ;
  assign n9325 = ( n1663 & n2618 ) | ( n1663 & n9324 ) | ( n2618 & n9324 ) ;
  assign n9326 = ( ~n487 & n2874 ) | ( ~n487 & n5581 ) | ( n2874 & n5581 ) ;
  assign n9327 = n872 & ~n6638 ;
  assign n9328 = n9327 ^ n5711 ^ n5170 ;
  assign n9329 = n9328 ^ n4566 ^ n4023 ;
  assign n9330 = n8083 | n9329 ;
  assign n9331 = n7284 | n9330 ;
  assign n9332 = ( ~x214 & n836 ) | ( ~x214 & n4526 ) | ( n836 & n4526 ) ;
  assign n9333 = n9332 ^ n8098 ^ n6634 ;
  assign n9334 = ( n310 & n6934 ) | ( n310 & n9333 ) | ( n6934 & n9333 ) ;
  assign n9335 = ( n814 & n1809 ) | ( n814 & ~n6776 ) | ( n1809 & ~n6776 ) ;
  assign n9336 = n7240 ^ n4932 ^ n1588 ;
  assign n9337 = ( n1098 & ~n9335 ) | ( n1098 & n9336 ) | ( ~n9335 & n9336 ) ;
  assign n9338 = ( n1510 & n9334 ) | ( n1510 & ~n9337 ) | ( n9334 & ~n9337 ) ;
  assign n9339 = ( n5403 & n9205 ) | ( n5403 & ~n9338 ) | ( n9205 & ~n9338 ) ;
  assign n9340 = n2218 ^ n365 ^ 1'b0 ;
  assign n9341 = ( n1267 & n6537 ) | ( n1267 & n9196 ) | ( n6537 & n9196 ) ;
  assign n9342 = ( n1521 & ~n5414 ) | ( n1521 & n9341 ) | ( ~n5414 & n9341 ) ;
  assign n9343 = n5283 ^ n1814 ^ x191 ;
  assign n9344 = n439 & n4594 ;
  assign n9345 = n781 | n9344 ;
  assign n9346 = n9343 | n9345 ;
  assign n9347 = ( n2855 & n6318 ) | ( n2855 & n8298 ) | ( n6318 & n8298 ) ;
  assign n9348 = ~n686 & n9347 ;
  assign n9349 = ~n4242 & n9348 ;
  assign n9350 = x210 & ~n2175 ;
  assign n9351 = ( x204 & n1564 ) | ( x204 & n8239 ) | ( n1564 & n8239 ) ;
  assign n9352 = ( n1107 & ~n9350 ) | ( n1107 & n9351 ) | ( ~n9350 & n9351 ) ;
  assign n9353 = n9352 ^ n1292 ^ 1'b0 ;
  assign n9354 = ( n9346 & ~n9349 ) | ( n9346 & n9353 ) | ( ~n9349 & n9353 ) ;
  assign n9359 = n3803 ^ n1891 ^ 1'b0 ;
  assign n9355 = n3486 ^ n1557 ^ x41 ;
  assign n9356 = n1730 & n3219 ;
  assign n9357 = n9356 ^ n1304 ^ 1'b0 ;
  assign n9358 = ( n277 & ~n9355 ) | ( n277 & n9357 ) | ( ~n9355 & n9357 ) ;
  assign n9360 = n9359 ^ n9358 ^ n491 ;
  assign n9362 = ( n1103 & n2046 ) | ( n1103 & n5930 ) | ( n2046 & n5930 ) ;
  assign n9361 = ( n2413 & n3118 ) | ( n2413 & ~n4440 ) | ( n3118 & ~n4440 ) ;
  assign n9363 = n9362 ^ n9361 ^ n2940 ;
  assign n9364 = ~n1678 & n2086 ;
  assign n9365 = ( n2317 & n3273 ) | ( n2317 & ~n9364 ) | ( n3273 & ~n9364 ) ;
  assign n9366 = n6335 ^ n3907 ^ n2799 ;
  assign n9367 = n5248 ^ n1532 ^ 1'b0 ;
  assign n9368 = n9366 & n9367 ;
  assign n9369 = ~n4604 & n5270 ;
  assign n9370 = n9368 & n9369 ;
  assign n9371 = ( x253 & ~n9365 ) | ( x253 & n9370 ) | ( ~n9365 & n9370 ) ;
  assign n9372 = n7335 ^ n823 ^ n773 ;
  assign n9373 = n6244 & ~n9372 ;
  assign n9374 = n9373 ^ n8980 ^ n3842 ;
  assign n9375 = n9374 ^ n2528 ^ n663 ;
  assign n9383 = n3731 | n4443 ;
  assign n9384 = n9383 ^ n2168 ^ n1187 ;
  assign n9376 = ~n6966 & n7745 ;
  assign n9377 = n1334 & n9376 ;
  assign n9378 = ( n1530 & n3374 ) | ( n1530 & n3573 ) | ( n3374 & n3573 ) ;
  assign n9379 = n9378 ^ n6172 ^ n1787 ;
  assign n9380 = ( n955 & n9377 ) | ( n955 & n9379 ) | ( n9377 & n9379 ) ;
  assign n9381 = ( n1624 & n3813 ) | ( n1624 & n8456 ) | ( n3813 & n8456 ) ;
  assign n9382 = ( n2042 & n9380 ) | ( n2042 & ~n9381 ) | ( n9380 & ~n9381 ) ;
  assign n9385 = n9384 ^ n9382 ^ n1338 ;
  assign n9386 = n2122 ^ n1886 ^ n904 ;
  assign n9387 = n950 & n4911 ;
  assign n9388 = ( n2920 & n9386 ) | ( n2920 & n9387 ) | ( n9386 & n9387 ) ;
  assign n9389 = n7112 ^ n1133 ^ n999 ;
  assign n9390 = ( n2117 & ~n7521 ) | ( n2117 & n9389 ) | ( ~n7521 & n9389 ) ;
  assign n9391 = ( ~n511 & n1418 ) | ( ~n511 & n3776 ) | ( n1418 & n3776 ) ;
  assign n9392 = ( ~n2012 & n6696 ) | ( ~n2012 & n9391 ) | ( n6696 & n9391 ) ;
  assign n9393 = ( n6025 & ~n9390 ) | ( n6025 & n9392 ) | ( ~n9390 & n9392 ) ;
  assign n9394 = n2340 ^ n2225 ^ n1207 ;
  assign n9395 = n5956 ^ n839 ^ 1'b0 ;
  assign n9396 = n9395 ^ n2314 ^ 1'b0 ;
  assign n9397 = n5426 & ~n9396 ;
  assign n9398 = n9397 ^ n8572 ^ n1701 ;
  assign n9399 = ( x190 & n3784 ) | ( x190 & n9398 ) | ( n3784 & n9398 ) ;
  assign n9400 = n4161 ^ n1814 ^ 1'b0 ;
  assign n9401 = n9399 & ~n9400 ;
  assign n9402 = ( n1612 & n9394 ) | ( n1612 & n9401 ) | ( n9394 & n9401 ) ;
  assign n9403 = n6202 | n7497 ;
  assign n9404 = n3713 | n9403 ;
  assign n9405 = ( ~n2230 & n6934 ) | ( ~n2230 & n9404 ) | ( n6934 & n9404 ) ;
  assign n9414 = ( ~n2570 & n7147 ) | ( ~n2570 & n9153 ) | ( n7147 & n9153 ) ;
  assign n9415 = ( ~n5045 & n6540 ) | ( ~n5045 & n9414 ) | ( n6540 & n9414 ) ;
  assign n9406 = ( x69 & n1433 ) | ( x69 & n2967 ) | ( n1433 & n2967 ) ;
  assign n9407 = n9406 ^ n8848 ^ n6375 ;
  assign n9408 = ( n517 & n2188 ) | ( n517 & ~n5581 ) | ( n2188 & ~n5581 ) ;
  assign n9409 = ( n933 & n5883 ) | ( n933 & n9408 ) | ( n5883 & n9408 ) ;
  assign n9410 = n9409 ^ n415 ^ 1'b0 ;
  assign n9411 = ( ~n8485 & n9407 ) | ( ~n8485 & n9410 ) | ( n9407 & n9410 ) ;
  assign n9412 = n7581 ^ n6037 ^ n3333 ;
  assign n9413 = n9411 & n9412 ;
  assign n9416 = n9415 ^ n9413 ^ 1'b0 ;
  assign n9417 = n9405 & ~n9416 ;
  assign n9418 = ~n6382 & n9417 ;
  assign n9419 = ( n3587 & ~n4688 ) | ( n3587 & n6574 ) | ( ~n4688 & n6574 ) ;
  assign n9422 = ( n1521 & n2237 ) | ( n1521 & n4452 ) | ( n2237 & n4452 ) ;
  assign n9421 = n3069 ^ n1432 ^ n1325 ;
  assign n9420 = ( n4986 & n8794 ) | ( n4986 & n8890 ) | ( n8794 & n8890 ) ;
  assign n9423 = n9422 ^ n9421 ^ n9420 ;
  assign n9424 = n9419 & n9423 ;
  assign n9425 = n9424 ^ n7416 ^ n1643 ;
  assign n9426 = n2025 ^ n1082 ^ 1'b0 ;
  assign n9427 = n7253 | n9426 ;
  assign n9428 = n9427 ^ n6951 ^ n5411 ;
  assign n9429 = n9428 ^ n3025 ^ n2250 ;
  assign n9430 = ( ~n1371 & n8690 ) | ( ~n1371 & n9429 ) | ( n8690 & n9429 ) ;
  assign n9431 = n9425 & ~n9430 ;
  assign n9432 = n6077 ^ n3510 ^ 1'b0 ;
  assign n9434 = n8876 ^ n1969 ^ n294 ;
  assign n9433 = ( n730 & ~n2084 ) | ( n730 & n9217 ) | ( ~n2084 & n9217 ) ;
  assign n9435 = n9434 ^ n9433 ^ n4176 ;
  assign n9436 = ~n9285 & n9435 ;
  assign n9437 = n9436 ^ n2063 ^ 1'b0 ;
  assign n9438 = n926 ^ n276 ^ 1'b0 ;
  assign n9439 = n9438 ^ n3433 ^ n1817 ;
  assign n9440 = ( n2332 & n6659 ) | ( n2332 & ~n7385 ) | ( n6659 & ~n7385 ) ;
  assign n9441 = ( n4445 & ~n6508 ) | ( n4445 & n9175 ) | ( ~n6508 & n9175 ) ;
  assign n9442 = n9441 ^ n3737 ^ x151 ;
  assign n9443 = ( n8357 & n9440 ) | ( n8357 & n9442 ) | ( n9440 & n9442 ) ;
  assign n9459 = ~n2105 & n8727 ;
  assign n9456 = n6021 ^ n6008 ^ 1'b0 ;
  assign n9457 = n2098 & n9456 ;
  assign n9458 = n9457 ^ n8112 ^ n953 ;
  assign n9460 = n9459 ^ n9458 ^ n7760 ;
  assign n9444 = n5499 ^ n345 ^ 1'b0 ;
  assign n9445 = n3201 ^ n489 ^ 1'b0 ;
  assign n9446 = n9445 ^ n371 ^ n281 ;
  assign n9447 = n9446 ^ n7163 ^ n4608 ;
  assign n9448 = ( n315 & ~n4091 ) | ( n315 & n6191 ) | ( ~n4091 & n6191 ) ;
  assign n9449 = ( ~n9444 & n9447 ) | ( ~n9444 & n9448 ) | ( n9447 & n9448 ) ;
  assign n9453 = n5222 ^ n5172 ^ n2845 ;
  assign n9450 = n6389 ^ n800 ^ 1'b0 ;
  assign n9451 = n1481 | n9450 ;
  assign n9452 = n1249 & ~n9451 ;
  assign n9454 = n9453 ^ n9452 ^ 1'b0 ;
  assign n9455 = ( ~x245 & n9449 ) | ( ~x245 & n9454 ) | ( n9449 & n9454 ) ;
  assign n9461 = n9460 ^ n9455 ^ 1'b0 ;
  assign n9465 = n4518 ^ n3888 ^ n957 ;
  assign n9466 = n9465 ^ n5008 ^ n4222 ;
  assign n9462 = ( ~x112 & x230 ) | ( ~x112 & n5499 ) | ( x230 & n5499 ) ;
  assign n9463 = ( ~n1880 & n4070 ) | ( ~n1880 & n9462 ) | ( n4070 & n9462 ) ;
  assign n9464 = ( n901 & n6335 ) | ( n901 & n9463 ) | ( n6335 & n9463 ) ;
  assign n9467 = n9466 ^ n9464 ^ n2507 ;
  assign n9468 = ( n470 & n1167 ) | ( n470 & n2530 ) | ( n1167 & n2530 ) ;
  assign n9469 = n8969 ^ n3213 ^ x229 ;
  assign n9470 = n4480 ^ n2796 ^ n547 ;
  assign n9471 = ( ~n2348 & n5366 ) | ( ~n2348 & n9470 ) | ( n5366 & n9470 ) ;
  assign n9472 = n7238 ^ n6976 ^ n5895 ;
  assign n9473 = ( ~n258 & n1320 ) | ( ~n258 & n9472 ) | ( n1320 & n9472 ) ;
  assign n9474 = n9473 ^ n2642 ^ 1'b0 ;
  assign n9475 = n9471 | n9474 ;
  assign n9476 = ( n7419 & ~n9469 ) | ( n7419 & n9475 ) | ( ~n9469 & n9475 ) ;
  assign n9477 = n6110 ^ n3416 ^ n1896 ;
  assign n9478 = n7817 & n8555 ;
  assign n9479 = n9477 & n9478 ;
  assign n9488 = ( ~n4617 & n5583 ) | ( ~n4617 & n9166 ) | ( n5583 & n9166 ) ;
  assign n9487 = n5090 ^ n4575 ^ x14 ;
  assign n9480 = n4229 ^ n1841 ^ n274 ;
  assign n9481 = ( n2198 & n2328 ) | ( n2198 & n8605 ) | ( n2328 & n8605 ) ;
  assign n9482 = n9481 ^ n3052 ^ n1695 ;
  assign n9483 = n4375 ^ n2272 ^ n1269 ;
  assign n9484 = ( n440 & n1056 ) | ( n440 & n9483 ) | ( n1056 & n9483 ) ;
  assign n9485 = ( n1290 & ~n9482 ) | ( n1290 & n9484 ) | ( ~n9482 & n9484 ) ;
  assign n9486 = ( n6494 & n9480 ) | ( n6494 & ~n9485 ) | ( n9480 & ~n9485 ) ;
  assign n9489 = n9488 ^ n9487 ^ n9486 ;
  assign n9490 = n9489 ^ n6871 ^ n3573 ;
  assign n9494 = n8795 ^ n2212 ^ n1278 ;
  assign n9491 = n2528 & ~n6269 ;
  assign n9492 = n9491 ^ n339 ^ 1'b0 ;
  assign n9493 = ( n1294 & ~n3482 ) | ( n1294 & n9492 ) | ( ~n3482 & n9492 ) ;
  assign n9495 = n9494 ^ n9493 ^ x165 ;
  assign n9496 = n3119 & n4332 ;
  assign n9498 = n3777 ^ n1240 ^ n792 ;
  assign n9499 = ( n1437 & n7441 ) | ( n1437 & n9498 ) | ( n7441 & n9498 ) ;
  assign n9500 = ( n1842 & ~n6867 ) | ( n1842 & n9499 ) | ( ~n6867 & n9499 ) ;
  assign n9497 = n6865 ^ n5288 ^ n1371 ;
  assign n9501 = n9500 ^ n9497 ^ n1468 ;
  assign n9502 = ( n263 & ~n6337 ) | ( n263 & n7142 ) | ( ~n6337 & n7142 ) ;
  assign n9503 = ( n9496 & n9501 ) | ( n9496 & n9502 ) | ( n9501 & n9502 ) ;
  assign n9504 = ( x75 & n1203 ) | ( x75 & ~n5499 ) | ( n1203 & ~n5499 ) ;
  assign n9505 = n9504 ^ n6532 ^ n593 ;
  assign n9506 = ( n1716 & n2225 ) | ( n1716 & ~n6451 ) | ( n2225 & ~n6451 ) ;
  assign n9507 = n6161 ^ n2003 ^ 1'b0 ;
  assign n9508 = ( n1643 & ~n3844 ) | ( n1643 & n6420 ) | ( ~n3844 & n6420 ) ;
  assign n9509 = ( n1752 & n1774 ) | ( n1752 & ~n9508 ) | ( n1774 & ~n9508 ) ;
  assign n9510 = ( n1394 & ~n9507 ) | ( n1394 & n9509 ) | ( ~n9507 & n9509 ) ;
  assign n9511 = ( ~x201 & n9506 ) | ( ~x201 & n9510 ) | ( n9506 & n9510 ) ;
  assign n9512 = ( n2890 & n3028 ) | ( n2890 & n3159 ) | ( n3028 & n3159 ) ;
  assign n9515 = n6356 ^ n1914 ^ n1656 ;
  assign n9513 = n8706 ^ n2464 ^ n1356 ;
  assign n9514 = ( n3547 & n4565 ) | ( n3547 & n9513 ) | ( n4565 & n9513 ) ;
  assign n9516 = n9515 ^ n9514 ^ n7165 ;
  assign n9517 = n6327 ^ n6323 ^ n3282 ;
  assign n9518 = ( n1362 & n2228 ) | ( n1362 & n3436 ) | ( n2228 & n3436 ) ;
  assign n9519 = ( ~n7037 & n9517 ) | ( ~n7037 & n9518 ) | ( n9517 & n9518 ) ;
  assign n9521 = n3749 ^ n3140 ^ n514 ;
  assign n9520 = n1682 ^ x29 ^ 1'b0 ;
  assign n9522 = n9521 ^ n9520 ^ 1'b0 ;
  assign n9523 = n9519 & ~n9522 ;
  assign n9524 = ( n1026 & ~n1535 ) | ( n1026 & n1662 ) | ( ~n1535 & n1662 ) ;
  assign n9525 = ( n1051 & ~n1914 ) | ( n1051 & n9524 ) | ( ~n1914 & n9524 ) ;
  assign n9526 = n9525 ^ x40 ^ 1'b0 ;
  assign n9527 = ~n9523 & n9526 ;
  assign n9528 = n9076 ^ n8011 ^ n2228 ;
  assign n9529 = n9528 ^ n2817 ^ 1'b0 ;
  assign n9530 = ( n1512 & n4094 ) | ( n1512 & n6838 ) | ( n4094 & n6838 ) ;
  assign n9531 = n9530 ^ n5501 ^ n5232 ;
  assign n9532 = n4288 ^ n306 ^ 1'b0 ;
  assign n9533 = n2771 | n9532 ;
  assign n9534 = n9533 ^ n4740 ^ n4643 ;
  assign n9542 = ( x177 & n2337 ) | ( x177 & ~n2847 ) | ( n2337 & ~n2847 ) ;
  assign n9543 = n3594 ^ n2583 ^ n1717 ;
  assign n9544 = ( n2688 & n9542 ) | ( n2688 & n9543 ) | ( n9542 & n9543 ) ;
  assign n9535 = n3474 ^ n3310 ^ n1109 ;
  assign n9537 = ( n772 & ~n2020 ) | ( n772 & n4308 ) | ( ~n2020 & n4308 ) ;
  assign n9536 = n5864 ^ n4725 ^ n4117 ;
  assign n9538 = n9537 ^ n9536 ^ n973 ;
  assign n9539 = ( ~n4237 & n8257 ) | ( ~n4237 & n9538 ) | ( n8257 & n9538 ) ;
  assign n9540 = n9539 ^ n4075 ^ 1'b0 ;
  assign n9541 = n9535 & ~n9540 ;
  assign n9545 = n9544 ^ n9541 ^ n2913 ;
  assign n9546 = n5760 ^ n5090 ^ x62 ;
  assign n9547 = n5865 & n9546 ;
  assign n9548 = n9547 ^ n2140 ^ 1'b0 ;
  assign n9550 = n7016 ^ n2813 ^ n621 ;
  assign n9549 = n3792 ^ n2683 ^ n2176 ;
  assign n9551 = n9550 ^ n9549 ^ n4764 ;
  assign n9552 = ( n2959 & n3945 ) | ( n2959 & ~n8712 ) | ( n3945 & ~n8712 ) ;
  assign n9553 = n3676 ^ n2036 ^ 1'b0 ;
  assign n9554 = n5361 | n9553 ;
  assign n9555 = ( n4382 & ~n5973 ) | ( n4382 & n9554 ) | ( ~n5973 & n9554 ) ;
  assign n9556 = n6966 ^ n333 ^ 1'b0 ;
  assign n9557 = ~n9555 & n9556 ;
  assign n9564 = n6608 ^ n3874 ^ n1515 ;
  assign n9565 = ( n4612 & ~n8709 ) | ( n4612 & n9564 ) | ( ~n8709 & n9564 ) ;
  assign n9558 = n3516 & ~n4903 ;
  assign n9559 = n2796 & n9558 ;
  assign n9560 = x153 & ~n3632 ;
  assign n9561 = ( n3957 & ~n9559 ) | ( n3957 & n9560 ) | ( ~n9559 & n9560 ) ;
  assign n9562 = n1670 & ~n9561 ;
  assign n9563 = n9562 ^ n4673 ^ 1'b0 ;
  assign n9566 = n9565 ^ n9563 ^ n4364 ;
  assign n9567 = ( ~x21 & n9557 ) | ( ~x21 & n9566 ) | ( n9557 & n9566 ) ;
  assign n9568 = ( n2277 & n4922 ) | ( n2277 & ~n7475 ) | ( n4922 & ~n7475 ) ;
  assign n9570 = n3294 ^ n1041 ^ n333 ;
  assign n9569 = ( n2728 & ~n3345 ) | ( n2728 & n7416 ) | ( ~n3345 & n7416 ) ;
  assign n9571 = n9570 ^ n9569 ^ 1'b0 ;
  assign n9572 = n7593 | n9571 ;
  assign n9573 = ( ~x48 & n1959 ) | ( ~x48 & n9572 ) | ( n1959 & n9572 ) ;
  assign n9574 = n9568 & n9573 ;
  assign n9575 = n9574 ^ n6929 ^ n3553 ;
  assign n9576 = ( ~n2098 & n2937 ) | ( ~n2098 & n6446 ) | ( n2937 & n6446 ) ;
  assign n9577 = n5763 ^ n3855 ^ n3819 ;
  assign n9578 = ( x12 & ~n3290 ) | ( x12 & n9577 ) | ( ~n3290 & n9577 ) ;
  assign n9579 = n9578 ^ n4238 ^ n3886 ;
  assign n9580 = ( n1828 & n9576 ) | ( n1828 & n9579 ) | ( n9576 & n9579 ) ;
  assign n9581 = n9580 ^ n9475 ^ n2247 ;
  assign n9582 = ( ~n6137 & n9575 ) | ( ~n6137 & n9581 ) | ( n9575 & n9581 ) ;
  assign n9585 = ( n4009 & ~n5422 ) | ( n4009 & n7745 ) | ( ~n5422 & n7745 ) ;
  assign n9586 = n6921 | n9585 ;
  assign n9587 = n9586 ^ n3681 ^ 1'b0 ;
  assign n9583 = n3836 | n4271 ;
  assign n9584 = n9583 ^ n1993 ^ 1'b0 ;
  assign n9588 = n9587 ^ n9584 ^ n5395 ;
  assign n9589 = n9588 ^ n8488 ^ n929 ;
  assign n9590 = n9070 ^ n7505 ^ n768 ;
  assign n9591 = n9590 ^ n1626 ^ n1317 ;
  assign n9592 = n9591 ^ n7055 ^ n6240 ;
  assign n9593 = n1953 ^ n511 ^ n398 ;
  assign n9594 = n9592 & ~n9593 ;
  assign n9595 = ( n3829 & ~n9589 ) | ( n3829 & n9594 ) | ( ~n9589 & n9594 ) ;
  assign n9596 = n2137 ^ n1546 ^ n1402 ;
  assign n9598 = n4357 ^ n1308 ^ 1'b0 ;
  assign n9597 = n6420 ^ n4472 ^ x241 ;
  assign n9599 = n9598 ^ n9597 ^ 1'b0 ;
  assign n9600 = ( n5576 & n9596 ) | ( n5576 & n9599 ) | ( n9596 & n9599 ) ;
  assign n9602 = n1654 | n7848 ;
  assign n9601 = ( n518 & n883 ) | ( n518 & ~n1576 ) | ( n883 & ~n1576 ) ;
  assign n9603 = n9602 ^ n9601 ^ n6859 ;
  assign n9604 = ( ~n5126 & n5312 ) | ( ~n5126 & n9603 ) | ( n5312 & n9603 ) ;
  assign n9605 = ( n613 & ~n6144 ) | ( n613 & n6805 ) | ( ~n6144 & n6805 ) ;
  assign n9606 = n6535 ^ n5030 ^ n4148 ;
  assign n9607 = ( ~n2346 & n5326 ) | ( ~n2346 & n9606 ) | ( n5326 & n9606 ) ;
  assign n9608 = ( n2603 & ~n7923 ) | ( n2603 & n9607 ) | ( ~n7923 & n9607 ) ;
  assign n9609 = ( ~n1211 & n5770 ) | ( ~n1211 & n9608 ) | ( n5770 & n9608 ) ;
  assign n9610 = n9605 & n9609 ;
  assign n9611 = ( ~n2656 & n9204 ) | ( ~n2656 & n9610 ) | ( n9204 & n9610 ) ;
  assign n9614 = n1276 ^ n1067 ^ n942 ;
  assign n9615 = n9614 ^ n4692 ^ n4644 ;
  assign n9612 = ~n5090 & n8698 ;
  assign n9613 = ~n8214 & n9612 ;
  assign n9616 = n9615 ^ n9613 ^ 1'b0 ;
  assign n9619 = n7014 ^ n5727 ^ n2945 ;
  assign n9617 = ( n437 & ~n5632 ) | ( n437 & n8006 ) | ( ~n5632 & n8006 ) ;
  assign n9618 = n9617 ^ n3086 ^ 1'b0 ;
  assign n9620 = n9619 ^ n9618 ^ n6831 ;
  assign n9627 = n9159 ^ n5245 ^ n893 ;
  assign n9628 = ( ~n546 & n3512 ) | ( ~n546 & n9627 ) | ( n3512 & n9627 ) ;
  assign n9629 = n9628 ^ n3049 ^ n2363 ;
  assign n9630 = ( n2483 & ~n7388 ) | ( n2483 & n9629 ) | ( ~n7388 & n9629 ) ;
  assign n9621 = n8768 ^ n2980 ^ n1358 ;
  assign n9622 = n3525 ^ n3273 ^ n1184 ;
  assign n9623 = n9622 ^ n3205 ^ 1'b0 ;
  assign n9624 = n9623 ^ n3178 ^ 1'b0 ;
  assign n9625 = ( n6681 & n9621 ) | ( n6681 & n9624 ) | ( n9621 & n9624 ) ;
  assign n9626 = ( n434 & ~n2397 ) | ( n434 & n9625 ) | ( ~n2397 & n9625 ) ;
  assign n9631 = n9630 ^ n9626 ^ 1'b0 ;
  assign n9650 = ( ~n1808 & n5615 ) | ( ~n1808 & n9513 ) | ( n5615 & n9513 ) ;
  assign n9635 = n3079 | n8782 ;
  assign n9632 = n4947 ^ n3074 ^ n1286 ;
  assign n9633 = n9632 ^ n3908 ^ n3755 ;
  assign n9634 = n9633 ^ n7702 ^ n4306 ;
  assign n9636 = n9635 ^ n9634 ^ n1613 ;
  assign n9637 = n1167 & n5766 ;
  assign n9638 = n9636 & n9637 ;
  assign n9642 = n3127 & n4892 ;
  assign n9643 = n4649 & n9642 ;
  assign n9644 = ( ~n2799 & n4922 ) | ( ~n2799 & n5800 ) | ( n4922 & n5800 ) ;
  assign n9645 = ( n5010 & n5177 ) | ( n5010 & n5704 ) | ( n5177 & n5704 ) ;
  assign n9646 = ( ~n3464 & n9644 ) | ( ~n3464 & n9645 ) | ( n9644 & n9645 ) ;
  assign n9647 = ( ~x51 & n9643 ) | ( ~x51 & n9646 ) | ( n9643 & n9646 ) ;
  assign n9639 = n9268 ^ n7208 ^ n1853 ;
  assign n9640 = n9639 ^ n5007 ^ n1498 ;
  assign n9641 = n9640 ^ n9279 ^ n3471 ;
  assign n9648 = n9647 ^ n9641 ^ 1'b0 ;
  assign n9649 = ~n9638 & n9648 ;
  assign n9651 = n9650 ^ n9649 ^ n8324 ;
  assign n9652 = n893 ^ n865 ^ n623 ;
  assign n9655 = ( n1312 & n2493 ) | ( n1312 & ~n2627 ) | ( n2493 & ~n2627 ) ;
  assign n9654 = n5391 ^ n1966 ^ 1'b0 ;
  assign n9656 = n9655 ^ n9654 ^ n4570 ;
  assign n9653 = n5121 | n6685 ;
  assign n9657 = n9656 ^ n9653 ^ 1'b0 ;
  assign n9658 = n1113 & ~n9657 ;
  assign n9659 = ( n8400 & n9652 ) | ( n8400 & n9658 ) | ( n9652 & n9658 ) ;
  assign n9660 = n6824 ^ n3191 ^ 1'b0 ;
  assign n9661 = n9659 & n9660 ;
  assign n9662 = n5249 ^ n4555 ^ n4446 ;
  assign n9663 = ( n3414 & ~n3622 ) | ( n3414 & n8141 ) | ( ~n3622 & n8141 ) ;
  assign n9664 = ( ~n2636 & n6186 ) | ( ~n2636 & n9663 ) | ( n6186 & n9663 ) ;
  assign n9665 = ( ~n2697 & n9662 ) | ( ~n2697 & n9664 ) | ( n9662 & n9664 ) ;
  assign n9666 = ~n1964 & n3293 ;
  assign n9667 = ~n4010 & n9666 ;
  assign n9668 = n5661 ^ n2271 ^ 1'b0 ;
  assign n9669 = n9668 ^ n7800 ^ n3002 ;
  assign n9670 = ( n4155 & n9667 ) | ( n4155 & n9669 ) | ( n9667 & n9669 ) ;
  assign n9671 = n9670 ^ n8970 ^ n8105 ;
  assign n9672 = n1209 & ~n2127 ;
  assign n9673 = n9672 ^ n9038 ^ 1'b0 ;
  assign n9674 = n9673 ^ n1217 ^ n268 ;
  assign n9675 = n7201 ^ n6748 ^ n4324 ;
  assign n9676 = ( n6352 & n9070 ) | ( n6352 & ~n9675 ) | ( n9070 & ~n9675 ) ;
  assign n9677 = n8495 ^ n7214 ^ n3807 ;
  assign n9678 = ( n4834 & ~n8041 ) | ( n4834 & n9677 ) | ( ~n8041 & n9677 ) ;
  assign n9686 = ( ~x217 & n8973 ) | ( ~x217 & n9346 ) | ( n8973 & n9346 ) ;
  assign n9687 = n6194 ^ n2851 ^ n780 ;
  assign n9688 = ( n4382 & n6576 ) | ( n4382 & n9076 ) | ( n6576 & n9076 ) ;
  assign n9689 = ( n3433 & n9687 ) | ( n3433 & ~n9688 ) | ( n9687 & ~n9688 ) ;
  assign n9690 = ( n915 & ~n9686 ) | ( n915 & n9689 ) | ( ~n9686 & n9689 ) ;
  assign n9679 = n8534 ^ n7553 ^ n3857 ;
  assign n9680 = n7722 ^ n5583 ^ n2813 ;
  assign n9681 = ( n3334 & n9679 ) | ( n3334 & n9680 ) | ( n9679 & n9680 ) ;
  assign n9682 = n6327 ^ n2398 ^ 1'b0 ;
  assign n9683 = ( n1506 & ~n2969 ) | ( n1506 & n4686 ) | ( ~n2969 & n4686 ) ;
  assign n9684 = n9682 | n9683 ;
  assign n9685 = n9681 | n9684 ;
  assign n9691 = n9690 ^ n9685 ^ n5734 ;
  assign n9692 = n525 ^ n489 ^ 1'b0 ;
  assign n9693 = ( n311 & ~n3424 ) | ( n311 & n5336 ) | ( ~n3424 & n5336 ) ;
  assign n9694 = n5193 & n9693 ;
  assign n9695 = ~n9692 & n9694 ;
  assign n9704 = ( n4234 & n4487 ) | ( n4234 & n5035 ) | ( n4487 & n5035 ) ;
  assign n9705 = n9704 ^ n6550 ^ 1'b0 ;
  assign n9706 = n4874 | n9705 ;
  assign n9707 = n5248 | n9706 ;
  assign n9699 = n7872 | n8669 ;
  assign n9700 = n1874 & ~n9699 ;
  assign n9701 = n9700 ^ n6650 ^ n2978 ;
  assign n9702 = ( ~n310 & n4817 ) | ( ~n310 & n5611 ) | ( n4817 & n5611 ) ;
  assign n9703 = ( n8844 & n9701 ) | ( n8844 & ~n9702 ) | ( n9701 & ~n9702 ) ;
  assign n9708 = n9707 ^ n9703 ^ n8122 ;
  assign n9714 = x154 & n5543 ;
  assign n9715 = n9714 ^ n7020 ^ 1'b0 ;
  assign n9716 = ( n2591 & ~n5314 ) | ( n2591 & n9715 ) | ( ~n5314 & n9715 ) ;
  assign n9717 = n9716 ^ n3458 ^ n2965 ;
  assign n9713 = ( ~n705 & n2757 ) | ( ~n705 & n6595 ) | ( n2757 & n6595 ) ;
  assign n9709 = n6256 & ~n6320 ;
  assign n9710 = ~x31 & n9709 ;
  assign n9711 = n9710 ^ n2984 ^ n2033 ;
  assign n9712 = n9711 ^ n8558 ^ n1838 ;
  assign n9718 = n9717 ^ n9713 ^ n9712 ;
  assign n9719 = n9718 ^ n5871 ^ n1178 ;
  assign n9720 = ( ~n4120 & n9708 ) | ( ~n4120 & n9719 ) | ( n9708 & n9719 ) ;
  assign n9721 = ( n4645 & ~n6876 ) | ( n4645 & n9720 ) | ( ~n6876 & n9720 ) ;
  assign n9696 = n3874 & ~n9279 ;
  assign n9697 = n9696 ^ n5571 ^ 1'b0 ;
  assign n9698 = x204 & n9697 ;
  assign n9722 = n9721 ^ n9698 ^ 1'b0 ;
  assign n9723 = ~n673 & n2184 ;
  assign n9724 = ( n370 & n1762 ) | ( n370 & n9723 ) | ( n1762 & n9723 ) ;
  assign n9725 = n9724 ^ n8030 ^ n7753 ;
  assign n9726 = ( n1512 & n5324 ) | ( n1512 & ~n7185 ) | ( n5324 & ~n7185 ) ;
  assign n9727 = n931 & ~n1531 ;
  assign n9728 = n9727 ^ n3080 ^ 1'b0 ;
  assign n9729 = n9728 ^ n7622 ^ n3129 ;
  assign n9730 = ( ~n591 & n2858 ) | ( ~n591 & n6307 ) | ( n2858 & n6307 ) ;
  assign n9731 = n9730 ^ n2583 ^ n1079 ;
  assign n9732 = ( ~n9726 & n9729 ) | ( ~n9726 & n9731 ) | ( n9729 & n9731 ) ;
  assign n9746 = ( ~n675 & n919 ) | ( ~n675 & n5889 ) | ( n919 & n5889 ) ;
  assign n9747 = ( n1283 & n1395 ) | ( n1283 & n3851 ) | ( n1395 & n3851 ) ;
  assign n9748 = ( n6056 & n9746 ) | ( n6056 & n9747 ) | ( n9746 & n9747 ) ;
  assign n9733 = ( n5633 & n6121 ) | ( n5633 & n7276 ) | ( n6121 & n7276 ) ;
  assign n9735 = n8336 | n8413 ;
  assign n9736 = n3003 & ~n9735 ;
  assign n9734 = n2492 | n4428 ;
  assign n9737 = n9736 ^ n9734 ^ 1'b0 ;
  assign n9738 = ( ~n5167 & n9733 ) | ( ~n5167 & n9737 ) | ( n9733 & n9737 ) ;
  assign n9741 = n7887 ^ n4914 ^ n875 ;
  assign n9739 = ( n1162 & n1537 ) | ( n1162 & n1738 ) | ( n1537 & n1738 ) ;
  assign n9740 = n9739 ^ n4141 ^ n1059 ;
  assign n9742 = n9741 ^ n9740 ^ n8984 ;
  assign n9743 = n9742 ^ n338 ^ 1'b0 ;
  assign n9744 = n7770 | n9743 ;
  assign n9745 = n9738 & ~n9744 ;
  assign n9749 = n9748 ^ n9745 ^ 1'b0 ;
  assign n9750 = n4959 ^ n4660 ^ n2803 ;
  assign n9751 = ( x16 & ~n1413 ) | ( x16 & n9750 ) | ( ~n1413 & n9750 ) ;
  assign n9752 = n8338 ^ n3450 ^ n2251 ;
  assign n9753 = ( ~n1829 & n3807 ) | ( ~n1829 & n9473 ) | ( n3807 & n9473 ) ;
  assign n9754 = ( n1795 & n9241 ) | ( n1795 & n9753 ) | ( n9241 & n9753 ) ;
  assign n9755 = n9754 ^ n6732 ^ 1'b0 ;
  assign n9756 = ( n7724 & ~n9752 ) | ( n7724 & n9755 ) | ( ~n9752 & n9755 ) ;
  assign n9757 = n5890 ^ n5309 ^ n3080 ;
  assign n9758 = ( n889 & ~n4370 ) | ( n889 & n9757 ) | ( ~n4370 & n9757 ) ;
  assign n9759 = n9758 ^ n2029 ^ 1'b0 ;
  assign n9760 = n9759 ^ n9166 ^ n4913 ;
  assign n9761 = n9760 ^ n4804 ^ n2473 ;
  assign n9762 = n3167 ^ n315 ^ x200 ;
  assign n9763 = ( n947 & n3222 ) | ( n947 & n7521 ) | ( n3222 & n7521 ) ;
  assign n9764 = n9763 ^ n4584 ^ n449 ;
  assign n9765 = n4375 ^ n3019 ^ 1'b0 ;
  assign n9766 = n3374 & n9765 ;
  assign n9767 = n9766 ^ n2097 ^ 1'b0 ;
  assign n9768 = ( n9762 & n9764 ) | ( n9762 & ~n9767 ) | ( n9764 & ~n9767 ) ;
  assign n9776 = n5662 ^ n2411 ^ 1'b0 ;
  assign n9775 = n2308 ^ n1404 ^ n865 ;
  assign n9777 = n9776 ^ n9775 ^ n4503 ;
  assign n9778 = n9777 ^ n5118 ^ n268 ;
  assign n9773 = ( n354 & n1896 ) | ( n354 & n2539 ) | ( n1896 & n2539 ) ;
  assign n9769 = n1502 | n3766 ;
  assign n9770 = n9769 ^ n4896 ^ 1'b0 ;
  assign n9771 = ( ~n515 & n840 ) | ( ~n515 & n9770 ) | ( n840 & n9770 ) ;
  assign n9772 = ( n2104 & n3264 ) | ( n2104 & n9771 ) | ( n3264 & n9771 ) ;
  assign n9774 = n9773 ^ n9772 ^ x37 ;
  assign n9779 = n9778 ^ n9774 ^ n2847 ;
  assign n9786 = ( n2058 & ~n2888 ) | ( n2058 & n7447 ) | ( ~n2888 & n7447 ) ;
  assign n9782 = ( n1777 & n1933 ) | ( n1777 & ~n5226 ) | ( n1933 & ~n5226 ) ;
  assign n9783 = ( n3960 & ~n5069 ) | ( n3960 & n9782 ) | ( ~n5069 & n9782 ) ;
  assign n9784 = n9783 ^ n3469 ^ 1'b0 ;
  assign n9785 = n9784 ^ n2986 ^ n2098 ;
  assign n9780 = n8256 ^ n3247 ^ n2552 ;
  assign n9781 = n9780 ^ n9475 ^ n7509 ;
  assign n9787 = n9786 ^ n9785 ^ n9781 ;
  assign n9788 = n7049 ^ n4867 ^ n3495 ;
  assign n9790 = ( n4085 & n4471 ) | ( n4085 & ~n8973 ) | ( n4471 & ~n8973 ) ;
  assign n9791 = n733 | n9790 ;
  assign n9792 = n9791 ^ n2541 ^ 1'b0 ;
  assign n9793 = n9792 ^ n7265 ^ n5559 ;
  assign n9789 = n7579 ^ n5593 ^ n3191 ;
  assign n9794 = n9793 ^ n9789 ^ 1'b0 ;
  assign n9802 = n2103 | n3837 ;
  assign n9803 = n7066 | n9802 ;
  assign n9798 = n2861 | n8785 ;
  assign n9799 = x91 | n9798 ;
  assign n9800 = n9799 ^ n6381 ^ n1567 ;
  assign n9801 = n9800 ^ n2750 ^ n1170 ;
  assign n9795 = n6801 ^ n5520 ^ n996 ;
  assign n9796 = ( ~x217 & n3621 ) | ( ~x217 & n9795 ) | ( n3621 & n9795 ) ;
  assign n9797 = ( n5918 & n6366 ) | ( n5918 & ~n9796 ) | ( n6366 & ~n9796 ) ;
  assign n9804 = n9803 ^ n9801 ^ n9797 ;
  assign n9818 = n9291 ^ n3514 ^ x241 ;
  assign n9819 = n9818 ^ n1475 ^ x93 ;
  assign n9815 = ( n496 & n3085 ) | ( n496 & ~n6038 ) | ( n3085 & ~n6038 ) ;
  assign n9816 = ( n1825 & ~n7352 ) | ( n1825 & n9815 ) | ( ~n7352 & n9815 ) ;
  assign n9811 = n7173 ^ n2436 ^ n2394 ;
  assign n9812 = n9811 ^ n5573 ^ n2715 ;
  assign n9813 = n9812 ^ n3147 ^ n706 ;
  assign n9814 = n4283 & ~n9813 ;
  assign n9817 = n9816 ^ n9814 ^ 1'b0 ;
  assign n9805 = ( n1033 & n1802 ) | ( n1033 & n1866 ) | ( n1802 & n1866 ) ;
  assign n9806 = ~n3376 & n9805 ;
  assign n9807 = ( ~n3197 & n3886 ) | ( ~n3197 & n9806 ) | ( n3886 & n9806 ) ;
  assign n9808 = ( n6748 & n7597 ) | ( n6748 & ~n9807 ) | ( n7597 & ~n9807 ) ;
  assign n9809 = ~n1009 & n6520 ;
  assign n9810 = ~n9808 & n9809 ;
  assign n9820 = n9819 ^ n9817 ^ n9810 ;
  assign n9821 = ( ~n2492 & n5763 ) | ( ~n2492 & n8222 ) | ( n5763 & n8222 ) ;
  assign n9822 = n9821 ^ n8626 ^ n7286 ;
  assign n9823 = n4889 ^ n3627 ^ n2492 ;
  assign n9825 = ( n701 & n1265 ) | ( n701 & n8113 ) | ( n1265 & n8113 ) ;
  assign n9826 = ( n1481 & ~n5667 ) | ( n1481 & n9825 ) | ( ~n5667 & n9825 ) ;
  assign n9824 = x71 & n7178 ;
  assign n9827 = n9826 ^ n9824 ^ 1'b0 ;
  assign n9828 = ( ~n9098 & n9823 ) | ( ~n9098 & n9827 ) | ( n9823 & n9827 ) ;
  assign n9834 = ( ~n1026 & n1618 ) | ( ~n1026 & n5586 ) | ( n1618 & n5586 ) ;
  assign n9835 = ( x149 & n3176 ) | ( x149 & ~n9834 ) | ( n3176 & ~n9834 ) ;
  assign n9829 = ( ~n763 & n2572 ) | ( ~n763 & n4126 ) | ( n2572 & n4126 ) ;
  assign n9830 = ~n1243 & n9829 ;
  assign n9831 = n9830 ^ n1469 ^ 1'b0 ;
  assign n9832 = ( ~n1868 & n6774 ) | ( ~n1868 & n9831 ) | ( n6774 & n9831 ) ;
  assign n9833 = ( n2634 & n9629 ) | ( n2634 & n9832 ) | ( n9629 & n9832 ) ;
  assign n9836 = n9835 ^ n9833 ^ n8223 ;
  assign n9837 = n2104 & ~n9836 ;
  assign n9838 = n5459 & ~n5750 ;
  assign n9839 = ~n8597 & n9838 ;
  assign n9851 = n814 | n2545 ;
  assign n9852 = n9851 ^ n1607 ^ 1'b0 ;
  assign n9850 = n5008 ^ n3464 ^ n2292 ;
  assign n9846 = ( x192 & n606 ) | ( x192 & n3594 ) | ( n606 & n3594 ) ;
  assign n9847 = n9846 ^ x174 ^ 1'b0 ;
  assign n9848 = n9847 ^ n5822 ^ 1'b0 ;
  assign n9844 = n4842 ^ n1506 ^ 1'b0 ;
  assign n9842 = n4855 ^ n1775 ^ 1'b0 ;
  assign n9843 = n1297 & ~n9842 ;
  assign n9840 = n5317 ^ n4521 ^ n2156 ;
  assign n9841 = ( ~n3701 & n6229 ) | ( ~n3701 & n9840 ) | ( n6229 & n9840 ) ;
  assign n9845 = n9844 ^ n9843 ^ n9841 ;
  assign n9849 = n9848 ^ n9845 ^ n3337 ;
  assign n9853 = n9852 ^ n9850 ^ n9849 ;
  assign n9854 = n1200 & ~n3727 ;
  assign n9855 = n9854 ^ n3829 ^ x70 ;
  assign n9856 = n9855 ^ n5615 ^ n2717 ;
  assign n9857 = n9856 ^ n5216 ^ n2828 ;
  assign n9858 = ( n7244 & n8036 ) | ( n7244 & ~n8974 ) | ( n8036 & ~n8974 ) ;
  assign n9859 = n9858 ^ n5203 ^ n2103 ;
  assign n9860 = ( n2575 & ~n6177 ) | ( n2575 & n6454 ) | ( ~n6177 & n6454 ) ;
  assign n9861 = n9860 ^ n7480 ^ x80 ;
  assign n9865 = ( n4147 & ~n5086 ) | ( n4147 & n5189 ) | ( ~n5086 & n5189 ) ;
  assign n9866 = n9865 ^ n3508 ^ n2421 ;
  assign n9867 = ( n2160 & n2309 ) | ( n2160 & ~n9866 ) | ( n2309 & ~n9866 ) ;
  assign n9868 = x74 | n9867 ;
  assign n9862 = n9597 ^ n8452 ^ n7822 ;
  assign n9863 = ( n489 & ~n2680 ) | ( n489 & n9862 ) | ( ~n2680 & n9862 ) ;
  assign n9864 = ( n6552 & n6780 ) | ( n6552 & n9863 ) | ( n6780 & n9863 ) ;
  assign n9869 = n9868 ^ n9864 ^ n6638 ;
  assign n9870 = ( ~n6750 & n8546 ) | ( ~n6750 & n9869 ) | ( n8546 & n9869 ) ;
  assign n9871 = ~n3242 & n9755 ;
  assign n9872 = ~n9870 & n9871 ;
  assign n9873 = ( n7469 & ~n9861 ) | ( n7469 & n9872 ) | ( ~n9861 & n9872 ) ;
  assign n9874 = x0 & n9873 ;
  assign n9877 = n7626 ^ n5897 ^ n3053 ;
  assign n9875 = n2732 ^ n1046 ^ 1'b0 ;
  assign n9876 = n7448 | n9875 ;
  assign n9878 = n9877 ^ n9876 ^ n4725 ;
  assign n9879 = n7685 ^ n2000 ^ n1231 ;
  assign n9883 = n6369 ^ n5283 ^ n2418 ;
  assign n9881 = ( ~x87 & n609 ) | ( ~x87 & n9776 ) | ( n609 & n9776 ) ;
  assign n9880 = n5822 ^ n3437 ^ n1810 ;
  assign n9882 = n9881 ^ n9880 ^ n5235 ;
  assign n9884 = n9883 ^ n9882 ^ n9797 ;
  assign n9885 = ( n6863 & n9879 ) | ( n6863 & n9884 ) | ( n9879 & n9884 ) ;
  assign n9893 = n3616 ^ n1136 ^ 1'b0 ;
  assign n9894 = n9893 ^ n9266 ^ n6373 ;
  assign n9895 = n9894 ^ n5691 ^ n2731 ;
  assign n9886 = n3279 ^ n2344 ^ n448 ;
  assign n9887 = n3810 | n4660 ;
  assign n9888 = n9886 | n9887 ;
  assign n9889 = n2475 & ~n9888 ;
  assign n9890 = n9889 ^ n1180 ^ 1'b0 ;
  assign n9891 = n6034 & n9890 ;
  assign n9892 = n9891 ^ n8407 ^ n7934 ;
  assign n9896 = n9895 ^ n9892 ^ n5110 ;
  assign n9897 = n7832 | n9896 ;
  assign n9898 = n2702 ^ n1700 ^ n710 ;
  assign n9899 = n9898 ^ n5185 ^ 1'b0 ;
  assign n9900 = n619 & n9899 ;
  assign n9901 = ( n1132 & ~n9897 ) | ( n1132 & n9900 ) | ( ~n9897 & n9900 ) ;
  assign n9902 = ( n4025 & ~n9885 ) | ( n4025 & n9901 ) | ( ~n9885 & n9901 ) ;
  assign n9903 = ~n7926 & n9855 ;
  assign n9904 = n9903 ^ n5090 ^ 1'b0 ;
  assign n9919 = ( n4429 & n4862 ) | ( n4429 & ~n8521 ) | ( n4862 & ~n8521 ) ;
  assign n9915 = ( n3743 & ~n4830 ) | ( n3743 & n4895 ) | ( ~n4830 & n4895 ) ;
  assign n9916 = n5900 | n9915 ;
  assign n9917 = n9916 ^ n6286 ^ 1'b0 ;
  assign n9918 = ( n5442 & n7703 ) | ( n5442 & n9917 ) | ( n7703 & n9917 ) ;
  assign n9920 = n9919 ^ n9918 ^ n2053 ;
  assign n9921 = n9920 ^ n4440 ^ n904 ;
  assign n9905 = n9268 ^ n8651 ^ n2986 ;
  assign n9906 = ~n413 & n5006 ;
  assign n9907 = n2480 & n9906 ;
  assign n9908 = n3515 | n6092 ;
  assign n9909 = n9908 ^ n6783 ^ 1'b0 ;
  assign n9910 = n9909 ^ n3245 ^ 1'b0 ;
  assign n9911 = n9907 | n9910 ;
  assign n9912 = ( n2344 & n9905 ) | ( n2344 & n9911 ) | ( n9905 & n9911 ) ;
  assign n9913 = ( n2724 & ~n8600 ) | ( n2724 & n9912 ) | ( ~n8600 & n9912 ) ;
  assign n9914 = ~n5148 & n9913 ;
  assign n9922 = n9921 ^ n9914 ^ 1'b0 ;
  assign n9923 = ( ~n3384 & n3560 ) | ( ~n3384 & n3827 ) | ( n3560 & n3827 ) ;
  assign n9928 = n5528 ^ n1477 ^ n629 ;
  assign n9927 = ( ~n2059 & n4948 ) | ( ~n2059 & n6768 ) | ( n4948 & n6768 ) ;
  assign n9925 = ( n1777 & n5512 ) | ( n1777 & ~n5624 ) | ( n5512 & ~n5624 ) ;
  assign n9924 = ~n4947 & n8085 ;
  assign n9926 = n9925 ^ n9924 ^ n8758 ;
  assign n9929 = n9928 ^ n9927 ^ n9926 ;
  assign n9930 = ( ~n1139 & n1762 ) | ( ~n1139 & n3168 ) | ( n1762 & n3168 ) ;
  assign n9931 = ( ~n565 & n2868 ) | ( ~n565 & n9930 ) | ( n2868 & n9930 ) ;
  assign n9932 = ( ~n2591 & n9099 ) | ( ~n2591 & n9931 ) | ( n9099 & n9931 ) ;
  assign n9933 = x25 & ~n1278 ;
  assign n9934 = n9933 ^ n2542 ^ 1'b0 ;
  assign n9935 = n9934 ^ n3225 ^ n2202 ;
  assign n9936 = ~n3680 & n7507 ;
  assign n9937 = n9935 & n9936 ;
  assign n9938 = n9932 & ~n9937 ;
  assign n9939 = n420 & n9938 ;
  assign n9940 = ( n9138 & ~n9555 ) | ( n9138 & n9939 ) | ( ~n9555 & n9939 ) ;
  assign n9941 = n3823 ^ n2957 ^ n1690 ;
  assign n9942 = n9941 ^ n1710 ^ n627 ;
  assign n9943 = n9942 ^ n4538 ^ n658 ;
  assign n9944 = n9940 & n9943 ;
  assign n9945 = ( ~n2969 & n6454 ) | ( ~n2969 & n9175 ) | ( n6454 & n9175 ) ;
  assign n9946 = ( n473 & ~n1989 ) | ( n473 & n4456 ) | ( ~n1989 & n4456 ) ;
  assign n9947 = n9946 ^ n2388 ^ 1'b0 ;
  assign n9963 = n5962 ^ n4404 ^ n3507 ;
  assign n9958 = ( n829 & n4121 ) | ( n829 & ~n4999 ) | ( n4121 & ~n4999 ) ;
  assign n9959 = n4802 ^ n3126 ^ n1134 ;
  assign n9960 = n9959 ^ n7505 ^ x245 ;
  assign n9961 = ( n3941 & ~n4282 ) | ( n3941 & n9960 ) | ( ~n4282 & n9960 ) ;
  assign n9962 = ( ~n2942 & n9958 ) | ( ~n2942 & n9961 ) | ( n9958 & n9961 ) ;
  assign n9964 = n9963 ^ n9962 ^ n2224 ;
  assign n9952 = n1590 ^ n964 ^ n519 ;
  assign n9953 = ~n4133 & n9952 ;
  assign n9948 = ( ~n3680 & n6581 ) | ( ~n3680 & n9250 ) | ( n6581 & n9250 ) ;
  assign n9949 = n9948 ^ n8116 ^ n6066 ;
  assign n9950 = ( n4377 & n7576 ) | ( n4377 & n9949 ) | ( n7576 & n9949 ) ;
  assign n9951 = ( n2656 & ~n7436 ) | ( n2656 & n9950 ) | ( ~n7436 & n9950 ) ;
  assign n9954 = n9953 ^ n9951 ^ n5558 ;
  assign n9955 = ( n3905 & n9746 ) | ( n3905 & n9954 ) | ( n9746 & n9954 ) ;
  assign n9956 = n9955 ^ n5608 ^ n491 ;
  assign n9957 = ~n6317 & n9956 ;
  assign n9965 = n9964 ^ n9957 ^ 1'b0 ;
  assign n9966 = ( n2861 & ~n3750 ) | ( n2861 & n6352 ) | ( ~n3750 & n6352 ) ;
  assign n9967 = n2706 & ~n9278 ;
  assign n9968 = n8208 & ~n9967 ;
  assign n9969 = n2234 & n9968 ;
  assign n9970 = ( ~n7511 & n9966 ) | ( ~n7511 & n9969 ) | ( n9966 & n9969 ) ;
  assign n9971 = n9970 ^ n8505 ^ n3153 ;
  assign n9972 = n927 & ~n2312 ;
  assign n9973 = ( n1551 & n9931 ) | ( n1551 & n9972 ) | ( n9931 & n9972 ) ;
  assign n9974 = n9973 ^ n7959 ^ n7248 ;
  assign n9975 = n9974 ^ n4145 ^ n3847 ;
  assign n9976 = n2634 | n2793 ;
  assign n9977 = n9976 ^ n9215 ^ 1'b0 ;
  assign n9979 = n1899 & n1977 ;
  assign n9980 = n9979 ^ n6396 ^ 1'b0 ;
  assign n9978 = ( n5647 & ~n6302 ) | ( n5647 & n9896 ) | ( ~n6302 & n9896 ) ;
  assign n9981 = n9980 ^ n9978 ^ n3630 ;
  assign n9982 = n9981 ^ n8055 ^ n5532 ;
  assign n9987 = n9457 ^ n814 ^ x51 ;
  assign n9988 = ( ~n1828 & n3094 ) | ( ~n1828 & n9987 ) | ( n3094 & n9987 ) ;
  assign n9983 = n4527 ^ n3964 ^ n2140 ;
  assign n9984 = ( n1725 & n3158 ) | ( n1725 & ~n4399 ) | ( n3158 & ~n4399 ) ;
  assign n9985 = n9984 ^ n4367 ^ n2188 ;
  assign n9986 = ( n974 & n9983 ) | ( n974 & n9985 ) | ( n9983 & n9985 ) ;
  assign n9989 = n9988 ^ n9986 ^ n2464 ;
  assign n9990 = ( n875 & ~n4220 ) | ( n875 & n8127 ) | ( ~n4220 & n8127 ) ;
  assign n9991 = n4536 ^ n3375 ^ n1910 ;
  assign n9992 = n3520 ^ n3103 ^ n777 ;
  assign n9993 = n8641 | n9992 ;
  assign n9994 = n9991 & ~n9993 ;
  assign n9999 = ( ~n3838 & n5135 ) | ( ~n3838 & n7567 ) | ( n5135 & n7567 ) ;
  assign n10000 = n2569 ^ x209 ^ 1'b0 ;
  assign n10001 = ~n9999 & n10000 ;
  assign n10002 = n6832 ^ n1064 ^ n1033 ;
  assign n10003 = ( n1786 & n10001 ) | ( n1786 & n10002 ) | ( n10001 & n10002 ) ;
  assign n9998 = n1909 ^ n1778 ^ n1238 ;
  assign n9995 = ~n2699 & n7824 ;
  assign n9996 = ( ~n3009 & n3018 ) | ( ~n3009 & n9995 ) | ( n3018 & n9995 ) ;
  assign n9997 = n9996 ^ n5647 ^ 1'b0 ;
  assign n10004 = n10003 ^ n9998 ^ n9997 ;
  assign n10005 = ( n3527 & n8448 ) | ( n3527 & ~n9525 ) | ( n8448 & ~n9525 ) ;
  assign n10006 = ( x147 & ~n9083 ) | ( x147 & n10005 ) | ( ~n9083 & n10005 ) ;
  assign n10012 = x37 & n3194 ;
  assign n10013 = ~n3866 & n10012 ;
  assign n10011 = n5953 ^ n2184 ^ n769 ;
  assign n10009 = ( n1624 & n4582 ) | ( n1624 & n4638 ) | ( n4582 & n4638 ) ;
  assign n10007 = n2990 | n6693 ;
  assign n10008 = x115 & ~n10007 ;
  assign n10010 = n10009 ^ n10008 ^ n4228 ;
  assign n10014 = n10013 ^ n10011 ^ n10010 ;
  assign n10015 = x141 & n1518 ;
  assign n10016 = n10015 ^ n8660 ^ 1'b0 ;
  assign n10017 = n10016 ^ n2697 ^ n2326 ;
  assign n10018 = ( n10006 & n10014 ) | ( n10006 & ~n10017 ) | ( n10014 & ~n10017 ) ;
  assign n10023 = ~n2675 & n3912 ;
  assign n10024 = n10023 ^ n6598 ^ 1'b0 ;
  assign n10022 = n2697 & n7262 ;
  assign n10020 = n7863 ^ n3793 ^ n2690 ;
  assign n10019 = n6040 ^ n2806 ^ n1188 ;
  assign n10021 = n10020 ^ n10019 ^ n5281 ;
  assign n10025 = n10024 ^ n10022 ^ n10021 ;
  assign n10026 = n10025 ^ n7652 ^ n4232 ;
  assign n10029 = n2078 ^ n1409 ^ 1'b0 ;
  assign n10030 = n3922 & ~n10029 ;
  assign n10027 = ~n1106 & n6952 ;
  assign n10028 = n10027 ^ n4488 ^ 1'b0 ;
  assign n10031 = n10030 ^ n10028 ^ n638 ;
  assign n10032 = ( n4120 & n5507 ) | ( n4120 & n10031 ) | ( n5507 & n10031 ) ;
  assign n10037 = n1119 & n6035 ;
  assign n10038 = n10037 ^ n3584 ^ 1'b0 ;
  assign n10033 = n8739 ^ n5611 ^ 1'b0 ;
  assign n10034 = n10033 ^ n6080 ^ n1226 ;
  assign n10035 = ( ~n1109 & n1345 ) | ( ~n1109 & n9995 ) | ( n1345 & n9995 ) ;
  assign n10036 = ( ~n6700 & n10034 ) | ( ~n6700 & n10035 ) | ( n10034 & n10035 ) ;
  assign n10039 = n10038 ^ n10036 ^ n8201 ;
  assign n10040 = ( n569 & n3503 ) | ( n569 & n10039 ) | ( n3503 & n10039 ) ;
  assign n10046 = ( ~n587 & n3744 ) | ( ~n587 & n5437 ) | ( n3744 & n5437 ) ;
  assign n10047 = n8260 & n10046 ;
  assign n10041 = n1990 & n2623 ;
  assign n10042 = n5417 & n10041 ;
  assign n10043 = ( n541 & n2299 ) | ( n541 & ~n10042 ) | ( n2299 & ~n10042 ) ;
  assign n10044 = ( n5804 & ~n9946 ) | ( n5804 & n10043 ) | ( ~n9946 & n10043 ) ;
  assign n10045 = n2641 & n10044 ;
  assign n10048 = n10047 ^ n10045 ^ 1'b0 ;
  assign n10049 = n4252 ^ n3635 ^ n2886 ;
  assign n10050 = n10049 ^ n9525 ^ n1347 ;
  assign n10051 = ~n4568 & n10050 ;
  assign n10052 = ~n4999 & n10051 ;
  assign n10053 = n7140 ^ n3816 ^ n2428 ;
  assign n10054 = ~n3407 & n8537 ;
  assign n10055 = n10054 ^ n2422 ^ n2277 ;
  assign n10056 = n8488 ^ n6127 ^ n2807 ;
  assign n10057 = n10056 ^ n9605 ^ n8515 ;
  assign n10058 = n2112 ^ n1132 ^ n1039 ;
  assign n10059 = ( ~n494 & n2265 ) | ( ~n494 & n3191 ) | ( n2265 & n3191 ) ;
  assign n10060 = ( ~x251 & n2867 ) | ( ~x251 & n10059 ) | ( n2867 & n10059 ) ;
  assign n10061 = n10058 & ~n10060 ;
  assign n10062 = ( n280 & n3305 ) | ( n280 & n5809 ) | ( n3305 & n5809 ) ;
  assign n10063 = n10062 ^ n4990 ^ n860 ;
  assign n10064 = n6915 ^ n4926 ^ 1'b0 ;
  assign n10065 = ~n1247 & n10064 ;
  assign n10066 = n10065 ^ n1806 ^ 1'b0 ;
  assign n10067 = n6158 & n10066 ;
  assign n10068 = ( n2267 & n10063 ) | ( n2267 & ~n10067 ) | ( n10063 & ~n10067 ) ;
  assign n10069 = n6768 ^ n685 ^ 1'b0 ;
  assign n10070 = n9821 ^ n7324 ^ n283 ;
  assign n10072 = n3090 ^ n1556 ^ 1'b0 ;
  assign n10071 = n8341 ^ n5090 ^ n2594 ;
  assign n10073 = n10072 ^ n10071 ^ n4940 ;
  assign n10074 = ( n3691 & ~n10070 ) | ( n3691 & n10073 ) | ( ~n10070 & n10073 ) ;
  assign n10083 = ( ~n524 & n1821 ) | ( ~n524 & n3317 ) | ( n1821 & n3317 ) ;
  assign n10081 = ( ~n3724 & n4082 ) | ( ~n3724 & n8412 ) | ( n4082 & n8412 ) ;
  assign n10082 = n10081 ^ n8857 ^ n5667 ;
  assign n10075 = n2775 ^ n2515 ^ n1613 ;
  assign n10076 = n10075 ^ n9559 ^ n4458 ;
  assign n10077 = n8473 ^ n3031 ^ n1322 ;
  assign n10078 = n10077 ^ n9022 ^ n2230 ;
  assign n10079 = n10078 ^ n9114 ^ n8057 ;
  assign n10080 = n10076 | n10079 ;
  assign n10084 = n10083 ^ n10082 ^ n10080 ;
  assign n10085 = ~n1587 & n6356 ;
  assign n10086 = n10085 ^ n3843 ^ 1'b0 ;
  assign n10095 = n4159 ^ n2429 ^ x162 ;
  assign n10096 = ( n739 & n1831 ) | ( n739 & ~n10095 ) | ( n1831 & ~n10095 ) ;
  assign n10097 = ( n579 & ~n715 ) | ( n579 & n10096 ) | ( ~n715 & n10096 ) ;
  assign n10098 = ( n2601 & ~n6395 ) | ( n2601 & n10097 ) | ( ~n6395 & n10097 ) ;
  assign n10094 = n9084 ^ n7196 ^ n6070 ;
  assign n10087 = n3942 ^ n3604 ^ x63 ;
  assign n10088 = ( ~n6245 & n8948 ) | ( ~n6245 & n10087 ) | ( n8948 & n10087 ) ;
  assign n10089 = ( n345 & n937 ) | ( n345 & n1470 ) | ( n937 & n1470 ) ;
  assign n10090 = n10089 ^ n6490 ^ 1'b0 ;
  assign n10091 = n2257 & n10090 ;
  assign n10092 = ~n10088 & n10091 ;
  assign n10093 = n10092 ^ n8035 ^ 1'b0 ;
  assign n10099 = n10098 ^ n10094 ^ n10093 ;
  assign n10100 = ( n7350 & n9606 ) | ( n7350 & ~n10099 ) | ( n9606 & ~n10099 ) ;
  assign n10116 = ( n1489 & n3772 ) | ( n1489 & ~n8277 ) | ( n3772 & ~n8277 ) ;
  assign n10104 = n3054 ^ n1225 ^ 1'b0 ;
  assign n10105 = n2117 | n10104 ;
  assign n10106 = n10105 ^ n5597 ^ n2036 ;
  assign n10107 = n6361 ^ n5386 ^ n3484 ;
  assign n10108 = ( ~n828 & n10106 ) | ( ~n828 & n10107 ) | ( n10106 & n10107 ) ;
  assign n10109 = n5461 ^ n2293 ^ 1'b0 ;
  assign n10110 = n2790 | n10109 ;
  assign n10111 = ( n820 & n3811 ) | ( n820 & ~n10110 ) | ( n3811 & ~n10110 ) ;
  assign n10112 = n10111 ^ n2401 ^ 1'b0 ;
  assign n10113 = n555 | n10112 ;
  assign n10114 = ( n3833 & ~n6321 ) | ( n3833 & n10113 ) | ( ~n6321 & n10113 ) ;
  assign n10115 = ( n5210 & n10108 ) | ( n5210 & ~n10114 ) | ( n10108 & ~n10114 ) ;
  assign n10101 = n3203 & n5422 ;
  assign n10102 = n10101 ^ n5843 ^ n1725 ;
  assign n10103 = n10102 ^ n4681 ^ n1195 ;
  assign n10117 = n10116 ^ n10115 ^ n10103 ;
  assign n10118 = ( n258 & ~n671 ) | ( n258 & n2867 ) | ( ~n671 & n2867 ) ;
  assign n10119 = n10118 ^ n2516 ^ n636 ;
  assign n10120 = ( ~n816 & n4893 ) | ( ~n816 & n10119 ) | ( n4893 & n10119 ) ;
  assign n10121 = n10120 ^ n5645 ^ n1567 ;
  assign n10122 = n10121 ^ n5379 ^ 1'b0 ;
  assign n10129 = n2100 ^ n1300 ^ n1099 ;
  assign n10130 = ( n5310 & n6122 ) | ( n5310 & ~n10129 ) | ( n6122 & ~n10129 ) ;
  assign n10131 = ( x82 & ~n8450 ) | ( x82 & n10130 ) | ( ~n8450 & n10130 ) ;
  assign n10133 = ( n1229 & n4855 ) | ( n1229 & n8534 ) | ( n4855 & n8534 ) ;
  assign n10132 = ( ~n812 & n2513 ) | ( ~n812 & n3710 ) | ( n2513 & n3710 ) ;
  assign n10134 = n10133 ^ n10132 ^ n6874 ;
  assign n10135 = n10134 ^ n5024 ^ n2963 ;
  assign n10136 = n9730 ^ n5605 ^ n1259 ;
  assign n10137 = ( n9885 & n10135 ) | ( n9885 & n10136 ) | ( n10135 & n10136 ) ;
  assign n10138 = n10131 | n10137 ;
  assign n10139 = n10138 ^ n6993 ^ 1'b0 ;
  assign n10124 = n9217 ^ n6415 ^ n442 ;
  assign n10125 = ~n1510 & n10124 ;
  assign n10126 = n3073 & n10125 ;
  assign n10123 = n5489 ^ n1219 ^ 1'b0 ;
  assign n10127 = n10126 ^ n10123 ^ n2385 ;
  assign n10128 = n3506 | n10127 ;
  assign n10140 = n10139 ^ n10128 ^ 1'b0 ;
  assign n10141 = ( n856 & ~n4048 ) | ( n856 & n10140 ) | ( ~n4048 & n10140 ) ;
  assign n10148 = n6238 ^ n2687 ^ 1'b0 ;
  assign n10149 = n10148 ^ n7128 ^ 1'b0 ;
  assign n10150 = n6318 & ~n10149 ;
  assign n10143 = ( n1495 & ~n1780 ) | ( n1495 & n4907 ) | ( ~n1780 & n4907 ) ;
  assign n10142 = n4458 ^ n2329 ^ 1'b0 ;
  assign n10144 = n10143 ^ n10142 ^ n1229 ;
  assign n10145 = ( n1108 & n2173 ) | ( n1108 & n10144 ) | ( n2173 & n10144 ) ;
  assign n10146 = n10145 ^ n3943 ^ n1464 ;
  assign n10147 = n10146 ^ n5914 ^ 1'b0 ;
  assign n10151 = n10150 ^ n10147 ^ n1008 ;
  assign n10152 = ( n1937 & n2102 ) | ( n1937 & n6580 ) | ( n2102 & n6580 ) ;
  assign n10153 = n8605 | n10152 ;
  assign n10172 = n6201 ^ n658 ^ 1'b0 ;
  assign n10173 = n8429 & n10172 ;
  assign n10170 = n6200 ^ n3185 ^ n655 ;
  assign n10158 = n3004 ^ n2231 ^ n1609 ;
  assign n10157 = n1944 & ~n7350 ;
  assign n10159 = n10158 ^ n10157 ^ 1'b0 ;
  assign n10160 = ( ~n5565 & n6010 ) | ( ~n5565 & n8426 ) | ( n6010 & n8426 ) ;
  assign n10166 = n7588 ^ n3294 ^ n3097 ;
  assign n10161 = n903 ^ n856 ^ n621 ;
  assign n10162 = ( n851 & ~n3201 ) | ( n851 & n10161 ) | ( ~n3201 & n10161 ) ;
  assign n10163 = n358 & n2305 ;
  assign n10164 = ( ~n3011 & n10162 ) | ( ~n3011 & n10163 ) | ( n10162 & n10163 ) ;
  assign n10165 = n10164 ^ n5938 ^ n3596 ;
  assign n10167 = n10166 ^ n10165 ^ n5709 ;
  assign n10168 = n10167 ^ n4687 ^ n379 ;
  assign n10169 = ( ~n10159 & n10160 ) | ( ~n10159 & n10168 ) | ( n10160 & n10168 ) ;
  assign n10154 = n7884 ^ n2147 ^ n1943 ;
  assign n10155 = n10154 ^ n2859 ^ n1161 ;
  assign n10156 = ( n7980 & n9961 ) | ( n7980 & ~n10155 ) | ( n9961 & ~n10155 ) ;
  assign n10171 = n10170 ^ n10169 ^ n10156 ;
  assign n10174 = n10173 ^ n10171 ^ n1171 ;
  assign n10175 = ( n578 & n2271 ) | ( n578 & ~n3107 ) | ( n2271 & ~n3107 ) ;
  assign n10176 = n9268 ^ n2084 ^ 1'b0 ;
  assign n10177 = n8005 | n10176 ;
  assign n10178 = ( n2913 & n10175 ) | ( n2913 & ~n10177 ) | ( n10175 & ~n10177 ) ;
  assign n10179 = ( n4915 & n8900 ) | ( n4915 & n10178 ) | ( n8900 & n10178 ) ;
  assign n10180 = ( ~n2991 & n10174 ) | ( ~n2991 & n10179 ) | ( n10174 & n10179 ) ;
  assign n10181 = ( x222 & ~n1130 ) | ( x222 & n6287 ) | ( ~n1130 & n6287 ) ;
  assign n10182 = ( ~n3234 & n5178 ) | ( ~n3234 & n9757 ) | ( n5178 & n9757 ) ;
  assign n10183 = ( n7846 & ~n10181 ) | ( n7846 & n10182 ) | ( ~n10181 & n10182 ) ;
  assign n10184 = n5762 & ~n9606 ;
  assign n10185 = n5040 & n10184 ;
  assign n10186 = ( n5458 & n5679 ) | ( n5458 & ~n8281 ) | ( n5679 & ~n8281 ) ;
  assign n10187 = ( n7545 & n10185 ) | ( n7545 & n10186 ) | ( n10185 & n10186 ) ;
  assign n10188 = ( ~n3841 & n10183 ) | ( ~n3841 & n10187 ) | ( n10183 & n10187 ) ;
  assign n10194 = n4732 ^ n2082 ^ 1'b0 ;
  assign n10189 = ( ~n631 & n1804 ) | ( ~n631 & n3031 ) | ( n1804 & n3031 ) ;
  assign n10190 = n3730 ^ n3043 ^ n1316 ;
  assign n10191 = ( n365 & n1425 ) | ( n365 & ~n10190 ) | ( n1425 & ~n10190 ) ;
  assign n10192 = ( n1211 & n10189 ) | ( n1211 & n10191 ) | ( n10189 & n10191 ) ;
  assign n10193 = n10192 ^ n8296 ^ n3307 ;
  assign n10195 = n10194 ^ n10193 ^ n9801 ;
  assign n10196 = ( ~n6529 & n10188 ) | ( ~n6529 & n10195 ) | ( n10188 & n10195 ) ;
  assign n10197 = n2422 | n4396 ;
  assign n10198 = ( n4344 & n9084 ) | ( n4344 & ~n10162 ) | ( n9084 & ~n10162 ) ;
  assign n10199 = ( n2019 & n10197 ) | ( n2019 & n10198 ) | ( n10197 & n10198 ) ;
  assign n10200 = n10199 ^ n6407 ^ n2713 ;
  assign n10201 = ( n3548 & n7117 ) | ( n3548 & ~n10200 ) | ( n7117 & ~n10200 ) ;
  assign n10205 = n6594 ^ n2984 ^ n1740 ;
  assign n10203 = ( n1758 & ~n3635 ) | ( n1758 & n6659 ) | ( ~n3635 & n6659 ) ;
  assign n10202 = ( ~n329 & n413 ) | ( ~n329 & n6137 ) | ( n413 & n6137 ) ;
  assign n10204 = n10203 ^ n10202 ^ n4679 ;
  assign n10206 = n10205 ^ n10204 ^ n5784 ;
  assign n10207 = n8938 ^ n8480 ^ n681 ;
  assign n10208 = n5329 ^ n3206 ^ 1'b0 ;
  assign n10209 = n1394 | n10208 ;
  assign n10210 = n10209 ^ n2745 ^ n866 ;
  assign n10211 = n10210 ^ n4356 ^ n2184 ;
  assign n10212 = ( ~n7236 & n10207 ) | ( ~n7236 & n10211 ) | ( n10207 & n10211 ) ;
  assign n10213 = n10212 ^ n3188 ^ n1891 ;
  assign n10214 = n400 & ~n681 ;
  assign n10215 = n10214 ^ n4502 ^ 1'b0 ;
  assign n10216 = n10215 ^ n3742 ^ n1595 ;
  assign n10217 = ( ~n1058 & n2252 ) | ( ~n1058 & n10216 ) | ( n2252 & n10216 ) ;
  assign n10218 = ( n1906 & ~n1935 ) | ( n1906 & n2151 ) | ( ~n1935 & n2151 ) ;
  assign n10219 = n10218 ^ n8430 ^ n3651 ;
  assign n10220 = ( n1665 & n2849 ) | ( n1665 & n10219 ) | ( n2849 & n10219 ) ;
  assign n10227 = ( x151 & n1755 ) | ( x151 & ~n3106 ) | ( n1755 & ~n3106 ) ;
  assign n10221 = ~n1971 & n9525 ;
  assign n10223 = n2481 ^ n996 ^ n701 ;
  assign n10224 = ( x38 & ~n1842 ) | ( x38 & n10223 ) | ( ~n1842 & n10223 ) ;
  assign n10222 = ( x250 & n4445 ) | ( x250 & ~n4833 ) | ( n4445 & ~n4833 ) ;
  assign n10225 = n10224 ^ n10222 ^ n7060 ;
  assign n10226 = ( n5695 & ~n10221 ) | ( n5695 & n10225 ) | ( ~n10221 & n10225 ) ;
  assign n10228 = n10227 ^ n10226 ^ n8876 ;
  assign n10229 = n10220 & n10228 ;
  assign n10230 = n10229 ^ n7156 ^ 1'b0 ;
  assign n10231 = n5710 & n10230 ;
  assign n10232 = ~n10217 & n10231 ;
  assign n10233 = n4911 ^ n2720 ^ 1'b0 ;
  assign n10234 = ( n3228 & n10071 ) | ( n3228 & ~n10233 ) | ( n10071 & ~n10233 ) ;
  assign n10235 = n4861 ^ n1188 ^ 1'b0 ;
  assign n10236 = n840 & n10235 ;
  assign n10237 = n9647 ^ n9142 ^ n1242 ;
  assign n10238 = ( n8821 & n10236 ) | ( n8821 & ~n10237 ) | ( n10236 & ~n10237 ) ;
  assign n10242 = n6197 ^ n6087 ^ n500 ;
  assign n10239 = n8964 ^ n5757 ^ n4213 ;
  assign n10240 = n2688 | n10239 ;
  assign n10241 = n10240 ^ n272 ^ 1'b0 ;
  assign n10243 = n10242 ^ n10241 ^ 1'b0 ;
  assign n10244 = ~n9088 & n10243 ;
  assign n10245 = ( n536 & n6359 ) | ( n536 & n10244 ) | ( n6359 & n10244 ) ;
  assign n10256 = n10226 ^ n3335 ^ n1147 ;
  assign n10257 = ( n5082 & n5742 ) | ( n5082 & ~n10256 ) | ( n5742 & ~n10256 ) ;
  assign n10255 = ( n2385 & n5444 ) | ( n2385 & n8971 ) | ( n5444 & n8971 ) ;
  assign n10258 = n10257 ^ n10255 ^ n5788 ;
  assign n10251 = n2606 ^ n2584 ^ n2006 ;
  assign n10247 = ( ~n903 & n1157 ) | ( ~n903 & n3432 ) | ( n1157 & n3432 ) ;
  assign n10246 = n8057 ^ n1796 ^ 1'b0 ;
  assign n10248 = n10247 ^ n10246 ^ n1830 ;
  assign n10249 = n10248 ^ n661 ^ x64 ;
  assign n10250 = n10249 ^ n1427 ^ n567 ;
  assign n10252 = n10251 ^ n10250 ^ n954 ;
  assign n10253 = ~n6720 & n10252 ;
  assign n10254 = n9961 | n10253 ;
  assign n10259 = n10258 ^ n10254 ^ 1'b0 ;
  assign n10260 = ( ~n1219 & n3980 ) | ( ~n1219 & n4713 ) | ( n3980 & n4713 ) ;
  assign n10261 = n10260 ^ n3443 ^ 1'b0 ;
  assign n10276 = x99 & n4404 ;
  assign n10277 = ~n403 & n10276 ;
  assign n10274 = n2994 ^ x237 ^ 1'b0 ;
  assign n10275 = n2063 & ~n10274 ;
  assign n10278 = n10277 ^ n10275 ^ n5736 ;
  assign n10271 = n903 & ~n1492 ;
  assign n10263 = x171 ^ x33 ^ 1'b0 ;
  assign n10270 = n5226 | n10263 ;
  assign n10272 = n10271 ^ n10270 ^ 1'b0 ;
  assign n10269 = n8366 ^ n3992 ^ n3640 ;
  assign n10262 = n2981 ^ n1001 ^ n300 ;
  assign n10264 = ( n1681 & ~n7090 ) | ( n1681 & n10263 ) | ( ~n7090 & n10263 ) ;
  assign n10265 = ~n5216 & n6883 ;
  assign n10266 = ~n9260 & n10265 ;
  assign n10267 = n10264 | n10266 ;
  assign n10268 = ( n1562 & ~n10262 ) | ( n1562 & n10267 ) | ( ~n10262 & n10267 ) ;
  assign n10273 = n10272 ^ n10269 ^ n10268 ;
  assign n10279 = n10278 ^ n10273 ^ n7749 ;
  assign n10281 = ( n1210 & n2767 ) | ( n1210 & n8131 ) | ( n2767 & n8131 ) ;
  assign n10282 = n10281 ^ n337 ^ 1'b0 ;
  assign n10280 = n7787 ^ n5768 ^ n5429 ;
  assign n10283 = n10282 ^ n10280 ^ 1'b0 ;
  assign n10284 = n5781 & n10283 ;
  assign n10285 = n9615 ^ n5397 ^ n448 ;
  assign n10286 = n4341 ^ n3525 ^ n682 ;
  assign n10287 = n10286 ^ n5259 ^ n3242 ;
  assign n10288 = ( n4709 & ~n10285 ) | ( n4709 & n10287 ) | ( ~n10285 & n10287 ) ;
  assign n10295 = n2447 ^ n2402 ^ n288 ;
  assign n10296 = ( n1838 & n6176 ) | ( n1838 & n10295 ) | ( n6176 & n10295 ) ;
  assign n10291 = n8857 ^ n4293 ^ n2385 ;
  assign n10292 = n10291 ^ n5993 ^ n5864 ;
  assign n10293 = ( ~n4070 & n9805 ) | ( ~n4070 & n10292 ) | ( n9805 & n10292 ) ;
  assign n10289 = n6195 ^ n5413 ^ n4039 ;
  assign n10290 = ( n411 & ~n1065 ) | ( n411 & n10289 ) | ( ~n1065 & n10289 ) ;
  assign n10294 = n10293 ^ n10290 ^ n9708 ;
  assign n10297 = n10296 ^ n10294 ^ n6254 ;
  assign n10298 = ( n2096 & n5196 ) | ( n2096 & ~n5286 ) | ( n5196 & ~n5286 ) ;
  assign n10299 = n10298 ^ n358 ^ 1'b0 ;
  assign n10301 = n5452 ^ n4113 ^ x214 ;
  assign n10300 = n9733 ^ n2214 ^ n632 ;
  assign n10302 = n10301 ^ n10300 ^ n7164 ;
  assign n10303 = n10302 ^ n6348 ^ n2237 ;
  assign n10317 = n5176 | n8500 ;
  assign n10318 = n10317 ^ n5964 ^ 1'b0 ;
  assign n10314 = n7253 ^ n4376 ^ n4038 ;
  assign n10315 = n10314 ^ n5401 ^ n554 ;
  assign n10316 = ( n540 & n1942 ) | ( n540 & n10315 ) | ( n1942 & n10315 ) ;
  assign n10319 = n10318 ^ n10316 ^ n9040 ;
  assign n10310 = n3346 ^ n1535 ^ 1'b0 ;
  assign n10311 = n10310 ^ n3751 ^ n1767 ;
  assign n10312 = n10311 ^ n2068 ^ x233 ;
  assign n10313 = n10312 ^ n6686 ^ n1928 ;
  assign n10320 = n10319 ^ n10313 ^ n4587 ;
  assign n10306 = ( n356 & ~n1812 ) | ( n356 & n4774 ) | ( ~n1812 & n4774 ) ;
  assign n10304 = ( n400 & n1212 ) | ( n400 & n2704 ) | ( n1212 & n2704 ) ;
  assign n10305 = n10304 ^ n7625 ^ n3515 ;
  assign n10307 = n10306 ^ n10305 ^ 1'b0 ;
  assign n10308 = ( n1171 & n8846 ) | ( n1171 & n10307 ) | ( n8846 & n10307 ) ;
  assign n10309 = ( n1389 & n1563 ) | ( n1389 & n10308 ) | ( n1563 & n10308 ) ;
  assign n10321 = n10320 ^ n10309 ^ n8052 ;
  assign n10323 = ( ~x162 & n2258 ) | ( ~x162 & n3194 ) | ( n2258 & n3194 ) ;
  assign n10322 = n9159 ^ n4520 ^ n3105 ;
  assign n10324 = n10323 ^ n10322 ^ n3057 ;
  assign n10329 = ( n1031 & ~n2803 ) | ( n1031 & n10030 ) | ( ~n2803 & n10030 ) ;
  assign n10330 = ( ~n561 & n6801 ) | ( ~n561 & n10329 ) | ( n6801 & n10329 ) ;
  assign n10325 = ~n1149 & n1156 ;
  assign n10326 = n10325 ^ n6396 ^ 1'b0 ;
  assign n10327 = n2255 ^ n2099 ^ n1356 ;
  assign n10328 = ( n4482 & ~n10326 ) | ( n4482 & n10327 ) | ( ~n10326 & n10327 ) ;
  assign n10331 = n10330 ^ n10328 ^ 1'b0 ;
  assign n10332 = n10331 ^ n8125 ^ n5039 ;
  assign n10333 = n5749 ^ n5194 ^ n1197 ;
  assign n10338 = n3900 ^ n3172 ^ n865 ;
  assign n10339 = ( n738 & n5459 ) | ( n738 & n10338 ) | ( n5459 & n10338 ) ;
  assign n10335 = n3703 ^ n1974 ^ n451 ;
  assign n10334 = n9654 ^ n875 ^ n629 ;
  assign n10336 = n10335 ^ n10334 ^ 1'b0 ;
  assign n10337 = n7313 & n10336 ;
  assign n10340 = n10339 ^ n10337 ^ n3005 ;
  assign n10341 = ( n992 & ~n2806 ) | ( n992 & n4760 ) | ( ~n2806 & n4760 ) ;
  assign n10342 = n10341 ^ n291 ^ 1'b0 ;
  assign n10344 = n4693 ^ n2758 ^ 1'b0 ;
  assign n10345 = n1880 & ~n10344 ;
  assign n10346 = ( x65 & n3115 ) | ( x65 & ~n10345 ) | ( n3115 & ~n10345 ) ;
  assign n10347 = ( ~n3790 & n7475 ) | ( ~n3790 & n10346 ) | ( n7475 & n10346 ) ;
  assign n10343 = n4470 & n8949 ;
  assign n10348 = n10347 ^ n10343 ^ 1'b0 ;
  assign n10349 = n3342 ^ n2292 ^ 1'b0 ;
  assign n10350 = ~n6180 & n10349 ;
  assign n10351 = ~n10348 & n10350 ;
  assign n10352 = n10351 ^ n1452 ^ 1'b0 ;
  assign n10353 = n10352 ^ n3885 ^ 1'b0 ;
  assign n10357 = n1986 ^ n1047 ^ n724 ;
  assign n10354 = n9496 ^ n9179 ^ n6996 ;
  assign n10355 = ( n3865 & ~n7799 ) | ( n3865 & n8753 ) | ( ~n7799 & n8753 ) ;
  assign n10356 = n10354 | n10355 ;
  assign n10358 = n10357 ^ n10356 ^ 1'b0 ;
  assign n10359 = n10358 ^ n9006 ^ n6056 ;
  assign n10360 = ~n1125 & n1829 ;
  assign n10361 = ~n3620 & n10360 ;
  assign n10362 = n9577 | n10361 ;
  assign n10363 = n1841 & ~n10362 ;
  assign n10364 = n4611 ^ n3670 ^ n1347 ;
  assign n10365 = n3947 & n8330 ;
  assign n10366 = ~n10364 & n10365 ;
  assign n10367 = n10366 ^ n7565 ^ n1259 ;
  assign n10368 = ( n4166 & n4971 ) | ( n4166 & ~n10367 ) | ( n4971 & ~n10367 ) ;
  assign n10369 = ( n1278 & n10363 ) | ( n1278 & ~n10368 ) | ( n10363 & ~n10368 ) ;
  assign n10370 = n4924 ^ n3878 ^ n1187 ;
  assign n10371 = n10370 ^ n7193 ^ 1'b0 ;
  assign n10372 = ~n9577 & n10371 ;
  assign n10373 = n10372 ^ n10298 ^ n8943 ;
  assign n10374 = n1686 | n8298 ;
  assign n10375 = n1497 | n10374 ;
  assign n10376 = n4078 | n10375 ;
  assign n10377 = n4009 ^ n3192 ^ 1'b0 ;
  assign n10378 = n10377 ^ n8693 ^ n8291 ;
  assign n10380 = ( n2399 & n3975 ) | ( n2399 & n5725 ) | ( n3975 & n5725 ) ;
  assign n10379 = n1844 ^ n1835 ^ n633 ;
  assign n10381 = n10380 ^ n10379 ^ 1'b0 ;
  assign n10382 = ~n4761 & n10381 ;
  assign n10383 = ( n8623 & ~n10378 ) | ( n8623 & n10382 ) | ( ~n10378 & n10382 ) ;
  assign n10384 = n2738 | n3542 ;
  assign n10385 = n4185 & ~n10384 ;
  assign n10386 = ( x83 & n1239 ) | ( x83 & n1243 ) | ( n1239 & n1243 ) ;
  assign n10387 = ( n1288 & n1943 ) | ( n1288 & n10386 ) | ( n1943 & n10386 ) ;
  assign n10389 = n6557 ^ n4765 ^ n3022 ;
  assign n10390 = ( n828 & n2122 ) | ( n828 & ~n10389 ) | ( n2122 & ~n10389 ) ;
  assign n10388 = n3580 | n6504 ;
  assign n10391 = n10390 ^ n10388 ^ 1'b0 ;
  assign n10392 = ( n906 & n9818 ) | ( n906 & ~n10391 ) | ( n9818 & ~n10391 ) ;
  assign n10393 = ( n1781 & n6528 ) | ( n1781 & ~n10392 ) | ( n6528 & ~n10392 ) ;
  assign n10395 = n6462 ^ n3930 ^ n2456 ;
  assign n10396 = n10395 ^ n4522 ^ n2829 ;
  assign n10394 = n5319 ^ n4099 ^ n2448 ;
  assign n10397 = n10396 ^ n10394 ^ n8141 ;
  assign n10398 = n10397 ^ n8842 ^ n6514 ;
  assign n10404 = ( n5053 & n5073 ) | ( n5053 & n6857 ) | ( n5073 & n6857 ) ;
  assign n10399 = n2963 ^ n2680 ^ n1905 ;
  assign n10400 = n7496 ^ n5203 ^ n3764 ;
  assign n10401 = ( n374 & ~n10399 ) | ( n374 & n10400 ) | ( ~n10399 & n10400 ) ;
  assign n10402 = ( n1231 & ~n7640 ) | ( n1231 & n10401 ) | ( ~n7640 & n10401 ) ;
  assign n10403 = n10402 ^ n4686 ^ n3490 ;
  assign n10405 = n10404 ^ n10403 ^ n5574 ;
  assign n10406 = n10405 ^ n8256 ^ n6900 ;
  assign n10407 = n7573 ^ n6454 ^ n2265 ;
  assign n10408 = ( n654 & ~n6079 ) | ( n654 & n10407 ) | ( ~n6079 & n10407 ) ;
  assign n10409 = n272 & ~n10408 ;
  assign n10411 = n6555 ^ n3372 ^ n2287 ;
  assign n10410 = ( n2541 & n5984 ) | ( n2541 & ~n10322 ) | ( n5984 & ~n10322 ) ;
  assign n10412 = n10411 ^ n10410 ^ 1'b0 ;
  assign n10413 = n5428 & ~n10412 ;
  assign n10414 = n3117 ^ n842 ^ 1'b0 ;
  assign n10415 = x230 & n10414 ;
  assign n10421 = ( n350 & ~n1651 ) | ( n350 & n5745 ) | ( ~n1651 & n5745 ) ;
  assign n10416 = n8803 ^ n638 ^ 1'b0 ;
  assign n10418 = n8113 ^ n2768 ^ n1030 ;
  assign n10417 = n4366 & ~n8170 ;
  assign n10419 = n10418 ^ n10417 ^ 1'b0 ;
  assign n10420 = ( ~n338 & n10416 ) | ( ~n338 & n10419 ) | ( n10416 & n10419 ) ;
  assign n10422 = n10421 ^ n10420 ^ n541 ;
  assign n10423 = ( ~n9269 & n10415 ) | ( ~n9269 & n10422 ) | ( n10415 & n10422 ) ;
  assign n10424 = n6313 ^ n5388 ^ n4736 ;
  assign n10425 = ( n3836 & n8817 ) | ( n3836 & ~n10424 ) | ( n8817 & ~n10424 ) ;
  assign n10426 = ( n655 & n1789 ) | ( n655 & n2786 ) | ( n1789 & n2786 ) ;
  assign n10427 = n10426 ^ n2695 ^ 1'b0 ;
  assign n10428 = n2942 & ~n10427 ;
  assign n10429 = ( n823 & ~n8473 ) | ( n823 & n10428 ) | ( ~n8473 & n10428 ) ;
  assign n10430 = n8450 ^ n7786 ^ n6572 ;
  assign n10431 = ( n6903 & n8772 ) | ( n6903 & ~n10430 ) | ( n8772 & ~n10430 ) ;
  assign n10432 = ( n4428 & n9759 ) | ( n4428 & n10431 ) | ( n9759 & n10431 ) ;
  assign n10433 = ( ~n7858 & n10429 ) | ( ~n7858 & n10432 ) | ( n10429 & n10432 ) ;
  assign n10434 = n10107 ^ n3526 ^ n3420 ;
  assign n10435 = ( n4041 & n5344 ) | ( n4041 & ~n5766 ) | ( n5344 & ~n5766 ) ;
  assign n10454 = n629 | n3499 ;
  assign n10450 = ( n2058 & n5302 ) | ( n2058 & ~n7794 ) | ( n5302 & ~n7794 ) ;
  assign n10451 = ( n1834 & n3580 ) | ( n1834 & n10450 ) | ( n3580 & n10450 ) ;
  assign n10452 = ( n5107 & ~n6557 ) | ( n5107 & n10451 ) | ( ~n6557 & n10451 ) ;
  assign n10453 = ( ~n3902 & n5204 ) | ( ~n3902 & n10452 ) | ( n5204 & n10452 ) ;
  assign n10455 = n10454 ^ n10453 ^ n6033 ;
  assign n10436 = n7625 ^ n1281 ^ x19 ;
  assign n10437 = n10436 ^ n6724 ^ 1'b0 ;
  assign n10438 = n3836 | n4570 ;
  assign n10439 = n10438 ^ n4984 ^ n2504 ;
  assign n10440 = n10439 ^ n6918 ^ n3717 ;
  assign n10441 = n6934 ^ n4892 ^ n4600 ;
  assign n10444 = n5178 ^ n5101 ^ n1183 ;
  assign n10442 = n8518 ^ n7725 ^ n5178 ;
  assign n10443 = n2778 & n10442 ;
  assign n10445 = n10444 ^ n10443 ^ 1'b0 ;
  assign n10446 = n677 & n3369 ;
  assign n10447 = n10446 ^ n275 ^ 1'b0 ;
  assign n10448 = ( n10441 & n10445 ) | ( n10441 & n10447 ) | ( n10445 & n10447 ) ;
  assign n10449 = ( ~n10437 & n10440 ) | ( ~n10437 & n10448 ) | ( n10440 & n10448 ) ;
  assign n10456 = n10455 ^ n10449 ^ n1335 ;
  assign n10457 = n5433 ^ n4474 ^ n4398 ;
  assign n10458 = n10331 ^ n9026 ^ n7332 ;
  assign n10459 = n5877 ^ n374 ^ 1'b0 ;
  assign n10460 = ( n10457 & n10458 ) | ( n10457 & ~n10459 ) | ( n10458 & ~n10459 ) ;
  assign n10463 = n6921 | n7753 ;
  assign n10464 = n3866 | n10463 ;
  assign n10465 = ( ~n826 & n2493 ) | ( ~n826 & n10464 ) | ( n2493 & n10464 ) ;
  assign n10461 = n5917 ^ n2485 ^ n1136 ;
  assign n10462 = n10461 ^ n7506 ^ n6238 ;
  assign n10466 = n10465 ^ n10462 ^ n3027 ;
  assign n10467 = ( n3845 & n4692 ) | ( n3845 & ~n10466 ) | ( n4692 & ~n10466 ) ;
  assign n10468 = n10277 ^ n6711 ^ 1'b0 ;
  assign n10469 = n2586 & ~n10468 ;
  assign n10470 = ( n2327 & n9329 ) | ( n2327 & ~n10469 ) | ( n9329 & ~n10469 ) ;
  assign n10471 = ( n2510 & n10467 ) | ( n2510 & ~n10470 ) | ( n10467 & ~n10470 ) ;
  assign n10472 = ( n6736 & n9503 ) | ( n6736 & n9560 ) | ( n9503 & n9560 ) ;
  assign n10473 = ( n2805 & ~n5334 ) | ( n2805 & n6660 ) | ( ~n5334 & n6660 ) ;
  assign n10483 = n1411 & ~n2668 ;
  assign n10484 = n10483 ^ n1350 ^ 1'b0 ;
  assign n10481 = n4819 | n6091 ;
  assign n10482 = n9841 & ~n10481 ;
  assign n10476 = ( ~x102 & n1267 ) | ( ~x102 & n1305 ) | ( n1267 & n1305 ) ;
  assign n10477 = ( n4013 & ~n8587 ) | ( n4013 & n9614 ) | ( ~n8587 & n9614 ) ;
  assign n10478 = n10477 ^ n6039 ^ x211 ;
  assign n10479 = ( n6215 & n10476 ) | ( n6215 & ~n10478 ) | ( n10476 & ~n10478 ) ;
  assign n10474 = n4456 ^ n2173 ^ n1599 ;
  assign n10475 = ( n2785 & n4656 ) | ( n2785 & ~n10474 ) | ( n4656 & ~n10474 ) ;
  assign n10480 = n10479 ^ n10475 ^ n8000 ;
  assign n10485 = n10484 ^ n10482 ^ n10480 ;
  assign n10486 = n10473 & n10485 ;
  assign n10487 = ( x79 & ~n1376 ) | ( x79 & n1382 ) | ( ~n1376 & n1382 ) ;
  assign n10488 = ( ~x92 & n2481 ) | ( ~x92 & n10487 ) | ( n2481 & n10487 ) ;
  assign n10489 = n8484 ^ n3564 ^ 1'b0 ;
  assign n10490 = ( n5140 & n10488 ) | ( n5140 & n10489 ) | ( n10488 & n10489 ) ;
  assign n10493 = n5848 & ~n8868 ;
  assign n10491 = ( ~n3887 & n7123 ) | ( ~n3887 & n7466 ) | ( n7123 & n7466 ) ;
  assign n10492 = n10491 ^ n10095 ^ n9995 ;
  assign n10494 = n10493 ^ n10492 ^ n3141 ;
  assign n10495 = ( ~n1929 & n4751 ) | ( ~n1929 & n8618 ) | ( n4751 & n8618 ) ;
  assign n10496 = n10495 ^ x102 ^ 1'b0 ;
  assign n10497 = n10494 | n10496 ;
  assign n10498 = n7451 ^ n2380 ^ 1'b0 ;
  assign n10499 = ( ~n1467 & n10497 ) | ( ~n1467 & n10498 ) | ( n10497 & n10498 ) ;
  assign n10500 = n10499 ^ n5966 ^ 1'b0 ;
  assign n10504 = ~n1583 & n2627 ;
  assign n10505 = n10504 ^ n7353 ^ n361 ;
  assign n10502 = ( ~x177 & n6092 ) | ( ~x177 & n6650 ) | ( n6092 & n6650 ) ;
  assign n10501 = n5790 ^ n5183 ^ n4002 ;
  assign n10503 = n10502 ^ n10501 ^ n9827 ;
  assign n10506 = n10505 ^ n10503 ^ n1528 ;
  assign n10507 = n10506 ^ n6715 ^ n6152 ;
  assign n10508 = n7980 ^ n7337 ^ n3979 ;
  assign n10512 = n2626 ^ n2463 ^ n1467 ;
  assign n10509 = ( ~n3819 & n6241 ) | ( ~n3819 & n7653 ) | ( n6241 & n7653 ) ;
  assign n10510 = n10509 ^ n2474 ^ n848 ;
  assign n10511 = n10510 ^ n9518 ^ n7202 ;
  assign n10513 = n10512 ^ n10511 ^ n371 ;
  assign n10514 = ( ~n5453 & n10508 ) | ( ~n5453 & n10513 ) | ( n10508 & n10513 ) ;
  assign n10515 = ( n2687 & ~n8803 ) | ( n2687 & n9991 ) | ( ~n8803 & n9991 ) ;
  assign n10516 = n10515 ^ n3615 ^ n3256 ;
  assign n10517 = ( n2381 & n4949 ) | ( n2381 & ~n10516 ) | ( n4949 & ~n10516 ) ;
  assign n10518 = x162 & n1356 ;
  assign n10519 = n2342 & n10518 ;
  assign n10520 = ( n763 & n4916 ) | ( n763 & n8293 ) | ( n4916 & n8293 ) ;
  assign n10521 = n10520 ^ n8858 ^ n340 ;
  assign n10522 = n1034 ^ n784 ^ n512 ;
  assign n10523 = ( x99 & n799 ) | ( x99 & n1112 ) | ( n799 & n1112 ) ;
  assign n10524 = ( n1896 & ~n10522 ) | ( n1896 & n10523 ) | ( ~n10522 & n10523 ) ;
  assign n10525 = ( n4826 & n9311 ) | ( n4826 & ~n10524 ) | ( n9311 & ~n10524 ) ;
  assign n10526 = ( ~n10519 & n10521 ) | ( ~n10519 & n10525 ) | ( n10521 & n10525 ) ;
  assign n10527 = n4869 ^ n3815 ^ n1051 ;
  assign n10528 = n4061 & n10386 ;
  assign n10529 = ( n8060 & ~n10527 ) | ( n8060 & n10528 ) | ( ~n10527 & n10528 ) ;
  assign n10530 = n10529 ^ n3414 ^ x245 ;
  assign n10531 = ( n718 & n1612 ) | ( n718 & n3891 ) | ( n1612 & n3891 ) ;
  assign n10532 = n4167 & n10531 ;
  assign n10533 = n1695 & n10532 ;
  assign n10534 = n10533 ^ n1599 ^ x174 ;
  assign n10541 = ( ~n276 & n2811 ) | ( ~n276 & n3779 ) | ( n2811 & n3779 ) ;
  assign n10535 = ( n519 & n1203 ) | ( n519 & n1454 ) | ( n1203 & n1454 ) ;
  assign n10536 = n10535 ^ n3559 ^ n3309 ;
  assign n10537 = n10536 ^ n3758 ^ 1'b0 ;
  assign n10538 = n379 & n10537 ;
  assign n10539 = n10538 ^ n4949 ^ n2017 ;
  assign n10540 = n10539 ^ n3732 ^ 1'b0 ;
  assign n10542 = n10541 ^ n10540 ^ x231 ;
  assign n10543 = ( ~n2682 & n10534 ) | ( ~n2682 & n10542 ) | ( n10534 & n10542 ) ;
  assign n10544 = n5219 ^ n4749 ^ n2738 ;
  assign n10545 = n4774 | n10544 ;
  assign n10546 = n8633 & ~n10545 ;
  assign n10547 = ( n3117 & ~n4882 ) | ( n3117 & n8558 ) | ( ~n4882 & n8558 ) ;
  assign n10548 = ( ~n6122 & n10189 ) | ( ~n6122 & n10547 ) | ( n10189 & n10547 ) ;
  assign n10549 = n10546 | n10548 ;
  assign n10550 = n4768 ^ n3183 ^ n2800 ;
  assign n10551 = ( n3887 & n8901 ) | ( n3887 & ~n10550 ) | ( n8901 & ~n10550 ) ;
  assign n10552 = ( n733 & n10549 ) | ( n733 & ~n10551 ) | ( n10549 & ~n10551 ) ;
  assign n10553 = ( n4553 & n8624 ) | ( n4553 & n10395 ) | ( n8624 & n10395 ) ;
  assign n10554 = ( n2631 & ~n6473 ) | ( n2631 & n9144 ) | ( ~n6473 & n9144 ) ;
  assign n10555 = n10554 ^ n1257 ^ n915 ;
  assign n10556 = ( n4015 & n6390 ) | ( n4015 & n10555 ) | ( n6390 & n10555 ) ;
  assign n10558 = ( n973 & n4908 ) | ( n973 & ~n8157 ) | ( n4908 & ~n8157 ) ;
  assign n10559 = n1565 & n10558 ;
  assign n10560 = n8165 & n10559 ;
  assign n10557 = ( n2563 & ~n3472 ) | ( n2563 & n8412 ) | ( ~n3472 & n8412 ) ;
  assign n10561 = n10560 ^ n10557 ^ n5585 ;
  assign n10562 = n6599 ^ n2835 ^ 1'b0 ;
  assign n10563 = n10562 ^ n8115 ^ n3845 ;
  assign n10564 = ( x21 & n2464 ) | ( x21 & ~n5863 ) | ( n2464 & ~n5863 ) ;
  assign n10565 = n10564 ^ n4915 ^ n4655 ;
  assign n10566 = ( n3278 & n6967 ) | ( n3278 & n10565 ) | ( n6967 & n10565 ) ;
  assign n10567 = ( n402 & n9280 ) | ( n402 & n10133 ) | ( n9280 & n10133 ) ;
  assign n10568 = ( n2213 & n5151 ) | ( n2213 & n10567 ) | ( n5151 & n10567 ) ;
  assign n10569 = ( n1303 & n10566 ) | ( n1303 & n10568 ) | ( n10566 & n10568 ) ;
  assign n10570 = ( n2885 & n3139 ) | ( n2885 & n3922 ) | ( n3139 & n3922 ) ;
  assign n10571 = n10570 ^ n9555 ^ n1690 ;
  assign n10572 = ( n3172 & n3496 ) | ( n3172 & n10571 ) | ( n3496 & n10571 ) ;
  assign n10574 = n3243 & ~n3582 ;
  assign n10575 = n10574 ^ n8257 ^ 1'b0 ;
  assign n10573 = ( x186 & n484 ) | ( x186 & ~n2647 ) | ( n484 & ~n2647 ) ;
  assign n10576 = n10575 ^ n10573 ^ n2860 ;
  assign n10577 = ( n3667 & ~n7793 ) | ( n3667 & n10407 ) | ( ~n7793 & n10407 ) ;
  assign n10578 = n4904 ^ n3943 ^ n2828 ;
  assign n10583 = n4774 ^ n3857 ^ n2824 ;
  assign n10584 = n10583 ^ n4663 ^ n1276 ;
  assign n10579 = n4338 ^ n2643 ^ n1419 ;
  assign n10580 = ( n2054 & n3127 ) | ( n2054 & ~n8414 ) | ( n3127 & ~n8414 ) ;
  assign n10581 = ~n3723 & n10580 ;
  assign n10582 = n10579 & n10581 ;
  assign n10585 = n10584 ^ n10582 ^ n7365 ;
  assign n10586 = n4490 & ~n7044 ;
  assign n10587 = n10585 & n10586 ;
  assign n10588 = ( n6293 & ~n10578 ) | ( n6293 & n10587 ) | ( ~n10578 & n10587 ) ;
  assign n10589 = ( x208 & n4482 ) | ( x208 & ~n5438 ) | ( n4482 & ~n5438 ) ;
  assign n10590 = ( n889 & n5940 ) | ( n889 & ~n10589 ) | ( n5940 & ~n10589 ) ;
  assign n10591 = ( n4150 & ~n4364 ) | ( n4150 & n10590 ) | ( ~n4364 & n10590 ) ;
  assign n10592 = ( n1379 & n3990 ) | ( n1379 & ~n5327 ) | ( n3990 & ~n5327 ) ;
  assign n10593 = ( n1788 & n2462 ) | ( n1788 & n9797 ) | ( n2462 & n9797 ) ;
  assign n10594 = ( n7671 & n10592 ) | ( n7671 & n10593 ) | ( n10592 & n10593 ) ;
  assign n10597 = n1640 | n7128 ;
  assign n10598 = n4054 | n10597 ;
  assign n10596 = ( n1044 & n1143 ) | ( n1044 & ~n8521 ) | ( n1143 & ~n8521 ) ;
  assign n10599 = n10598 ^ n10596 ^ n5128 ;
  assign n10595 = ( n3898 & n5686 ) | ( n3898 & ~n6243 ) | ( n5686 & ~n6243 ) ;
  assign n10600 = n10599 ^ n10595 ^ n870 ;
  assign n10601 = n479 & ~n1431 ;
  assign n10602 = n10601 ^ n1439 ^ 1'b0 ;
  assign n10603 = n1760 ^ n907 ^ n847 ;
  assign n10604 = ~n1064 & n10603 ;
  assign n10605 = n2468 & n10604 ;
  assign n10606 = ( n2141 & n5148 ) | ( n2141 & ~n10605 ) | ( n5148 & ~n10605 ) ;
  assign n10607 = ~n10602 & n10606 ;
  assign n10608 = ( n10594 & n10600 ) | ( n10594 & n10607 ) | ( n10600 & n10607 ) ;
  assign n10609 = n4662 ^ n3526 ^ 1'b0 ;
  assign n10610 = n7869 & ~n10609 ;
  assign n10611 = n6742 ^ n5836 ^ n1600 ;
  assign n10612 = n1809 | n1870 ;
  assign n10613 = n10612 ^ n8237 ^ 1'b0 ;
  assign n10614 = ( ~n387 & n1836 ) | ( ~n387 & n1928 ) | ( n1836 & n1928 ) ;
  assign n10615 = n10614 ^ n8573 ^ 1'b0 ;
  assign n10616 = ( ~n10611 & n10613 ) | ( ~n10611 & n10615 ) | ( n10613 & n10615 ) ;
  assign n10617 = n9177 ^ n2888 ^ 1'b0 ;
  assign n10618 = n10617 ^ n4320 ^ n2212 ;
  assign n10619 = ( ~n3576 & n5122 ) | ( ~n3576 & n10618 ) | ( n5122 & n10618 ) ;
  assign n10620 = n3365 | n8978 ;
  assign n10621 = ( ~n3124 & n7790 ) | ( ~n3124 & n10620 ) | ( n7790 & n10620 ) ;
  assign n10622 = n10621 ^ n6583 ^ n4363 ;
  assign n10623 = ( n4453 & ~n7833 ) | ( n4453 & n9433 ) | ( ~n7833 & n9433 ) ;
  assign n10624 = ( ~n1888 & n4082 ) | ( ~n1888 & n6237 ) | ( n4082 & n6237 ) ;
  assign n10625 = n10624 ^ n6640 ^ n5289 ;
  assign n10626 = ( n1283 & ~n2062 ) | ( n1283 & n5228 ) | ( ~n2062 & n5228 ) ;
  assign n10627 = n1392 & n1828 ;
  assign n10628 = n10626 & n10627 ;
  assign n10629 = n10628 ^ n6257 ^ n3429 ;
  assign n10630 = n10629 ^ x238 ^ 1'b0 ;
  assign n10631 = n3105 & ~n10630 ;
  assign n10632 = n895 & n2126 ;
  assign n10633 = n10632 ^ n4148 ^ 1'b0 ;
  assign n10634 = n10633 ^ n2640 ^ x137 ;
  assign n10635 = ( n3436 & n3489 ) | ( n3436 & ~n10634 ) | ( n3489 & ~n10634 ) ;
  assign n10636 = ( n4743 & n6388 ) | ( n4743 & ~n10635 ) | ( n6388 & ~n10635 ) ;
  assign n10637 = ( x66 & n7254 ) | ( x66 & ~n10636 ) | ( n7254 & ~n10636 ) ;
  assign n10638 = ( ~n10625 & n10631 ) | ( ~n10625 & n10637 ) | ( n10631 & n10637 ) ;
  assign n10639 = n3427 & ~n4700 ;
  assign n10640 = n10639 ^ n3502 ^ 1'b0 ;
  assign n10641 = ( n8358 & ~n9931 ) | ( n8358 & n10640 ) | ( ~n9931 & n10640 ) ;
  assign n10642 = n10641 ^ n5886 ^ n2515 ;
  assign n10643 = ( n1969 & n8281 ) | ( n1969 & ~n9741 ) | ( n8281 & ~n9741 ) ;
  assign n10644 = n7860 ^ n5649 ^ n5225 ;
  assign n10645 = n10643 & n10644 ;
  assign n10646 = n10642 & n10645 ;
  assign n10647 = n10646 ^ n9256 ^ n4430 ;
  assign n10648 = ( ~n5368 & n8844 ) | ( ~n5368 & n10647 ) | ( n8844 & n10647 ) ;
  assign n10649 = n10648 ^ n426 ^ x149 ;
  assign n10650 = ( n1513 & n2838 ) | ( n1513 & ~n4220 ) | ( n2838 & ~n4220 ) ;
  assign n10651 = n10650 ^ n10306 ^ n8699 ;
  assign n10652 = n10651 ^ n6144 ^ n3139 ;
  assign n10653 = ( n2630 & n6512 ) | ( n2630 & ~n9308 ) | ( n6512 & ~n9308 ) ;
  assign n10654 = ( ~n4391 & n4484 ) | ( ~n4391 & n10653 ) | ( n4484 & n10653 ) ;
  assign n10655 = ( ~n737 & n10652 ) | ( ~n737 & n10654 ) | ( n10652 & n10654 ) ;
  assign n10656 = x66 & ~n4629 ;
  assign n10657 = n10656 ^ n4390 ^ 1'b0 ;
  assign n10658 = n10657 ^ n9258 ^ n2514 ;
  assign n10659 = n393 & n8290 ;
  assign n10660 = ( n8447 & ~n10658 ) | ( n8447 & n10659 ) | ( ~n10658 & n10659 ) ;
  assign n10661 = n10660 ^ n6074 ^ n1182 ;
  assign n10669 = n5245 ^ n2275 ^ n1261 ;
  assign n10666 = ~n504 & n8221 ;
  assign n10667 = ~n3975 & n10666 ;
  assign n10668 = ( n495 & n1589 ) | ( n495 & ~n10667 ) | ( n1589 & ~n10667 ) ;
  assign n10662 = n2654 | n9424 ;
  assign n10663 = n10662 ^ n4529 ^ 1'b0 ;
  assign n10664 = n6466 | n10663 ;
  assign n10665 = n10664 ^ n6761 ^ 1'b0 ;
  assign n10670 = n10669 ^ n10668 ^ n10665 ;
  assign n10671 = ( n1213 & n2140 ) | ( n1213 & n4361 ) | ( n2140 & n4361 ) ;
  assign n10672 = n10671 ^ n1535 ^ n1450 ;
  assign n10673 = n6513 & n10672 ;
  assign n10682 = n6829 ^ n3864 ^ n2658 ;
  assign n10680 = n6124 ^ n4629 ^ n1219 ;
  assign n10681 = n10680 ^ n3558 ^ n3265 ;
  assign n10683 = n10682 ^ n10681 ^ n979 ;
  assign n10674 = ( x62 & ~n2396 ) | ( x62 & n3484 ) | ( ~n2396 & n3484 ) ;
  assign n10675 = ( n6480 & n7436 ) | ( n6480 & n10674 ) | ( n7436 & n10674 ) ;
  assign n10676 = n10675 ^ n5930 ^ n2308 ;
  assign n10677 = n9292 ^ n3195 ^ n1944 ;
  assign n10678 = ( n5496 & ~n10676 ) | ( n5496 & n10677 ) | ( ~n10676 & n10677 ) ;
  assign n10679 = n10678 ^ n9177 ^ n3403 ;
  assign n10684 = n10683 ^ n10679 ^ n3098 ;
  assign n10685 = ( n9372 & ~n9420 ) | ( n9372 & n10684 ) | ( ~n9420 & n10684 ) ;
  assign n10686 = n8440 ^ n5800 ^ n1055 ;
  assign n10687 = n820 & ~n8429 ;
  assign n10688 = ( ~n663 & n5782 ) | ( ~n663 & n10687 ) | ( n5782 & n10687 ) ;
  assign n10689 = n10633 ^ n2839 ^ n1526 ;
  assign n10690 = ( n10686 & ~n10688 ) | ( n10686 & n10689 ) | ( ~n10688 & n10689 ) ;
  assign n10691 = ~n5892 & n10681 ;
  assign n10692 = ~n10690 & n10691 ;
  assign n10693 = n1125 & n7696 ;
  assign n10696 = n5169 ^ n1182 ^ 1'b0 ;
  assign n10697 = ~n2813 & n10696 ;
  assign n10694 = n5663 & ~n6991 ;
  assign n10695 = n10694 ^ n2542 ^ n1431 ;
  assign n10698 = n10697 ^ n10695 ^ n5860 ;
  assign n10708 = ( n601 & n651 ) | ( n601 & ~n849 ) | ( n651 & ~n849 ) ;
  assign n10709 = ( ~n962 & n2018 ) | ( ~n962 & n10708 ) | ( n2018 & n10708 ) ;
  assign n10710 = ( ~n736 & n1212 ) | ( ~n736 & n1440 ) | ( n1212 & n1440 ) ;
  assign n10711 = ( x9 & n6185 ) | ( x9 & ~n10710 ) | ( n6185 & ~n10710 ) ;
  assign n10712 = ( n4319 & n10709 ) | ( n4319 & n10711 ) | ( n10709 & n10711 ) ;
  assign n10713 = ( n3209 & n5061 ) | ( n3209 & ~n10712 ) | ( n5061 & ~n10712 ) ;
  assign n10707 = n2553 ^ n698 ^ 1'b0 ;
  assign n10714 = n10713 ^ n10707 ^ n8945 ;
  assign n10699 = n4668 & n8044 ;
  assign n10700 = n10699 ^ n3764 ^ 1'b0 ;
  assign n10703 = n284 & n1299 ;
  assign n10704 = ~x118 & n10703 ;
  assign n10701 = n1648 ^ n1067 ^ n439 ;
  assign n10702 = ( ~n659 & n6084 ) | ( ~n659 & n10701 ) | ( n6084 & n10701 ) ;
  assign n10705 = n10704 ^ n10702 ^ n4999 ;
  assign n10706 = ( ~n5837 & n10700 ) | ( ~n5837 & n10705 ) | ( n10700 & n10705 ) ;
  assign n10715 = n10714 ^ n10706 ^ n10488 ;
  assign n10716 = n7154 & n8284 ;
  assign n10717 = n2100 & n10716 ;
  assign n10718 = ~n301 & n10717 ;
  assign n10719 = n10718 ^ n7046 ^ n2952 ;
  assign n10720 = n9564 ^ n9420 ^ n2842 ;
  assign n10721 = ( ~n258 & n8939 ) | ( ~n258 & n9291 ) | ( n8939 & n9291 ) ;
  assign n10722 = ( ~n7396 & n8627 ) | ( ~n7396 & n10721 ) | ( n8627 & n10721 ) ;
  assign n10723 = ( n10719 & n10720 ) | ( n10719 & ~n10722 ) | ( n10720 & ~n10722 ) ;
  assign n10724 = ( n856 & n1084 ) | ( n856 & n9537 ) | ( n1084 & n9537 ) ;
  assign n10725 = ( x181 & n2240 ) | ( x181 & ~n4792 ) | ( n2240 & ~n4792 ) ;
  assign n10726 = n10725 ^ n1927 ^ n1694 ;
  assign n10727 = n10726 ^ n5308 ^ n287 ;
  assign n10728 = n5178 ^ n1372 ^ 1'b0 ;
  assign n10729 = n7444 & ~n10728 ;
  assign n10730 = ( n6994 & ~n8335 ) | ( n6994 & n10729 ) | ( ~n8335 & n10729 ) ;
  assign n10731 = n10730 ^ n7953 ^ n7882 ;
  assign n10732 = ( n6807 & n10727 ) | ( n6807 & ~n10731 ) | ( n10727 & ~n10731 ) ;
  assign n10733 = ( ~n3317 & n10724 ) | ( ~n3317 & n10732 ) | ( n10724 & n10732 ) ;
  assign n10734 = n8006 ^ n3468 ^ n2314 ;
  assign n10735 = n10734 ^ n2134 ^ n831 ;
  assign n10737 = n6967 ^ n2602 ^ n389 ;
  assign n10738 = ( ~n1176 & n4842 ) | ( ~n1176 & n7510 ) | ( n4842 & n7510 ) ;
  assign n10739 = n10737 & ~n10738 ;
  assign n10740 = n10739 ^ n3797 ^ 1'b0 ;
  assign n10741 = n10584 ^ n6851 ^ n595 ;
  assign n10742 = ( n2563 & n10740 ) | ( n2563 & ~n10741 ) | ( n10740 & ~n10741 ) ;
  assign n10736 = n3831 ^ n2020 ^ n1683 ;
  assign n10743 = n10742 ^ n10736 ^ n5866 ;
  assign n10744 = ( n8634 & n9641 ) | ( n8634 & ~n10063 ) | ( n9641 & ~n10063 ) ;
  assign n10745 = ( n10735 & n10743 ) | ( n10735 & n10744 ) | ( n10743 & n10744 ) ;
  assign n10746 = n5439 ^ n2856 ^ n1653 ;
  assign n10747 = n8152 & ~n10746 ;
  assign n10748 = n10745 & n10747 ;
  assign n10749 = ( ~n1364 & n6884 ) | ( ~n1364 & n9503 ) | ( n6884 & n9503 ) ;
  assign n10750 = n1033 & n7529 ;
  assign n10751 = n4584 & ~n7980 ;
  assign n10752 = n10751 ^ n5225 ^ n903 ;
  assign n10753 = n10752 ^ n327 ^ 1'b0 ;
  assign n10754 = n10753 ^ n7519 ^ n541 ;
  assign n10755 = n8045 ^ x157 ^ 1'b0 ;
  assign n10756 = ~n5210 & n10755 ;
  assign n10757 = n1175 & n10756 ;
  assign n10758 = n10757 ^ n5416 ^ 1'b0 ;
  assign n10759 = n10758 ^ n7129 ^ n5296 ;
  assign n10760 = ( x60 & ~n435 ) | ( x60 & n10759 ) | ( ~n435 & n10759 ) ;
  assign n10761 = n10760 ^ n5262 ^ n1130 ;
  assign n10762 = ( ~n683 & n883 ) | ( ~n683 & n1344 ) | ( n883 & n1344 ) ;
  assign n10763 = ( n838 & n2762 ) | ( n838 & ~n5475 ) | ( n2762 & ~n5475 ) ;
  assign n10764 = n10763 ^ n2645 ^ n433 ;
  assign n10765 = n3523 ^ n3103 ^ 1'b0 ;
  assign n10766 = ( n10762 & ~n10764 ) | ( n10762 & n10765 ) | ( ~n10764 & n10765 ) ;
  assign n10767 = n10766 ^ n1469 ^ 1'b0 ;
  assign n10768 = ( n3569 & ~n3602 ) | ( n3569 & n10767 ) | ( ~n3602 & n10767 ) ;
  assign n10769 = n4214 ^ n3385 ^ n1461 ;
  assign n10770 = n10769 ^ n8620 ^ n2286 ;
  assign n10774 = ( n2999 & ~n3743 ) | ( n2999 & n4448 ) | ( ~n3743 & n4448 ) ;
  assign n10775 = n4495 ^ n2949 ^ n1515 ;
  assign n10776 = n10775 ^ n5691 ^ n1562 ;
  assign n10777 = n10776 ^ n3383 ^ 1'b0 ;
  assign n10778 = ( n1158 & n10774 ) | ( n1158 & ~n10777 ) | ( n10774 & ~n10777 ) ;
  assign n10771 = n10633 ^ n1897 ^ 1'b0 ;
  assign n10772 = n8592 & ~n10771 ;
  assign n10773 = ( ~n1656 & n10167 ) | ( ~n1656 & n10772 ) | ( n10167 & n10772 ) ;
  assign n10779 = n10778 ^ n10773 ^ n4150 ;
  assign n10780 = ( n2126 & n10770 ) | ( n2126 & ~n10779 ) | ( n10770 & ~n10779 ) ;
  assign n10787 = n1788 & n5397 ;
  assign n10788 = n3883 & n10787 ;
  assign n10782 = ( n1067 & n1437 ) | ( n1067 & ~n6253 ) | ( n1437 & ~n6253 ) ;
  assign n10781 = n8277 ^ n4390 ^ n4058 ;
  assign n10783 = n10782 ^ n10781 ^ n6082 ;
  assign n10784 = ( n6086 & ~n6200 ) | ( n6086 & n10783 ) | ( ~n6200 & n10783 ) ;
  assign n10785 = n10784 ^ n9521 ^ n5232 ;
  assign n10786 = n10785 ^ n10131 ^ x176 ;
  assign n10789 = n10788 ^ n10786 ^ n9041 ;
  assign n10790 = n5532 ^ n314 ^ 1'b0 ;
  assign n10791 = ( n2517 & n4571 ) | ( n2517 & ~n10593 ) | ( n4571 & ~n10593 ) ;
  assign n10792 = ( n6493 & ~n8784 ) | ( n6493 & n10791 ) | ( ~n8784 & n10791 ) ;
  assign n10793 = ( ~n2206 & n10790 ) | ( ~n2206 & n10792 ) | ( n10790 & n10792 ) ;
  assign n10795 = n3830 ^ n2244 ^ 1'b0 ;
  assign n10794 = ( x136 & n1930 ) | ( x136 & n3602 ) | ( n1930 & n3602 ) ;
  assign n10796 = n10795 ^ n10794 ^ n3712 ;
  assign n10797 = n7539 ^ n7024 ^ n1630 ;
  assign n10798 = ( n7820 & n9263 ) | ( n7820 & n10797 ) | ( n9263 & n10797 ) ;
  assign n10799 = n943 ^ n538 ^ n530 ;
  assign n10800 = n10799 ^ n8696 ^ 1'b0 ;
  assign n10801 = n10800 ^ n9086 ^ 1'b0 ;
  assign n10802 = n10801 ^ n4216 ^ 1'b0 ;
  assign n10803 = n7923 ^ n4022 ^ n2521 ;
  assign n10804 = n6681 & ~n10803 ;
  assign n10808 = n4877 ^ n4876 ^ n1167 ;
  assign n10809 = ( ~n2576 & n3622 ) | ( ~n2576 & n10808 ) | ( n3622 & n10808 ) ;
  assign n10805 = n10418 ^ n10400 ^ n4337 ;
  assign n10806 = ( ~n2833 & n10216 ) | ( ~n2833 & n10805 ) | ( n10216 & n10805 ) ;
  assign n10807 = ( n3670 & ~n7525 ) | ( n3670 & n10806 ) | ( ~n7525 & n10806 ) ;
  assign n10810 = n10809 ^ n10807 ^ n10225 ;
  assign n10811 = ( n1136 & n3343 ) | ( n1136 & ~n10810 ) | ( n3343 & ~n10810 ) ;
  assign n10812 = ( n10260 & ~n10804 ) | ( n10260 & n10811 ) | ( ~n10804 & n10811 ) ;
  assign n10813 = n7905 ^ n2852 ^ n2573 ;
  assign n10815 = n5836 & ~n6733 ;
  assign n10814 = n9268 ^ n7083 ^ n1737 ;
  assign n10816 = n10815 ^ n10814 ^ n7346 ;
  assign n10820 = n7188 ^ n6827 ^ n4988 ;
  assign n10818 = n8152 ^ n5285 ^ n1881 ;
  assign n10819 = n10818 ^ n9139 ^ n760 ;
  assign n10817 = n8054 ^ n5994 ^ 1'b0 ;
  assign n10821 = n10820 ^ n10819 ^ n10817 ;
  assign n10822 = ( n3374 & n9897 ) | ( n3374 & n10821 ) | ( n9897 & n10821 ) ;
  assign n10823 = ( n8429 & ~n10816 ) | ( n8429 & n10822 ) | ( ~n10816 & n10822 ) ;
  assign n10829 = n7489 ^ n3306 ^ x222 ;
  assign n10826 = n465 & ~n2076 ;
  assign n10825 = ( ~n1362 & n3050 ) | ( ~n1362 & n5580 ) | ( n3050 & n5580 ) ;
  assign n10827 = n10826 ^ n10825 ^ n1611 ;
  assign n10828 = n10827 ^ n733 ^ 1'b0 ;
  assign n10824 = n6938 ^ n3655 ^ 1'b0 ;
  assign n10830 = n10829 ^ n10828 ^ n10824 ;
  assign n10831 = ( n874 & ~n1166 ) | ( n874 & n6914 ) | ( ~n1166 & n6914 ) ;
  assign n10832 = ( ~n5548 & n7225 ) | ( ~n5548 & n10831 ) | ( n7225 & n10831 ) ;
  assign n10833 = n10832 ^ n10225 ^ n6273 ;
  assign n10834 = n10833 ^ n10442 ^ n3075 ;
  assign n10838 = n6815 ^ n6736 ^ n1204 ;
  assign n10839 = ( n520 & n2907 ) | ( n520 & ~n10838 ) | ( n2907 & ~n10838 ) ;
  assign n10835 = n3125 ^ n1607 ^ x120 ;
  assign n10836 = n4751 & n10835 ;
  assign n10837 = ( x124 & ~n5309 ) | ( x124 & n10836 ) | ( ~n5309 & n10836 ) ;
  assign n10840 = n10839 ^ n10837 ^ 1'b0 ;
  assign n10841 = n6187 ^ n5209 ^ n369 ;
  assign n10842 = ( n2200 & ~n2268 ) | ( n2200 & n2598 ) | ( ~n2268 & n2598 ) ;
  assign n10843 = n10842 ^ n4080 ^ n846 ;
  assign n10844 = n10709 ^ n10614 ^ n9972 ;
  assign n10845 = ~n10843 & n10844 ;
  assign n10846 = n10845 ^ n8302 ^ n1700 ;
  assign n10847 = ( n10840 & n10841 ) | ( n10840 & n10846 ) | ( n10841 & n10846 ) ;
  assign n10848 = n2691 ^ n2071 ^ n1007 ;
  assign n10849 = n10848 ^ n666 ^ 1'b0 ;
  assign n10850 = n10849 ^ n9758 ^ n8268 ;
  assign n10851 = n2195 | n10850 ;
  assign n10852 = n10315 | n10851 ;
  assign n10853 = n6014 ^ n4487 ^ n1111 ;
  assign n10854 = n10853 ^ n1899 ^ 1'b0 ;
  assign n10855 = n8725 ^ n3620 ^ n3118 ;
  assign n10856 = n10770 ^ x219 ^ 1'b0 ;
  assign n10857 = n4729 & ~n10856 ;
  assign n10858 = n10857 ^ n2963 ^ n949 ;
  assign n10859 = n5374 ^ n5368 ^ 1'b0 ;
  assign n10860 = n6526 & n10859 ;
  assign n10861 = n3417 ^ n1897 ^ x44 ;
  assign n10862 = n10861 ^ n2797 ^ n1619 ;
  assign n10865 = ( n1387 & n2462 ) | ( n1387 & n7605 ) | ( n2462 & n7605 ) ;
  assign n10863 = ~n1095 & n1295 ;
  assign n10864 = ~n5680 & n10863 ;
  assign n10866 = n10865 ^ n10864 ^ n8653 ;
  assign n10867 = ( ~n256 & n10862 ) | ( ~n256 & n10866 ) | ( n10862 & n10866 ) ;
  assign n10868 = n10867 ^ n10646 ^ n5540 ;
  assign n10869 = ( ~n1741 & n2345 ) | ( ~n1741 & n5499 ) | ( n2345 & n5499 ) ;
  assign n10870 = n1055 ^ n807 ^ x117 ;
  assign n10871 = n10870 ^ n4629 ^ n2389 ;
  assign n10872 = n10869 | n10871 ;
  assign n10873 = n4908 | n10872 ;
  assign n10874 = ( n1000 & n3866 ) | ( n1000 & ~n7496 ) | ( n3866 & ~n7496 ) ;
  assign n10875 = n7295 ^ n7090 ^ n5980 ;
  assign n10876 = ( n5796 & n10874 ) | ( n5796 & ~n10875 ) | ( n10874 & ~n10875 ) ;
  assign n10877 = n6177 ^ n2605 ^ n288 ;
  assign n10878 = ( n6443 & n7097 ) | ( n6443 & n10635 ) | ( n7097 & n10635 ) ;
  assign n10879 = ( n885 & n10482 ) | ( n885 & ~n10878 ) | ( n10482 & ~n10878 ) ;
  assign n10880 = ( n2572 & ~n10877 ) | ( n2572 & n10879 ) | ( ~n10877 & n10879 ) ;
  assign n10882 = n5831 ^ n4654 ^ n1724 ;
  assign n10883 = ( ~n4935 & n8440 ) | ( ~n4935 & n10882 ) | ( n8440 & n10882 ) ;
  assign n10881 = n8158 ^ n4165 ^ n3938 ;
  assign n10884 = n10883 ^ n10881 ^ n3643 ;
  assign n10885 = n10884 ^ n7259 ^ n6993 ;
  assign n10886 = ( n4864 & n10880 ) | ( n4864 & ~n10885 ) | ( n10880 & ~n10885 ) ;
  assign n10887 = n5567 ^ n3185 ^ n1697 ;
  assign n10893 = n8974 ^ n7962 ^ n3110 ;
  assign n10888 = n4316 | n7753 ;
  assign n10889 = n3729 | n10888 ;
  assign n10890 = n6548 & n10889 ;
  assign n10891 = ~n4058 & n10890 ;
  assign n10892 = ( ~n3195 & n6172 ) | ( ~n3195 & n10891 ) | ( n6172 & n10891 ) ;
  assign n10894 = n10893 ^ n10892 ^ n10226 ;
  assign n10909 = n9677 ^ n8897 ^ n3784 ;
  assign n10904 = n3479 ^ n2643 ^ n1478 ;
  assign n10905 = n750 & ~n2824 ;
  assign n10906 = n1390 & n10905 ;
  assign n10907 = ( n651 & ~n10904 ) | ( n651 & n10906 ) | ( ~n10904 & n10906 ) ;
  assign n10899 = ~n1078 & n1683 ;
  assign n10900 = n10899 ^ n1911 ^ n1030 ;
  assign n10901 = ( n836 & ~n2543 ) | ( n836 & n10900 ) | ( ~n2543 & n10900 ) ;
  assign n10902 = n10901 ^ n5536 ^ n2256 ;
  assign n10903 = n10902 ^ n8946 ^ n8277 ;
  assign n10908 = n10907 ^ n10903 ^ n10165 ;
  assign n10910 = n10909 ^ n10908 ^ 1'b0 ;
  assign n10895 = n7432 ^ n1593 ^ n1584 ;
  assign n10896 = ( n4396 & ~n4932 ) | ( n4396 & n10895 ) | ( ~n4932 & n10895 ) ;
  assign n10897 = n7339 ^ n6484 ^ n929 ;
  assign n10898 = n10896 & n10897 ;
  assign n10911 = n10910 ^ n10898 ^ 1'b0 ;
  assign n10912 = n1695 | n8285 ;
  assign n10913 = n10912 ^ n3768 ^ 1'b0 ;
  assign n10914 = n10913 ^ n10538 ^ n3514 ;
  assign n10915 = ( n295 & ~n1601 ) | ( n295 & n8321 ) | ( ~n1601 & n8321 ) ;
  assign n10916 = ( n1223 & n6143 ) | ( n1223 & ~n10915 ) | ( n6143 & ~n10915 ) ;
  assign n10917 = n10916 ^ n1859 ^ x63 ;
  assign n10918 = n1176 & n10917 ;
  assign n10919 = n10918 ^ n10394 ^ 1'b0 ;
  assign n10920 = ( n10466 & ~n10914 ) | ( n10466 & n10919 ) | ( ~n10914 & n10919 ) ;
  assign n10921 = ( n1424 & ~n2240 ) | ( n1424 & n5344 ) | ( ~n2240 & n5344 ) ;
  assign n10922 = ( n759 & n3816 ) | ( n759 & n10921 ) | ( n3816 & n10921 ) ;
  assign n10923 = n4698 | n8165 ;
  assign n10924 = n10923 ^ n4708 ^ x70 ;
  assign n10925 = ( n9536 & n10922 ) | ( n9536 & n10924 ) | ( n10922 & n10924 ) ;
  assign n10926 = ~n8281 & n10925 ;
  assign n10927 = ~n2828 & n10926 ;
  assign n10928 = n4490 & ~n10927 ;
  assign n10929 = n10928 ^ n2902 ^ 1'b0 ;
  assign n10930 = n8521 ^ n1628 ^ n988 ;
  assign n10931 = n10930 ^ n4969 ^ 1'b0 ;
  assign n10932 = ( n2535 & n6018 ) | ( n2535 & ~n6908 ) | ( n6018 & ~n6908 ) ;
  assign n10933 = n2980 | n10932 ;
  assign n10934 = n1132 ^ n693 ^ 1'b0 ;
  assign n10935 = n8892 ^ n4398 ^ x196 ;
  assign n10936 = ( n3533 & ~n10934 ) | ( n3533 & n10935 ) | ( ~n10934 & n10935 ) ;
  assign n10937 = n8464 ^ n6668 ^ n2637 ;
  assign n10938 = ( n2844 & n3838 ) | ( n2844 & ~n10937 ) | ( n3838 & ~n10937 ) ;
  assign n10939 = ( n1912 & ~n2412 ) | ( n1912 & n10938 ) | ( ~n2412 & n10938 ) ;
  assign n10940 = ( n4852 & n5587 ) | ( n4852 & n10939 ) | ( n5587 & n10939 ) ;
  assign n10941 = ( ~n1485 & n3503 ) | ( ~n1485 & n8924 ) | ( n3503 & n8924 ) ;
  assign n10942 = n10941 ^ n4381 ^ n855 ;
  assign n10943 = n10940 | n10942 ;
  assign n10944 = n10943 ^ n9177 ^ 1'b0 ;
  assign n10945 = ~n929 & n6777 ;
  assign n10946 = n10945 ^ n6208 ^ 1'b0 ;
  assign n10947 = ( n8793 & ~n9940 ) | ( n8793 & n10946 ) | ( ~n9940 & n10946 ) ;
  assign n10952 = n2974 ^ n2105 ^ n1962 ;
  assign n10953 = n10952 ^ n8466 ^ n1442 ;
  assign n10948 = n8016 ^ n6598 ^ n264 ;
  assign n10949 = n10948 ^ n4487 ^ n3498 ;
  assign n10950 = n10949 ^ n3675 ^ n575 ;
  assign n10951 = ( n4368 & ~n7367 ) | ( n4368 & n10950 ) | ( ~n7367 & n10950 ) ;
  assign n10954 = n10953 ^ n10951 ^ n1906 ;
  assign n10955 = ( n1387 & ~n1901 ) | ( n1387 & n4941 ) | ( ~n1901 & n4941 ) ;
  assign n10956 = ~n3693 & n10955 ;
  assign n10957 = n10956 ^ n4038 ^ n871 ;
  assign n10958 = n9587 ^ n7150 ^ 1'b0 ;
  assign n10959 = ~n4427 & n10958 ;
  assign n10960 = ( ~n1804 & n2541 ) | ( ~n1804 & n10554 ) | ( n2541 & n10554 ) ;
  assign n10961 = ( n10957 & ~n10959 ) | ( n10957 & n10960 ) | ( ~n10959 & n10960 ) ;
  assign n10965 = n4804 & n8852 ;
  assign n10963 = n4823 ^ n3714 ^ n2362 ;
  assign n10962 = ( n4525 & n8586 ) | ( n4525 & ~n10848 ) | ( n8586 & ~n10848 ) ;
  assign n10964 = n10963 ^ n10962 ^ n1634 ;
  assign n10966 = n10965 ^ n10964 ^ n8849 ;
  assign n10967 = n3255 ^ n3105 ^ n871 ;
  assign n10968 = ( n7545 & n9829 ) | ( n7545 & n10967 ) | ( n9829 & n10967 ) ;
  assign n10969 = n4755 ^ n1924 ^ n380 ;
  assign n10970 = n10969 ^ n9104 ^ 1'b0 ;
  assign n10971 = n7619 ^ n4402 ^ n3154 ;
  assign n10972 = n4092 ^ n1817 ^ 1'b0 ;
  assign n10973 = n6272 ^ n3810 ^ n2447 ;
  assign n10974 = n1950 & ~n7667 ;
  assign n10975 = ( ~n6905 & n10973 ) | ( ~n6905 & n10974 ) | ( n10973 & n10974 ) ;
  assign n10976 = ( n9097 & n10972 ) | ( n9097 & ~n10975 ) | ( n10972 & ~n10975 ) ;
  assign n10977 = ( n623 & n5113 ) | ( n623 & ~n6362 ) | ( n5113 & ~n6362 ) ;
  assign n10979 = ( n724 & n1307 ) | ( n724 & n1368 ) | ( n1307 & n1368 ) ;
  assign n10978 = ( n693 & n1976 ) | ( n693 & ~n7250 ) | ( n1976 & ~n7250 ) ;
  assign n10980 = n10979 ^ n10978 ^ n4873 ;
  assign n10981 = ~n10977 & n10980 ;
  assign n10982 = n10976 & n10981 ;
  assign n10986 = n4187 ^ n2814 ^ n1741 ;
  assign n10985 = ( ~n741 & n4052 ) | ( ~n741 & n8776 ) | ( n4052 & n8776 ) ;
  assign n10983 = ( ~n2091 & n3870 ) | ( ~n2091 & n7171 ) | ( n3870 & n7171 ) ;
  assign n10984 = n10983 ^ n4112 ^ 1'b0 ;
  assign n10987 = n10986 ^ n10985 ^ n10984 ;
  assign n10988 = n8013 ^ n2967 ^ 1'b0 ;
  assign n10989 = n10988 ^ n1762 ^ 1'b0 ;
  assign n10990 = ~n6864 & n10989 ;
  assign n10991 = ( n3011 & ~n5593 ) | ( n3011 & n10990 ) | ( ~n5593 & n10990 ) ;
  assign n10992 = ( ~n3034 & n9554 ) | ( ~n3034 & n10991 ) | ( n9554 & n10991 ) ;
  assign n10993 = n6655 ^ n3354 ^ n3076 ;
  assign n10994 = ( n1780 & n7215 ) | ( n1780 & ~n10271 ) | ( n7215 & ~n10271 ) ;
  assign n10995 = ( n2936 & ~n10993 ) | ( n2936 & n10994 ) | ( ~n10993 & n10994 ) ;
  assign n10996 = ( n383 & n9183 ) | ( n383 & n10995 ) | ( n9183 & n10995 ) ;
  assign n11000 = ( x59 & ~n2077 ) | ( x59 & n5609 ) | ( ~n2077 & n5609 ) ;
  assign n10997 = ( n1013 & ~n1689 ) | ( n1013 & n2505 ) | ( ~n1689 & n2505 ) ;
  assign n10998 = n820 & ~n10997 ;
  assign n10999 = n10998 ^ n4869 ^ 1'b0 ;
  assign n11001 = n11000 ^ n10999 ^ 1'b0 ;
  assign n11002 = n11001 ^ n9164 ^ n1220 ;
  assign n11003 = n11002 ^ n6532 ^ x0 ;
  assign n11004 = ( n7756 & n8418 ) | ( n7756 & ~n11003 ) | ( n8418 & ~n11003 ) ;
  assign n11005 = n9052 ^ n8320 ^ n6940 ;
  assign n11006 = ( n1370 & ~n5244 ) | ( n1370 & n11005 ) | ( ~n5244 & n11005 ) ;
  assign n11007 = n2562 & ~n11006 ;
  assign n11008 = ( n5121 & n10042 ) | ( n5121 & n11007 ) | ( n10042 & n11007 ) ;
  assign n11009 = ( ~n627 & n4262 ) | ( ~n627 & n11008 ) | ( n4262 & n11008 ) ;
  assign n11010 = n10073 | n11009 ;
  assign n11011 = n10110 ^ n7764 ^ n1827 ;
  assign n11012 = n6443 ^ n967 ^ 1'b0 ;
  assign n11013 = ( n6543 & n6581 ) | ( n6543 & n7597 ) | ( n6581 & n7597 ) ;
  assign n11014 = ( n2549 & ~n6574 ) | ( n2549 & n11013 ) | ( ~n6574 & n11013 ) ;
  assign n11015 = n4235 ^ n3887 ^ n417 ;
  assign n11016 = n3269 & ~n11015 ;
  assign n11017 = n11016 ^ n5981 ^ n3921 ;
  assign n11018 = n727 & ~n11017 ;
  assign n11019 = n10218 | n11018 ;
  assign n11020 = n6138 & ~n11019 ;
  assign n11021 = n11020 ^ n10348 ^ n2821 ;
  assign n11022 = ( n5556 & n11014 ) | ( n5556 & n11021 ) | ( n11014 & n11021 ) ;
  assign n11023 = ( n7242 & ~n8232 ) | ( n7242 & n11022 ) | ( ~n8232 & n11022 ) ;
  assign n11024 = n1627 | n11023 ;
  assign n11025 = n11012 & ~n11024 ;
  assign n11026 = n989 & n8292 ;
  assign n11027 = ~x128 & n11026 ;
  assign n11028 = n5203 | n11027 ;
  assign n11029 = n6957 | n11028 ;
  assign n11030 = n11029 ^ n9480 ^ n2316 ;
  assign n11031 = ~n1254 & n11030 ;
  assign n11032 = n11031 ^ n1457 ^ 1'b0 ;
  assign n11033 = n11032 ^ n8639 ^ 1'b0 ;
  assign n11037 = ~n3352 & n6406 ;
  assign n11034 = ( n2790 & n7802 ) | ( n2790 & ~n10614 ) | ( n7802 & ~n10614 ) ;
  assign n11035 = ( n3621 & n8466 ) | ( n3621 & n11034 ) | ( n8466 & n11034 ) ;
  assign n11036 = n11035 ^ n8523 ^ n3124 ;
  assign n11038 = n11037 ^ n11036 ^ n3268 ;
  assign n11040 = ( ~x185 & n2152 ) | ( ~x185 & n4275 ) | ( n2152 & n4275 ) ;
  assign n11039 = n5470 ^ n1968 ^ n1266 ;
  assign n11041 = n11040 ^ n11039 ^ n10719 ;
  assign n11042 = n11041 ^ n10418 ^ n5255 ;
  assign n11043 = ( n688 & n3522 ) | ( n688 & n9549 ) | ( n3522 & n9549 ) ;
  assign n11044 = ( n7375 & n8107 ) | ( n7375 & ~n11043 ) | ( n8107 & ~n11043 ) ;
  assign n11052 = ( ~n809 & n2402 ) | ( ~n809 & n7132 ) | ( n2402 & n7132 ) ;
  assign n11051 = ( n2997 & n3577 ) | ( n2997 & ~n4936 ) | ( n3577 & ~n4936 ) ;
  assign n11045 = n9190 ^ n726 ^ n684 ;
  assign n11046 = n763 & ~n11045 ;
  assign n11047 = ( n4129 & n5030 ) | ( n4129 & ~n11046 ) | ( n5030 & ~n11046 ) ;
  assign n11048 = ( x104 & n2375 ) | ( x104 & ~n4602 ) | ( n2375 & ~n4602 ) ;
  assign n11049 = ( n4351 & n10063 ) | ( n4351 & n11048 ) | ( n10063 & n11048 ) ;
  assign n11050 = ( ~n8227 & n11047 ) | ( ~n8227 & n11049 ) | ( n11047 & n11049 ) ;
  assign n11053 = n11052 ^ n11051 ^ n11050 ;
  assign n11054 = ( n1485 & n3984 ) | ( n1485 & n4364 ) | ( n3984 & n4364 ) ;
  assign n11055 = n4310 & ~n9609 ;
  assign n11056 = n11054 & n11055 ;
  assign n11057 = n7176 ^ n654 ^ 1'b0 ;
  assign n11058 = ( n5713 & n8232 ) | ( n5713 & n11057 ) | ( n8232 & n11057 ) ;
  assign n11059 = n11058 ^ n9021 ^ x229 ;
  assign n11060 = ( ~n2443 & n6645 ) | ( ~n2443 & n11059 ) | ( n6645 & n11059 ) ;
  assign n11061 = ( n4160 & ~n11056 ) | ( n4160 & n11060 ) | ( ~n11056 & n11060 ) ;
  assign n11062 = ( n11044 & ~n11053 ) | ( n11044 & n11061 ) | ( ~n11053 & n11061 ) ;
  assign n11064 = n9533 ^ n4925 ^ n1749 ;
  assign n11063 = n6985 ^ n6618 ^ n4829 ;
  assign n11065 = n11064 ^ n11063 ^ x169 ;
  assign n11066 = n11065 ^ n8201 ^ n4229 ;
  assign n11067 = n4458 ^ n2473 ^ n595 ;
  assign n11068 = ( n5444 & ~n7086 ) | ( n5444 & n8237 ) | ( ~n7086 & n8237 ) ;
  assign n11069 = ( n9218 & n9733 ) | ( n9218 & n11068 ) | ( n9733 & n11068 ) ;
  assign n11070 = ( ~n9555 & n11067 ) | ( ~n9555 & n11069 ) | ( n11067 & n11069 ) ;
  assign n11071 = n11066 & ~n11070 ;
  assign n11072 = n11071 ^ n9964 ^ 1'b0 ;
  assign n11081 = n3273 ^ n3019 ^ n1391 ;
  assign n11078 = n10531 ^ n4918 ^ n1487 ;
  assign n11079 = n2615 & ~n11078 ;
  assign n11080 = ( n3823 & ~n7526 ) | ( n3823 & n11079 ) | ( ~n7526 & n11079 ) ;
  assign n11073 = ( n3337 & ~n3464 ) | ( n3337 & n5179 ) | ( ~n3464 & n5179 ) ;
  assign n11074 = n9015 ^ n6025 ^ 1'b0 ;
  assign n11075 = n6599 ^ n4051 ^ n2593 ;
  assign n11076 = ( ~n11073 & n11074 ) | ( ~n11073 & n11075 ) | ( n11074 & n11075 ) ;
  assign n11077 = n11076 ^ n5656 ^ n3146 ;
  assign n11082 = n11081 ^ n11080 ^ n11077 ;
  assign n11083 = n8555 ^ n7076 ^ n4096 ;
  assign n11084 = ( n8842 & n11074 ) | ( n8842 & ~n11083 ) | ( n11074 & ~n11083 ) ;
  assign n11085 = n11084 ^ n5058 ^ 1'b0 ;
  assign n11086 = ~n2051 & n11085 ;
  assign n11087 = ( n722 & n4271 ) | ( n722 & ~n9570 ) | ( n4271 & ~n9570 ) ;
  assign n11088 = ( ~n3011 & n3172 ) | ( ~n3011 & n5206 ) | ( n3172 & n5206 ) ;
  assign n11089 = n5944 ^ n4833 ^ n1952 ;
  assign n11090 = ~n1745 & n11089 ;
  assign n11091 = n11090 ^ n3452 ^ n2523 ;
  assign n11092 = ( n2080 & n11088 ) | ( n2080 & n11091 ) | ( n11088 & n11091 ) ;
  assign n11093 = ( n2422 & n11087 ) | ( n2422 & n11092 ) | ( n11087 & n11092 ) ;
  assign n11094 = n8587 ^ n3974 ^ n3461 ;
  assign n11095 = ( ~n2216 & n7055 ) | ( ~n2216 & n8822 ) | ( n7055 & n8822 ) ;
  assign n11096 = ( ~x4 & n11094 ) | ( ~x4 & n11095 ) | ( n11094 & n11095 ) ;
  assign n11102 = ( n539 & ~n596 ) | ( n539 & n897 ) | ( ~n596 & n897 ) ;
  assign n11100 = ( ~n1678 & n1816 ) | ( ~n1678 & n4791 ) | ( n1816 & n4791 ) ;
  assign n11099 = n7882 ^ n2708 ^ n489 ;
  assign n11101 = n11100 ^ n11099 ^ n2852 ;
  assign n11103 = n11102 ^ n11101 ^ n7237 ;
  assign n11097 = ( n1454 & n2769 ) | ( n1454 & ~n3866 ) | ( n2769 & ~n3866 ) ;
  assign n11098 = n11097 ^ n4390 ^ 1'b0 ;
  assign n11104 = n11103 ^ n11098 ^ n7057 ;
  assign n11105 = n11104 ^ n8938 ^ n1571 ;
  assign n11106 = ( n719 & ~n2526 ) | ( n719 & n2949 ) | ( ~n2526 & n2949 ) ;
  assign n11107 = ( ~n288 & n10408 ) | ( ~n288 & n11106 ) | ( n10408 & n11106 ) ;
  assign n11121 = ( n1033 & n5769 ) | ( n1033 & ~n7510 ) | ( n5769 & ~n7510 ) ;
  assign n11122 = n11121 ^ n10628 ^ n8916 ;
  assign n11120 = n2585 & ~n9662 ;
  assign n11118 = n8267 ^ n2593 ^ x173 ;
  assign n11113 = n5993 ^ n5870 ^ n4277 ;
  assign n11114 = n11113 ^ n7067 ^ n683 ;
  assign n11115 = n11114 ^ n8380 ^ n5855 ;
  assign n11108 = x204 & ~n4802 ;
  assign n11109 = n11108 ^ n971 ^ 1'b0 ;
  assign n11110 = ( n1601 & n2776 ) | ( n1601 & ~n11109 ) | ( n2776 & ~n11109 ) ;
  assign n11111 = n11110 ^ n8632 ^ 1'b0 ;
  assign n11112 = n6975 & n11111 ;
  assign n11116 = n11115 ^ n11112 ^ n860 ;
  assign n11117 = n11116 ^ n6863 ^ 1'b0 ;
  assign n11119 = n11118 ^ n11117 ^ n10697 ;
  assign n11123 = n11122 ^ n11120 ^ n11119 ;
  assign n11124 = ( x103 & ~x223 ) | ( x103 & n4676 ) | ( ~x223 & n4676 ) ;
  assign n11125 = ( ~n1689 & n8160 ) | ( ~n1689 & n11124 ) | ( n8160 & n11124 ) ;
  assign n11126 = n11125 ^ n8628 ^ n7953 ;
  assign n11127 = ~n901 & n4858 ;
  assign n11128 = n3198 & n11127 ;
  assign n11129 = ( n3194 & n8066 ) | ( n3194 & n11128 ) | ( n8066 & n11128 ) ;
  assign n11130 = n11129 ^ n9241 ^ n3206 ;
  assign n11131 = ( n2517 & n11126 ) | ( n2517 & n11130 ) | ( n11126 & n11130 ) ;
  assign n11132 = n3782 & n11131 ;
  assign n11140 = ~n2551 & n2850 ;
  assign n11138 = n1130 & ~n8608 ;
  assign n11139 = n11138 ^ n4955 ^ 1'b0 ;
  assign n11141 = n11140 ^ n11139 ^ n10711 ;
  assign n11134 = ( n678 & ~n2713 ) | ( n678 & n5359 ) | ( ~n2713 & n5359 ) ;
  assign n11135 = n11134 ^ n3777 ^ n2306 ;
  assign n11136 = n10437 ^ n6482 ^ 1'b0 ;
  assign n11137 = ( n4732 & n11135 ) | ( n4732 & n11136 ) | ( n11135 & n11136 ) ;
  assign n11133 = ( n5722 & n10065 ) | ( n5722 & ~n10103 ) | ( n10065 & ~n10103 ) ;
  assign n11142 = n11141 ^ n11137 ^ n11133 ;
  assign n11143 = n11142 ^ n9780 ^ n7457 ;
  assign n11144 = n5308 ^ n3849 ^ n1952 ;
  assign n11145 = n4859 & n11144 ;
  assign n11146 = ( n4505 & n8302 ) | ( n4505 & n11145 ) | ( n8302 & n11145 ) ;
  assign n11147 = n2388 & ~n4835 ;
  assign n11148 = n11147 ^ n7665 ^ n5611 ;
  assign n11149 = n6396 ^ n5142 ^ n1637 ;
  assign n11150 = ( n2925 & n11148 ) | ( n2925 & n11149 ) | ( n11148 & n11149 ) ;
  assign n11151 = ( n3575 & n5645 ) | ( n3575 & ~n11150 ) | ( n5645 & ~n11150 ) ;
  assign n11153 = n8668 ^ n6468 ^ n3228 ;
  assign n11154 = n11153 ^ n1298 ^ 1'b0 ;
  assign n11152 = n6684 ^ n3516 ^ n2200 ;
  assign n11155 = n11154 ^ n11152 ^ n9298 ;
  assign n11164 = n6476 ^ n3342 ^ n668 ;
  assign n11159 = ( n529 & n2100 ) | ( n529 & n2456 ) | ( n2100 & n2456 ) ;
  assign n11160 = ( x237 & n406 ) | ( x237 & ~n3922 ) | ( n406 & ~n3922 ) ;
  assign n11161 = n355 & ~n11160 ;
  assign n11162 = ~n11159 & n11161 ;
  assign n11163 = n11162 ^ n9079 ^ n4910 ;
  assign n11156 = n3943 ^ n3592 ^ n2985 ;
  assign n11157 = ( n2778 & n5956 ) | ( n2778 & ~n11156 ) | ( n5956 & ~n11156 ) ;
  assign n11158 = n11157 ^ n3527 ^ n1226 ;
  assign n11165 = n11164 ^ n11163 ^ n11158 ;
  assign n11166 = ( n2747 & n11155 ) | ( n2747 & ~n11165 ) | ( n11155 & ~n11165 ) ;
  assign n11186 = n6567 ^ n4823 ^ 1'b0 ;
  assign n11182 = n6573 ^ n2884 ^ n1170 ;
  assign n11183 = n11182 ^ n4441 ^ n1510 ;
  assign n11184 = ( n5503 & n7455 ) | ( n5503 & ~n11183 ) | ( n7455 & ~n11183 ) ;
  assign n11175 = n2292 ^ n926 ^ n318 ;
  assign n11176 = n5182 | n5201 ;
  assign n11177 = n11176 ^ n437 ^ 1'b0 ;
  assign n11178 = ( n6361 & n9022 ) | ( n6361 & n11177 ) | ( n9022 & n11177 ) ;
  assign n11179 = n3228 | n11178 ;
  assign n11180 = n4676 & ~n11179 ;
  assign n11181 = ( n7093 & n11175 ) | ( n7093 & n11180 ) | ( n11175 & n11180 ) ;
  assign n11185 = n11184 ^ n11181 ^ n3227 ;
  assign n11167 = n4011 ^ n879 ^ n582 ;
  assign n11170 = n4320 ^ n3636 ^ n1211 ;
  assign n11171 = ( ~n1044 & n8822 ) | ( ~n1044 & n11170 ) | ( n8822 & n11170 ) ;
  assign n11168 = n10598 ^ n10118 ^ n5124 ;
  assign n11169 = ( ~n5565 & n6121 ) | ( ~n5565 & n11168 ) | ( n6121 & n11168 ) ;
  assign n11172 = n11171 ^ n11169 ^ n10838 ;
  assign n11173 = n4326 & ~n11172 ;
  assign n11174 = ~n11167 & n11173 ;
  assign n11187 = n11186 ^ n11185 ^ n11174 ;
  assign n11188 = n7771 ^ n6238 ^ 1'b0 ;
  assign n11189 = n6826 & ~n11188 ;
  assign n11190 = n3581 | n4151 ;
  assign n11191 = n11190 ^ n7186 ^ 1'b0 ;
  assign n11192 = ( n4085 & n11189 ) | ( n4085 & n11191 ) | ( n11189 & n11191 ) ;
  assign n11193 = ~n1514 & n5675 ;
  assign n11194 = n11193 ^ n2677 ^ 1'b0 ;
  assign n11195 = ( n1884 & ~n3577 ) | ( n1884 & n11194 ) | ( ~n3577 & n11194 ) ;
  assign n11196 = ( n2992 & ~n5309 ) | ( n2992 & n10135 ) | ( ~n5309 & n10135 ) ;
  assign n11197 = ( ~n6493 & n9316 ) | ( ~n6493 & n11196 ) | ( n9316 & n11196 ) ;
  assign n11198 = ( n1664 & ~n2114 ) | ( n1664 & n11197 ) | ( ~n2114 & n11197 ) ;
  assign n11199 = ( x71 & n1786 ) | ( x71 & ~n2305 ) | ( n1786 & ~n2305 ) ;
  assign n11200 = n11199 ^ n6357 ^ 1'b0 ;
  assign n11201 = n10323 ^ n4472 ^ n2689 ;
  assign n11202 = ( ~n9385 & n11200 ) | ( ~n9385 & n11201 ) | ( n11200 & n11201 ) ;
  assign n11203 = ( n11195 & n11198 ) | ( n11195 & n11202 ) | ( n11198 & n11202 ) ;
  assign n11204 = ( x0 & n4625 ) | ( x0 & n10215 ) | ( n4625 & n10215 ) ;
  assign n11205 = ( n1275 & ~n1663 ) | ( n1275 & n11204 ) | ( ~n1663 & n11204 ) ;
  assign n11206 = ( n558 & n3180 ) | ( n558 & n11205 ) | ( n3180 & n11205 ) ;
  assign n11207 = n5176 ^ n2728 ^ x205 ;
  assign n11208 = ( n870 & ~n4580 ) | ( n870 & n11207 ) | ( ~n4580 & n11207 ) ;
  assign n11209 = n4403 ^ n3590 ^ 1'b0 ;
  assign n11210 = ( n4036 & ~n11208 ) | ( n4036 & n11209 ) | ( ~n11208 & n11209 ) ;
  assign n11216 = ~n972 & n1219 ;
  assign n11214 = n4422 ^ n3645 ^ n2614 ;
  assign n11213 = ( n3015 & ~n4219 ) | ( n3015 & n5171 ) | ( ~n4219 & n5171 ) ;
  assign n11211 = n10220 ^ n8737 ^ n7804 ;
  assign n11212 = n11211 ^ n8535 ^ n736 ;
  assign n11215 = n11214 ^ n11213 ^ n11212 ;
  assign n11217 = n11216 ^ n11215 ^ n4739 ;
  assign n11218 = ( ~n11206 & n11210 ) | ( ~n11206 & n11217 ) | ( n11210 & n11217 ) ;
  assign n11219 = ( n1906 & ~n4031 ) | ( n1906 & n8849 ) | ( ~n4031 & n8849 ) ;
  assign n11220 = ( n1622 & n2333 ) | ( n1622 & ~n8122 ) | ( n2333 & ~n8122 ) ;
  assign n11224 = n8509 ^ n5700 ^ n424 ;
  assign n11225 = ( n1030 & n7239 ) | ( n1030 & n11224 ) | ( n7239 & n11224 ) ;
  assign n11221 = n3347 ^ n3153 ^ n1505 ;
  assign n11222 = n11221 ^ x40 ^ 1'b0 ;
  assign n11223 = n1622 | n11222 ;
  assign n11226 = n11225 ^ n11223 ^ n10640 ;
  assign n11227 = n875 | n11226 ;
  assign n11228 = n10900 & ~n11227 ;
  assign n11229 = ( n11219 & n11220 ) | ( n11219 & n11228 ) | ( n11220 & n11228 ) ;
  assign n11233 = n10612 ^ n9241 ^ n1272 ;
  assign n11234 = ( n742 & n10658 ) | ( n742 & ~n11233 ) | ( n10658 & ~n11233 ) ;
  assign n11230 = ( n3702 & ~n4242 ) | ( n3702 & n10059 ) | ( ~n4242 & n10059 ) ;
  assign n11231 = ( ~n5843 & n7113 ) | ( ~n5843 & n11230 ) | ( n7113 & n11230 ) ;
  assign n11232 = n11231 ^ n10308 ^ n1384 ;
  assign n11235 = n11234 ^ n11232 ^ n5540 ;
  assign n11236 = n11235 ^ n10917 ^ n10909 ;
  assign n11237 = ( x66 & ~n1046 ) | ( x66 & n6643 ) | ( ~n1046 & n6643 ) ;
  assign n11238 = ( n1777 & n3181 ) | ( n1777 & n3573 ) | ( n3181 & n3573 ) ;
  assign n11239 = n11238 ^ n9082 ^ n681 ;
  assign n11240 = n11237 & ~n11239 ;
  assign n11255 = n5600 & ~n10504 ;
  assign n11251 = n4885 ^ n2086 ^ 1'b0 ;
  assign n11252 = n10973 | n11251 ;
  assign n11253 = n5263 ^ n1467 ^ 1'b0 ;
  assign n11254 = n11252 | n11253 ;
  assign n11256 = n11255 ^ n11254 ^ n872 ;
  assign n11249 = n5160 ^ n2012 ^ 1'b0 ;
  assign n11250 = n9338 | n11249 ;
  assign n11257 = n11256 ^ n11250 ^ 1'b0 ;
  assign n11247 = ( x120 & n2286 ) | ( x120 & n2692 ) | ( n2286 & n2692 ) ;
  assign n11241 = n8472 ^ n5759 ^ n2017 ;
  assign n11242 = ( n561 & n5148 ) | ( n561 & n11241 ) | ( n5148 & n11241 ) ;
  assign n11243 = n4599 | n8488 ;
  assign n11244 = n2302 | n11243 ;
  assign n11245 = n11244 ^ n2507 ^ x76 ;
  assign n11246 = n11242 & ~n11245 ;
  assign n11248 = n11247 ^ n11246 ^ 1'b0 ;
  assign n11258 = n11257 ^ n11248 ^ 1'b0 ;
  assign n11259 = ( n6849 & n10512 ) | ( n6849 & n11258 ) | ( n10512 & n11258 ) ;
  assign n11260 = n8810 ^ n2689 ^ x95 ;
  assign n11263 = ( n365 & n2205 ) | ( n365 & ~n10504 ) | ( n2205 & ~n10504 ) ;
  assign n11261 = n574 & ~n4245 ;
  assign n11262 = n6906 & n11261 ;
  assign n11264 = n11263 ^ n11262 ^ n491 ;
  assign n11265 = n11264 ^ n3255 ^ 1'b0 ;
  assign n11266 = n11265 ^ n6353 ^ n3786 ;
  assign n11267 = ( ~n5475 & n10658 ) | ( ~n5475 & n10941 ) | ( n10658 & n10941 ) ;
  assign n11268 = ( n9006 & ~n11266 ) | ( n9006 & n11267 ) | ( ~n11266 & n11267 ) ;
  assign n11269 = ( ~n4436 & n6316 ) | ( ~n4436 & n11268 ) | ( n6316 & n11268 ) ;
  assign n11270 = n6145 & ~n11269 ;
  assign n11271 = n11270 ^ n9615 ^ n2749 ;
  assign n11272 = ( n1158 & n3382 ) | ( n1158 & n3779 ) | ( n3382 & n3779 ) ;
  assign n11273 = n585 | n11272 ;
  assign n11274 = n4366 | n11273 ;
  assign n11275 = ( n7073 & n10882 ) | ( n7073 & ~n11274 ) | ( n10882 & ~n11274 ) ;
  assign n11276 = n9846 ^ n4728 ^ n4111 ;
  assign n11277 = n11276 ^ n7135 ^ 1'b0 ;
  assign n11278 = ~n912 & n8053 ;
  assign n11279 = n7206 & n11278 ;
  assign n11280 = ( n2747 & n8104 ) | ( n2747 & n11279 ) | ( n8104 & n11279 ) ;
  assign n11281 = n5530 ^ n4231 ^ x120 ;
  assign n11282 = n6848 ^ n2307 ^ x203 ;
  assign n11283 = n11282 ^ n1934 ^ n1539 ;
  assign n11284 = ( n11280 & n11281 ) | ( n11280 & ~n11283 ) | ( n11281 & ~n11283 ) ;
  assign n11285 = ( n11275 & n11277 ) | ( n11275 & ~n11284 ) | ( n11277 & ~n11284 ) ;
  assign n11287 = n1835 & n6369 ;
  assign n11288 = ( n1170 & ~n6791 ) | ( n1170 & n11287 ) | ( ~n6791 & n11287 ) ;
  assign n11289 = ( ~n476 & n8269 ) | ( ~n476 & n11288 ) | ( n8269 & n11288 ) ;
  assign n11286 = n3847 ^ n1523 ^ x155 ;
  assign n11290 = n11289 ^ n11286 ^ n9279 ;
  assign n11291 = ~n548 & n1965 ;
  assign n11292 = n11291 ^ n4981 ^ n3090 ;
  assign n11293 = ( x10 & n4636 ) | ( x10 & n6491 ) | ( n4636 & n6491 ) ;
  assign n11294 = n11293 ^ n2016 ^ 1'b0 ;
  assign n11295 = n11292 & n11294 ;
  assign n11296 = n8372 ^ n2243 ^ x92 ;
  assign n11297 = ( ~n6045 & n8632 ) | ( ~n6045 & n11296 ) | ( n8632 & n11296 ) ;
  assign n11300 = n1312 & ~n1582 ;
  assign n11298 = n9398 ^ n5386 ^ n2331 ;
  assign n11299 = n11298 ^ n1988 ^ n1690 ;
  assign n11301 = n11300 ^ n11299 ^ 1'b0 ;
  assign n11302 = ( ~n8140 & n11297 ) | ( ~n8140 & n11301 ) | ( n11297 & n11301 ) ;
  assign n11303 = ( x148 & ~n3243 ) | ( x148 & n9542 ) | ( ~n3243 & n9542 ) ;
  assign n11304 = n9597 ^ n5743 ^ n4180 ;
  assign n11306 = ( n574 & n1423 ) | ( n574 & n2881 ) | ( n1423 & n2881 ) ;
  assign n11305 = x236 & ~n7249 ;
  assign n11307 = n11306 ^ n11305 ^ 1'b0 ;
  assign n11308 = ( n10819 & n11304 ) | ( n10819 & n11307 ) | ( n11304 & n11307 ) ;
  assign n11309 = n11303 & ~n11308 ;
  assign n11318 = n3123 ^ n3000 ^ n1175 ;
  assign n11312 = ~n4729 & n8619 ;
  assign n11313 = x28 & ~n8256 ;
  assign n11314 = n11313 ^ n4950 ^ 1'b0 ;
  assign n11315 = n11314 ^ n2893 ^ n1924 ;
  assign n11316 = ~n11312 & n11315 ;
  assign n11317 = n288 & n11316 ;
  assign n11310 = n8776 ^ n5417 ^ 1'b0 ;
  assign n11311 = n11310 ^ n9900 ^ n8880 ;
  assign n11319 = n11318 ^ n11317 ^ n11311 ;
  assign n11320 = ( ~x137 & n9693 ) | ( ~x137 & n11319 ) | ( n9693 & n11319 ) ;
  assign n11327 = n7527 ^ n4100 ^ n2198 ;
  assign n11328 = ( n1553 & n4018 ) | ( n1553 & n11327 ) | ( n4018 & n11327 ) ;
  assign n11322 = n8372 ^ n2125 ^ n2058 ;
  assign n11323 = ( n2067 & n10515 ) | ( n2067 & n11322 ) | ( n10515 & n11322 ) ;
  assign n11324 = ~n5067 & n11323 ;
  assign n11325 = n1503 & n11324 ;
  assign n11321 = n4122 | n7815 ;
  assign n11326 = n11325 ^ n11321 ^ n7472 ;
  assign n11329 = n11328 ^ n11326 ^ n6008 ;
  assign n11330 = ( ~n3688 & n4027 ) | ( ~n3688 & n11329 ) | ( n4027 & n11329 ) ;
  assign n11331 = n10377 ^ n9496 ^ n2508 ;
  assign n11332 = ( n904 & ~n6417 ) | ( n904 & n7290 ) | ( ~n6417 & n7290 ) ;
  assign n11333 = n11332 ^ n8220 ^ n6735 ;
  assign n11341 = ( n743 & n6378 ) | ( n743 & ~n9072 ) | ( n6378 & ~n9072 ) ;
  assign n11342 = n5479 ^ n857 ^ n772 ;
  assign n11343 = n11342 ^ n2316 ^ n904 ;
  assign n11344 = ( ~n1822 & n11341 ) | ( ~n1822 & n11343 ) | ( n11341 & n11343 ) ;
  assign n11337 = n2001 ^ n485 ^ x44 ;
  assign n11338 = ( ~n1165 & n1385 ) | ( ~n1165 & n11337 ) | ( n1385 & n11337 ) ;
  assign n11335 = n10442 ^ n7219 ^ n3207 ;
  assign n11336 = n11335 ^ n7484 ^ n6013 ;
  assign n11334 = n6690 ^ n4551 ^ n4223 ;
  assign n11339 = n11338 ^ n11336 ^ n11334 ;
  assign n11340 = ( n4390 & n8674 ) | ( n4390 & ~n11339 ) | ( n8674 & ~n11339 ) ;
  assign n11345 = n11344 ^ n11340 ^ n9453 ;
  assign n11350 = n6298 ^ n935 ^ n736 ;
  assign n11351 = n5255 ^ n901 ^ 1'b0 ;
  assign n11352 = n11350 & ~n11351 ;
  assign n11353 = ( n5635 & n6240 ) | ( n5635 & n11352 ) | ( n6240 & n11352 ) ;
  assign n11348 = ( n2747 & n4031 ) | ( n2747 & ~n4370 ) | ( n4031 & ~n4370 ) ;
  assign n11346 = n11054 ^ n4738 ^ 1'b0 ;
  assign n11347 = ( n7513 & ~n8707 ) | ( n7513 & n11346 ) | ( ~n8707 & n11346 ) ;
  assign n11349 = n11348 ^ n11347 ^ n1992 ;
  assign n11354 = n11353 ^ n11349 ^ x92 ;
  assign n11355 = ( n974 & n11345 ) | ( n974 & n11354 ) | ( n11345 & n11354 ) ;
  assign n11356 = n4834 ^ n4037 ^ n854 ;
  assign n11357 = n11356 ^ n6415 ^ n1836 ;
  assign n11358 = ( n636 & n9465 ) | ( n636 & n10113 ) | ( n9465 & n10113 ) ;
  assign n11363 = n5122 ^ n1531 ^ n828 ;
  assign n11362 = ( n438 & ~n3013 ) | ( n438 & n3569 ) | ( ~n3013 & n3569 ) ;
  assign n11364 = n11363 ^ n11362 ^ n1060 ;
  assign n11365 = n11364 ^ n10144 ^ n1776 ;
  assign n11359 = ( n4308 & n5066 ) | ( n4308 & n11195 ) | ( n5066 & n11195 ) ;
  assign n11360 = ( n5935 & ~n8739 ) | ( n5935 & n11359 ) | ( ~n8739 & n11359 ) ;
  assign n11361 = n11360 ^ n7610 ^ n5923 ;
  assign n11366 = n11365 ^ n11361 ^ 1'b0 ;
  assign n11367 = ~n11358 & n11366 ;
  assign n11368 = ( x85 & n11357 ) | ( x85 & n11367 ) | ( n11357 & n11367 ) ;
  assign n11369 = n3249 & ~n8560 ;
  assign n11370 = ~n4908 & n11369 ;
  assign n11371 = n9779 ^ n4750 ^ 1'b0 ;
  assign n11372 = ~n11370 & n11371 ;
  assign n11375 = ( ~n1252 & n3008 ) | ( ~n1252 & n5113 ) | ( n3008 & n5113 ) ;
  assign n11376 = n11375 ^ n10251 ^ n9433 ;
  assign n11373 = n8315 & n8818 ;
  assign n11374 = n11373 ^ n3015 ^ n2843 ;
  assign n11377 = n11376 ^ n11374 ^ n6333 ;
  assign n11378 = n2438 ^ n1704 ^ 1'b0 ;
  assign n11379 = n3213 & n11378 ;
  assign n11380 = n3073 ^ n2160 ^ 1'b0 ;
  assign n11381 = ( n371 & n1823 ) | ( n371 & n3779 ) | ( n1823 & n3779 ) ;
  assign n11382 = ( n4516 & n11380 ) | ( n4516 & n11381 ) | ( n11380 & n11381 ) ;
  assign n11383 = ( n3127 & n10487 ) | ( n3127 & ~n11382 ) | ( n10487 & ~n11382 ) ;
  assign n11384 = n7835 ^ n4956 ^ 1'b0 ;
  assign n11385 = ( n11379 & n11383 ) | ( n11379 & n11384 ) | ( n11383 & n11384 ) ;
  assign n11386 = ( n4379 & n11377 ) | ( n4379 & n11385 ) | ( n11377 & n11385 ) ;
  assign n11387 = n2152 ^ n851 ^ 1'b0 ;
  assign n11388 = ~n534 & n11387 ;
  assign n11389 = n11388 ^ n4680 ^ n530 ;
  assign n11394 = ~n2081 & n5907 ;
  assign n11395 = ~n773 & n11394 ;
  assign n11396 = ( n1521 & n4636 ) | ( n1521 & ~n8037 ) | ( n4636 & ~n8037 ) ;
  assign n11397 = ( n5983 & n11395 ) | ( n5983 & ~n11396 ) | ( n11395 & ~n11396 ) ;
  assign n11392 = n10640 ^ n2273 ^ n1563 ;
  assign n11390 = n1510 & ~n5791 ;
  assign n11391 = n7290 | n11390 ;
  assign n11393 = n11392 ^ n11391 ^ n2595 ;
  assign n11398 = n11397 ^ n11393 ^ n4520 ;
  assign n11399 = ( n7551 & n11389 ) | ( n7551 & ~n11398 ) | ( n11389 & ~n11398 ) ;
  assign n11407 = ( x39 & n5175 ) | ( x39 & ~n6451 ) | ( n5175 & ~n6451 ) ;
  assign n11408 = ( ~x230 & n835 ) | ( ~x230 & n11407 ) | ( n835 & n11407 ) ;
  assign n11401 = n5073 ^ n896 ^ n632 ;
  assign n11402 = ( n1264 & ~n10842 ) | ( n1264 & n11401 ) | ( ~n10842 & n11401 ) ;
  assign n11403 = ~n823 & n11402 ;
  assign n11404 = n11403 ^ n340 ^ 1'b0 ;
  assign n11400 = n7609 ^ n3960 ^ n2962 ;
  assign n11405 = n11404 ^ n11400 ^ n2975 ;
  assign n11406 = n11405 ^ n8088 ^ n5691 ;
  assign n11409 = n11408 ^ n11406 ^ n4309 ;
  assign n11410 = n6757 ^ n4001 ^ n1537 ;
  assign n11411 = ~n4343 & n4932 ;
  assign n11412 = ( n1446 & n11410 ) | ( n1446 & ~n11411 ) | ( n11410 & ~n11411 ) ;
  assign n11413 = n4177 ^ n4074 ^ n2911 ;
  assign n11414 = n11413 ^ n11238 ^ 1'b0 ;
  assign n11415 = n3238 & n11414 ;
  assign n11416 = ( n2624 & n7020 ) | ( n2624 & ~n7650 ) | ( n7020 & ~n7650 ) ;
  assign n11417 = n11415 & n11416 ;
  assign n11420 = n9627 ^ n5767 ^ n2497 ;
  assign n11418 = n469 | n7411 ;
  assign n11419 = n3948 & ~n11418 ;
  assign n11421 = n11420 ^ n11419 ^ n5621 ;
  assign n11422 = n4271 ^ n640 ^ x237 ;
  assign n11423 = n1540 ^ n720 ^ 1'b0 ;
  assign n11424 = ~n1033 & n11423 ;
  assign n11425 = n11424 ^ n3454 ^ n2347 ;
  assign n11426 = ( n8854 & ~n11422 ) | ( n8854 & n11425 ) | ( ~n11422 & n11425 ) ;
  assign n11427 = ( ~n5150 & n5470 ) | ( ~n5150 & n11426 ) | ( n5470 & n11426 ) ;
  assign n11428 = n4897 ^ n1613 ^ 1'b0 ;
  assign n11438 = ( n2211 & n3866 ) | ( n2211 & ~n8031 ) | ( n3866 & ~n8031 ) ;
  assign n11437 = n10708 ^ n5586 ^ n2408 ;
  assign n11429 = n3908 ^ n431 ^ 1'b0 ;
  assign n11430 = ( ~n266 & n3307 ) | ( ~n266 & n6669 ) | ( n3307 & n6669 ) ;
  assign n11431 = n2196 ^ n1419 ^ n332 ;
  assign n11432 = n11430 & n11431 ;
  assign n11433 = ~n11429 & n11432 ;
  assign n11434 = n11433 ^ n7400 ^ n3983 ;
  assign n11435 = n11434 ^ n5135 ^ 1'b0 ;
  assign n11436 = x185 & n11435 ;
  assign n11439 = n11438 ^ n11437 ^ n11436 ;
  assign n11440 = ( ~n11427 & n11428 ) | ( ~n11427 & n11439 ) | ( n11428 & n11439 ) ;
  assign n11442 = n1153 | n1609 ;
  assign n11443 = n11442 ^ n10641 ^ n5149 ;
  assign n11441 = ( n1881 & n4078 ) | ( n1881 & ~n4309 ) | ( n4078 & ~n4309 ) ;
  assign n11444 = n11443 ^ n11441 ^ n11264 ;
  assign n11445 = n11444 ^ n10579 ^ n4324 ;
  assign n11446 = n8880 ^ n7007 ^ n6388 ;
  assign n11447 = n4509 & ~n11446 ;
  assign n11448 = n11447 ^ n11077 ^ 1'b0 ;
  assign n11449 = n11448 ^ n9224 ^ n1944 ;
  assign n11450 = n6079 ^ n3820 ^ n3297 ;
  assign n11451 = ( n4010 & ~n4748 ) | ( n4010 & n11450 ) | ( ~n4748 & n11450 ) ;
  assign n11454 = n8429 ^ n3981 ^ n1182 ;
  assign n11452 = n9428 ^ n5536 ^ n1603 ;
  assign n11453 = ( ~n1084 & n10354 ) | ( ~n1084 & n11452 ) | ( n10354 & n11452 ) ;
  assign n11455 = n11454 ^ n11453 ^ 1'b0 ;
  assign n11456 = n11451 & ~n11455 ;
  assign n11457 = n11247 ^ n10152 ^ n1856 ;
  assign n11458 = ( n6292 & n10179 ) | ( n6292 & n11457 ) | ( n10179 & n11457 ) ;
  assign n11460 = n9287 ^ n8531 ^ n7540 ;
  assign n11459 = n791 & ~n5303 ;
  assign n11461 = n11460 ^ n11459 ^ 1'b0 ;
  assign n11462 = ( n691 & ~n2767 ) | ( n691 & n3103 ) | ( ~n2767 & n3103 ) ;
  assign n11463 = n11462 ^ n8219 ^ 1'b0 ;
  assign n11464 = n3753 ^ n2992 ^ n1961 ;
  assign n11465 = ( n1232 & ~n9888 ) | ( n1232 & n11464 ) | ( ~n9888 & n11464 ) ;
  assign n11466 = n11465 ^ n11286 ^ n5142 ;
  assign n11471 = ( ~n1111 & n3635 ) | ( ~n1111 & n4680 ) | ( n3635 & n4680 ) ;
  assign n11470 = n639 | n6095 ;
  assign n11467 = x227 & n947 ;
  assign n11468 = n11467 ^ x157 ^ 1'b0 ;
  assign n11469 = n11468 ^ n5960 ^ n2244 ;
  assign n11472 = n11471 ^ n11470 ^ n11469 ;
  assign n11477 = n7955 ^ n6238 ^ n2935 ;
  assign n11473 = ( n593 & n1124 ) | ( n593 & n1271 ) | ( n1124 & n1271 ) ;
  assign n11474 = n2027 ^ n1666 ^ 1'b0 ;
  assign n11475 = n1416 & n11474 ;
  assign n11476 = n11473 & ~n11475 ;
  assign n11478 = n11477 ^ n11476 ^ 1'b0 ;
  assign n11479 = ( ~n6002 & n6558 ) | ( ~n6002 & n10973 ) | ( n6558 & n10973 ) ;
  assign n11480 = n6782 & ~n11479 ;
  assign n11481 = n11480 ^ n6980 ^ 1'b0 ;
  assign n11482 = ( n4245 & n7574 ) | ( n4245 & n11481 ) | ( n7574 & n11481 ) ;
  assign n11483 = ( ~n6027 & n6865 ) | ( ~n6027 & n6867 ) | ( n6865 & n6867 ) ;
  assign n11484 = ( ~n1077 & n1469 ) | ( ~n1077 & n3468 ) | ( n1469 & n3468 ) ;
  assign n11485 = ( n1446 & ~n2588 ) | ( n1446 & n11484 ) | ( ~n2588 & n11484 ) ;
  assign n11486 = x8 & n539 ;
  assign n11487 = n5895 & n11486 ;
  assign n11488 = ( n1838 & n6793 ) | ( n1838 & n7373 ) | ( n6793 & n7373 ) ;
  assign n11489 = n11488 ^ n6897 ^ 1'b0 ;
  assign n11490 = n11487 | n11489 ;
  assign n11491 = ( ~n11483 & n11485 ) | ( ~n11483 & n11490 ) | ( n11485 & n11490 ) ;
  assign n11492 = ( n4897 & ~n11482 ) | ( n4897 & n11491 ) | ( ~n11482 & n11491 ) ;
  assign n11493 = n11492 ^ n9060 ^ n5735 ;
  assign n11494 = n11493 ^ n4611 ^ n2846 ;
  assign n11495 = n11494 ^ n9063 ^ 1'b0 ;
  assign n11496 = n11478 | n11495 ;
  assign n11497 = ( n395 & n1959 ) | ( n395 & n8070 ) | ( n1959 & n8070 ) ;
  assign n11498 = ( ~n6565 & n8660 ) | ( ~n6565 & n11497 ) | ( n8660 & n11497 ) ;
  assign n11499 = n4608 ^ n3045 ^ n2250 ;
  assign n11500 = ( ~n1494 & n5710 ) | ( ~n1494 & n11499 ) | ( n5710 & n11499 ) ;
  assign n11501 = ( n1677 & n10465 ) | ( n1677 & ~n11500 ) | ( n10465 & ~n11500 ) ;
  assign n11502 = ( n2264 & ~n3022 ) | ( n2264 & n11501 ) | ( ~n3022 & n11501 ) ;
  assign n11503 = ( n760 & n11498 ) | ( n760 & ~n11502 ) | ( n11498 & ~n11502 ) ;
  assign n11504 = n10133 | n11503 ;
  assign n11505 = ~n3116 & n3160 ;
  assign n11506 = n3282 ^ n2220 ^ 1'b0 ;
  assign n11507 = ( n4816 & n6216 ) | ( n4816 & n11506 ) | ( n6216 & n11506 ) ;
  assign n11508 = n9466 ^ n7476 ^ n1219 ;
  assign n11509 = n5014 & ~n11508 ;
  assign n11510 = n11507 & n11509 ;
  assign n11511 = ( ~n6439 & n11505 ) | ( ~n6439 & n11510 ) | ( n11505 & n11510 ) ;
  assign n11512 = n11511 ^ n2099 ^ n1739 ;
  assign n11516 = ( ~n4061 & n4133 ) | ( ~n4061 & n6420 ) | ( n4133 & n6420 ) ;
  assign n11513 = n1100 & n8112 ;
  assign n11514 = n11513 ^ n11481 ^ 1'b0 ;
  assign n11515 = ( n885 & n5004 ) | ( n885 & n11514 ) | ( n5004 & n11514 ) ;
  assign n11517 = n11516 ^ n11515 ^ n1195 ;
  assign n11518 = n10625 & n11517 ;
  assign n11519 = n3887 & n9251 ;
  assign n11526 = n7496 ^ n6607 ^ n5441 ;
  assign n11527 = n1074 | n5115 ;
  assign n11528 = n11527 ^ n445 ^ 1'b0 ;
  assign n11529 = ( n832 & ~n3820 ) | ( n832 & n11528 ) | ( ~n3820 & n11528 ) ;
  assign n11530 = n11529 ^ n10602 ^ 1'b0 ;
  assign n11531 = ( n7914 & n11526 ) | ( n7914 & n11530 ) | ( n11526 & n11530 ) ;
  assign n11520 = n2692 ^ n1587 ^ n435 ;
  assign n11521 = n5050 ^ n400 ^ 1'b0 ;
  assign n11522 = n11521 ^ n2614 ^ n1289 ;
  assign n11523 = ( n11464 & n11520 ) | ( n11464 & ~n11522 ) | ( n11520 & ~n11522 ) ;
  assign n11524 = n11523 ^ n9850 ^ n6071 ;
  assign n11525 = ( n2429 & n3205 ) | ( n2429 & ~n11524 ) | ( n3205 & ~n11524 ) ;
  assign n11532 = n11531 ^ n11525 ^ 1'b0 ;
  assign n11533 = n7859 | n11532 ;
  assign n11534 = n6905 | n10160 ;
  assign n11535 = n11534 ^ n1153 ^ 1'b0 ;
  assign n11536 = n11535 ^ n9812 ^ n2353 ;
  assign n11537 = n10107 ^ n6316 ^ n1059 ;
  assign n11538 = ( n990 & n2817 ) | ( n990 & ~n6581 ) | ( n2817 & ~n6581 ) ;
  assign n11539 = n10277 ^ n4198 ^ n1647 ;
  assign n11540 = ( ~n2130 & n11538 ) | ( ~n2130 & n11539 ) | ( n11538 & n11539 ) ;
  assign n11541 = ~n5319 & n8378 ;
  assign n11542 = n7468 & n11541 ;
  assign n11543 = n11542 ^ n10392 ^ n2649 ;
  assign n11544 = ( n2714 & ~n4293 ) | ( n2714 & n11543 ) | ( ~n4293 & n11543 ) ;
  assign n11546 = ( n4210 & n4336 ) | ( n4210 & ~n6327 ) | ( n4336 & ~n6327 ) ;
  assign n11545 = ~n758 & n3886 ;
  assign n11547 = n11546 ^ n11545 ^ 1'b0 ;
  assign n11548 = ( n3147 & ~n5596 ) | ( n3147 & n10721 ) | ( ~n5596 & n10721 ) ;
  assign n11549 = n7524 ^ n4439 ^ n376 ;
  assign n11550 = ~n590 & n5298 ;
  assign n11551 = n11550 ^ n3335 ^ 1'b0 ;
  assign n11552 = n11551 ^ n5836 ^ n5216 ;
  assign n11553 = n4939 ^ n3183 ^ n921 ;
  assign n11554 = ( n2944 & n5387 ) | ( n2944 & n10538 ) | ( n5387 & n10538 ) ;
  assign n11555 = ( n11552 & n11553 ) | ( n11552 & n11554 ) | ( n11553 & n11554 ) ;
  assign n11557 = n8345 ^ n3227 ^ n2694 ;
  assign n11556 = n9143 ^ n6270 ^ x4 ;
  assign n11558 = n11557 ^ n11556 ^ n5091 ;
  assign n11559 = n11558 ^ n7397 ^ n5098 ;
  assign n11560 = ( n11549 & ~n11555 ) | ( n11549 & n11559 ) | ( ~n11555 & n11559 ) ;
  assign n11561 = n7637 ^ n1476 ^ n359 ;
  assign n11562 = ( n2360 & n2641 ) | ( n2360 & ~n8098 ) | ( n2641 & ~n8098 ) ;
  assign n11563 = n5930 & n8119 ;
  assign n11564 = n11563 ^ n6484 ^ x92 ;
  assign n11565 = n11562 & n11564 ;
  assign n11569 = ( x11 & ~n5134 ) | ( x11 & n7910 ) | ( ~n5134 & n7910 ) ;
  assign n11568 = ( ~n5559 & n8669 ) | ( ~n5559 & n10105 ) | ( n8669 & n10105 ) ;
  assign n11566 = ( n907 & n1750 ) | ( n907 & ~n7110 ) | ( n1750 & ~n7110 ) ;
  assign n11567 = n11566 ^ n3948 ^ n3588 ;
  assign n11570 = n11569 ^ n11568 ^ n11567 ;
  assign n11571 = ( n497 & ~n1983 ) | ( n497 & n3578 ) | ( ~n1983 & n3578 ) ;
  assign n11572 = ( n582 & n11516 ) | ( n582 & n11571 ) | ( n11516 & n11571 ) ;
  assign n11578 = ( ~n317 & n5652 ) | ( ~n317 & n6261 ) | ( n5652 & n6261 ) ;
  assign n11574 = n6148 ^ n2385 ^ n2336 ;
  assign n11575 = n11574 ^ n5091 ^ n3479 ;
  assign n11576 = n11575 ^ n6938 ^ n5734 ;
  assign n11577 = ( n2872 & ~n7576 ) | ( n2872 & n11576 ) | ( ~n7576 & n11576 ) ;
  assign n11579 = n11578 ^ n11577 ^ n6318 ;
  assign n11580 = ~n11147 & n11579 ;
  assign n11573 = ( n6244 & n6667 ) | ( n6244 & n10815 ) | ( n6667 & n10815 ) ;
  assign n11581 = n11580 ^ n11573 ^ n713 ;
  assign n11582 = n4582 ^ n4487 ^ n1993 ;
  assign n11583 = n11582 ^ n9937 ^ n2338 ;
  assign n11584 = n11583 ^ n6244 ^ n5799 ;
  assign n11585 = n7473 ^ n3659 ^ x221 ;
  assign n11586 = n11585 ^ n3307 ^ n2369 ;
  assign n11587 = n9366 ^ n4536 ^ n2410 ;
  assign n11588 = n2682 ^ n2564 ^ n937 ;
  assign n11589 = n1622 ^ n1443 ^ n1248 ;
  assign n11590 = ( n1945 & ~n3757 ) | ( n1945 & n11589 ) | ( ~n3757 & n11589 ) ;
  assign n11591 = ( n1000 & n11588 ) | ( n1000 & ~n11590 ) | ( n11588 & ~n11590 ) ;
  assign n11592 = ( n8059 & ~n11587 ) | ( n8059 & n11591 ) | ( ~n11587 & n11591 ) ;
  assign n11593 = n11592 ^ n11304 ^ 1'b0 ;
  assign n11594 = n11586 | n11593 ;
  assign n11596 = n6573 ^ n590 ^ n372 ;
  assign n11595 = ( ~n448 & n5731 ) | ( ~n448 & n7438 ) | ( n5731 & n7438 ) ;
  assign n11597 = n11596 ^ n11595 ^ n8425 ;
  assign n11598 = n11597 ^ n8842 ^ 1'b0 ;
  assign n11599 = n299 | n11007 ;
  assign n11600 = ( n2468 & n6741 ) | ( n2468 & n11599 ) | ( n6741 & n11599 ) ;
  assign n11601 = n7438 | n11600 ;
  assign n11602 = n11601 ^ n5175 ^ 1'b0 ;
  assign n11603 = n3488 & n11087 ;
  assign n11604 = n11603 ^ x69 ^ 1'b0 ;
  assign n11605 = n8293 ^ n2826 ^ 1'b0 ;
  assign n11606 = ( n7398 & n7615 ) | ( n7398 & n11557 ) | ( n7615 & n11557 ) ;
  assign n11607 = ( n4038 & n11605 ) | ( n4038 & n11606 ) | ( n11605 & n11606 ) ;
  assign n11608 = n11604 | n11607 ;
  assign n11609 = n11602 & ~n11608 ;
  assign n11614 = n10921 ^ n8140 ^ n2201 ;
  assign n11612 = n5126 & n10782 ;
  assign n11613 = n11612 ^ n10772 ^ n3090 ;
  assign n11615 = n11614 ^ n11613 ^ n954 ;
  assign n11610 = ( n431 & n2804 ) | ( n431 & ~n8928 ) | ( n2804 & ~n8928 ) ;
  assign n11611 = n11610 ^ n6522 ^ n3898 ;
  assign n11616 = n11615 ^ n11611 ^ n2398 ;
  assign n11621 = n5503 | n8563 ;
  assign n11622 = n11621 ^ n4459 ^ 1'b0 ;
  assign n11617 = ( n5028 & ~n8742 ) | ( n5028 & n9188 ) | ( ~n8742 & n9188 ) ;
  assign n11618 = n11617 ^ n1309 ^ n817 ;
  assign n11619 = ( ~n5314 & n6552 ) | ( ~n5314 & n11291 ) | ( n6552 & n11291 ) ;
  assign n11620 = ( n8667 & ~n11618 ) | ( n8667 & n11619 ) | ( ~n11618 & n11619 ) ;
  assign n11623 = n11622 ^ n11620 ^ n8931 ;
  assign n11624 = ( n893 & n1370 ) | ( n893 & n2098 ) | ( n1370 & n2098 ) ;
  assign n11625 = ( n3598 & n5819 ) | ( n3598 & n6244 ) | ( n5819 & n6244 ) ;
  assign n11626 = n11624 & n11625 ;
  assign n11629 = n10713 ^ n1415 ^ 1'b0 ;
  assign n11630 = n2528 & ~n11629 ;
  assign n11627 = n6211 ^ n6119 ^ n6115 ;
  assign n11628 = n7166 & ~n11627 ;
  assign n11631 = n11630 ^ n11628 ^ 1'b0 ;
  assign n11632 = n4905 & n7790 ;
  assign n11633 = n11632 ^ n2576 ^ n667 ;
  assign n11634 = ( ~n2367 & n5675 ) | ( ~n2367 & n8011 ) | ( n5675 & n8011 ) ;
  assign n11635 = n11634 ^ n10181 ^ n6694 ;
  assign n11636 = n8682 & ~n11635 ;
  assign n11637 = ( x68 & ~n1373 ) | ( x68 & n11636 ) | ( ~n1373 & n11636 ) ;
  assign n11638 = ( n1809 & ~n11633 ) | ( n1809 & n11637 ) | ( ~n11633 & n11637 ) ;
  assign n11639 = n6520 ^ n5782 ^ n5131 ;
  assign n11640 = ( ~n4970 & n6907 ) | ( ~n4970 & n9190 ) | ( n6907 & n9190 ) ;
  assign n11641 = n11640 ^ n721 ^ 1'b0 ;
  assign n11642 = n11641 ^ n918 ^ 1'b0 ;
  assign n11643 = ~n5591 & n11642 ;
  assign n11644 = ~n11639 & n11643 ;
  assign n11650 = n7672 ^ n3818 ^ n1839 ;
  assign n11645 = ( n4691 & n5069 ) | ( n4691 & ~n10477 ) | ( n5069 & ~n10477 ) ;
  assign n11646 = ( x206 & n4107 ) | ( x206 & ~n11645 ) | ( n4107 & ~n11645 ) ;
  assign n11647 = ( n3997 & ~n5027 ) | ( n3997 & n7350 ) | ( ~n5027 & n7350 ) ;
  assign n11648 = ( n1834 & ~n11646 ) | ( n1834 & n11647 ) | ( ~n11646 & n11647 ) ;
  assign n11649 = n11648 ^ n5516 ^ n1955 ;
  assign n11651 = n11650 ^ n11649 ^ n7368 ;
  assign n11652 = ( x201 & n1005 ) | ( x201 & n8283 ) | ( n1005 & n8283 ) ;
  assign n11653 = n11652 ^ n354 ^ 1'b0 ;
  assign n11654 = ( n4319 & n6199 ) | ( n4319 & ~n11653 ) | ( n6199 & ~n11653 ) ;
  assign n11655 = ( ~n1998 & n5428 ) | ( ~n1998 & n11654 ) | ( n5428 & n11654 ) ;
  assign n11656 = ( n3829 & ~n6289 ) | ( n3829 & n11655 ) | ( ~n6289 & n11655 ) ;
  assign n11658 = n1531 ^ n493 ^ 1'b0 ;
  assign n11659 = n1182 | n11658 ;
  assign n11660 = ( ~n5790 & n7481 ) | ( ~n5790 & n11659 ) | ( n7481 & n11659 ) ;
  assign n11657 = n1976 & n9524 ;
  assign n11661 = n11660 ^ n11657 ^ 1'b0 ;
  assign n11667 = n2212 ^ n1576 ^ n743 ;
  assign n11665 = n1388 | n3034 ;
  assign n11666 = n9391 & ~n11665 ;
  assign n11668 = n11667 ^ n11666 ^ n11450 ;
  assign n11662 = ( ~n1077 & n3061 ) | ( ~n1077 & n3479 ) | ( n3061 & n3479 ) ;
  assign n11663 = n11662 ^ n5597 ^ 1'b0 ;
  assign n11664 = ( ~n1482 & n2592 ) | ( ~n1482 & n11663 ) | ( n2592 & n11663 ) ;
  assign n11669 = n11668 ^ n11664 ^ n2622 ;
  assign n11670 = n11661 | n11669 ;
  assign n11677 = ( x232 & n2687 ) | ( x232 & n4239 ) | ( n2687 & n4239 ) ;
  assign n11678 = n11677 ^ n11659 ^ n8112 ;
  assign n11674 = n1396 ^ n334 ^ x180 ;
  assign n11671 = ( ~x186 & n2382 ) | ( ~x186 & n5006 ) | ( n2382 & n5006 ) ;
  assign n11672 = ( ~n1654 & n8573 ) | ( ~n1654 & n11671 ) | ( n8573 & n11671 ) ;
  assign n11673 = ( n4282 & n9248 ) | ( n4282 & n11672 ) | ( n9248 & n11672 ) ;
  assign n11675 = n11674 ^ n11673 ^ n678 ;
  assign n11676 = n11675 ^ n8816 ^ n2955 ;
  assign n11679 = n11678 ^ n11676 ^ n10009 ;
  assign n11683 = n6689 ^ n3768 ^ x124 ;
  assign n11682 = n11499 ^ n7240 ^ n3594 ;
  assign n11680 = ( n571 & ~n7433 ) | ( n571 & n7981 ) | ( ~n7433 & n7981 ) ;
  assign n11681 = n11680 ^ n1619 ^ n438 ;
  assign n11684 = n11683 ^ n11682 ^ n11681 ;
  assign n11691 = n3379 ^ n2759 ^ 1'b0 ;
  assign n11692 = ~n3316 & n11691 ;
  assign n11693 = n9644 ^ n6874 ^ n4564 ;
  assign n11694 = ( n3464 & n6833 ) | ( n3464 & ~n11693 ) | ( n6833 & ~n11693 ) ;
  assign n11695 = n11694 ^ n4458 ^ n1471 ;
  assign n11696 = ( n4012 & ~n11692 ) | ( n4012 & n11695 ) | ( ~n11692 & n11695 ) ;
  assign n11688 = n4439 ^ n4189 ^ n1301 ;
  assign n11689 = ( n1315 & ~n3297 ) | ( n1315 & n11688 ) | ( ~n3297 & n11688 ) ;
  assign n11685 = n1181 & ~n2380 ;
  assign n11686 = n11685 ^ n9464 ^ 1'b0 ;
  assign n11687 = n11686 ^ n9909 ^ n6452 ;
  assign n11690 = n11689 ^ n11687 ^ n10326 ;
  assign n11697 = n11696 ^ n11690 ^ n2237 ;
  assign n11699 = ( n721 & n3858 ) | ( n721 & ~n4187 ) | ( n3858 & ~n4187 ) ;
  assign n11700 = ( n3343 & ~n6669 ) | ( n3343 & n11699 ) | ( ~n6669 & n11699 ) ;
  assign n11701 = n11700 ^ n3347 ^ n761 ;
  assign n11698 = n3881 ^ n2121 ^ n1132 ;
  assign n11702 = n11701 ^ n11698 ^ n1406 ;
  assign n11703 = ( ~n3058 & n5437 ) | ( ~n3058 & n11336 ) | ( n5437 & n11336 ) ;
  assign n11704 = n11703 ^ n2646 ^ n689 ;
  assign n11705 = n11704 ^ n6133 ^ x46 ;
  assign n11706 = n5324 & ~n11705 ;
  assign n11707 = n11706 ^ n8140 ^ n7571 ;
  assign n11708 = n4155 ^ n2251 ^ 1'b0 ;
  assign n11710 = ( n2767 & ~n3348 ) | ( n2767 & n5329 ) | ( ~n3348 & n5329 ) ;
  assign n11709 = n8084 ^ n705 ^ n383 ;
  assign n11711 = n11710 ^ n11709 ^ n8716 ;
  assign n11712 = n1807 ^ n1671 ^ 1'b0 ;
  assign n11713 = n5458 & n7771 ;
  assign n11714 = ( ~n5573 & n11712 ) | ( ~n5573 & n11713 ) | ( n11712 & n11713 ) ;
  assign n11724 = n5374 ^ n5296 ^ n2316 ;
  assign n11725 = n11724 ^ n5749 ^ x19 ;
  assign n11723 = n7265 ^ n5304 ^ n1887 ;
  assign n11720 = n11596 ^ n9153 ^ n4817 ;
  assign n11718 = ( n1839 & n4604 ) | ( n1839 & ~n10218 ) | ( n4604 & ~n10218 ) ;
  assign n11719 = n11718 ^ n1734 ^ n1567 ;
  assign n11721 = n11720 ^ n11719 ^ n2189 ;
  assign n11716 = n2440 ^ n1601 ^ n1417 ;
  assign n11717 = n11716 ^ n7936 ^ n6737 ;
  assign n11722 = n11721 ^ n11717 ^ n1286 ;
  assign n11726 = n11725 ^ n11723 ^ n11722 ;
  assign n11715 = n9852 ^ n6458 ^ n3673 ;
  assign n11727 = n11726 ^ n11715 ^ n2383 ;
  assign n11728 = n11714 | n11727 ;
  assign n11729 = n11711 | n11728 ;
  assign n11730 = n3887 ^ n2237 ^ 1'b0 ;
  assign n11731 = n4198 ^ n3100 ^ n2710 ;
  assign n11732 = n7710 ^ n6177 ^ 1'b0 ;
  assign n11733 = ~n11731 & n11732 ;
  assign n11734 = n11733 ^ n973 ^ n779 ;
  assign n11735 = ( ~n4299 & n6263 ) | ( ~n4299 & n6979 ) | ( n6263 & n6979 ) ;
  assign n11736 = ( n358 & n4768 ) | ( n358 & n5626 ) | ( n4768 & n5626 ) ;
  assign n11737 = ~n11735 & n11736 ;
  assign n11738 = n11737 ^ n6147 ^ 1'b0 ;
  assign n11741 = n4381 ^ n742 ^ 1'b0 ;
  assign n11742 = n11741 ^ n6894 ^ n4390 ;
  assign n11739 = ( n629 & n1744 ) | ( n629 & ~n10997 ) | ( n1744 & ~n10997 ) ;
  assign n11740 = ( n3236 & n6377 ) | ( n3236 & ~n11739 ) | ( n6377 & ~n11739 ) ;
  assign n11743 = n11742 ^ n11740 ^ n2580 ;
  assign n11746 = ( n1537 & ~n3476 ) | ( n1537 & n4742 ) | ( ~n3476 & n4742 ) ;
  assign n11744 = ( n857 & n1315 ) | ( n857 & n1861 ) | ( n1315 & n1861 ) ;
  assign n11745 = ( x22 & ~n6675 ) | ( x22 & n11744 ) | ( ~n6675 & n11744 ) ;
  assign n11747 = n11746 ^ n11745 ^ n868 ;
  assign n11748 = ( ~n5915 & n6056 ) | ( ~n5915 & n9291 ) | ( n6056 & n9291 ) ;
  assign n11749 = ( n2098 & n2113 ) | ( n2098 & n11748 ) | ( n2113 & n11748 ) ;
  assign n11750 = n4700 ^ n4568 ^ n3688 ;
  assign n11751 = ( n1025 & n1874 ) | ( n1025 & n11750 ) | ( n1874 & n11750 ) ;
  assign n11752 = ( n2328 & n3992 ) | ( n2328 & n9780 ) | ( n3992 & n9780 ) ;
  assign n11753 = x229 & ~n11752 ;
  assign n11754 = ~n3765 & n11753 ;
  assign n11755 = n4031 | n7358 ;
  assign n11756 = n11754 & ~n11755 ;
  assign n11757 = ( n10009 & ~n10841 ) | ( n10009 & n11756 ) | ( ~n10841 & n11756 ) ;
  assign n11758 = ( n1224 & ~n1422 ) | ( n1224 & n4300 ) | ( ~n1422 & n4300 ) ;
  assign n11759 = ( n1744 & n6680 ) | ( n1744 & ~n11758 ) | ( n6680 & ~n11758 ) ;
  assign n11760 = ( n11751 & n11757 ) | ( n11751 & ~n11759 ) | ( n11757 & ~n11759 ) ;
  assign n11761 = n11749 | n11760 ;
  assign n11762 = n7011 & ~n11761 ;
  assign n11766 = ~n9862 & n10307 ;
  assign n11767 = ~n556 & n11766 ;
  assign n11763 = n3040 ^ n1756 ^ 1'b0 ;
  assign n11764 = n6233 | n11763 ;
  assign n11765 = n11764 ^ n2953 ^ 1'b0 ;
  assign n11768 = n11767 ^ n11765 ^ n6171 ;
  assign n11769 = n7188 ^ n3137 ^ n1375 ;
  assign n11770 = n11769 ^ n10795 ^ n1435 ;
  assign n11771 = ( n6987 & ~n11569 ) | ( n6987 & n11770 ) | ( ~n11569 & n11770 ) ;
  assign n11772 = n11771 ^ n4358 ^ 1'b0 ;
  assign n11773 = n5327 | n11772 ;
  assign n11774 = ~n3780 & n11773 ;
  assign n11775 = n4098 ^ n1640 ^ 1'b0 ;
  assign n11776 = n11775 ^ n2717 ^ n644 ;
  assign n11777 = n11776 ^ n4796 ^ n2085 ;
  assign n11778 = n9790 | n11777 ;
  assign n11779 = ( ~n292 & n1367 ) | ( ~n292 & n10478 ) | ( n1367 & n10478 ) ;
  assign n11780 = n11779 ^ n7948 ^ n3393 ;
  assign n11781 = n2667 ^ n284 ^ 1'b0 ;
  assign n11782 = n9728 ^ n6596 ^ n4238 ;
  assign n11783 = n11782 ^ n3369 ^ n1589 ;
  assign n11785 = n7837 ^ n2138 ^ 1'b0 ;
  assign n11784 = n3014 & ~n8136 ;
  assign n11786 = n11785 ^ n11784 ^ 1'b0 ;
  assign n11787 = ~n11783 & n11786 ;
  assign n11788 = ~n11781 & n11787 ;
  assign n11789 = n7544 ^ n6502 ^ n4837 ;
  assign n11790 = ( n2163 & ~n4842 ) | ( n2163 & n4891 ) | ( ~n4842 & n4891 ) ;
  assign n11795 = ( n523 & n3703 ) | ( n523 & n9006 ) | ( n3703 & n9006 ) ;
  assign n11796 = n11795 ^ n10963 ^ n8661 ;
  assign n11791 = ( n815 & ~n2953 ) | ( n815 & n4023 ) | ( ~n2953 & n4023 ) ;
  assign n11792 = n11791 ^ n2706 ^ 1'b0 ;
  assign n11793 = n9462 ^ n3871 ^ 1'b0 ;
  assign n11794 = n11792 & ~n11793 ;
  assign n11797 = n11796 ^ n11794 ^ n5785 ;
  assign n11798 = ( ~n2002 & n6967 ) | ( ~n2002 & n7519 ) | ( n6967 & n7519 ) ;
  assign n11799 = ( n4985 & n8172 ) | ( n4985 & ~n11798 ) | ( n8172 & ~n11798 ) ;
  assign n11800 = n11513 ^ n10536 ^ n1800 ;
  assign n11801 = n11800 ^ n6884 ^ 1'b0 ;
  assign n11806 = n4180 ^ n2697 ^ n1612 ;
  assign n11807 = n2448 & ~n11806 ;
  assign n11803 = ( ~n722 & n1294 ) | ( ~n722 & n6913 ) | ( n1294 & n6913 ) ;
  assign n11804 = ( x139 & n6279 ) | ( x139 & n11803 ) | ( n6279 & n11803 ) ;
  assign n11805 = ( n5005 & n5764 ) | ( n5005 & n11804 ) | ( n5764 & n11804 ) ;
  assign n11802 = n1131 & n8092 ;
  assign n11808 = n11807 ^ n11805 ^ n11802 ;
  assign n11809 = n11808 ^ n5393 ^ n3616 ;
  assign n11820 = n5147 ^ n2926 ^ x111 ;
  assign n11813 = n3384 | n6639 ;
  assign n11814 = n4134 | n11813 ;
  assign n11815 = ( ~n365 & n3749 ) | ( ~n365 & n4467 ) | ( n3749 & n4467 ) ;
  assign n11816 = ( x193 & ~n3009 ) | ( x193 & n11815 ) | ( ~n3009 & n11815 ) ;
  assign n11817 = ( n2338 & ~n11814 ) | ( n2338 & n11816 ) | ( ~n11814 & n11816 ) ;
  assign n11818 = n11817 ^ n8518 ^ n8152 ;
  assign n11819 = ~n7549 & n11818 ;
  assign n11821 = n11820 ^ n11819 ^ 1'b0 ;
  assign n11822 = n7368 & n11821 ;
  assign n11810 = n10557 ^ n4260 ^ n2430 ;
  assign n11811 = n11810 ^ n11016 ^ n10866 ;
  assign n11812 = n11811 ^ n5450 ^ n2693 ;
  assign n11823 = n11822 ^ n11812 ^ n10508 ;
  assign n11824 = n3342 ^ n1800 ^ x75 ;
  assign n11825 = ~x158 & n4532 ;
  assign n11826 = n11825 ^ n3543 ^ 1'b0 ;
  assign n11827 = ( n784 & n1031 ) | ( n784 & n11742 ) | ( n1031 & n11742 ) ;
  assign n11828 = n1267 | n11827 ;
  assign n11829 = n3419 | n11828 ;
  assign n11830 = n11829 ^ n8217 ^ 1'b0 ;
  assign n11831 = n4922 & ~n11830 ;
  assign n11832 = n4910 | n11831 ;
  assign n11833 = ( n10401 & n11826 ) | ( n10401 & n11832 ) | ( n11826 & n11832 ) ;
  assign n11834 = ( n979 & n11824 ) | ( n979 & n11833 ) | ( n11824 & n11833 ) ;
  assign n11835 = ( n1911 & ~n2309 ) | ( n1911 & n10567 ) | ( ~n2309 & n10567 ) ;
  assign n11836 = n11835 ^ n8787 ^ n2387 ;
  assign n11837 = n11836 ^ n9111 ^ n801 ;
  assign n11838 = n9726 ^ n8233 ^ n2213 ;
  assign n11839 = n10002 ^ n7492 ^ n4086 ;
  assign n11840 = n11021 ^ n6334 ^ n3092 ;
  assign n11841 = ( ~n1148 & n9101 ) | ( ~n1148 & n11840 ) | ( n9101 & n11840 ) ;
  assign n11842 = ( n4693 & n11839 ) | ( n4693 & ~n11841 ) | ( n11839 & ~n11841 ) ;
  assign n11843 = ( n6133 & n10680 ) | ( n6133 & n10999 ) | ( n10680 & n10999 ) ;
  assign n11844 = n11843 ^ n3094 ^ n327 ;
  assign n11847 = n11363 ^ n3893 ^ n3656 ;
  assign n11848 = ( n3890 & n4902 ) | ( n3890 & ~n11847 ) | ( n4902 & ~n11847 ) ;
  assign n11849 = n3999 | n11848 ;
  assign n11850 = n11849 ^ n2351 ^ 1'b0 ;
  assign n11845 = n6359 ^ n3885 ^ n3345 ;
  assign n11846 = n8032 & n11845 ;
  assign n11851 = n11850 ^ n11846 ^ 1'b0 ;
  assign n11852 = ( n4237 & n11844 ) | ( n4237 & ~n11851 ) | ( n11844 & ~n11851 ) ;
  assign n11853 = n2959 ^ n2578 ^ x166 ;
  assign n11854 = n2529 ^ n2254 ^ n1118 ;
  assign n11855 = ( n3676 & n5185 ) | ( n3676 & n7905 ) | ( n5185 & n7905 ) ;
  assign n11856 = n1026 & ~n1515 ;
  assign n11857 = n7270 ^ n4611 ^ 1'b0 ;
  assign n11858 = ~n11856 & n11857 ;
  assign n11859 = ( n11854 & ~n11855 ) | ( n11854 & n11858 ) | ( ~n11855 & n11858 ) ;
  assign n11860 = n11853 & n11859 ;
  assign n11861 = n11824 ^ n626 ^ x153 ;
  assign n11867 = n4986 ^ n1250 ^ x80 ;
  assign n11862 = ~n3752 & n6417 ;
  assign n11863 = n6774 & n11862 ;
  assign n11864 = n11863 ^ n5571 ^ n5083 ;
  assign n11865 = n11864 ^ n8090 ^ n883 ;
  assign n11866 = ( ~n885 & n1605 ) | ( ~n885 & n11865 ) | ( n1605 & n11865 ) ;
  assign n11868 = n11867 ^ n11866 ^ n1073 ;
  assign n11869 = n2649 ^ n2345 ^ n676 ;
  assign n11870 = n2595 ^ n1474 ^ 1'b0 ;
  assign n11871 = n1906 & n11870 ;
  assign n11872 = n6238 ^ n1388 ^ 1'b0 ;
  assign n11873 = n11872 ^ n5504 ^ n3782 ;
  assign n11874 = n11871 & ~n11873 ;
  assign n11875 = n11874 ^ n9383 ^ 1'b0 ;
  assign n11876 = n7385 ^ n4758 ^ n4565 ;
  assign n11877 = n11876 ^ n3353 ^ 1'b0 ;
  assign n11878 = n11877 ^ n11720 ^ 1'b0 ;
  assign n11879 = ( ~n11869 & n11875 ) | ( ~n11869 & n11878 ) | ( n11875 & n11878 ) ;
  assign n11884 = n4016 & ~n5972 ;
  assign n11885 = ~n1509 & n11884 ;
  assign n11880 = n3162 & ~n8283 ;
  assign n11881 = ~n8853 & n11880 ;
  assign n11882 = n11881 ^ n3550 ^ 1'b0 ;
  assign n11883 = n5646 | n11882 ;
  assign n11886 = n11885 ^ n11883 ^ n4263 ;
  assign n11887 = n7362 ^ n1567 ^ n808 ;
  assign n11888 = ( n9083 & n11886 ) | ( n9083 & ~n11887 ) | ( n11886 & ~n11887 ) ;
  assign n11889 = ( ~n1007 & n4122 ) | ( ~n1007 & n6601 ) | ( n4122 & n6601 ) ;
  assign n11890 = ( ~n8078 & n9440 ) | ( ~n8078 & n11889 ) | ( n9440 & n11889 ) ;
  assign n11891 = ( x90 & ~n2395 ) | ( x90 & n5876 ) | ( ~n2395 & n5876 ) ;
  assign n11892 = ( n5845 & ~n10431 ) | ( n5845 & n11891 ) | ( ~n10431 & n11891 ) ;
  assign n11893 = ( n2645 & n6889 ) | ( n2645 & n8006 ) | ( n6889 & n8006 ) ;
  assign n11894 = ( x199 & n11892 ) | ( x199 & n11893 ) | ( n11892 & n11893 ) ;
  assign n11901 = ( n1088 & n5976 ) | ( n1088 & ~n6288 ) | ( n5976 & ~n6288 ) ;
  assign n11902 = n11901 ^ n9114 ^ n6976 ;
  assign n11897 = ( ~x145 & n2250 ) | ( ~x145 & n5245 ) | ( n2250 & n5245 ) ;
  assign n11898 = ( ~n3386 & n11182 ) | ( ~n3386 & n11897 ) | ( n11182 & n11897 ) ;
  assign n11899 = ~n5022 & n11898 ;
  assign n11900 = n11899 ^ n11677 ^ n6109 ;
  assign n11895 = ( ~n2925 & n4184 ) | ( ~n2925 & n5177 ) | ( n4184 & n5177 ) ;
  assign n11896 = ( ~n2171 & n10488 ) | ( ~n2171 & n11895 ) | ( n10488 & n11895 ) ;
  assign n11903 = n11902 ^ n11900 ^ n11896 ;
  assign n11904 = n10113 ^ n2476 ^ n975 ;
  assign n11905 = ( n1719 & n4689 ) | ( n1719 & n11904 ) | ( n4689 & n11904 ) ;
  assign n11906 = n11856 ^ n8141 ^ n2317 ;
  assign n11907 = n11906 ^ n9850 ^ n3785 ;
  assign n11908 = n11907 ^ n11283 ^ n8622 ;
  assign n11909 = ( n9408 & n11905 ) | ( n9408 & n11908 ) | ( n11905 & n11908 ) ;
  assign n11911 = ~n1374 & n2960 ;
  assign n11912 = n11911 ^ n7201 ^ 1'b0 ;
  assign n11910 = ( ~n3561 & n4788 ) | ( ~n3561 & n11566 ) | ( n4788 & n11566 ) ;
  assign n11913 = n11912 ^ n11910 ^ n6698 ;
  assign n11914 = n11913 ^ n6075 ^ n4545 ;
  assign n11915 = n4943 ^ n3357 ^ n1449 ;
  assign n11916 = n2711 & ~n11915 ;
  assign n11917 = ( n8380 & n9160 ) | ( n8380 & ~n9726 ) | ( n9160 & ~n9726 ) ;
  assign n11918 = ( ~n11914 & n11916 ) | ( ~n11914 & n11917 ) | ( n11916 & n11917 ) ;
  assign n11919 = n11918 ^ n7167 ^ n3445 ;
  assign n11920 = ( ~n1881 & n7393 ) | ( ~n1881 & n11919 ) | ( n7393 & n11919 ) ;
  assign n11921 = n6828 ^ n6297 ^ n2076 ;
  assign n11924 = n8884 ^ n3759 ^ n1395 ;
  assign n11925 = n11924 ^ n6428 ^ n3752 ;
  assign n11926 = n8141 ^ n633 ^ n598 ;
  assign n11927 = n11926 ^ n3714 ^ 1'b0 ;
  assign n11928 = n8494 & ~n11927 ;
  assign n11929 = ( ~n1472 & n6607 ) | ( ~n1472 & n11928 ) | ( n6607 & n11928 ) ;
  assign n11930 = n11925 & ~n11929 ;
  assign n11922 = ( x225 & n2303 ) | ( x225 & n7646 ) | ( n2303 & n7646 ) ;
  assign n11923 = n9194 | n11922 ;
  assign n11931 = n11930 ^ n11923 ^ n11116 ;
  assign n11932 = ( n1319 & ~n3765 ) | ( n1319 & n11147 ) | ( ~n3765 & n11147 ) ;
  assign n11940 = n8673 ^ n6775 ^ n679 ;
  assign n11941 = n11940 ^ n4873 ^ n4811 ;
  assign n11942 = n1846 & n11941 ;
  assign n11943 = ~n8618 & n11942 ;
  assign n11945 = n9025 ^ n6659 ^ n1385 ;
  assign n11944 = n3811 | n6063 ;
  assign n11946 = n11945 ^ n11944 ^ 1'b0 ;
  assign n11947 = n11946 ^ n1955 ^ 1'b0 ;
  assign n11948 = n11943 | n11947 ;
  assign n11938 = n6746 ^ n3393 ^ n851 ;
  assign n11935 = ~n979 & n8044 ;
  assign n11936 = ~n6178 & n11935 ;
  assign n11937 = n7070 | n11936 ;
  assign n11933 = ( n3472 & ~n3887 ) | ( n3472 & n11337 ) | ( ~n3887 & n11337 ) ;
  assign n11934 = n11933 ^ n6925 ^ n6439 ;
  assign n11939 = n11938 ^ n11937 ^ n11934 ;
  assign n11949 = n11948 ^ n11939 ^ 1'b0 ;
  assign n11950 = ~n11932 & n11949 ;
  assign n11951 = ( n6304 & ~n6414 ) | ( n6304 & n9073 ) | ( ~n6414 & n9073 ) ;
  assign n11952 = n11951 ^ n10398 ^ n3831 ;
  assign n11955 = ( ~n2154 & n7888 ) | ( ~n2154 & n8695 ) | ( n7888 & n8695 ) ;
  assign n11953 = ~n5109 & n9961 ;
  assign n11954 = n11953 ^ n3920 ^ n333 ;
  assign n11956 = n11955 ^ n11954 ^ n10146 ;
  assign n11957 = n4164 ^ n3926 ^ 1'b0 ;
  assign n11958 = n7666 | n11957 ;
  assign n11959 = n11958 ^ n6373 ^ n1154 ;
  assign n11960 = ( n4125 & n8771 ) | ( n4125 & n11959 ) | ( n8771 & n11959 ) ;
  assign n11969 = ( n1731 & ~n5966 ) | ( n1731 & n6917 ) | ( ~n5966 & n6917 ) ;
  assign n11970 = ( n5756 & n7708 ) | ( n5756 & n11969 ) | ( n7708 & n11969 ) ;
  assign n11968 = n5507 ^ n5270 ^ n3958 ;
  assign n11962 = n8171 & n9265 ;
  assign n11963 = ( n1021 & n4147 ) | ( n1021 & ~n10009 ) | ( n4147 & ~n10009 ) ;
  assign n11964 = n11963 ^ n5611 ^ 1'b0 ;
  assign n11965 = n11962 & ~n11964 ;
  assign n11966 = ( n651 & n7959 ) | ( n651 & n11965 ) | ( n7959 & n11965 ) ;
  assign n11961 = n7115 ^ n6066 ^ n1817 ;
  assign n11967 = n11966 ^ n11961 ^ n6513 ;
  assign n11971 = n11970 ^ n11968 ^ n11967 ;
  assign n11973 = n11177 ^ n6360 ^ n4412 ;
  assign n11974 = ( n1839 & n3237 ) | ( n1839 & ~n11973 ) | ( n3237 & ~n11973 ) ;
  assign n11972 = n8593 ^ n1089 ^ n721 ;
  assign n11975 = n11974 ^ n11972 ^ n719 ;
  assign n11976 = n11975 ^ n8031 ^ n461 ;
  assign n11977 = n2564 & n11976 ;
  assign n11981 = n5498 ^ n2241 ^ 1'b0 ;
  assign n11982 = n11981 ^ n11914 ^ n5383 ;
  assign n11978 = n7858 & n8783 ;
  assign n11979 = n11978 ^ n4921 ^ 1'b0 ;
  assign n11980 = ( n7403 & n9030 ) | ( n7403 & ~n11979 ) | ( n9030 & ~n11979 ) ;
  assign n11983 = n11982 ^ n11980 ^ n987 ;
  assign n11997 = n9948 ^ n7201 ^ 1'b0 ;
  assign n11998 = n4129 | n11997 ;
  assign n11999 = n11998 ^ n1325 ^ 1'b0 ;
  assign n12000 = n6929 & ~n11999 ;
  assign n11984 = ( ~n4755 & n5885 ) | ( ~n4755 & n7497 ) | ( n5885 & n7497 ) ;
  assign n11986 = ( ~n351 & n521 ) | ( ~n351 & n1181 ) | ( n521 & n1181 ) ;
  assign n11987 = ( n536 & n10323 ) | ( n536 & n11986 ) | ( n10323 & n11986 ) ;
  assign n11988 = ( n4304 & n4885 ) | ( n4304 & ~n11987 ) | ( n4885 & ~n11987 ) ;
  assign n11989 = n11988 ^ n5628 ^ 1'b0 ;
  assign n11985 = ( ~n1160 & n4445 ) | ( ~n1160 & n5296 ) | ( n4445 & n5296 ) ;
  assign n11990 = n11989 ^ n11985 ^ n1895 ;
  assign n11993 = ~x109 & n3814 ;
  assign n11994 = ( n2533 & n3916 ) | ( n2533 & n11993 ) | ( n3916 & n11993 ) ;
  assign n11991 = n8735 ^ n8475 ^ n5505 ;
  assign n11992 = n11991 ^ n3755 ^ n1964 ;
  assign n11995 = n11994 ^ n11992 ^ n3012 ;
  assign n11996 = ( n11984 & n11990 ) | ( n11984 & n11995 ) | ( n11990 & n11995 ) ;
  assign n12001 = n12000 ^ n11996 ^ n6971 ;
  assign n12002 = n6245 ^ n5178 ^ n3352 ;
  assign n12003 = n12002 ^ n5140 ^ n2012 ;
  assign n12004 = ( ~n6231 & n8386 ) | ( ~n6231 & n12003 ) | ( n8386 & n12003 ) ;
  assign n12005 = n834 & ~n12004 ;
  assign n12007 = ( n5944 & n8336 ) | ( n5944 & ~n11538 ) | ( n8336 & ~n11538 ) ;
  assign n12008 = n12007 ^ n9523 ^ n1524 ;
  assign n12006 = ( n1549 & ~n2811 ) | ( n1549 & n9253 ) | ( ~n2811 & n9253 ) ;
  assign n12009 = n12008 ^ n12006 ^ n6707 ;
  assign n12010 = ( n7524 & n12005 ) | ( n7524 & n12009 ) | ( n12005 & n12009 ) ;
  assign n12017 = ( n1288 & n5840 ) | ( n1288 & n11254 ) | ( n5840 & n11254 ) ;
  assign n12015 = n8974 ^ n3004 ^ n2096 ;
  assign n12012 = ( n5954 & n8146 ) | ( n5954 & ~n10580 ) | ( n8146 & ~n10580 ) ;
  assign n12013 = n12012 ^ n3719 ^ n1677 ;
  assign n12011 = ~n4082 & n11539 ;
  assign n12014 = n12013 ^ n12011 ^ 1'b0 ;
  assign n12016 = n12015 ^ n12014 ^ n1149 ;
  assign n12018 = n12017 ^ n12016 ^ n11715 ;
  assign n12021 = ( n418 & n1914 ) | ( n418 & ~n5395 ) | ( n1914 & ~n5395 ) ;
  assign n12022 = ( n5568 & ~n10985 ) | ( n5568 & n12021 ) | ( ~n10985 & n12021 ) ;
  assign n12019 = ( n559 & ~n6218 ) | ( n559 & n7024 ) | ( ~n6218 & n7024 ) ;
  assign n12020 = n12019 ^ n10568 ^ n931 ;
  assign n12023 = n12022 ^ n12020 ^ n3319 ;
  assign n12024 = n2100 | n3143 ;
  assign n12025 = n9251 & ~n12024 ;
  assign n12026 = n3777 & n8829 ;
  assign n12027 = n12026 ^ n1657 ^ 1'b0 ;
  assign n12028 = ( n2567 & ~n8627 ) | ( n2567 & n12027 ) | ( ~n8627 & n12027 ) ;
  assign n12030 = ( ~n1744 & n2195 ) | ( ~n1744 & n4501 ) | ( n2195 & n4501 ) ;
  assign n12029 = n6911 ^ n3312 ^ n1239 ;
  assign n12031 = n12030 ^ n12029 ^ n1471 ;
  assign n12032 = ( n465 & ~n12028 ) | ( n465 & n12031 ) | ( ~n12028 & n12031 ) ;
  assign n12042 = n2546 ^ n1345 ^ n897 ;
  assign n12034 = n2078 & n6608 ;
  assign n12035 = n12034 ^ x209 ^ 1'b0 ;
  assign n12036 = n12035 ^ n2229 ^ x185 ;
  assign n12037 = ( ~n3267 & n6786 ) | ( ~n3267 & n12036 ) | ( n6786 & n12036 ) ;
  assign n12033 = n3070 | n9860 ;
  assign n12038 = n12037 ^ n12033 ^ 1'b0 ;
  assign n12039 = x40 & n7872 ;
  assign n12040 = n12039 ^ n8919 ^ 1'b0 ;
  assign n12041 = n12038 & n12040 ;
  assign n12043 = n12042 ^ n12041 ^ n11168 ;
  assign n12044 = ( ~n2474 & n10781 ) | ( ~n2474 & n11775 ) | ( n10781 & n11775 ) ;
  assign n12045 = ( n2019 & n4615 ) | ( n2019 & n12044 ) | ( n4615 & n12044 ) ;
  assign n12046 = ( x216 & n8161 ) | ( x216 & ~n12045 ) | ( n8161 & ~n12045 ) ;
  assign n12047 = n2421 ^ n2054 ^ n1403 ;
  assign n12048 = n4417 ^ n1497 ^ n1133 ;
  assign n12049 = ( ~x9 & n4430 ) | ( ~x9 & n12048 ) | ( n4430 & n12048 ) ;
  assign n12050 = ( ~n4415 & n7379 ) | ( ~n4415 & n12049 ) | ( n7379 & n12049 ) ;
  assign n12051 = ( n8011 & n12047 ) | ( n8011 & ~n12050 ) | ( n12047 & ~n12050 ) ;
  assign n12052 = n1771 & n7642 ;
  assign n12053 = n12052 ^ n9052 ^ 1'b0 ;
  assign n12054 = ~n8725 & n12053 ;
  assign n12055 = n5002 & ~n8234 ;
  assign n12056 = ( ~x73 & n3432 ) | ( ~x73 & n9244 ) | ( n3432 & n9244 ) ;
  assign n12057 = n12056 ^ n9447 ^ n5075 ;
  assign n12058 = n11988 ^ n9041 ^ 1'b0 ;
  assign n12059 = n12057 & n12058 ;
  assign n12060 = n9987 ^ n9421 ^ n481 ;
  assign n12061 = ~n3211 & n6189 ;
  assign n12062 = n3950 & n12061 ;
  assign n12063 = ~n12060 & n12062 ;
  assign n12064 = ( ~x7 & n2594 ) | ( ~x7 & n8472 ) | ( n2594 & n8472 ) ;
  assign n12065 = ( x160 & n2042 ) | ( x160 & ~n2375 ) | ( n2042 & ~n2375 ) ;
  assign n12066 = n8281 ^ n3623 ^ n2708 ;
  assign n12067 = ( ~n862 & n12065 ) | ( ~n862 & n12066 ) | ( n12065 & n12066 ) ;
  assign n12068 = ( n5560 & n5784 ) | ( n5560 & n12067 ) | ( n5784 & n12067 ) ;
  assign n12069 = ( n9261 & ~n12064 ) | ( n9261 & n12068 ) | ( ~n12064 & n12068 ) ;
  assign n12070 = n4459 ^ n4385 ^ n3608 ;
  assign n12071 = n12070 ^ n11735 ^ n7442 ;
  assign n12072 = n2347 & n9263 ;
  assign n12073 = n499 & n12072 ;
  assign n12074 = n8478 ^ n1722 ^ 1'b0 ;
  assign n12075 = ( ~n7945 & n10224 ) | ( ~n7945 & n12074 ) | ( n10224 & n12074 ) ;
  assign n12076 = n8767 ^ n5841 ^ 1'b0 ;
  assign n12077 = n5373 & n12076 ;
  assign n12078 = n2126 & ~n8485 ;
  assign n12079 = ( n964 & n3535 ) | ( n964 & ~n8156 ) | ( n3535 & ~n8156 ) ;
  assign n12080 = ( n12077 & n12078 ) | ( n12077 & ~n12079 ) | ( n12078 & ~n12079 ) ;
  assign n12081 = ( n3363 & n4625 ) | ( n3363 & ~n12080 ) | ( n4625 & ~n12080 ) ;
  assign n12090 = n3991 ^ x252 ^ 1'b0 ;
  assign n12091 = n12090 ^ n4116 ^ n2275 ;
  assign n12082 = ( n968 & ~n4925 ) | ( n968 & n5767 ) | ( ~n4925 & n5767 ) ;
  assign n12084 = ( n2521 & ~n3696 ) | ( n2521 & n6482 ) | ( ~n3696 & n6482 ) ;
  assign n12085 = n12084 ^ n8498 ^ 1'b0 ;
  assign n12083 = n1761 & n5520 ;
  assign n12086 = n12085 ^ n12083 ^ 1'b0 ;
  assign n12087 = n7543 & n12086 ;
  assign n12088 = n12087 ^ n4240 ^ 1'b0 ;
  assign n12089 = ( n11528 & ~n12082 ) | ( n11528 & n12088 ) | ( ~n12082 & n12088 ) ;
  assign n12092 = n12091 ^ n12089 ^ 1'b0 ;
  assign n12093 = n7111 & n12092 ;
  assign n12098 = n2917 & n3814 ;
  assign n12096 = n5738 ^ n5116 ^ n2389 ;
  assign n12094 = ( n3323 & ~n5213 ) | ( n3323 & n6907 ) | ( ~n5213 & n6907 ) ;
  assign n12095 = n10166 & ~n12094 ;
  assign n12097 = n12096 ^ n12095 ^ 1'b0 ;
  assign n12099 = n12098 ^ n12097 ^ n5208 ;
  assign n12100 = ( ~n1841 & n7714 ) | ( ~n1841 & n12099 ) | ( n7714 & n12099 ) ;
  assign n12101 = n1930 & n4598 ;
  assign n12102 = n12101 ^ n8257 ^ 1'b0 ;
  assign n12103 = ( x242 & n2542 ) | ( x242 & n12102 ) | ( n2542 & n12102 ) ;
  assign n12104 = ( ~n1779 & n10997 ) | ( ~n1779 & n12103 ) | ( n10997 & n12103 ) ;
  assign n12105 = n12104 ^ n10547 ^ n1819 ;
  assign n12106 = n5859 ^ n5212 ^ n4128 ;
  assign n12107 = n9420 ^ n3818 ^ n1704 ;
  assign n12108 = n3576 ^ n1519 ^ 1'b0 ;
  assign n12109 = n12108 ^ n8358 ^ x185 ;
  assign n12110 = ( n848 & ~n1277 ) | ( n848 & n7103 ) | ( ~n1277 & n7103 ) ;
  assign n12111 = n12110 ^ n8928 ^ 1'b0 ;
  assign n12112 = ( n415 & ~n12109 ) | ( n415 & n12111 ) | ( ~n12109 & n12111 ) ;
  assign n12113 = n12112 ^ n7205 ^ n1633 ;
  assign n12115 = n5713 ^ n5178 ^ n2290 ;
  assign n12116 = n12115 ^ n5491 ^ 1'b0 ;
  assign n12114 = n7725 ^ n5388 ^ n2837 ;
  assign n12117 = n12116 ^ n12114 ^ n3251 ;
  assign n12118 = ( n12042 & n12113 ) | ( n12042 & n12117 ) | ( n12113 & n12117 ) ;
  assign n12119 = ( ~x176 & n1883 ) | ( ~x176 & n3272 ) | ( n1883 & n3272 ) ;
  assign n12120 = ( x61 & ~n310 ) | ( x61 & n783 ) | ( ~n310 & n783 ) ;
  assign n12121 = n4774 ^ n3598 ^ n2157 ;
  assign n12122 = ( n1055 & ~n12120 ) | ( n1055 & n12121 ) | ( ~n12120 & n12121 ) ;
  assign n12123 = ( n4560 & n6828 ) | ( n4560 & n12122 ) | ( n6828 & n12122 ) ;
  assign n12124 = ( n5553 & n12119 ) | ( n5553 & n12123 ) | ( n12119 & n12123 ) ;
  assign n12130 = n4165 ^ n2577 ^ x209 ;
  assign n12131 = ( ~n1028 & n7338 ) | ( ~n1028 & n12130 ) | ( n7338 & n12130 ) ;
  assign n12132 = ( n925 & n3406 ) | ( n925 & n12131 ) | ( n3406 & n12131 ) ;
  assign n12126 = ( ~n5033 & n5083 ) | ( ~n5033 & n11442 ) | ( n5083 & n11442 ) ;
  assign n12125 = n8204 ^ n643 ^ 1'b0 ;
  assign n12127 = n12126 ^ n12125 ^ n6243 ;
  assign n12128 = n1602 ^ n767 ^ 1'b0 ;
  assign n12129 = n12127 | n12128 ;
  assign n12133 = n12132 ^ n12129 ^ 1'b0 ;
  assign n12134 = n12124 & n12133 ;
  assign n12135 = ( n6241 & n7426 ) | ( n6241 & n9325 ) | ( n7426 & n9325 ) ;
  assign n12136 = n12135 ^ n4042 ^ x56 ;
  assign n12137 = n7487 & ~n7650 ;
  assign n12141 = n820 & n1052 ;
  assign n12142 = n12141 ^ n3932 ^ 1'b0 ;
  assign n12143 = n12142 ^ n12080 ^ n8340 ;
  assign n12144 = n12143 ^ n9885 ^ n9357 ;
  assign n12138 = n5437 ^ n2955 ^ n1320 ;
  assign n12139 = n12138 ^ n6824 ^ 1'b0 ;
  assign n12140 = ( n6187 & n6567 ) | ( n6187 & n12139 ) | ( n6567 & n12139 ) ;
  assign n12145 = n12144 ^ n12140 ^ 1'b0 ;
  assign n12146 = n6694 ^ n6214 ^ n1512 ;
  assign n12147 = n11792 & ~n12146 ;
  assign n12148 = n12147 ^ n2919 ^ 1'b0 ;
  assign n12149 = n3602 | n4676 ;
  assign n12150 = n12149 ^ n5226 ^ 1'b0 ;
  assign n12152 = n10602 ^ n2432 ^ 1'b0 ;
  assign n12151 = ( n1646 & n3471 ) | ( n1646 & n4426 ) | ( n3471 & n4426 ) ;
  assign n12153 = n12152 ^ n12151 ^ n4167 ;
  assign n12164 = ( n628 & ~n711 ) | ( n628 & n6995 ) | ( ~n711 & n6995 ) ;
  assign n12161 = ( n842 & n6610 ) | ( n842 & n8378 ) | ( n6610 & n8378 ) ;
  assign n12162 = ( n502 & ~n5953 ) | ( n502 & n12161 ) | ( ~n5953 & n12161 ) ;
  assign n12163 = n12162 ^ n11212 ^ n6148 ;
  assign n12158 = n9564 ^ n4174 ^ n3709 ;
  assign n12159 = n12158 ^ n3256 ^ n2673 ;
  assign n12157 = n11539 ^ n4852 ^ 1'b0 ;
  assign n12156 = n8468 ^ n7509 ^ n7051 ;
  assign n12160 = n12159 ^ n12157 ^ n12156 ;
  assign n12165 = n12164 ^ n12163 ^ n12160 ;
  assign n12154 = n6308 ^ n2715 ^ x237 ;
  assign n12155 = n8313 | n12154 ;
  assign n12166 = n12165 ^ n12155 ^ 1'b0 ;
  assign n12167 = ( n12150 & ~n12153 ) | ( n12150 & n12166 ) | ( ~n12153 & n12166 ) ;
  assign n12168 = n5456 & n10291 ;
  assign n12169 = n5417 ^ n3255 ^ n2753 ;
  assign n12170 = ( n4038 & ~n12168 ) | ( n4038 & n12169 ) | ( ~n12168 & n12169 ) ;
  assign n12171 = ( ~n2534 & n9139 ) | ( ~n2534 & n10431 ) | ( n9139 & n10431 ) ;
  assign n12172 = ( n3422 & ~n12170 ) | ( n3422 & n12171 ) | ( ~n12170 & n12171 ) ;
  assign n12173 = ( ~x146 & n11746 ) | ( ~x146 & n12172 ) | ( n11746 & n12172 ) ;
  assign n12174 = n10044 ^ n8895 ^ n486 ;
  assign n12175 = n9552 ^ n6837 ^ n2230 ;
  assign n12176 = n4221 & n7581 ;
  assign n12177 = n4929 & ~n12176 ;
  assign n12178 = ~n7578 & n12177 ;
  assign n12179 = ( n681 & n7667 ) | ( n681 & ~n12178 ) | ( n7667 & ~n12178 ) ;
  assign n12180 = ( n2108 & ~n10397 ) | ( n2108 & n12179 ) | ( ~n10397 & n12179 ) ;
  assign n12184 = n9919 ^ n5124 ^ 1'b0 ;
  assign n12181 = n2499 ^ n1991 ^ 1'b0 ;
  assign n12182 = n9035 & n12181 ;
  assign n12183 = ( n6229 & n10479 ) | ( n6229 & ~n12182 ) | ( n10479 & ~n12182 ) ;
  assign n12185 = n12184 ^ n12183 ^ n4592 ;
  assign n12186 = n4787 ^ n1973 ^ n1394 ;
  assign n12187 = n8080 ^ n5287 ^ 1'b0 ;
  assign n12188 = ~n12186 & n12187 ;
  assign n12192 = ( n6627 & ~n7247 ) | ( n6627 & n7329 ) | ( ~n7247 & n7329 ) ;
  assign n12190 = n7484 ^ n5344 ^ n3200 ;
  assign n12191 = ( n11314 & ~n11497 ) | ( n11314 & n12190 ) | ( ~n11497 & n12190 ) ;
  assign n12193 = n12192 ^ n12191 ^ 1'b0 ;
  assign n12194 = n11040 & n12193 ;
  assign n12189 = ~n1512 & n9258 ;
  assign n12195 = n12194 ^ n12189 ^ 1'b0 ;
  assign n12196 = ( n12185 & n12188 ) | ( n12185 & ~n12195 ) | ( n12188 & ~n12195 ) ;
  assign n12197 = n3941 & ~n9762 ;
  assign n12198 = n6029 & n12197 ;
  assign n12199 = ( ~n6750 & n9681 ) | ( ~n6750 & n12198 ) | ( n9681 & n12198 ) ;
  assign n12200 = ( ~n426 & n1670 ) | ( ~n426 & n5219 ) | ( n1670 & n5219 ) ;
  assign n12201 = ( n5141 & ~n5422 ) | ( n5141 & n12200 ) | ( ~n5422 & n12200 ) ;
  assign n12202 = ( n5749 & n7688 ) | ( n5749 & n12201 ) | ( n7688 & n12201 ) ;
  assign n12203 = ( ~n2435 & n6815 ) | ( ~n2435 & n9217 ) | ( n6815 & n9217 ) ;
  assign n12204 = n12203 ^ n5132 ^ n456 ;
  assign n12205 = n12204 ^ n5273 ^ n4812 ;
  assign n12206 = ( ~n12199 & n12202 ) | ( ~n12199 & n12205 ) | ( n12202 & n12205 ) ;
  assign n12207 = n7721 ^ n6805 ^ n3133 ;
  assign n12208 = ( ~n7616 & n11267 ) | ( ~n7616 & n12207 ) | ( n11267 & n12207 ) ;
  assign n12209 = n4187 | n8007 ;
  assign n12210 = n12209 ^ n4890 ^ 1'b0 ;
  assign n12211 = n9811 ^ n8025 ^ n3711 ;
  assign n12212 = n12211 ^ n9568 ^ n2564 ;
  assign n12213 = ( ~n2309 & n12210 ) | ( ~n2309 & n12212 ) | ( n12210 & n12212 ) ;
  assign n12214 = ( ~n4742 & n7014 ) | ( ~n4742 & n9457 ) | ( n7014 & n9457 ) ;
  assign n12215 = ( n4750 & n4994 ) | ( n4750 & ~n11180 ) | ( n4994 & ~n11180 ) ;
  assign n12216 = ( n473 & n12214 ) | ( n473 & ~n12215 ) | ( n12214 & ~n12215 ) ;
  assign n12217 = n4285 & ~n12216 ;
  assign n12218 = ( n4509 & ~n6678 ) | ( n4509 & n10711 ) | ( ~n6678 & n10711 ) ;
  assign n12219 = n5790 & ~n9762 ;
  assign n12220 = ( n4351 & ~n5413 ) | ( n4351 & n7405 ) | ( ~n5413 & n7405 ) ;
  assign n12221 = ( ~n288 & n4778 ) | ( ~n288 & n12220 ) | ( n4778 & n12220 ) ;
  assign n12222 = n9843 ^ n9155 ^ n3638 ;
  assign n12223 = ( n685 & n3901 ) | ( n685 & n12222 ) | ( n3901 & n12222 ) ;
  assign n12224 = ( n12219 & n12221 ) | ( n12219 & ~n12223 ) | ( n12221 & ~n12223 ) ;
  assign n12225 = ( ~n10507 & n12218 ) | ( ~n10507 & n12224 ) | ( n12218 & n12224 ) ;
  assign n12226 = ( ~n652 & n3114 ) | ( ~n652 & n3558 ) | ( n3114 & n3558 ) ;
  assign n12227 = n11867 | n12226 ;
  assign n12228 = n8174 & ~n12227 ;
  assign n12229 = ( n3990 & n4446 ) | ( n3990 & ~n12228 ) | ( n4446 & ~n12228 ) ;
  assign n12230 = n3708 ^ n3627 ^ n660 ;
  assign n12231 = n12230 ^ n9160 ^ n2336 ;
  assign n12232 = ~n9406 & n10111 ;
  assign n12233 = ( n8498 & n12231 ) | ( n8498 & n12232 ) | ( n12231 & n12232 ) ;
  assign n12234 = n3068 | n9784 ;
  assign n12235 = n12234 ^ n1708 ^ 1'b0 ;
  assign n12236 = n2993 | n10105 ;
  assign n12237 = n1217 | n12236 ;
  assign n12238 = n6683 & ~n12237 ;
  assign n12239 = ( n1035 & n1449 ) | ( n1035 & ~n6967 ) | ( n1449 & ~n6967 ) ;
  assign n12240 = n12239 ^ n6832 ^ n5328 ;
  assign n12241 = ~n12238 & n12240 ;
  assign n12242 = ~n12235 & n12241 ;
  assign n12249 = n4584 ^ n1744 ^ 1'b0 ;
  assign n12250 = ( n6451 & ~n9176 ) | ( n6451 & n12249 ) | ( ~n9176 & n12249 ) ;
  assign n12243 = n1445 ^ n757 ^ n653 ;
  assign n12244 = ( n924 & n10076 ) | ( n924 & ~n12243 ) | ( n10076 & ~n12243 ) ;
  assign n12245 = n12244 ^ n5944 ^ n578 ;
  assign n12246 = n4981 ^ n2458 ^ 1'b0 ;
  assign n12247 = ( n4401 & n5669 ) | ( n4401 & ~n12246 ) | ( n5669 & ~n12246 ) ;
  assign n12248 = ( n6161 & ~n12245 ) | ( n6161 & n12247 ) | ( ~n12245 & n12247 ) ;
  assign n12251 = n12250 ^ n12248 ^ n3837 ;
  assign n12252 = ~n4802 & n12251 ;
  assign n12253 = n12242 & n12252 ;
  assign n12269 = n5210 ^ n1911 ^ n722 ;
  assign n12267 = ( ~x223 & n3398 ) | ( ~x223 & n6799 ) | ( n3398 & n6799 ) ;
  assign n12268 = n12267 ^ n12203 ^ n3641 ;
  assign n12270 = n12269 ^ n12268 ^ n3976 ;
  assign n12258 = n1431 | n7497 ;
  assign n12259 = n12258 ^ n2374 ^ 1'b0 ;
  assign n12257 = ( n1261 & n5058 ) | ( n1261 & ~n5480 ) | ( n5058 & ~n5480 ) ;
  assign n12256 = n11856 ^ n8189 ^ n5184 ;
  assign n12260 = n12259 ^ n12257 ^ n12256 ;
  assign n12254 = n4389 ^ n4036 ^ n3849 ;
  assign n12255 = n10969 | n12254 ;
  assign n12261 = n12260 ^ n12255 ^ 1'b0 ;
  assign n12262 = ( n294 & n3005 ) | ( n294 & ~n4042 ) | ( n3005 & ~n4042 ) ;
  assign n12263 = n5259 & ~n12262 ;
  assign n12264 = n12263 ^ n1712 ^ 1'b0 ;
  assign n12265 = n265 & n12264 ;
  assign n12266 = n12261 & n12265 ;
  assign n12271 = n12270 ^ n12266 ^ n454 ;
  assign n12272 = ( ~n3403 & n7224 ) | ( ~n3403 & n8014 ) | ( n7224 & n8014 ) ;
  assign n12273 = ~n4778 & n12272 ;
  assign n12274 = n7735 ^ n5941 ^ n2748 ;
  assign n12275 = ( n7449 & n9578 ) | ( n7449 & ~n12274 ) | ( n9578 & ~n12274 ) ;
  assign n12276 = ( n7548 & n12273 ) | ( n7548 & n12275 ) | ( n12273 & n12275 ) ;
  assign n12277 = n3206 & ~n8525 ;
  assign n12278 = ( n4475 & n10250 ) | ( n4475 & ~n12277 ) | ( n10250 & ~n12277 ) ;
  assign n12279 = ( ~x171 & n9230 ) | ( ~x171 & n9606 ) | ( n9230 & n9606 ) ;
  assign n12280 = ( n3198 & ~n7454 ) | ( n3198 & n12279 ) | ( ~n7454 & n12279 ) ;
  assign n12281 = ~n12278 & n12280 ;
  assign n12282 = n1783 & n1889 ;
  assign n12283 = ~n3661 & n12282 ;
  assign n12284 = n4876 | n11744 ;
  assign n12285 = n12284 ^ x123 ^ 1'b0 ;
  assign n12286 = n3526 | n12285 ;
  assign n12287 = n8894 ^ n5470 ^ 1'b0 ;
  assign n12288 = n12286 & n12287 ;
  assign n12289 = ~n6253 & n12288 ;
  assign n12290 = n12283 & n12289 ;
  assign n12291 = ( n2492 & n3195 ) | ( n2492 & n12290 ) | ( n3195 & n12290 ) ;
  assign n12293 = ( n827 & n8273 ) | ( n827 & ~n11615 ) | ( n8273 & ~n11615 ) ;
  assign n12292 = n10239 ^ n8678 ^ n6069 ;
  assign n12294 = n12293 ^ n12292 ^ n3238 ;
  assign n12295 = n10969 ^ n4643 ^ n663 ;
  assign n12303 = n6319 & n11006 ;
  assign n12304 = n12303 ^ n515 ^ 1'b0 ;
  assign n12296 = n10493 ^ n9864 ^ 1'b0 ;
  assign n12297 = ~n1581 & n4935 ;
  assign n12298 = n12297 ^ n3641 ^ n855 ;
  assign n12299 = n12298 ^ n10582 ^ 1'b0 ;
  assign n12300 = n12296 & ~n12299 ;
  assign n12301 = n766 & n12300 ;
  assign n12302 = ~n5002 & n12301 ;
  assign n12305 = n12304 ^ n12302 ^ n7870 ;
  assign n12306 = ( ~n4770 & n12295 ) | ( ~n4770 & n12305 ) | ( n12295 & n12305 ) ;
  assign n12307 = n12306 ^ n10631 ^ n10519 ;
  assign n12308 = n1552 & ~n5029 ;
  assign n12309 = n1519 | n12308 ;
  assign n12310 = n1106 & ~n12309 ;
  assign n12311 = n12310 ^ n2544 ^ n519 ;
  assign n12312 = ( n3476 & ~n6729 ) | ( n3476 & n11118 ) | ( ~n6729 & n11118 ) ;
  assign n12313 = n3632 ^ x190 ^ 1'b0 ;
  assign n12314 = n1298 & ~n7279 ;
  assign n12315 = ~n12313 & n12314 ;
  assign n12316 = n7417 | n12315 ;
  assign n12317 = ( n3390 & n12312 ) | ( n3390 & n12316 ) | ( n12312 & n12316 ) ;
  assign n12318 = ( n6328 & n12311 ) | ( n6328 & ~n12317 ) | ( n12311 & ~n12317 ) ;
  assign n12319 = ( n1776 & n2514 ) | ( n1776 & ~n3345 ) | ( n2514 & ~n3345 ) ;
  assign n12320 = n12319 ^ n3002 ^ 1'b0 ;
  assign n12326 = ( ~n313 & n3168 ) | ( ~n313 & n9924 ) | ( n3168 & n9924 ) ;
  assign n12327 = n12326 ^ n2760 ^ n2293 ;
  assign n12323 = n11897 ^ n11895 ^ n6301 ;
  assign n12321 = n2368 ^ x27 ^ 1'b0 ;
  assign n12322 = n12321 ^ n6230 ^ n2768 ;
  assign n12324 = n12323 ^ n12322 ^ n6022 ;
  assign n12325 = n12324 ^ n9032 ^ n1841 ;
  assign n12328 = n12327 ^ n12325 ^ 1'b0 ;
  assign n12329 = n8376 & ~n12328 ;
  assign n12330 = ( n2306 & ~n2424 ) | ( n2306 & n3669 ) | ( ~n2424 & n3669 ) ;
  assign n12331 = ( n3942 & ~n6465 ) | ( n3942 & n12330 ) | ( ~n6465 & n12330 ) ;
  assign n12332 = ( n10313 & ~n12329 ) | ( n10313 & n12331 ) | ( ~n12329 & n12331 ) ;
  assign n12333 = ( n1279 & n1499 ) | ( n1279 & ~n12332 ) | ( n1499 & ~n12332 ) ;
  assign n12334 = ( n1425 & ~n12320 ) | ( n1425 & n12333 ) | ( ~n12320 & n12333 ) ;
  assign n12338 = n2588 ^ n2080 ^ x17 ;
  assign n12339 = n269 | n9434 ;
  assign n12340 = n2429 | n12339 ;
  assign n12341 = ( n1060 & ~n8561 ) | ( n1060 & n12340 ) | ( ~n8561 & n12340 ) ;
  assign n12342 = ( ~n3612 & n5878 ) | ( ~n3612 & n6759 ) | ( n5878 & n6759 ) ;
  assign n12343 = ( n3672 & ~n12341 ) | ( n3672 & n12342 ) | ( ~n12341 & n12342 ) ;
  assign n12344 = ( n6208 & n12338 ) | ( n6208 & ~n12343 ) | ( n12338 & ~n12343 ) ;
  assign n12335 = n5010 ^ n1469 ^ n750 ;
  assign n12336 = ( n1686 & n9444 ) | ( n1686 & ~n10072 ) | ( n9444 & ~n10072 ) ;
  assign n12337 = ( ~n2932 & n12335 ) | ( ~n2932 & n12336 ) | ( n12335 & n12336 ) ;
  assign n12345 = n12344 ^ n12337 ^ n4676 ;
  assign n12349 = n1730 & n2176 ;
  assign n12350 = n7923 & n12349 ;
  assign n12346 = n7745 ^ n486 ^ x2 ;
  assign n12347 = n12065 & n12346 ;
  assign n12348 = ( n1663 & n6371 ) | ( n1663 & ~n12347 ) | ( n6371 & ~n12347 ) ;
  assign n12351 = n12350 ^ n12348 ^ n4457 ;
  assign n12352 = n3272 & n10290 ;
  assign n12353 = n12352 ^ n10224 ^ 1'b0 ;
  assign n12354 = ( n2006 & n2506 ) | ( n2006 & ~n6717 ) | ( n2506 & ~n6717 ) ;
  assign n12355 = n11627 ^ n10990 ^ n5714 ;
  assign n12359 = ( n4648 & n5706 ) | ( n4648 & ~n6254 ) | ( n5706 & ~n6254 ) ;
  assign n12360 = ( ~n3864 & n5213 ) | ( ~n3864 & n7734 ) | ( n5213 & n7734 ) ;
  assign n12361 = ( n12011 & n12359 ) | ( n12011 & n12360 ) | ( n12359 & n12360 ) ;
  assign n12362 = n12361 ^ n11068 ^ n5650 ;
  assign n12356 = ( n9268 & n9301 ) | ( n9268 & ~n11275 ) | ( n9301 & ~n11275 ) ;
  assign n12357 = ( n501 & n4600 ) | ( n501 & ~n12356 ) | ( n4600 & ~n12356 ) ;
  assign n12358 = n12357 ^ n4433 ^ n1473 ;
  assign n12363 = n12362 ^ n12358 ^ 1'b0 ;
  assign n12364 = n12355 & n12363 ;
  assign n12365 = n2592 & n12364 ;
  assign n12366 = n1807 & n2797 ;
  assign n12367 = n12366 ^ n10633 ^ n5626 ;
  assign n12368 = n12367 ^ n9492 ^ n8269 ;
  assign n12369 = ( n430 & n867 ) | ( n430 & n7020 ) | ( n867 & n7020 ) ;
  assign n12370 = ( ~n8665 & n9750 ) | ( ~n8665 & n12369 ) | ( n9750 & n12369 ) ;
  assign n12371 = ( n2858 & n3580 ) | ( n2858 & n5223 ) | ( n3580 & n5223 ) ;
  assign n12372 = n5289 ^ n4863 ^ n1955 ;
  assign n12373 = ( n6279 & ~n12371 ) | ( n6279 & n12372 ) | ( ~n12371 & n12372 ) ;
  assign n12374 = n10719 ^ n3019 ^ n2211 ;
  assign n12375 = n12374 ^ n12321 ^ x39 ;
  assign n12376 = ( n5893 & ~n12373 ) | ( n5893 & n12375 ) | ( ~n12373 & n12375 ) ;
  assign n12377 = ( ~n3381 & n12370 ) | ( ~n3381 & n12376 ) | ( n12370 & n12376 ) ;
  assign n12380 = n5774 ^ n3148 ^ 1'b0 ;
  assign n12381 = ( n2457 & n6593 ) | ( n2457 & n12380 ) | ( n6593 & n12380 ) ;
  assign n12378 = n5099 ^ n4235 ^ n291 ;
  assign n12379 = n4115 | n12378 ;
  assign n12382 = n12381 ^ n12379 ^ 1'b0 ;
  assign n12390 = n11429 ^ n11021 ^ n5650 ;
  assign n12391 = n5597 | n12390 ;
  assign n12392 = n12391 ^ n4171 ^ 1'b0 ;
  assign n12387 = n6768 ^ n6502 ^ n4456 ;
  assign n12388 = n12387 ^ n5088 ^ n2714 ;
  assign n12384 = ( n640 & n1424 ) | ( n640 & ~n6038 ) | ( n1424 & ~n6038 ) ;
  assign n12385 = n12384 ^ n7743 ^ n269 ;
  assign n12386 = n12385 ^ n10707 ^ n6972 ;
  assign n12389 = n12388 ^ n12386 ^ n2711 ;
  assign n12383 = n6951 ^ n6757 ^ n5832 ;
  assign n12393 = n12392 ^ n12389 ^ n12383 ;
  assign n12394 = ( n3976 & n7780 ) | ( n3976 & n12393 ) | ( n7780 & n12393 ) ;
  assign n12401 = ( n991 & n2890 ) | ( n991 & ~n7063 ) | ( n2890 & ~n7063 ) ;
  assign n12397 = n7593 ^ n3037 ^ n1974 ;
  assign n12398 = n10765 | n12397 ;
  assign n12399 = x242 | n12398 ;
  assign n12395 = ( n1594 & n2916 ) | ( n1594 & n5345 ) | ( n2916 & n5345 ) ;
  assign n12396 = n12395 ^ n3637 ^ 1'b0 ;
  assign n12400 = n12399 ^ n12396 ^ n665 ;
  assign n12402 = n12401 ^ n12400 ^ n8548 ;
  assign n12403 = n7606 ^ n6148 ^ n579 ;
  assign n12404 = ( ~n431 & n2340 ) | ( ~n431 & n9864 ) | ( n2340 & n9864 ) ;
  assign n12405 = ( ~n11876 & n12403 ) | ( ~n11876 & n12404 ) | ( n12403 & n12404 ) ;
  assign n12406 = ( n787 & ~n7211 ) | ( n787 & n12405 ) | ( ~n7211 & n12405 ) ;
  assign n12409 = ( x59 & n3991 ) | ( x59 & ~n4316 ) | ( n3991 & ~n4316 ) ;
  assign n12410 = n1779 & ~n2207 ;
  assign n12411 = ~n12409 & n12410 ;
  assign n12407 = n5505 ^ n5134 ^ n2001 ;
  assign n12408 = ( n2151 & n6554 ) | ( n2151 & ~n12407 ) | ( n6554 & ~n12407 ) ;
  assign n12412 = n12411 ^ n12408 ^ 1'b0 ;
  assign n12413 = n9109 ^ n3205 ^ n626 ;
  assign n12414 = n12413 ^ n11083 ^ n4748 ;
  assign n12415 = ( x135 & n6029 ) | ( x135 & ~n12414 ) | ( n6029 & ~n12414 ) ;
  assign n12416 = n12415 ^ n8297 ^ 1'b0 ;
  assign n12417 = n7802 ^ n7203 ^ 1'b0 ;
  assign n12418 = n6239 & n12417 ;
  assign n12419 = n12418 ^ n9028 ^ n1122 ;
  assign n12420 = n8760 ^ n4394 ^ x61 ;
  assign n12421 = ( n2330 & ~n3897 ) | ( n2330 & n4645 ) | ( ~n3897 & n4645 ) ;
  assign n12422 = ( n7260 & n12420 ) | ( n7260 & n12421 ) | ( n12420 & n12421 ) ;
  assign n12423 = ( n2166 & n2626 ) | ( n2166 & ~n12422 ) | ( n2626 & ~n12422 ) ;
  assign n12427 = ( n3353 & ~n5662 ) | ( n3353 & n10596 ) | ( ~n5662 & n10596 ) ;
  assign n12428 = n2455 ^ n581 ^ 1'b0 ;
  assign n12429 = ~n12427 & n12428 ;
  assign n12424 = ( n4110 & n5228 ) | ( n4110 & n10838 ) | ( n5228 & n10838 ) ;
  assign n12425 = ( n1674 & ~n6507 ) | ( n1674 & n12424 ) | ( ~n6507 & n12424 ) ;
  assign n12426 = n5515 & n12425 ;
  assign n12430 = n12429 ^ n12426 ^ 1'b0 ;
  assign n12431 = n8425 ^ n1007 ^ n533 ;
  assign n12437 = n10107 ^ n8454 ^ x91 ;
  assign n12432 = n289 | n1257 ;
  assign n12433 = n7810 ^ n4638 ^ x97 ;
  assign n12434 = n10323 & ~n12433 ;
  assign n12435 = ~n8201 & n12434 ;
  assign n12436 = ( n472 & n12432 ) | ( n472 & n12435 ) | ( n12432 & n12435 ) ;
  assign n12438 = n12437 ^ n12436 ^ 1'b0 ;
  assign n12439 = n4856 & ~n12438 ;
  assign n12440 = ( ~n6783 & n10148 ) | ( ~n6783 & n11256 ) | ( n10148 & n11256 ) ;
  assign n12448 = ( n2431 & n3002 ) | ( n2431 & n8101 ) | ( n3002 & n8101 ) ;
  assign n12445 = ( n5455 & n6765 ) | ( n5455 & ~n9473 ) | ( n6765 & ~n9473 ) ;
  assign n12446 = ( n2268 & ~n11233 ) | ( n2268 & n12445 ) | ( ~n11233 & n12445 ) ;
  assign n12447 = ( n6155 & n8615 ) | ( n6155 & ~n12446 ) | ( n8615 & ~n12446 ) ;
  assign n12443 = n7139 ^ n1948 ^ x193 ;
  assign n12441 = n9806 ^ n9368 ^ n774 ;
  assign n12442 = n12441 ^ n9920 ^ n4579 ;
  assign n12444 = n12443 ^ n12442 ^ n6262 ;
  assign n12449 = n12448 ^ n12447 ^ n12444 ;
  assign n12450 = ( ~n12439 & n12440 ) | ( ~n12439 & n12449 ) | ( n12440 & n12449 ) ;
  assign n12451 = n8555 ^ n1112 ^ 1'b0 ;
  assign n12452 = n12451 ^ n9566 ^ n6014 ;
  assign n12462 = n8827 ^ n2157 ^ n1283 ;
  assign n12463 = n12462 ^ n5848 ^ 1'b0 ;
  assign n12464 = n7903 ^ n930 ^ 1'b0 ;
  assign n12465 = n10512 & n12464 ;
  assign n12466 = ( n5183 & n7022 ) | ( n5183 & n12465 ) | ( n7022 & n12465 ) ;
  assign n12467 = ~n4319 & n12466 ;
  assign n12468 = ( n7034 & n12463 ) | ( n7034 & ~n12467 ) | ( n12463 & ~n12467 ) ;
  assign n12458 = n2458 ^ n2060 ^ n556 ;
  assign n12455 = n6685 ^ n2628 ^ n1332 ;
  assign n12456 = ( n3988 & ~n6669 ) | ( n3988 & n12455 ) | ( ~n6669 & n12455 ) ;
  assign n12457 = ( ~n3508 & n7417 ) | ( ~n3508 & n12456 ) | ( n7417 & n12456 ) ;
  assign n12459 = n12458 ^ n12457 ^ n2824 ;
  assign n12453 = n2356 ^ n1197 ^ x154 ;
  assign n12454 = n12453 ^ n5882 ^ n2528 ;
  assign n12460 = n12459 ^ n12454 ^ n4650 ;
  assign n12461 = ( n4215 & n6508 ) | ( n4215 & ~n12460 ) | ( n6508 & ~n12460 ) ;
  assign n12469 = n12468 ^ n12461 ^ n4070 ;
  assign n12474 = ( x244 & n1762 ) | ( x244 & ~n5312 ) | ( n1762 & ~n5312 ) ;
  assign n12473 = n4319 ^ n3426 ^ n2071 ;
  assign n12470 = ( n3502 & n5462 ) | ( n3502 & n5880 ) | ( n5462 & n5880 ) ;
  assign n12471 = n10126 ^ n7520 ^ 1'b0 ;
  assign n12472 = ( n3968 & n12470 ) | ( n3968 & n12471 ) | ( n12470 & n12471 ) ;
  assign n12475 = n12474 ^ n12473 ^ n12472 ;
  assign n12476 = n6516 ^ n2279 ^ 1'b0 ;
  assign n12477 = ( n4557 & ~n6357 ) | ( n4557 & n12476 ) | ( ~n6357 & n12476 ) ;
  assign n12478 = ( ~n3934 & n8990 ) | ( ~n3934 & n12477 ) | ( n8990 & n12477 ) ;
  assign n12479 = n12478 ^ n11736 ^ 1'b0 ;
  assign n12480 = n12479 ^ n12399 ^ n8609 ;
  assign n12487 = ( x119 & ~x183 ) | ( x119 & n4447 ) | ( ~x183 & n4447 ) ;
  assign n12481 = ( n4213 & n6287 ) | ( n4213 & ~n7947 ) | ( n6287 & ~n7947 ) ;
  assign n12482 = ( ~n4065 & n4558 ) | ( ~n4065 & n11451 ) | ( n4558 & n11451 ) ;
  assign n12484 = ( n4122 & n8844 ) | ( n4122 & ~n10377 ) | ( n8844 & ~n10377 ) ;
  assign n12483 = n10729 & ~n10838 ;
  assign n12485 = n12484 ^ n12483 ^ 1'b0 ;
  assign n12486 = ( n12481 & n12482 ) | ( n12481 & n12485 ) | ( n12482 & n12485 ) ;
  assign n12488 = n12487 ^ n12486 ^ n5709 ;
  assign n12491 = ( n1424 & ~n2344 ) | ( n1424 & n2761 ) | ( ~n2344 & n2761 ) ;
  assign n12489 = ( x144 & ~n6752 ) | ( x144 & n10438 ) | ( ~n6752 & n10438 ) ;
  assign n12490 = ( n1629 & n1968 ) | ( n1629 & n12489 ) | ( n1968 & n12489 ) ;
  assign n12492 = n12491 ^ n12490 ^ n2230 ;
  assign n12493 = ( n4289 & n6654 ) | ( n4289 & n11160 ) | ( n6654 & n11160 ) ;
  assign n12494 = n12493 ^ n9268 ^ n5507 ;
  assign n12495 = n2778 ^ n2403 ^ n721 ;
  assign n12496 = n7424 ^ n1709 ^ 1'b0 ;
  assign n12497 = ( ~n12494 & n12495 ) | ( ~n12494 & n12496 ) | ( n12495 & n12496 ) ;
  assign n12498 = n12497 ^ n5192 ^ n4033 ;
  assign n12499 = ( n11815 & ~n12492 ) | ( n11815 & n12498 ) | ( ~n12492 & n12498 ) ;
  assign n12500 = n11875 ^ n8311 ^ n3425 ;
  assign n12501 = ~n284 & n865 ;
  assign n12502 = n11232 ^ n5635 ^ 1'b0 ;
  assign n12503 = ( n3332 & ~n3507 ) | ( n3332 & n12502 ) | ( ~n3507 & n12502 ) ;
  assign n12510 = ( n2899 & ~n8430 ) | ( n2899 & n8679 ) | ( ~n8430 & n8679 ) ;
  assign n12508 = ( n3088 & n5688 ) | ( n3088 & ~n5907 ) | ( n5688 & ~n5907 ) ;
  assign n12504 = n404 & n1667 ;
  assign n12505 = n12504 ^ n8140 ^ 1'b0 ;
  assign n12506 = ( n590 & n1588 ) | ( n590 & ~n12505 ) | ( n1588 & ~n12505 ) ;
  assign n12507 = n12506 ^ n453 ^ x1 ;
  assign n12509 = n12508 ^ n12507 ^ n7524 ;
  assign n12511 = n12510 ^ n12509 ^ n9241 ;
  assign n12512 = n6335 ^ n3586 ^ n1281 ;
  assign n12513 = ( n415 & n2396 ) | ( n415 & n12512 ) | ( n2396 & n12512 ) ;
  assign n12514 = n12513 ^ n7654 ^ n933 ;
  assign n12515 = n12514 ^ n6061 ^ n1888 ;
  assign n12516 = ( n876 & n1527 ) | ( n876 & ~n7198 ) | ( n1527 & ~n7198 ) ;
  assign n12517 = ( n1551 & ~n9192 ) | ( n1551 & n12516 ) | ( ~n9192 & n12516 ) ;
  assign n12518 = ~x45 & n12517 ;
  assign n12528 = n6574 ^ n2445 ^ n1281 ;
  assign n12529 = n12528 ^ n8698 ^ n5908 ;
  assign n12519 = n5543 ^ n1371 ^ n806 ;
  assign n12520 = n12519 ^ n5505 ^ n2403 ;
  assign n12521 = ( ~n4015 & n7293 ) | ( ~n4015 & n12520 ) | ( n7293 & n12520 ) ;
  assign n12522 = n4770 | n12521 ;
  assign n12523 = n6099 | n12522 ;
  assign n12524 = n9162 ^ n8378 ^ 1'b0 ;
  assign n12525 = n12524 ^ n12321 ^ n2387 ;
  assign n12526 = n12523 & n12525 ;
  assign n12527 = n12526 ^ n3811 ^ 1'b0 ;
  assign n12530 = n12529 ^ n12527 ^ n12145 ;
  assign n12532 = n10720 | n12042 ;
  assign n12533 = n7225 | n12532 ;
  assign n12531 = n1051 | n10976 ;
  assign n12534 = n12533 ^ n12531 ^ 1'b0 ;
  assign n12538 = n1749 & n5970 ;
  assign n12539 = ( n3278 & n11959 ) | ( n3278 & ~n12538 ) | ( n11959 & ~n12538 ) ;
  assign n12536 = n3062 ^ n2172 ^ n1828 ;
  assign n12537 = ( n3255 & n6082 ) | ( n3255 & n12536 ) | ( n6082 & n12536 ) ;
  assign n12540 = n12539 ^ n12537 ^ n7853 ;
  assign n12541 = n8392 ^ n7264 ^ n2639 ;
  assign n12542 = ( x166 & n3035 ) | ( x166 & ~n3744 ) | ( n3035 & ~n3744 ) ;
  assign n12543 = n12542 ^ n5910 ^ n2347 ;
  assign n12544 = n11710 ^ n3298 ^ n2534 ;
  assign n12545 = ( ~n7418 & n12543 ) | ( ~n7418 & n12544 ) | ( n12543 & n12544 ) ;
  assign n12546 = n11473 ^ n9549 ^ n4468 ;
  assign n12547 = ( n12541 & n12545 ) | ( n12541 & n12546 ) | ( n12545 & n12546 ) ;
  assign n12548 = ( ~n5465 & n12540 ) | ( ~n5465 & n12547 ) | ( n12540 & n12547 ) ;
  assign n12535 = ( n2274 & n3767 ) | ( n2274 & n8342 ) | ( n3767 & n8342 ) ;
  assign n12549 = n12548 ^ n12535 ^ n5271 ;
  assign n12550 = ( n2430 & ~n4293 ) | ( n2430 & n7373 ) | ( ~n4293 & n7373 ) ;
  assign n12551 = ( ~n8066 & n9335 ) | ( ~n8066 & n9459 ) | ( n9335 & n9459 ) ;
  assign n12552 = n12551 ^ n4772 ^ n2956 ;
  assign n12553 = ( ~n7256 & n11840 ) | ( ~n7256 & n12552 ) | ( n11840 & n12552 ) ;
  assign n12554 = ( n10753 & ~n12550 ) | ( n10753 & n12553 ) | ( ~n12550 & n12553 ) ;
  assign n12555 = n4560 ^ n2521 ^ n728 ;
  assign n12556 = ( ~n5224 & n10821 ) | ( ~n5224 & n12555 ) | ( n10821 & n12555 ) ;
  assign n12557 = ( n4221 & ~n12017 ) | ( n4221 & n12556 ) | ( ~n12017 & n12556 ) ;
  assign n12558 = ( n1899 & n2437 ) | ( n1899 & ~n2785 ) | ( n2437 & ~n2785 ) ;
  assign n12559 = n12558 ^ n12203 ^ n814 ;
  assign n12560 = n12559 ^ n7070 ^ n3322 ;
  assign n12561 = n12560 ^ n10178 ^ n5881 ;
  assign n12562 = n12561 ^ n817 ^ 1'b0 ;
  assign n12563 = ( n2130 & n5644 ) | ( n2130 & n7018 ) | ( n5644 & n7018 ) ;
  assign n12565 = ( n692 & n4775 ) | ( n692 & ~n10345 ) | ( n4775 & ~n10345 ) ;
  assign n12566 = ( n276 & n1111 ) | ( n276 & ~n12565 ) | ( n1111 & ~n12565 ) ;
  assign n12564 = n3283 ^ n2780 ^ n868 ;
  assign n12567 = n12566 ^ n12564 ^ n7992 ;
  assign n12568 = ( ~n5334 & n10773 ) | ( ~n5334 & n12567 ) | ( n10773 & n12567 ) ;
  assign n12569 = n673 | n7952 ;
  assign n12570 = n7690 | n12569 ;
  assign n12571 = n12570 ^ n11922 ^ n2630 ;
  assign n12572 = n2856 & n12571 ;
  assign n12573 = n12572 ^ n6269 ^ 1'b0 ;
  assign n12574 = ( ~n3941 & n6197 ) | ( ~n3941 & n7370 ) | ( n6197 & n7370 ) ;
  assign n12575 = x168 & n4019 ;
  assign n12576 = n12524 & n12575 ;
  assign n12577 = ( n1828 & ~n5181 ) | ( n1828 & n8291 ) | ( ~n5181 & n8291 ) ;
  assign n12578 = n7029 ^ n6905 ^ n1879 ;
  assign n12579 = n5148 & ~n6928 ;
  assign n12580 = n12579 ^ n11815 ^ 1'b0 ;
  assign n12581 = ( ~n12577 & n12578 ) | ( ~n12577 & n12580 ) | ( n12578 & n12580 ) ;
  assign n12582 = ( ~n3300 & n5253 ) | ( ~n3300 & n6534 ) | ( n5253 & n6534 ) ;
  assign n12583 = n12582 ^ n7139 ^ n663 ;
  assign n12584 = ( ~n1424 & n2860 ) | ( ~n1424 & n10494 ) | ( n2860 & n10494 ) ;
  assign n12585 = n2681 ^ n1937 ^ n1046 ;
  assign n12586 = ( n12583 & n12584 ) | ( n12583 & ~n12585 ) | ( n12584 & ~n12585 ) ;
  assign n12587 = n6763 ^ n4259 ^ n2813 ;
  assign n12588 = n12587 ^ n6520 ^ n5746 ;
  assign n12589 = n7977 ^ n4936 ^ 1'b0 ;
  assign n12590 = n4016 & n12589 ;
  assign n12591 = ( n1771 & n7238 ) | ( n1771 & n12590 ) | ( n7238 & n12590 ) ;
  assign n12592 = ( ~n5050 & n12588 ) | ( ~n5050 & n12591 ) | ( n12588 & n12591 ) ;
  assign n12593 = n12019 ^ x228 ^ 1'b0 ;
  assign n12594 = n12593 ^ n4640 ^ 1'b0 ;
  assign n12595 = ( ~n3286 & n5670 ) | ( ~n3286 & n12594 ) | ( n5670 & n12594 ) ;
  assign n12596 = ( n1494 & n1927 ) | ( n1494 & ~n12595 ) | ( n1927 & ~n12595 ) ;
  assign n12597 = ( n1141 & ~n12493 ) | ( n1141 & n12565 ) | ( ~n12493 & n12565 ) ;
  assign n12598 = n12597 ^ n3492 ^ 1'b0 ;
  assign n12599 = n6844 & n12598 ;
  assign n12600 = n4100 ^ n1005 ^ 1'b0 ;
  assign n12601 = ~n8463 & n9775 ;
  assign n12602 = n10146 ^ n4390 ^ 1'b0 ;
  assign n12603 = n12601 | n12602 ;
  assign n12604 = n12603 ^ n9263 ^ n3219 ;
  assign n12605 = ( n5768 & n9686 ) | ( n5768 & ~n9997 ) | ( n9686 & ~n9997 ) ;
  assign n12613 = n6260 | n6803 ;
  assign n12607 = ~n2096 & n3812 ;
  assign n12608 = n4122 & ~n9465 ;
  assign n12609 = ~n12607 & n12608 ;
  assign n12610 = n10772 & ~n12609 ;
  assign n12611 = n12610 ^ n9880 ^ 1'b0 ;
  assign n12606 = n3153 | n4390 ;
  assign n12612 = n12611 ^ n12606 ^ 1'b0 ;
  assign n12614 = n12613 ^ n12612 ^ n6395 ;
  assign n12615 = ~n12605 & n12614 ;
  assign n12616 = n12615 ^ n9658 ^ n6230 ;
  assign n12617 = n11700 ^ n7234 ^ n4127 ;
  assign n12618 = n6786 & ~n11384 ;
  assign n12619 = n12618 ^ n7727 ^ 1'b0 ;
  assign n12620 = n5044 ^ n3083 ^ n1209 ;
  assign n12622 = n7526 & ~n8776 ;
  assign n12623 = n12622 ^ n6428 ^ 1'b0 ;
  assign n12621 = n5360 ^ n4305 ^ n3927 ;
  assign n12624 = n12623 ^ n12621 ^ n2874 ;
  assign n12627 = ( ~n1937 & n2439 ) | ( ~n1937 & n5163 ) | ( n2439 & n5163 ) ;
  assign n12628 = n12627 ^ n291 ^ 1'b0 ;
  assign n12625 = n9826 ^ n3307 ^ n1527 ;
  assign n12626 = n12625 ^ n11620 ^ n662 ;
  assign n12629 = n12628 ^ n12626 ^ n6308 ;
  assign n12630 = ( ~n4400 & n7265 ) | ( ~n4400 & n10956 ) | ( n7265 & n10956 ) ;
  assign n12631 = n4602 & ~n7740 ;
  assign n12632 = ( n1684 & n3885 ) | ( n1684 & n7795 ) | ( n3885 & n7795 ) ;
  assign n12633 = n12632 ^ n4417 ^ n389 ;
  assign n12634 = ( ~n926 & n3400 ) | ( ~n926 & n11191 ) | ( n3400 & n11191 ) ;
  assign n12635 = n12634 ^ n3319 ^ n1705 ;
  assign n12636 = ( ~n6979 & n12633 ) | ( ~n6979 & n12635 ) | ( n12633 & n12635 ) ;
  assign n12637 = ( n464 & n8377 ) | ( n464 & ~n8488 ) | ( n8377 & ~n8488 ) ;
  assign n12643 = ( n773 & n5228 ) | ( n773 & n11588 ) | ( n5228 & n11588 ) ;
  assign n12644 = n12643 ^ n5884 ^ n2935 ;
  assign n12638 = ( ~n759 & n1610 ) | ( ~n759 & n3209 ) | ( n1610 & n3209 ) ;
  assign n12639 = n12638 ^ n7150 ^ n1588 ;
  assign n12640 = n546 | n5328 ;
  assign n12641 = ( n7127 & ~n12639 ) | ( n7127 & n12640 ) | ( ~n12639 & n12640 ) ;
  assign n12642 = ( ~n3579 & n9196 ) | ( ~n3579 & n12641 ) | ( n9196 & n12641 ) ;
  assign n12645 = n12644 ^ n12642 ^ n7543 ;
  assign n12646 = n12645 ^ n10600 ^ n4555 ;
  assign n12647 = n10227 ^ n2074 ^ 1'b0 ;
  assign n12648 = ( n1260 & ~n9617 ) | ( n1260 & n12647 ) | ( ~n9617 & n12647 ) ;
  assign n12649 = ( n8824 & ~n9034 ) | ( n8824 & n12648 ) | ( ~n9034 & n12648 ) ;
  assign n12650 = n12649 ^ n5351 ^ x244 ;
  assign n12651 = n9298 ^ n4579 ^ n685 ;
  assign n12652 = ( n396 & ~n4096 ) | ( n396 & n12651 ) | ( ~n4096 & n12651 ) ;
  assign n12653 = n11803 ^ n6859 ^ n5704 ;
  assign n12654 = ( n3064 & n8621 ) | ( n3064 & ~n12653 ) | ( n8621 & ~n12653 ) ;
  assign n12655 = ( ~n5170 & n12652 ) | ( ~n5170 & n12654 ) | ( n12652 & n12654 ) ;
  assign n12656 = ( n1324 & ~n6139 ) | ( n1324 & n12655 ) | ( ~n6139 & n12655 ) ;
  assign n12657 = ( n1545 & n3185 ) | ( n1545 & ~n3219 ) | ( n3185 & ~n3219 ) ;
  assign n12658 = n1155 & ~n11869 ;
  assign n12659 = n12658 ^ n2637 ^ 1'b0 ;
  assign n12660 = ( n12142 & n12657 ) | ( n12142 & ~n12659 ) | ( n12657 & ~n12659 ) ;
  assign n12661 = ( n2735 & ~n6129 ) | ( n2735 & n12660 ) | ( ~n6129 & n12660 ) ;
  assign n12662 = ( n2621 & n2654 ) | ( n2621 & ~n3191 ) | ( n2654 & ~n3191 ) ;
  assign n12663 = n6286 ^ n4301 ^ 1'b0 ;
  assign n12664 = ( ~n6186 & n12662 ) | ( ~n6186 & n12663 ) | ( n12662 & n12663 ) ;
  assign n12665 = n12664 ^ n3823 ^ x28 ;
  assign n12666 = ( n6988 & ~n8131 ) | ( n6988 & n12665 ) | ( ~n8131 & n12665 ) ;
  assign n12668 = ~n524 & n6028 ;
  assign n12667 = ( ~n5743 & n6137 ) | ( ~n5743 & n8098 ) | ( n6137 & n8098 ) ;
  assign n12669 = n12668 ^ n12667 ^ n8179 ;
  assign n12670 = ( n4279 & n5553 ) | ( n4279 & n6804 ) | ( n5553 & n6804 ) ;
  assign n12671 = n546 | n11099 ;
  assign n12672 = n12671 ^ n1973 ^ 1'b0 ;
  assign n12674 = ( ~n903 & n2261 ) | ( ~n903 & n4184 ) | ( n2261 & n4184 ) ;
  assign n12675 = n11853 ^ n5635 ^ 1'b0 ;
  assign n12676 = ~n12674 & n12675 ;
  assign n12673 = n12296 ^ n2541 ^ n1957 ;
  assign n12677 = n12676 ^ n12673 ^ n736 ;
  assign n12678 = ( ~n2093 & n12672 ) | ( ~n2093 & n12677 ) | ( n12672 & n12677 ) ;
  assign n12679 = n7591 & ~n7650 ;
  assign n12680 = n12679 ^ n6202 ^ 1'b0 ;
  assign n12681 = n1416 | n1772 ;
  assign n12682 = n10129 & ~n12681 ;
  assign n12683 = n8345 ^ n1897 ^ 1'b0 ;
  assign n12684 = ~n8484 & n12683 ;
  assign n12685 = n12684 ^ n10046 ^ n964 ;
  assign n12686 = ( ~n12680 & n12682 ) | ( ~n12680 & n12685 ) | ( n12682 & n12685 ) ;
  assign n12687 = ( ~n345 & n2844 ) | ( ~n345 & n5399 ) | ( n2844 & n5399 ) ;
  assign n12688 = n1501 & ~n12687 ;
  assign n12689 = n10168 ^ n6203 ^ n1388 ;
  assign n12690 = ( n4152 & ~n12688 ) | ( n4152 & n12689 ) | ( ~n12688 & n12689 ) ;
  assign n12691 = n4625 ^ n3816 ^ 1'b0 ;
  assign n12692 = ~n8876 & n12691 ;
  assign n12695 = n11898 ^ n1501 ^ 1'b0 ;
  assign n12693 = ( ~n2981 & n4122 ) | ( ~n2981 & n9607 ) | ( n4122 & n9607 ) ;
  assign n12694 = n12693 ^ n7846 ^ n653 ;
  assign n12696 = n12695 ^ n12694 ^ n298 ;
  assign n12697 = n7882 ^ n5029 ^ n1035 ;
  assign n12698 = n12697 ^ n8106 ^ n3455 ;
  assign n12699 = n2180 & n3250 ;
  assign n12700 = n949 & n12699 ;
  assign n12701 = n8309 ^ n6085 ^ 1'b0 ;
  assign n12702 = ( ~n10806 & n12700 ) | ( ~n10806 & n12701 ) | ( n12700 & n12701 ) ;
  assign n12703 = ( n2971 & n12698 ) | ( n2971 & ~n12702 ) | ( n12698 & ~n12702 ) ;
  assign n12707 = ( ~n756 & n1075 ) | ( ~n756 & n1354 ) | ( n1075 & n1354 ) ;
  assign n12708 = ( ~n6023 & n6799 ) | ( ~n6023 & n12707 ) | ( n6799 & n12707 ) ;
  assign n12705 = n7525 | n8505 ;
  assign n12704 = ( n4366 & ~n11574 ) | ( n4366 & n11981 ) | ( ~n11574 & n11981 ) ;
  assign n12706 = n12705 ^ n12704 ^ n2389 ;
  assign n12709 = n12708 ^ n12706 ^ n4713 ;
  assign n12710 = n7338 ^ n6638 ^ n1019 ;
  assign n12711 = n6433 ^ n4167 ^ 1'b0 ;
  assign n12712 = n1308 | n12711 ;
  assign n12713 = ( n1137 & ~n4331 ) | ( n1137 & n4836 ) | ( ~n4331 & n4836 ) ;
  assign n12714 = n12713 ^ n10588 ^ n9424 ;
  assign n12715 = ( ~n12710 & n12712 ) | ( ~n12710 & n12714 ) | ( n12712 & n12714 ) ;
  assign n12721 = n3729 ^ n3380 ^ x121 ;
  assign n12716 = n8456 ^ n4656 ^ x53 ;
  assign n12717 = ( n2351 & n11219 ) | ( n2351 & n12716 ) | ( n11219 & n12716 ) ;
  assign n12718 = n12717 ^ n6639 ^ n1381 ;
  assign n12719 = n3719 & ~n11617 ;
  assign n12720 = n12718 & n12719 ;
  assign n12722 = n12721 ^ n12720 ^ n9867 ;
  assign n12723 = ~n1643 & n5392 ;
  assign n12724 = n1618 & n12723 ;
  assign n12725 = n10310 ^ n8645 ^ 1'b0 ;
  assign n12726 = n12725 ^ n859 ^ 1'b0 ;
  assign n12727 = n12724 | n12726 ;
  assign n12728 = n7444 & n12727 ;
  assign n12729 = n7980 ^ n5984 ^ n430 ;
  assign n12730 = ( n3914 & ~n10672 ) | ( n3914 & n12729 ) | ( ~n10672 & n12729 ) ;
  assign n12735 = ( n1181 & n4012 ) | ( n1181 & ~n5619 ) | ( n4012 & ~n5619 ) ;
  assign n12736 = n12735 ^ n11299 ^ n6162 ;
  assign n12731 = ( ~n1697 & n6952 ) | ( ~n1697 & n10729 ) | ( n6952 & n10729 ) ;
  assign n12732 = n12731 ^ n9421 ^ n6733 ;
  assign n12733 = n12732 ^ n8688 ^ n4636 ;
  assign n12734 = n9738 & n12733 ;
  assign n12737 = n12736 ^ n12734 ^ 1'b0 ;
  assign n12738 = ( n5179 & n11549 ) | ( n5179 & ~n11962 ) | ( n11549 & ~n11962 ) ;
  assign n12739 = n12738 ^ n12158 ^ n359 ;
  assign n12740 = n12739 ^ n10839 ^ 1'b0 ;
  assign n12741 = n5704 | n12740 ;
  assign n12742 = n7087 & n11298 ;
  assign n12743 = ( n624 & n1673 ) | ( n624 & n2662 ) | ( n1673 & n2662 ) ;
  assign n12744 = n12743 ^ n8022 ^ n2686 ;
  assign n12745 = n2027 & n12744 ;
  assign n12746 = n6882 & n12745 ;
  assign n12747 = n11400 ^ n8337 ^ n6938 ;
  assign n12749 = ( ~n1435 & n2049 ) | ( ~n1435 & n2377 ) | ( n2049 & n2377 ) ;
  assign n12750 = n2137 & n12749 ;
  assign n12751 = ~n11634 & n12750 ;
  assign n12748 = ( x6 & ~n2589 ) | ( x6 & n9365 ) | ( ~n2589 & n9365 ) ;
  assign n12752 = n12751 ^ n12748 ^ n11303 ;
  assign n12753 = n12752 ^ n489 ^ n420 ;
  assign n12758 = n7905 ^ n733 ^ n365 ;
  assign n12759 = ~n10669 & n12638 ;
  assign n12760 = n12758 & n12759 ;
  assign n12754 = ( n371 & ~n1650 ) | ( n371 & n2967 ) | ( ~n1650 & n2967 ) ;
  assign n12755 = n12754 ^ n5549 ^ n2523 ;
  assign n12756 = n5571 | n12755 ;
  assign n12757 = n8916 | n12756 ;
  assign n12761 = n12760 ^ n12757 ^ n313 ;
  assign n12762 = ( n4470 & ~n7522 ) | ( n4470 & n12761 ) | ( ~n7522 & n12761 ) ;
  assign n12763 = ( n2945 & n12753 ) | ( n2945 & n12762 ) | ( n12753 & n12762 ) ;
  assign n12764 = ~n12747 & n12763 ;
  assign n12765 = ( ~n4406 & n6570 ) | ( ~n4406 & n6752 ) | ( n6570 & n6752 ) ;
  assign n12766 = n6091 ^ n2035 ^ 1'b0 ;
  assign n12767 = n12766 ^ n2897 ^ n1714 ;
  assign n12768 = n1810 & ~n11688 ;
  assign n12769 = n1939 & n12768 ;
  assign n12770 = n1874 | n12769 ;
  assign n12771 = n12767 | n12770 ;
  assign n12772 = ( n8004 & n12765 ) | ( n8004 & ~n12771 ) | ( n12765 & ~n12771 ) ;
  assign n12773 = n12772 ^ n1811 ^ 1'b0 ;
  assign n12774 = ( ~n3980 & n7092 ) | ( ~n3980 & n12773 ) | ( n7092 & n12773 ) ;
  assign n12775 = n5991 ^ n2949 ^ n346 ;
  assign n12776 = n12775 ^ n3614 ^ n2661 ;
  assign n12777 = ( n1180 & n3085 ) | ( n1180 & n11505 ) | ( n3085 & n11505 ) ;
  assign n12778 = n12777 ^ n5882 ^ n828 ;
  assign n12779 = n6917 ^ n5979 ^ n257 ;
  assign n12780 = n922 ^ n544 ^ x73 ;
  assign n12781 = n4110 ^ n3443 ^ n2587 ;
  assign n12782 = ( n1607 & n12780 ) | ( n1607 & n12781 ) | ( n12780 & n12781 ) ;
  assign n12783 = ( n1662 & ~n12779 ) | ( n1662 & n12782 ) | ( ~n12779 & n12782 ) ;
  assign n12784 = ( n1403 & ~n1788 ) | ( n1403 & n9217 ) | ( ~n1788 & n9217 ) ;
  assign n12785 = ( x231 & ~n6650 ) | ( x231 & n12784 ) | ( ~n6650 & n12784 ) ;
  assign n12786 = ( n10688 & n12783 ) | ( n10688 & n12785 ) | ( n12783 & n12785 ) ;
  assign n12789 = ( n7428 & ~n8761 ) | ( n7428 & n11488 ) | ( ~n8761 & n11488 ) ;
  assign n12787 = ( n2994 & ~n4382 ) | ( n2994 & n6880 ) | ( ~n4382 & n6880 ) ;
  assign n12788 = n12787 ^ n9874 ^ n6819 ;
  assign n12790 = n12789 ^ n12788 ^ n4904 ;
  assign n12792 = ( ~n3532 & n7521 ) | ( ~n3532 & n9704 ) | ( n7521 & n9704 ) ;
  assign n12793 = ( n7698 & n12705 ) | ( n7698 & n12792 ) | ( n12705 & n12792 ) ;
  assign n12791 = n12462 ^ n9761 ^ x123 ;
  assign n12794 = n12793 ^ n12791 ^ n6583 ;
  assign n12795 = ( n3374 & n4921 ) | ( n3374 & ~n7252 ) | ( n4921 & ~n7252 ) ;
  assign n12796 = n4935 & ~n8336 ;
  assign n12797 = n12796 ^ n9716 ^ 1'b0 ;
  assign n12798 = ( x23 & ~n9265 ) | ( x23 & n12797 ) | ( ~n9265 & n12797 ) ;
  assign n12799 = n12798 ^ n1621 ^ x209 ;
  assign n12800 = ( n6803 & n12795 ) | ( n6803 & n12799 ) | ( n12795 & n12799 ) ;
  assign n12801 = n6524 ^ n3233 ^ n1745 ;
  assign n12802 = n7681 | n12801 ;
  assign n12803 = n12802 ^ n10418 ^ 1'b0 ;
  assign n12804 = ~n6263 & n12803 ;
  assign n12805 = n10774 ^ n6458 ^ n1345 ;
  assign n12808 = n11839 ^ n11709 ^ n1750 ;
  assign n12806 = ( n5128 & n5201 ) | ( n5128 & ~n11213 ) | ( n5201 & ~n11213 ) ;
  assign n12807 = n12806 ^ n7446 ^ n3522 ;
  assign n12809 = n12808 ^ n12807 ^ n11389 ;
  assign n12810 = ( n1543 & ~n4088 ) | ( n1543 & n4375 ) | ( ~n4088 & n4375 ) ;
  assign n12811 = x192 & n669 ;
  assign n12812 = n12811 ^ n1771 ^ 1'b0 ;
  assign n12813 = n409 | n2383 ;
  assign n12814 = n1578 & ~n12813 ;
  assign n12815 = ( n1649 & n5309 ) | ( n1649 & n12814 ) | ( n5309 & n12814 ) ;
  assign n12816 = n3566 ^ n2770 ^ n1636 ;
  assign n12817 = n12815 & ~n12816 ;
  assign n12818 = n12812 & n12817 ;
  assign n12819 = ( ~n618 & n623 ) | ( ~n618 & n1313 ) | ( n623 & n1313 ) ;
  assign n12820 = ~n12818 & n12819 ;
  assign n12821 = n12810 & n12820 ;
  assign n12822 = ( x26 & n3706 ) | ( x26 & n5730 ) | ( n3706 & n5730 ) ;
  assign n12823 = n12822 ^ n9471 ^ 1'b0 ;
  assign n12824 = n5244 ^ n4691 ^ n368 ;
  assign n12825 = ( n2826 & ~n12823 ) | ( n2826 & n12824 ) | ( ~n12823 & n12824 ) ;
  assign n12826 = ( n5321 & ~n12821 ) | ( n5321 & n12825 ) | ( ~n12821 & n12825 ) ;
  assign n12834 = n9390 ^ n6457 ^ n1732 ;
  assign n12835 = n12834 ^ n7525 ^ n430 ;
  assign n12836 = n12835 ^ n6907 ^ n6835 ;
  assign n12827 = ( n3443 & n4357 ) | ( n3443 & ~n4447 ) | ( n4357 & ~n4447 ) ;
  assign n12828 = ( ~n4428 & n10164 ) | ( ~n4428 & n12827 ) | ( n10164 & n12827 ) ;
  assign n12829 = n2953 & ~n3848 ;
  assign n12830 = n12829 ^ n9894 ^ 1'b0 ;
  assign n12831 = ( n1955 & ~n12828 ) | ( n1955 & n12830 ) | ( ~n12828 & n12830 ) ;
  assign n12832 = ( n2990 & n8221 ) | ( n2990 & ~n12831 ) | ( n8221 & ~n12831 ) ;
  assign n12833 = ( ~n897 & n10893 ) | ( ~n897 & n12832 ) | ( n10893 & n12832 ) ;
  assign n12837 = n12836 ^ n12833 ^ n3300 ;
  assign n12838 = n12837 ^ n8982 ^ x95 ;
  assign n12839 = ( ~n1422 & n1688 ) | ( ~n1422 & n5148 ) | ( n1688 & n5148 ) ;
  assign n12840 = ( n3415 & ~n6224 ) | ( n3415 & n12839 ) | ( ~n6224 & n12839 ) ;
  assign n12841 = ( n617 & n5680 ) | ( n617 & ~n12840 ) | ( n5680 & ~n12840 ) ;
  assign n12842 = ( n998 & n2493 ) | ( n998 & n12841 ) | ( n2493 & n12841 ) ;
  assign n12843 = n529 | n12017 ;
  assign n12844 = ~n12842 & n12843 ;
  assign n12845 = ~n1915 & n12844 ;
  assign n12846 = ( n1439 & n2384 ) | ( n1439 & ~n11521 ) | ( n2384 & ~n11521 ) ;
  assign n12847 = ( n1307 & ~n2922 ) | ( n1307 & n7545 ) | ( ~n2922 & n7545 ) ;
  assign n12848 = ( ~n9477 & n10531 ) | ( ~n9477 & n12847 ) | ( n10531 & n12847 ) ;
  assign n12849 = ( n480 & ~n5930 ) | ( n480 & n8600 ) | ( ~n5930 & n8600 ) ;
  assign n12850 = n12849 ^ n3664 ^ n2839 ;
  assign n12851 = x115 & n4680 ;
  assign n12852 = n333 & n12851 ;
  assign n12853 = ( n12848 & n12850 ) | ( n12848 & n12852 ) | ( n12850 & n12852 ) ;
  assign n12863 = ( n4382 & n5757 ) | ( n4382 & ~n9394 ) | ( n5757 & ~n9394 ) ;
  assign n12860 = n8463 ^ n3759 ^ 1'b0 ;
  assign n12861 = n5460 & ~n12860 ;
  assign n12862 = n12861 ^ n10482 ^ n10136 ;
  assign n12864 = n12863 ^ n12862 ^ n7053 ;
  assign n12856 = n7508 ^ n4661 ^ 1'b0 ;
  assign n12857 = n12084 | n12856 ;
  assign n12858 = n12857 ^ n6346 ^ n1474 ;
  assign n12854 = n5543 ^ n918 ^ 1'b0 ;
  assign n12855 = ( n1398 & n7786 ) | ( n1398 & n12854 ) | ( n7786 & n12854 ) ;
  assign n12859 = n12858 ^ n12855 ^ n11287 ;
  assign n12865 = n12864 ^ n12859 ^ n9293 ;
  assign n12866 = n12210 ^ n5474 ^ n2237 ;
  assign n12867 = ( ~n734 & n4259 ) | ( ~n734 & n4880 ) | ( n4259 & n4880 ) ;
  assign n12868 = ( ~n7615 & n9282 ) | ( ~n7615 & n12044 ) | ( n9282 & n12044 ) ;
  assign n12869 = ( ~n3473 & n12867 ) | ( ~n3473 & n12868 ) | ( n12867 & n12868 ) ;
  assign n12870 = ( n3625 & ~n12866 ) | ( n3625 & n12869 ) | ( ~n12866 & n12869 ) ;
  assign n12884 = n4582 ^ n1967 ^ n1756 ;
  assign n12881 = n3080 ^ n2821 ^ n397 ;
  assign n12882 = ( n905 & ~n8673 ) | ( n905 & n12881 ) | ( ~n8673 & n12881 ) ;
  assign n12879 = n4475 ^ n2684 ^ 1'b0 ;
  assign n12876 = n8876 ^ n3153 ^ n1939 ;
  assign n12877 = ~n10379 & n12876 ;
  assign n12878 = n12877 ^ n3135 ^ 1'b0 ;
  assign n12880 = n12879 ^ n12878 ^ n4658 ;
  assign n12883 = n12882 ^ n12880 ^ n2484 ;
  assign n12872 = ~n1296 & n2171 ;
  assign n12873 = n653 & n12872 ;
  assign n12871 = ( n917 & n5849 ) | ( n917 & ~n6721 ) | ( n5849 & ~n6721 ) ;
  assign n12874 = n12873 ^ n12871 ^ n5896 ;
  assign n12875 = n12874 ^ n2400 ^ 1'b0 ;
  assign n12885 = n12884 ^ n12883 ^ n12875 ;
  assign n12886 = n8150 ^ n2268 ^ 1'b0 ;
  assign n12891 = n11566 ^ n9069 ^ n2239 ;
  assign n12892 = ( x35 & n2934 ) | ( x35 & ~n12891 ) | ( n2934 & ~n12891 ) ;
  assign n12889 = n2927 ^ n1118 ^ n319 ;
  assign n12890 = n12889 ^ n12341 ^ n6339 ;
  assign n12887 = n7257 & n8530 ;
  assign n12888 = n12887 ^ n1336 ^ 1'b0 ;
  assign n12893 = n12892 ^ n12890 ^ n12888 ;
  assign n12895 = n6131 ^ n4726 ^ n4427 ;
  assign n12894 = n8630 & n8750 ;
  assign n12896 = n12895 ^ n12894 ^ 1'b0 ;
  assign n12897 = ( n2268 & n5450 ) | ( n2268 & ~n12896 ) | ( n5450 & ~n12896 ) ;
  assign n12898 = ( ~n11570 & n12893 ) | ( ~n11570 & n12897 ) | ( n12893 & n12897 ) ;
  assign n12899 = n1342 & n2599 ;
  assign n12900 = n3625 & n12899 ;
  assign n12901 = ( x24 & n5948 ) | ( x24 & n12900 ) | ( n5948 & n12900 ) ;
  assign n12902 = ( ~n2055 & n5445 ) | ( ~n2055 & n12901 ) | ( n5445 & n12901 ) ;
  assign n12903 = n12902 ^ n11451 ^ n7752 ;
  assign n12904 = ( n4333 & ~n5055 ) | ( n4333 & n10531 ) | ( ~n5055 & n10531 ) ;
  assign n12907 = n3567 ^ n1528 ^ n917 ;
  assign n12905 = ~n8195 & n9697 ;
  assign n12906 = n4079 & n12905 ;
  assign n12908 = n12907 ^ n12906 ^ 1'b0 ;
  assign n12909 = n12904 & ~n12908 ;
  assign n12910 = ( n8554 & n12903 ) | ( n8554 & ~n12909 ) | ( n12903 & ~n12909 ) ;
  assign n12911 = n3764 & n8040 ;
  assign n12912 = n12471 ^ n5290 ^ n1660 ;
  assign n12915 = ( n1607 & n4103 ) | ( n1607 & ~n10708 ) | ( n4103 & ~n10708 ) ;
  assign n12913 = n1974 ^ n1910 ^ n1401 ;
  assign n12914 = n12913 ^ n2178 ^ n2077 ;
  assign n12916 = n12915 ^ n12914 ^ n9664 ;
  assign n12917 = ( n12911 & n12912 ) | ( n12911 & ~n12916 ) | ( n12912 & ~n12916 ) ;
  assign n12918 = n6708 ^ n3274 ^ 1'b0 ;
  assign n12919 = x10 & n12918 ;
  assign n12920 = n1080 & n12919 ;
  assign n12921 = ( n4173 & n4269 ) | ( n4173 & n7987 ) | ( n4269 & n7987 ) ;
  assign n12922 = n12921 ^ n2244 ^ 1'b0 ;
  assign n12923 = n3670 & n12922 ;
  assign n12924 = n5029 & n12923 ;
  assign n12937 = n8407 ^ n993 ^ 1'b0 ;
  assign n12938 = ( ~n7740 & n9063 ) | ( ~n7740 & n12937 ) | ( n9063 & n12937 ) ;
  assign n12929 = n1553 ^ n781 ^ n548 ;
  assign n12930 = n12929 ^ n11300 ^ n4597 ;
  assign n12931 = n12930 ^ n9465 ^ n4937 ;
  assign n12932 = ( ~n1195 & n3225 ) | ( ~n1195 & n3713 ) | ( n3225 & n3713 ) ;
  assign n12933 = n12932 ^ n5814 ^ n4136 ;
  assign n12934 = n12933 ^ n11672 ^ 1'b0 ;
  assign n12935 = n3461 & ~n12934 ;
  assign n12936 = ( n6219 & n12931 ) | ( n6219 & n12935 ) | ( n12931 & n12935 ) ;
  assign n12927 = ( n7795 & n9310 ) | ( n7795 & ~n11156 ) | ( n9310 & ~n11156 ) ;
  assign n12925 = ~n6330 & n11986 ;
  assign n12926 = ( ~x127 & n5980 ) | ( ~x127 & n12925 ) | ( n5980 & n12925 ) ;
  assign n12928 = n12927 ^ n12926 ^ n7358 ;
  assign n12939 = n12938 ^ n12936 ^ n12928 ;
  assign n12940 = ( ~n755 & n4627 ) | ( ~n755 & n7066 ) | ( n4627 & n7066 ) ;
  assign n12941 = ( n9508 & ~n11097 ) | ( n9508 & n11863 ) | ( ~n11097 & n11863 ) ;
  assign n12942 = n12941 ^ n3184 ^ 1'b0 ;
  assign n12943 = ( n2785 & n4271 ) | ( n2785 & n11901 ) | ( n4271 & n11901 ) ;
  assign n12944 = n12943 ^ n5977 ^ n882 ;
  assign n12945 = ( n12940 & n12942 ) | ( n12940 & ~n12944 ) | ( n12942 & ~n12944 ) ;
  assign n12958 = n4098 | n8312 ;
  assign n12949 = n7278 ^ n4582 ^ x87 ;
  assign n12950 = n12949 ^ n6433 ^ n1970 ;
  assign n12951 = n12950 ^ n6957 ^ n1452 ;
  assign n12952 = ( ~n417 & n3279 ) | ( ~n417 & n3652 ) | ( n3279 & n3652 ) ;
  assign n12953 = n6251 | n12952 ;
  assign n12954 = n12953 ^ n8802 ^ 1'b0 ;
  assign n12955 = ( n5969 & n12951 ) | ( n5969 & n12954 ) | ( n12951 & n12954 ) ;
  assign n12946 = n4755 ^ n4308 ^ n2864 ;
  assign n12947 = ( n10635 & ~n11064 ) | ( n10635 & n12946 ) | ( ~n11064 & n12946 ) ;
  assign n12948 = n12947 ^ n11578 ^ 1'b0 ;
  assign n12956 = n12955 ^ n12948 ^ n4856 ;
  assign n12957 = ~n2342 & n12956 ;
  assign n12959 = n12958 ^ n12957 ^ n6695 ;
  assign n12966 = n12626 ^ n12395 ^ n6396 ;
  assign n12967 = n12966 ^ n10337 ^ n4197 ;
  assign n12960 = n7980 ^ n2320 ^ 1'b0 ;
  assign n12961 = n2704 | n8603 ;
  assign n12962 = ( n1072 & ~n2819 ) | ( n1072 & n12961 ) | ( ~n2819 & n12961 ) ;
  assign n12963 = ( n7290 & ~n7294 ) | ( n7290 & n12962 ) | ( ~n7294 & n12962 ) ;
  assign n12964 = n12963 ^ n10329 ^ n6484 ;
  assign n12965 = ( n10183 & n12960 ) | ( n10183 & ~n12964 ) | ( n12960 & ~n12964 ) ;
  assign n12968 = n12967 ^ n12965 ^ n1979 ;
  assign n12969 = n11100 ^ n9844 ^ n6557 ;
  assign n12970 = n12969 ^ n11260 ^ n1912 ;
  assign n12975 = n8758 ^ n4357 ^ n2664 ;
  assign n12973 = ( n2214 & n2799 ) | ( n2214 & ~n5282 ) | ( n2799 & ~n5282 ) ;
  assign n12972 = n4273 ^ n2600 ^ x133 ;
  assign n12971 = ( n427 & n7669 ) | ( n427 & n10444 ) | ( n7669 & n10444 ) ;
  assign n12974 = n12973 ^ n12972 ^ n12971 ;
  assign n12976 = n12975 ^ n12974 ^ n1865 ;
  assign n12979 = ( n2715 & n4520 ) | ( n2715 & ~n8221 ) | ( n4520 & ~n8221 ) ;
  assign n12978 = ( n4352 & n5821 ) | ( n4352 & ~n8201 ) | ( n5821 & ~n8201 ) ;
  assign n12980 = n12979 ^ n12978 ^ n9278 ;
  assign n12977 = n3056 & n11643 ;
  assign n12981 = n12980 ^ n12977 ^ n5796 ;
  assign n12984 = ( n2411 & n3692 ) | ( n2411 & ~n12662 ) | ( n3692 & ~n12662 ) ;
  assign n12982 = n8788 ^ n5667 ^ 1'b0 ;
  assign n12983 = n3999 | n12982 ;
  assign n12985 = n12984 ^ n12983 ^ n11099 ;
  assign n12994 = ~n2428 & n5725 ;
  assign n12995 = ( n8738 & n8802 ) | ( n8738 & n12994 ) | ( n8802 & n12994 ) ;
  assign n12988 = ( x75 & n4588 ) | ( x75 & ~n5286 ) | ( n4588 & ~n5286 ) ;
  assign n12989 = ( ~n2022 & n3780 ) | ( ~n2022 & n5017 ) | ( n3780 & n5017 ) ;
  assign n12990 = ( n1281 & n12988 ) | ( n1281 & ~n12989 ) | ( n12988 & ~n12989 ) ;
  assign n12987 = n5195 | n7206 ;
  assign n12991 = n12990 ^ n12987 ^ 1'b0 ;
  assign n12992 = n12991 ^ n3126 ^ 1'b0 ;
  assign n12986 = ( ~n2421 & n6659 ) | ( ~n2421 & n8640 ) | ( n6659 & n8640 ) ;
  assign n12993 = n12992 ^ n12986 ^ n2853 ;
  assign n12996 = n12995 ^ n12993 ^ n11956 ;
  assign n12997 = ( n1614 & n12985 ) | ( n1614 & n12996 ) | ( n12985 & n12996 ) ;
  assign n12998 = n7088 ^ n4542 ^ x48 ;
  assign n12999 = ( n6347 & n9778 ) | ( n6347 & n10057 ) | ( n9778 & n10057 ) ;
  assign n13000 = ~n12998 & n12999 ;
  assign n13001 = n8003 ^ n3941 ^ n3928 ;
  assign n13006 = n11451 ^ n3042 ^ n973 ;
  assign n13007 = n13006 ^ n7867 ^ 1'b0 ;
  assign n13002 = ( n2508 & n3630 ) | ( n2508 & ~n5560 ) | ( n3630 & ~n5560 ) ;
  assign n13003 = ( n2851 & ~n11014 ) | ( n2851 & n13002 ) | ( ~n11014 & n13002 ) ;
  assign n13004 = ( ~n1705 & n9593 ) | ( ~n1705 & n13003 ) | ( n9593 & n13003 ) ;
  assign n13005 = n13004 ^ n6121 ^ n3002 ;
  assign n13008 = n13007 ^ n13005 ^ n3209 ;
  assign n13009 = n12510 ^ n11100 ^ n3333 ;
  assign n13010 = ( ~n3572 & n5756 ) | ( ~n3572 & n7328 ) | ( n5756 & n7328 ) ;
  assign n13011 = ( n2941 & n12919 ) | ( n2941 & ~n13010 ) | ( n12919 & ~n13010 ) ;
  assign n13020 = ( n3260 & ~n6467 ) | ( n3260 & n6951 ) | ( ~n6467 & n6951 ) ;
  assign n13012 = n3272 ^ n1155 ^ 1'b0 ;
  assign n13013 = n10580 ^ n4075 ^ 1'b0 ;
  assign n13014 = n13012 & ~n13013 ;
  assign n13015 = n4828 ^ x104 ^ x101 ;
  assign n13016 = n13015 ^ n1986 ^ n641 ;
  assign n13017 = ( x110 & n2535 ) | ( x110 & ~n13016 ) | ( n2535 & ~n13016 ) ;
  assign n13018 = n10965 & ~n13017 ;
  assign n13019 = ~n13014 & n13018 ;
  assign n13021 = n13020 ^ n13019 ^ 1'b0 ;
  assign n13025 = n12330 ^ n4819 ^ 1'b0 ;
  assign n13022 = ~n3562 & n8639 ;
  assign n13023 = ~n11864 & n13022 ;
  assign n13024 = n681 | n13023 ;
  assign n13026 = n13025 ^ n13024 ^ 1'b0 ;
  assign n13027 = ~n6375 & n13026 ;
  assign n13028 = n13027 ^ n1471 ^ 1'b0 ;
  assign n13029 = ( n800 & n2532 ) | ( n800 & ~n10509 ) | ( n2532 & ~n10509 ) ;
  assign n13030 = n12182 ^ n7378 ^ n5301 ;
  assign n13031 = n13030 ^ n7722 ^ n4420 ;
  assign n13032 = ( n7702 & n9128 ) | ( n7702 & ~n13031 ) | ( n9128 & ~n13031 ) ;
  assign n13033 = n10701 ^ n3050 ^ n2360 ;
  assign n13040 = n4403 ^ n4342 ^ n3905 ;
  assign n13038 = x234 & n8947 ;
  assign n13039 = n2384 & n13038 ;
  assign n13034 = n6039 ^ n5746 ^ n895 ;
  assign n13035 = n13034 ^ n9985 ^ n4402 ;
  assign n13036 = n7279 ^ n6884 ^ n3800 ;
  assign n13037 = ( n6947 & ~n13035 ) | ( n6947 & n13036 ) | ( ~n13035 & n13036 ) ;
  assign n13041 = n13040 ^ n13039 ^ n13037 ;
  assign n13047 = n3526 ^ n2225 ^ n1157 ;
  assign n13048 = ( n4423 & n10993 ) | ( n4423 & n13047 ) | ( n10993 & n13047 ) ;
  assign n13049 = ( n652 & n4033 ) | ( n652 & ~n13048 ) | ( n4033 & ~n13048 ) ;
  assign n13042 = ( ~n1014 & n1340 ) | ( ~n1014 & n1861 ) | ( n1340 & n1861 ) ;
  assign n13043 = ( n2360 & n3153 ) | ( n2360 & n4583 ) | ( n3153 & n4583 ) ;
  assign n13044 = n13042 | n13043 ;
  assign n13045 = n13044 ^ n9381 ^ n7732 ;
  assign n13046 = n13045 ^ n12892 ^ n7225 ;
  assign n13050 = n13049 ^ n13046 ^ n12080 ;
  assign n13051 = ( n1985 & n6617 ) | ( n1985 & ~n8171 ) | ( n6617 & ~n8171 ) ;
  assign n13052 = n13051 ^ n1866 ^ n1599 ;
  assign n13053 = ( n467 & ~n3735 ) | ( n467 & n10549 ) | ( ~n3735 & n10549 ) ;
  assign n13054 = ( n6094 & n13052 ) | ( n6094 & ~n13053 ) | ( n13052 & ~n13053 ) ;
  assign n13055 = n13054 ^ n5308 ^ n2039 ;
  assign n13059 = ( n3698 & ~n6200 ) | ( n3698 & n6565 ) | ( ~n6200 & n6565 ) ;
  assign n13058 = ( n1968 & n5983 ) | ( n1968 & n6261 ) | ( n5983 & n6261 ) ;
  assign n13060 = n13059 ^ n13058 ^ 1'b0 ;
  assign n13056 = n1517 | n10185 ;
  assign n13057 = n13056 ^ n5480 ^ 1'b0 ;
  assign n13061 = n13060 ^ n13057 ^ n10358 ;
  assign n13062 = ( n4733 & n8220 ) | ( n4733 & ~n12388 ) | ( n8220 & ~n12388 ) ;
  assign n13063 = n5550 ^ n1833 ^ n560 ;
  assign n13067 = ( x192 & n2332 ) | ( x192 & n9299 ) | ( n2332 & n9299 ) ;
  assign n13068 = n13067 ^ n7019 ^ n3770 ;
  assign n13064 = n6501 ^ n5005 ^ n451 ;
  assign n13065 = ( n2744 & n8469 ) | ( n2744 & ~n13064 ) | ( n8469 & ~n13064 ) ;
  assign n13066 = n10852 & ~n13065 ;
  assign n13069 = n13068 ^ n13066 ^ 1'b0 ;
  assign n13070 = ( n9042 & n13063 ) | ( n9042 & ~n13069 ) | ( n13063 & ~n13069 ) ;
  assign n13078 = n453 & ~n1648 ;
  assign n13079 = n13078 ^ n6147 ^ n2625 ;
  assign n13071 = ( x239 & n1447 ) | ( x239 & n2391 ) | ( n1447 & n2391 ) ;
  assign n13072 = n10523 & ~n11007 ;
  assign n13073 = n13071 & n13072 ;
  assign n13074 = n13073 ^ n5369 ^ 1'b0 ;
  assign n13075 = ~n12682 & n13074 ;
  assign n13076 = ( n1406 & n6394 ) | ( n1406 & ~n11610 ) | ( n6394 & ~n11610 ) ;
  assign n13077 = ( n3353 & n13075 ) | ( n3353 & n13076 ) | ( n13075 & n13076 ) ;
  assign n13080 = n13079 ^ n13077 ^ n7560 ;
  assign n13081 = ( n2872 & ~n3861 ) | ( n2872 & n4361 ) | ( ~n3861 & n4361 ) ;
  assign n13082 = ( n3095 & n5017 ) | ( n3095 & n13081 ) | ( n5017 & n13081 ) ;
  assign n13083 = n13082 ^ n7902 ^ n2125 ;
  assign n13084 = n10364 ^ n9826 ^ n276 ;
  assign n13087 = n10667 ^ n10598 ^ n3209 ;
  assign n13085 = n7753 ^ n5170 ^ x47 ;
  assign n13086 = ( n1517 & n8207 ) | ( n1517 & n13085 ) | ( n8207 & n13085 ) ;
  assign n13088 = n13087 ^ n13086 ^ n8673 ;
  assign n13089 = n13084 | n13088 ;
  assign n13090 = n9154 | n13089 ;
  assign n13091 = n13090 ^ n3475 ^ n478 ;
  assign n13092 = n12259 ^ n9919 ^ n3514 ;
  assign n13093 = n13092 ^ n11299 ^ n10355 ;
  assign n13094 = n13093 ^ n1188 ^ n410 ;
  assign n13095 = ( n3734 & n4856 ) | ( n3734 & ~n8772 ) | ( n4856 & ~n8772 ) ;
  assign n13096 = ( n3224 & n10251 ) | ( n3224 & ~n13095 ) | ( n10251 & ~n13095 ) ;
  assign n13097 = ( n1702 & ~n5814 ) | ( n1702 & n13096 ) | ( ~n5814 & n13096 ) ;
  assign n13098 = ( n5679 & n13086 ) | ( n5679 & n13097 ) | ( n13086 & n13097 ) ;
  assign n13099 = n13098 ^ n7683 ^ n7332 ;
  assign n13100 = ( n2799 & ~n8271 ) | ( n2799 & n13099 ) | ( ~n8271 & n13099 ) ;
  assign n13101 = n10324 | n13100 ;
  assign n13102 = x34 | n13101 ;
  assign n13103 = n7790 ^ n5843 ^ 1'b0 ;
  assign n13104 = ( n1187 & n1974 ) | ( n1187 & n2200 ) | ( n1974 & n2200 ) ;
  assign n13105 = ( n3073 & ~n3891 ) | ( n3073 & n13104 ) | ( ~n3891 & n13104 ) ;
  assign n13106 = n13105 ^ n9100 ^ 1'b0 ;
  assign n13107 = n13103 & n13106 ;
  assign n13108 = n13107 ^ n5997 ^ 1'b0 ;
  assign n13109 = n13108 ^ n7727 ^ n4786 ;
  assign n13124 = n6172 ^ n5267 ^ n357 ;
  assign n13110 = n10410 ^ n7250 ^ n5474 ;
  assign n13111 = n4516 ^ n4273 ^ 1'b0 ;
  assign n13112 = ~n4246 & n13111 ;
  assign n13113 = n3801 ^ n3082 ^ x248 ;
  assign n13114 = n12285 ^ n3116 ^ n1998 ;
  assign n13115 = ~n6252 & n13114 ;
  assign n13116 = ~n13113 & n13115 ;
  assign n13117 = ( ~n13110 & n13112 ) | ( ~n13110 & n13116 ) | ( n13112 & n13116 ) ;
  assign n13118 = n11529 ^ n8585 ^ n5053 ;
  assign n13119 = ( n3297 & n3751 ) | ( n3297 & ~n4208 ) | ( n3751 & ~n4208 ) ;
  assign n13120 = ( n10260 & n13118 ) | ( n10260 & ~n13119 ) | ( n13118 & ~n13119 ) ;
  assign n13121 = n10143 ^ n2387 ^ n1196 ;
  assign n13122 = ( n13117 & ~n13120 ) | ( n13117 & n13121 ) | ( ~n13120 & n13121 ) ;
  assign n13123 = n13122 ^ n6554 ^ 1'b0 ;
  assign n13125 = n13124 ^ n13123 ^ n6672 ;
  assign n13126 = n8625 ^ n3403 ^ n851 ;
  assign n13127 = ( ~x156 & n305 ) | ( ~x156 & n1831 ) | ( n305 & n1831 ) ;
  assign n13128 = ( n678 & n3282 ) | ( n678 & ~n4287 ) | ( n3282 & ~n4287 ) ;
  assign n13129 = ( n8502 & ~n13127 ) | ( n8502 & n13128 ) | ( ~n13127 & n13128 ) ;
  assign n13130 = ( ~x120 & n3635 ) | ( ~x120 & n13129 ) | ( n3635 & n13129 ) ;
  assign n13131 = n13130 ^ n11781 ^ n8300 ;
  assign n13132 = ( n3585 & ~n4331 ) | ( n3585 & n5319 ) | ( ~n4331 & n5319 ) ;
  assign n13140 = n2243 ^ n2122 ^ n940 ;
  assign n13141 = n13140 ^ n4145 ^ n1714 ;
  assign n13142 = n6123 & n13141 ;
  assign n13143 = n1954 & n13142 ;
  assign n13144 = n13143 ^ n3056 ^ n2948 ;
  assign n13145 = n13144 ^ n3895 ^ 1'b0 ;
  assign n13146 = n11254 | n13145 ;
  assign n13137 = x31 & ~n6985 ;
  assign n13138 = n13137 ^ n1579 ^ 1'b0 ;
  assign n13133 = n5855 ^ n5033 ^ n3823 ;
  assign n13134 = n13133 ^ n8159 ^ n5106 ;
  assign n13135 = ( n4825 & n12783 ) | ( n4825 & ~n13134 ) | ( n12783 & ~n13134 ) ;
  assign n13136 = n13135 ^ n8065 ^ n6435 ;
  assign n13139 = n13138 ^ n13136 ^ n4702 ;
  assign n13147 = n13146 ^ n13139 ^ n9587 ;
  assign n13148 = ( n12688 & n13132 ) | ( n12688 & ~n13147 ) | ( n13132 & ~n13147 ) ;
  assign n13149 = ( ~x210 & n2549 ) | ( ~x210 & n12512 ) | ( n2549 & n12512 ) ;
  assign n13150 = n13149 ^ n8821 ^ n1082 ;
  assign n13151 = n2397 ^ n2038 ^ n829 ;
  assign n13152 = n13151 ^ n6557 ^ n4177 ;
  assign n13153 = n2552 ^ n522 ^ x106 ;
  assign n13154 = ( ~n10354 & n12731 ) | ( ~n10354 & n13153 ) | ( n12731 & n13153 ) ;
  assign n13155 = ( n12331 & n13152 ) | ( n12331 & n13154 ) | ( n13152 & n13154 ) ;
  assign n13156 = ( n6454 & n9389 ) | ( n6454 & n13155 ) | ( n9389 & n13155 ) ;
  assign n13160 = ( n3325 & n6819 ) | ( n3325 & ~n8553 ) | ( n6819 & ~n8553 ) ;
  assign n13157 = n7889 ^ n6021 ^ n2296 ;
  assign n13158 = ( n1302 & n2074 ) | ( n1302 & ~n12991 ) | ( n2074 & ~n12991 ) ;
  assign n13159 = ( n2682 & ~n13157 ) | ( n2682 & n13158 ) | ( ~n13157 & n13158 ) ;
  assign n13161 = n13160 ^ n13159 ^ n13048 ;
  assign n13163 = n7743 ^ n5477 ^ n4141 ;
  assign n13164 = n13163 ^ n8930 ^ n2340 ;
  assign n13162 = ( n1612 & ~n6045 ) | ( n1612 & n12411 ) | ( ~n6045 & n12411 ) ;
  assign n13165 = n13164 ^ n13162 ^ 1'b0 ;
  assign n13166 = ~n955 & n13165 ;
  assign n13167 = n13166 ^ n9970 ^ 1'b0 ;
  assign n13168 = ~n12715 & n13167 ;
  assign n13169 = ( x249 & n6822 ) | ( x249 & n10570 ) | ( n6822 & n10570 ) ;
  assign n13170 = n5679 & ~n7103 ;
  assign n13171 = ~n13169 & n13170 ;
  assign n13172 = ( n5870 & n12594 ) | ( n5870 & n13171 ) | ( n12594 & n13171 ) ;
  assign n13173 = n11835 ^ n4082 ^ x80 ;
  assign n13174 = n13173 ^ n9907 ^ n6385 ;
  assign n13175 = ( n1397 & n1512 ) | ( n1397 & ~n2237 ) | ( n1512 & ~n2237 ) ;
  assign n13176 = n11075 & ~n13175 ;
  assign n13177 = ( n9032 & n11097 ) | ( n9032 & ~n13176 ) | ( n11097 & ~n13176 ) ;
  assign n13178 = n13177 ^ n6326 ^ n5422 ;
  assign n13179 = n13118 ^ n5625 ^ n5392 ;
  assign n13180 = n13179 ^ n11382 ^ n9055 ;
  assign n13181 = ( n3259 & n10746 ) | ( n3259 & n13180 ) | ( n10746 & n13180 ) ;
  assign n13182 = ( n5678 & n11340 ) | ( n5678 & n13181 ) | ( n11340 & n13181 ) ;
  assign n13183 = ( ~n1695 & n13178 ) | ( ~n1695 & n13182 ) | ( n13178 & n13182 ) ;
  assign n13191 = n2752 & n3904 ;
  assign n13192 = n13191 ^ n4464 ^ 1'b0 ;
  assign n13185 = n4961 ^ n3469 ^ n361 ;
  assign n13186 = n13185 ^ n9597 ^ n6244 ;
  assign n13187 = ( n1465 & n4617 ) | ( n1465 & n13186 ) | ( n4617 & n13186 ) ;
  assign n13188 = n5575 & ~n13187 ;
  assign n13189 = n13188 ^ n6368 ^ 1'b0 ;
  assign n13184 = n7387 ^ n3509 ^ 1'b0 ;
  assign n13190 = n13189 ^ n13184 ^ n1416 ;
  assign n13193 = n13192 ^ n13190 ^ n7511 ;
  assign n13196 = n10346 ^ n3653 ^ n1718 ;
  assign n13194 = x75 & n8335 ;
  assign n13195 = n2983 & n13194 ;
  assign n13197 = n13196 ^ n13195 ^ n4615 ;
  assign n13198 = ( n3736 & n4224 ) | ( n3736 & n4511 ) | ( n4224 & n4511 ) ;
  assign n13199 = n3787 ^ n1734 ^ 1'b0 ;
  assign n13200 = ~n13198 & n13199 ;
  assign n13204 = n4729 ^ n3489 ^ x105 ;
  assign n13203 = n8740 ^ n1489 ^ 1'b0 ;
  assign n13201 = ( n5997 & n11114 ) | ( n5997 & n11562 ) | ( n11114 & n11562 ) ;
  assign n13202 = n13201 ^ n5511 ^ n536 ;
  assign n13205 = n13204 ^ n13203 ^ n13202 ;
  assign n13210 = n12441 ^ n12350 ^ n7473 ;
  assign n13208 = ~n2184 & n3916 ;
  assign n13209 = ( ~n2389 & n8588 ) | ( ~n2389 & n13208 ) | ( n8588 & n13208 ) ;
  assign n13206 = n3804 ^ n2479 ^ n1217 ;
  assign n13207 = n13206 ^ n11215 ^ n7103 ;
  assign n13211 = n13210 ^ n13209 ^ n13207 ;
  assign n13219 = n6676 ^ n2844 ^ n433 ;
  assign n13220 = ( n9882 & ~n10134 ) | ( n9882 & n13219 ) | ( ~n10134 & n13219 ) ;
  assign n13217 = n7956 ^ n3038 ^ n809 ;
  assign n13216 = n12932 ^ n7658 ^ 1'b0 ;
  assign n13218 = n13217 ^ n13216 ^ n5198 ;
  assign n13212 = n4433 ^ n2449 ^ n2025 ;
  assign n13213 = ( n1409 & n2843 ) | ( n1409 & n9934 ) | ( n2843 & n9934 ) ;
  assign n13214 = n9865 & ~n13213 ;
  assign n13215 = ( n8902 & ~n13212 ) | ( n8902 & n13214 ) | ( ~n13212 & n13214 ) ;
  assign n13221 = n13220 ^ n13218 ^ n13215 ;
  assign n13222 = n10820 ^ n6367 ^ n4544 ;
  assign n13223 = ~n4772 & n8248 ;
  assign n13224 = n13223 ^ n3837 ^ n1698 ;
  assign n13225 = ( n5479 & ~n9499 ) | ( n5479 & n13224 ) | ( ~n9499 & n13224 ) ;
  assign n13226 = n13225 ^ n9412 ^ n1484 ;
  assign n13227 = ~n10326 & n13226 ;
  assign n13228 = ( n3608 & ~n13222 ) | ( n3608 & n13227 ) | ( ~n13222 & n13227 ) ;
  assign n13229 = n10643 ^ n7286 ^ n496 ;
  assign n13230 = n6141 | n13229 ;
  assign n13231 = n13230 ^ n9521 ^ 1'b0 ;
  assign n13232 = ( x92 & n654 ) | ( x92 & ~n969 ) | ( n654 & ~n969 ) ;
  assign n13233 = n12674 ^ n4651 ^ n2235 ;
  assign n13234 = n8398 ^ n7771 ^ 1'b0 ;
  assign n13235 = n13233 | n13234 ;
  assign n13236 = ( n5121 & n13232 ) | ( n5121 & ~n13235 ) | ( n13232 & ~n13235 ) ;
  assign n13237 = ( n9399 & ~n13231 ) | ( n9399 & n13236 ) | ( ~n13231 & n13236 ) ;
  assign n13238 = n5818 & n10442 ;
  assign n13239 = n2158 & n13238 ;
  assign n13240 = ( n7299 & n10058 ) | ( n7299 & ~n13239 ) | ( n10058 & ~n13239 ) ;
  assign n13241 = n13240 ^ n10651 ^ n5391 ;
  assign n13242 = n6084 ^ n5719 ^ n2061 ;
  assign n13243 = n5850 ^ n1647 ^ 1'b0 ;
  assign n13244 = n4774 | n13243 ;
  assign n13245 = ( ~n518 & n13242 ) | ( ~n518 & n13244 ) | ( n13242 & n13244 ) ;
  assign n13246 = ( n7764 & ~n7962 ) | ( n7764 & n13245 ) | ( ~n7962 & n13245 ) ;
  assign n13247 = n13246 ^ n4095 ^ 1'b0 ;
  assign n13248 = n2341 & n13247 ;
  assign n13249 = ~n10266 & n13248 ;
  assign n13250 = n13249 ^ n10646 ^ 1'b0 ;
  assign n13252 = n2034 ^ n1741 ^ n1184 ;
  assign n13251 = ( n3493 & n11256 ) | ( n3493 & n12220 ) | ( n11256 & n12220 ) ;
  assign n13253 = n13252 ^ n13251 ^ n6085 ;
  assign n13254 = ( n2385 & ~n6334 ) | ( n2385 & n13253 ) | ( ~n6334 & n13253 ) ;
  assign n13256 = n5907 ^ n5730 ^ n1729 ;
  assign n13257 = ( n602 & n1838 ) | ( n602 & ~n13256 ) | ( n1838 & ~n13256 ) ;
  assign n13258 = ( n3849 & n4029 ) | ( n3849 & n13257 ) | ( n4029 & n13257 ) ;
  assign n13255 = n8838 & n12528 ;
  assign n13259 = n13258 ^ n13255 ^ 1'b0 ;
  assign n13260 = ( n2561 & n8468 ) | ( n2561 & n8546 ) | ( n8468 & n8546 ) ;
  assign n13261 = n13260 ^ n10071 ^ n3025 ;
  assign n13262 = ( x201 & n5324 ) | ( x201 & n13261 ) | ( n5324 & n13261 ) ;
  assign n13263 = ( n12577 & n13259 ) | ( n12577 & ~n13262 ) | ( n13259 & ~n13262 ) ;
  assign n13264 = ( ~n1503 & n2793 ) | ( ~n1503 & n4945 ) | ( n2793 & n4945 ) ;
  assign n13265 = n13264 ^ n5403 ^ n5093 ;
  assign n13266 = ( ~n3808 & n6855 ) | ( ~n3808 & n12245 ) | ( n6855 & n12245 ) ;
  assign n13267 = n2104 | n13266 ;
  assign n13268 = n1339 ^ x169 ^ 1'b0 ;
  assign n13269 = ( n6527 & ~n10260 ) | ( n6527 & n12336 ) | ( ~n10260 & n12336 ) ;
  assign n13270 = ( n2122 & n12625 ) | ( n2122 & ~n13269 ) | ( n12625 & ~n13269 ) ;
  assign n13271 = ( ~n3554 & n4740 ) | ( ~n3554 & n12674 ) | ( n4740 & n12674 ) ;
  assign n13272 = n11254 ^ n3064 ^ x131 ;
  assign n13273 = n6435 & n13272 ;
  assign n13274 = ~n9958 & n13273 ;
  assign n13275 = n4143 ^ n2818 ^ n846 ;
  assign n13276 = ( ~n3782 & n13274 ) | ( ~n3782 & n13275 ) | ( n13274 & n13275 ) ;
  assign n13277 = ( ~n4863 & n13271 ) | ( ~n4863 & n13276 ) | ( n13271 & n13276 ) ;
  assign n13278 = n7817 ^ n7807 ^ 1'b0 ;
  assign n13279 = ( ~n2521 & n5738 ) | ( ~n2521 & n9048 ) | ( n5738 & n9048 ) ;
  assign n13280 = n13222 ^ n8854 ^ n8536 ;
  assign n13285 = n8536 ^ n1603 ^ n623 ;
  assign n13281 = n11557 ^ n3266 ^ n1490 ;
  assign n13282 = n13281 ^ n476 ^ 1'b0 ;
  assign n13283 = n2614 ^ n2412 ^ n1283 ;
  assign n13284 = ( ~n4148 & n13282 ) | ( ~n4148 & n13283 ) | ( n13282 & n13283 ) ;
  assign n13286 = n13285 ^ n13284 ^ n12570 ;
  assign n13287 = ~x74 & n4214 ;
  assign n13288 = ( n3691 & n5240 ) | ( n3691 & n13287 ) | ( n5240 & n13287 ) ;
  assign n13289 = n13288 ^ n1544 ^ 1'b0 ;
  assign n13290 = ( ~n3776 & n6477 ) | ( ~n3776 & n12841 ) | ( n6477 & n12841 ) ;
  assign n13291 = n9677 ^ n3862 ^ x64 ;
  assign n13292 = n13291 ^ n13164 ^ n5386 ;
  assign n13293 = n13292 ^ n12038 ^ n7609 ;
  assign n13294 = n13293 ^ n8223 ^ n6898 ;
  assign n13295 = ( ~n3499 & n12229 ) | ( ~n3499 & n13294 ) | ( n12229 & n13294 ) ;
  assign n13302 = ( n561 & ~n5238 ) | ( n561 & n9389 ) | ( ~n5238 & n9389 ) ;
  assign n13300 = n4401 ^ n4160 ^ n1698 ;
  assign n13299 = ( ~n1056 & n6455 ) | ( ~n1056 & n7921 ) | ( n6455 & n7921 ) ;
  assign n13296 = ( ~n10170 & n10603 ) | ( ~n10170 & n13176 ) | ( n10603 & n13176 ) ;
  assign n13297 = ~n11848 & n13296 ;
  assign n13298 = ~n11263 & n13297 ;
  assign n13301 = n13300 ^ n13299 ^ n13298 ;
  assign n13303 = n13302 ^ n13301 ^ n12242 ;
  assign n13304 = n6958 ^ n5135 ^ x155 ;
  assign n13305 = ( n8699 & n12900 ) | ( n8699 & n13304 ) | ( n12900 & n13304 ) ;
  assign n13306 = n5400 ^ n1623 ^ 1'b0 ;
  assign n13309 = ~n3870 & n7044 ;
  assign n13310 = n725 & ~n13309 ;
  assign n13311 = n13310 ^ n12716 ^ 1'b0 ;
  assign n13307 = ( n1751 & ~n2643 ) | ( n1751 & n8103 ) | ( ~n2643 & n8103 ) ;
  assign n13308 = ( n1270 & n5885 ) | ( n1270 & n13307 ) | ( n5885 & n13307 ) ;
  assign n13312 = n13311 ^ n13308 ^ 1'b0 ;
  assign n13313 = ( n6154 & n9032 ) | ( n6154 & ~n13312 ) | ( n9032 & ~n13312 ) ;
  assign n13314 = n3581 ^ x58 ^ 1'b0 ;
  assign n13315 = n4387 | n13314 ;
  assign n13316 = n13315 ^ n3471 ^ 1'b0 ;
  assign n13319 = ( ~n1987 & n2087 ) | ( ~n1987 & n6164 ) | ( n2087 & n6164 ) ;
  assign n13320 = n3731 | n13319 ;
  assign n13321 = n13320 ^ n422 ^ 1'b0 ;
  assign n13322 = n13321 ^ n4245 ^ 1'b0 ;
  assign n13317 = n5804 ^ n3751 ^ 1'b0 ;
  assign n13318 = n13052 & ~n13317 ;
  assign n13323 = n13322 ^ n13318 ^ n8857 ;
  assign n13324 = ( n13313 & ~n13316 ) | ( n13313 & n13323 ) | ( ~n13316 & n13323 ) ;
  assign n13325 = n8660 & ~n13324 ;
  assign n13326 = ~n881 & n13325 ;
  assign n13327 = ( n3410 & n5452 ) | ( n3410 & n8412 ) | ( n5452 & n8412 ) ;
  assign n13330 = ( x107 & n1154 ) | ( x107 & ~n2464 ) | ( n1154 & ~n2464 ) ;
  assign n13331 = n13330 ^ n4653 ^ n1487 ;
  assign n13328 = ( n1435 & ~n9939 ) | ( n1435 & n10296 ) | ( ~n9939 & n10296 ) ;
  assign n13329 = ( n5740 & ~n12384 ) | ( n5740 & n13328 ) | ( ~n12384 & n13328 ) ;
  assign n13332 = n13331 ^ n13329 ^ n9272 ;
  assign n13334 = ( n3290 & n4864 ) | ( n3290 & n10770 ) | ( n4864 & n10770 ) ;
  assign n13335 = n13334 ^ n3339 ^ n2822 ;
  assign n13333 = n1264 & n3690 ;
  assign n13336 = n13335 ^ n13333 ^ 1'b0 ;
  assign n13337 = n5237 ^ n1734 ^ n1165 ;
  assign n13338 = n1507 | n5152 ;
  assign n13339 = n13337 & ~n13338 ;
  assign n13340 = ( ~n411 & n2278 ) | ( ~n411 & n4402 ) | ( n2278 & n4402 ) ;
  assign n13341 = ( ~n857 & n1097 ) | ( ~n857 & n6347 ) | ( n1097 & n6347 ) ;
  assign n13342 = ( n534 & ~n11272 ) | ( n534 & n13341 ) | ( ~n11272 & n13341 ) ;
  assign n13343 = n9741 ^ n1009 ^ 1'b0 ;
  assign n13344 = n13342 & n13343 ;
  assign n13348 = x165 & ~n6894 ;
  assign n13345 = ( ~n1623 & n8302 ) | ( ~n1623 & n9279 ) | ( n8302 & n9279 ) ;
  assign n13346 = ~n1851 & n3307 ;
  assign n13347 = n13345 & n13346 ;
  assign n13349 = n13348 ^ n13347 ^ n9616 ;
  assign n13350 = ( n13340 & ~n13344 ) | ( n13340 & n13349 ) | ( ~n13344 & n13349 ) ;
  assign n13352 = ( n6665 & ~n7251 ) | ( n6665 & n8158 ) | ( ~n7251 & n8158 ) ;
  assign n13351 = ( n1594 & n3921 ) | ( n1594 & ~n7634 ) | ( n3921 & ~n7634 ) ;
  assign n13353 = n13352 ^ n13351 ^ 1'b0 ;
  assign n13357 = n7737 ^ n5739 ^ x109 ;
  assign n13358 = n13357 ^ n13034 ^ n3983 ;
  assign n13359 = n7791 & ~n13358 ;
  assign n13354 = ( ~n1420 & n1684 ) | ( ~n1420 & n6029 ) | ( n1684 & n6029 ) ;
  assign n13355 = n13354 ^ n4473 ^ 1'b0 ;
  assign n13356 = ~n5134 & n13355 ;
  assign n13360 = n13359 ^ n13356 ^ n3535 ;
  assign n13361 = ( n12302 & ~n13353 ) | ( n12302 & n13360 ) | ( ~n13353 & n13360 ) ;
  assign n13362 = ( n8769 & n11775 ) | ( n8769 & ~n13361 ) | ( n11775 & ~n13361 ) ;
  assign n13363 = ( n5570 & n6834 ) | ( n5570 & n11030 ) | ( n6834 & n11030 ) ;
  assign n13369 = ( n2113 & n6273 ) | ( n2113 & n7725 ) | ( n6273 & n7725 ) ;
  assign n13370 = ( ~n3790 & n5452 ) | ( ~n3790 & n13369 ) | ( n5452 & n13369 ) ;
  assign n13366 = ~n7977 & n10862 ;
  assign n13367 = n13366 ^ n675 ^ 1'b0 ;
  assign n13364 = n2583 | n3790 ;
  assign n13365 = n13364 ^ n11683 ^ x12 ;
  assign n13368 = n13367 ^ n13365 ^ n3711 ;
  assign n13371 = n13370 ^ n13368 ^ n8666 ;
  assign n13372 = n13363 | n13371 ;
  assign n13373 = n8232 & ~n13372 ;
  assign n13374 = n8159 | n13373 ;
  assign n13375 = n13374 ^ n10205 ^ 1'b0 ;
  assign n13378 = n4784 ^ n4292 ^ n370 ;
  assign n13376 = n7333 | n9268 ;
  assign n13377 = ( n2759 & n12903 ) | ( n2759 & n13376 ) | ( n12903 & n13376 ) ;
  assign n13379 = n13378 ^ n13377 ^ n4295 ;
  assign n13380 = n13379 ^ n5969 ^ n991 ;
  assign n13381 = ~n6572 & n6714 ;
  assign n13382 = ( n2234 & n11731 ) | ( n2234 & ~n13381 ) | ( n11731 & ~n13381 ) ;
  assign n13383 = ( n343 & n8293 ) | ( n343 & ~n8344 ) | ( n8293 & ~n8344 ) ;
  assign n13384 = n13383 ^ n9535 ^ n3934 ;
  assign n13386 = n2253 & n2645 ;
  assign n13385 = n1856 & ~n7721 ;
  assign n13387 = n13386 ^ n13385 ^ n1230 ;
  assign n13401 = n11897 ^ n596 ^ n557 ;
  assign n13399 = ( n1989 & n6276 ) | ( n1989 & n7886 ) | ( n6276 & n7886 ) ;
  assign n13400 = n13399 ^ n6055 ^ 1'b0 ;
  assign n13395 = n11959 ^ n5242 ^ n5022 ;
  assign n13388 = ( n5143 & n7259 ) | ( n5143 & n10674 ) | ( n7259 & n10674 ) ;
  assign n13389 = ~n3607 & n11219 ;
  assign n13390 = n13389 ^ n6750 ^ n1026 ;
  assign n13391 = n11205 ^ n7685 ^ n2803 ;
  assign n13392 = n13391 ^ n268 ^ 1'b0 ;
  assign n13393 = n13392 ^ n8162 ^ n4922 ;
  assign n13394 = ( ~n13388 & n13390 ) | ( ~n13388 & n13393 ) | ( n13390 & n13393 ) ;
  assign n13396 = n13395 ^ n13394 ^ n8918 ;
  assign n13397 = n269 | n13396 ;
  assign n13398 = n8655 & ~n13397 ;
  assign n13402 = n13401 ^ n13400 ^ n13398 ;
  assign n13403 = ( n13384 & ~n13387 ) | ( n13384 & n13402 ) | ( ~n13387 & n13402 ) ;
  assign n13404 = ( n4058 & ~n12694 ) | ( n4058 & n13403 ) | ( ~n12694 & n13403 ) ;
  assign n13405 = n3696 ^ n2421 ^ n2185 ;
  assign n13406 = ( n1284 & n5148 ) | ( n1284 & n13405 ) | ( n5148 & n13405 ) ;
  assign n13407 = ( ~n2804 & n8388 ) | ( ~n2804 & n9569 ) | ( n8388 & n9569 ) ;
  assign n13408 = n3818 & n7818 ;
  assign n13409 = n13408 ^ n900 ^ 1'b0 ;
  assign n13410 = n5352 & n13409 ;
  assign n13411 = n13410 ^ n5615 ^ 1'b0 ;
  assign n13412 = n10734 ^ n1696 ^ 1'b0 ;
  assign n13413 = ( n3494 & n12766 ) | ( n3494 & n13412 ) | ( n12766 & n13412 ) ;
  assign n13414 = ( n13407 & n13411 ) | ( n13407 & ~n13413 ) | ( n13411 & ~n13413 ) ;
  assign n13418 = n3027 & n3565 ;
  assign n13419 = ( n3619 & n5208 ) | ( n3619 & ~n13418 ) | ( n5208 & ~n13418 ) ;
  assign n13420 = n13419 ^ n9934 ^ n7753 ;
  assign n13415 = ( n1269 & n2925 ) | ( n1269 & n12901 ) | ( n2925 & n12901 ) ;
  assign n13416 = n10521 & ~n13415 ;
  assign n13417 = ~n3498 & n13416 ;
  assign n13421 = n13420 ^ n13417 ^ 1'b0 ;
  assign n13425 = ( ~x133 & n1133 ) | ( ~x133 & n12952 ) | ( n1133 & n12952 ) ;
  assign n13422 = n3972 ^ n3667 ^ 1'b0 ;
  assign n13423 = n13422 ^ n13245 ^ n1067 ;
  assign n13424 = n13423 ^ n10743 ^ n9066 ;
  assign n13426 = n13425 ^ n13424 ^ n6494 ;
  assign n13427 = n4817 ^ n3984 ^ n2528 ;
  assign n13428 = ( n3656 & n3766 ) | ( n3656 & n13427 ) | ( n3766 & n13427 ) ;
  assign n13429 = n2006 & ~n2358 ;
  assign n13430 = n10323 ^ n2743 ^ n990 ;
  assign n13431 = n13430 ^ n4869 ^ 1'b0 ;
  assign n13432 = ~n13429 & n13431 ;
  assign n13433 = ( x176 & n905 ) | ( x176 & n13432 ) | ( n905 & n13432 ) ;
  assign n13447 = ( x105 & ~n2589 ) | ( x105 & n3384 ) | ( ~n2589 & n3384 ) ;
  assign n13448 = n10674 ^ n1949 ^ n1732 ;
  assign n13449 = ( ~n7120 & n13447 ) | ( ~n7120 & n13448 ) | ( n13447 & n13448 ) ;
  assign n13443 = ( n2231 & ~n5262 ) | ( n2231 & n7753 ) | ( ~n5262 & n7753 ) ;
  assign n13444 = ( n2249 & n2532 ) | ( n2249 & n13443 ) | ( n2532 & n13443 ) ;
  assign n13441 = ( n394 & n3528 ) | ( n394 & ~n8658 ) | ( n3528 & ~n8658 ) ;
  assign n13442 = ( n2147 & n4238 ) | ( n2147 & n13441 ) | ( n4238 & n13441 ) ;
  assign n13445 = n13444 ^ n13442 ^ n7846 ;
  assign n13446 = ( n1786 & n12162 ) | ( n1786 & ~n13445 ) | ( n12162 & ~n13445 ) ;
  assign n13450 = n13449 ^ n13446 ^ n12839 ;
  assign n13434 = ( n1069 & n6570 ) | ( n1069 & ~n10072 ) | ( n6570 & ~n10072 ) ;
  assign n13435 = ( ~n2819 & n12743 ) | ( ~n2819 & n13434 ) | ( n12743 & n13434 ) ;
  assign n13436 = n13435 ^ n4950 ^ n3737 ;
  assign n13437 = ( ~n1666 & n3040 ) | ( ~n1666 & n13436 ) | ( n3040 & n13436 ) ;
  assign n13438 = n1527 ^ n1266 ^ n897 ;
  assign n13439 = ( n6413 & ~n10906 ) | ( n6413 & n13438 ) | ( ~n10906 & n13438 ) ;
  assign n13440 = ( n7178 & ~n13437 ) | ( n7178 & n13439 ) | ( ~n13437 & n13439 ) ;
  assign n13451 = n13450 ^ n13440 ^ n13019 ;
  assign n13452 = n7592 ^ n6502 ^ n1295 ;
  assign n13453 = ( n3638 & n7169 ) | ( n3638 & n8336 ) | ( n7169 & n8336 ) ;
  assign n13454 = n3512 | n6705 ;
  assign n13455 = n13454 ^ n7748 ^ 1'b0 ;
  assign n13456 = n4077 & n13455 ;
  assign n13457 = ( n320 & n4110 ) | ( n320 & ~n13386 ) | ( n4110 & ~n13386 ) ;
  assign n13460 = ( n580 & n2168 ) | ( n580 & n8536 ) | ( n2168 & n8536 ) ;
  assign n13458 = ( ~n3165 & n4871 ) | ( ~n3165 & n8714 ) | ( n4871 & n8714 ) ;
  assign n13459 = n13458 ^ n638 ^ 1'b0 ;
  assign n13461 = n13460 ^ n13459 ^ n11657 ;
  assign n13462 = n1571 & ~n8447 ;
  assign n13463 = n13462 ^ x43 ^ 1'b0 ;
  assign n13464 = n715 | n13463 ;
  assign n13465 = n13464 ^ n6846 ^ 1'b0 ;
  assign n13466 = ~n4271 & n13465 ;
  assign n13469 = n11392 ^ n11391 ^ n5235 ;
  assign n13470 = ( ~n3460 & n7509 ) | ( ~n3460 & n13469 ) | ( n7509 & n13469 ) ;
  assign n13467 = ( n3889 & n5414 ) | ( n3889 & n7296 ) | ( n5414 & n7296 ) ;
  assign n13468 = n13467 ^ n9327 ^ n5474 ;
  assign n13471 = n13470 ^ n13468 ^ x160 ;
  assign n13472 = n9555 ^ n8841 ^ n3449 ;
  assign n13473 = ( n779 & ~n2757 ) | ( n779 & n10690 ) | ( ~n2757 & n10690 ) ;
  assign n13474 = ( n7514 & ~n13472 ) | ( n7514 & n13473 ) | ( ~n13472 & n13473 ) ;
  assign n13475 = n13474 ^ n10730 ^ n333 ;
  assign n13478 = ( n1300 & n2599 ) | ( n1300 & n3474 ) | ( n2599 & n3474 ) ;
  assign n13479 = n4227 | n13478 ;
  assign n13476 = n9643 ^ n3335 ^ n964 ;
  assign n13477 = n13476 ^ n10880 ^ n2074 ;
  assign n13480 = n13479 ^ n13477 ^ n8111 ;
  assign n13481 = n9601 ^ n5152 ^ n2758 ;
  assign n13482 = n6091 ^ n2965 ^ 1'b0 ;
  assign n13483 = n3819 | n13482 ;
  assign n13484 = ( n393 & ~n2643 ) | ( n393 & n13483 ) | ( ~n2643 & n13483 ) ;
  assign n13485 = n13484 ^ n11666 ^ n8985 ;
  assign n13486 = n6488 ^ n5106 ^ n4943 ;
  assign n13488 = ( n1634 & n8009 ) | ( n1634 & n8143 ) | ( n8009 & n8143 ) ;
  assign n13487 = ( ~n4573 & n4637 ) | ( ~n4573 & n8714 ) | ( n4637 & n8714 ) ;
  assign n13489 = n13488 ^ n13487 ^ n13097 ;
  assign n13490 = n13486 | n13489 ;
  assign n13491 = n5895 & ~n13490 ;
  assign n13492 = ( n2065 & n4051 ) | ( n2065 & ~n10564 ) | ( n4051 & ~n10564 ) ;
  assign n13493 = n13492 ^ n11095 ^ n7214 ;
  assign n13494 = n13493 ^ n1178 ^ n644 ;
  assign n13495 = n13494 ^ n6554 ^ 1'b0 ;
  assign n13496 = n13491 | n13495 ;
  assign n13497 = ( n13481 & n13485 ) | ( n13481 & n13496 ) | ( n13485 & n13496 ) ;
  assign n13498 = n4400 ^ n1491 ^ x62 ;
  assign n13499 = n13498 ^ n7247 ^ 1'b0 ;
  assign n13500 = n6057 & n13499 ;
  assign n13501 = n10331 ^ n7253 ^ x9 ;
  assign n13509 = ( ~n3677 & n3992 ) | ( ~n3677 & n5580 ) | ( n3992 & n5580 ) ;
  assign n13506 = ( n2856 & n4581 ) | ( n2856 & ~n8772 ) | ( n4581 & ~n8772 ) ;
  assign n13507 = ( ~x197 & n8246 ) | ( ~x197 & n13506 ) | ( n8246 & n13506 ) ;
  assign n13505 = ( ~n2577 & n3927 ) | ( ~n2577 & n11186 ) | ( n3927 & n11186 ) ;
  assign n13508 = n13507 ^ n13505 ^ n5148 ;
  assign n13510 = n13509 ^ n13508 ^ 1'b0 ;
  assign n13511 = n1621 & ~n13510 ;
  assign n13512 = ( n2860 & n10257 ) | ( n2860 & n13511 ) | ( n10257 & n13511 ) ;
  assign n13502 = n10438 ^ n756 ^ 1'b0 ;
  assign n13503 = n8454 | n13502 ;
  assign n13504 = n13503 ^ n7668 ^ n5655 ;
  assign n13513 = n13512 ^ n13504 ^ 1'b0 ;
  assign n13514 = ( n13500 & ~n13501 ) | ( n13500 & n13513 ) | ( ~n13501 & n13513 ) ;
  assign n13515 = ( n1425 & n3727 ) | ( n1425 & n7071 ) | ( n3727 & n7071 ) ;
  assign n13516 = n13515 ^ n3449 ^ 1'b0 ;
  assign n13517 = n5761 | n13516 ;
  assign n13518 = n13517 ^ n11865 ^ n11610 ;
  assign n13519 = n9613 ^ n7425 ^ 1'b0 ;
  assign n13520 = ( n2392 & n7347 ) | ( n2392 & n13519 ) | ( n7347 & n13519 ) ;
  assign n13521 = ( n4156 & ~n5194 ) | ( n4156 & n10407 ) | ( ~n5194 & n10407 ) ;
  assign n13522 = ( n1613 & n6019 ) | ( n1613 & ~n13521 ) | ( n6019 & ~n13521 ) ;
  assign n13523 = n13522 ^ n8356 ^ n7642 ;
  assign n13524 = ( n657 & n13520 ) | ( n657 & ~n13523 ) | ( n13520 & ~n13523 ) ;
  assign n13539 = n2479 ^ n1822 ^ n430 ;
  assign n13528 = ( x113 & n1896 ) | ( x113 & ~n10118 ) | ( n1896 & ~n10118 ) ;
  assign n13525 = n7140 & n7319 ;
  assign n13526 = n13525 ^ n4057 ^ 1'b0 ;
  assign n13527 = n13526 ^ n5198 ^ n5196 ;
  assign n13529 = n13528 ^ n13527 ^ n5728 ;
  assign n13530 = n13529 ^ n13103 ^ n6263 ;
  assign n13531 = ( n885 & ~n4142 ) | ( n885 & n13530 ) | ( ~n4142 & n13530 ) ;
  assign n13534 = ~n2085 & n2619 ;
  assign n13535 = ( x135 & n1284 ) | ( x135 & ~n3788 ) | ( n1284 & ~n3788 ) ;
  assign n13536 = ( ~n533 & n13534 ) | ( ~n533 & n13535 ) | ( n13534 & n13535 ) ;
  assign n13532 = ( ~n1518 & n6324 ) | ( ~n1518 & n9232 ) | ( n6324 & n9232 ) ;
  assign n13533 = ( ~n851 & n6747 ) | ( ~n851 & n13532 ) | ( n6747 & n13532 ) ;
  assign n13537 = n13536 ^ n13533 ^ n4581 ;
  assign n13538 = ( n11178 & n13531 ) | ( n11178 & n13537 ) | ( n13531 & n13537 ) ;
  assign n13540 = n13539 ^ n13538 ^ n4525 ;
  assign n13541 = n8962 ^ n5510 ^ n3836 ;
  assign n13542 = ( n2878 & n6689 ) | ( n2878 & ~n7139 ) | ( n6689 & ~n7139 ) ;
  assign n13543 = ( n9707 & n13541 ) | ( n9707 & ~n13542 ) | ( n13541 & ~n13542 ) ;
  assign n13547 = ( n569 & n3066 ) | ( n569 & ~n5955 ) | ( n3066 & ~n5955 ) ;
  assign n13545 = ~n682 & n11818 ;
  assign n13544 = ~n850 & n10372 ;
  assign n13546 = n13545 ^ n13544 ^ 1'b0 ;
  assign n13548 = n13547 ^ n13546 ^ n2917 ;
  assign n13550 = ( ~n1327 & n2293 ) | ( ~n1327 & n9308 ) | ( n2293 & n9308 ) ;
  assign n13551 = ( ~n4366 & n11562 ) | ( ~n4366 & n13550 ) | ( n11562 & n13550 ) ;
  assign n13549 = ( n7303 & n9581 ) | ( n7303 & n12544 ) | ( n9581 & n12544 ) ;
  assign n13552 = n13551 ^ n13549 ^ n12550 ;
  assign n13553 = ( n2139 & ~n3904 ) | ( n2139 & n10181 ) | ( ~n3904 & n10181 ) ;
  assign n13554 = n12028 ^ n3638 ^ n2197 ;
  assign n13555 = ( n10422 & n13553 ) | ( n10422 & n13554 ) | ( n13553 & n13554 ) ;
  assign n13556 = ( n8997 & ~n9627 ) | ( n8997 & n11700 ) | ( ~n9627 & n11700 ) ;
  assign n13558 = n6915 ^ n3903 ^ 1'b0 ;
  assign n13559 = n5218 & ~n13558 ;
  assign n13560 = n13559 ^ n7029 ^ n2006 ;
  assign n13557 = n6983 ^ n4674 ^ n3658 ;
  assign n13561 = n13560 ^ n13557 ^ n12631 ;
  assign n13562 = n3451 ^ n636 ^ 1'b0 ;
  assign n13563 = ~n326 & n13562 ;
  assign n13564 = n13563 ^ n5393 ^ n1842 ;
  assign n13565 = n13564 ^ n6214 ^ n4302 ;
  assign n13566 = n1539 & ~n3865 ;
  assign n13567 = ( n1756 & ~n12582 ) | ( n1756 & n13566 ) | ( ~n12582 & n13566 ) ;
  assign n13568 = n13567 ^ n7449 ^ n7112 ;
  assign n13569 = n857 & n13568 ;
  assign n13570 = n1691 & n13569 ;
  assign n13571 = ( n7844 & n13565 ) | ( n7844 & ~n13570 ) | ( n13565 & ~n13570 ) ;
  assign n13589 = n683 & n3402 ;
  assign n13573 = ~n5891 & n11350 ;
  assign n13574 = n13573 ^ n3645 ^ 1'b0 ;
  assign n13575 = n6356 ^ n3443 ^ n2535 ;
  assign n13576 = x73 & n9265 ;
  assign n13577 = n13576 ^ n3649 ^ 1'b0 ;
  assign n13578 = ( x192 & ~n1527 ) | ( x192 & n3133 ) | ( ~n1527 & n3133 ) ;
  assign n13579 = n13578 ^ n11596 ^ n2679 ;
  assign n13580 = n3207 | n13579 ;
  assign n13581 = n13577 | n13580 ;
  assign n13582 = ( n470 & n3708 ) | ( n470 & ~n5490 ) | ( n3708 & ~n5490 ) ;
  assign n13583 = n13582 ^ n1088 ^ n464 ;
  assign n13584 = n9072 | n10657 ;
  assign n13585 = n13584 ^ n2410 ^ n957 ;
  assign n13586 = ( n8760 & ~n13583 ) | ( n8760 & n13585 ) | ( ~n13583 & n13585 ) ;
  assign n13587 = ( n949 & ~n13581 ) | ( n949 & n13586 ) | ( ~n13581 & n13586 ) ;
  assign n13588 = ( n13574 & ~n13575 ) | ( n13574 & n13587 ) | ( ~n13575 & n13587 ) ;
  assign n13572 = ( n4565 & ~n6713 ) | ( n4565 & n9205 ) | ( ~n6713 & n9205 ) ;
  assign n13590 = n13589 ^ n13588 ^ n13572 ;
  assign n13591 = ( n2853 & n6723 ) | ( n2853 & ~n13590 ) | ( n6723 & ~n13590 ) ;
  assign n13592 = ( n2028 & n8060 ) | ( n2028 & n12308 ) | ( n8060 & n12308 ) ;
  assign n13593 = n11500 ^ n4102 ^ n3526 ;
  assign n13594 = ( ~n3455 & n13592 ) | ( ~n3455 & n13593 ) | ( n13592 & n13593 ) ;
  assign n13595 = n9946 ^ n3449 ^ n1396 ;
  assign n13596 = n13595 ^ n9463 ^ n4451 ;
  assign n13597 = ( n8553 & ~n10848 ) | ( n8553 & n13596 ) | ( ~n10848 & n13596 ) ;
  assign n13598 = n13597 ^ n6080 ^ n2513 ;
  assign n13602 = n12519 ^ n3891 ^ n2691 ;
  assign n13603 = ( n1563 & n2897 ) | ( n1563 & ~n13602 ) | ( n2897 & ~n13602 ) ;
  assign n13599 = n13015 ^ n3979 ^ n2498 ;
  assign n13600 = n6122 & ~n13599 ;
  assign n13601 = ( n643 & n6834 ) | ( n643 & ~n13600 ) | ( n6834 & ~n13600 ) ;
  assign n13604 = n13603 ^ n13601 ^ n1701 ;
  assign n13606 = ( ~n333 & n415 ) | ( ~n333 & n782 ) | ( n415 & n782 ) ;
  assign n13607 = n13606 ^ n9860 ^ n6475 ;
  assign n13605 = n12267 ^ n8811 ^ n3716 ;
  assign n13608 = n13607 ^ n13605 ^ 1'b0 ;
  assign n13609 = n3945 | n13608 ;
  assign n13610 = ( n744 & n12950 ) | ( n744 & ~n13609 ) | ( n12950 & ~n13609 ) ;
  assign n13611 = n13610 ^ n12646 ^ n2623 ;
  assign n13612 = ( n1993 & n5138 ) | ( n1993 & n10519 ) | ( n5138 & n10519 ) ;
  assign n13613 = ( n5335 & n8317 ) | ( n5335 & ~n13612 ) | ( n8317 & ~n13612 ) ;
  assign n13614 = n5969 ^ n5807 ^ n3541 ;
  assign n13616 = n2295 | n8170 ;
  assign n13617 = ( ~n939 & n5422 ) | ( ~n939 & n13616 ) | ( n5422 & n13616 ) ;
  assign n13618 = n13617 ^ n4621 ^ 1'b0 ;
  assign n13619 = x25 & ~n13618 ;
  assign n13615 = n7772 ^ n4201 ^ n1485 ;
  assign n13620 = n13619 ^ n13615 ^ 1'b0 ;
  assign n13621 = n13614 & ~n13620 ;
  assign n13622 = n9338 ^ n3820 ^ 1'b0 ;
  assign n13623 = ( n5244 & ~n9133 ) | ( n5244 & n13622 ) | ( ~n9133 & n13622 ) ;
  assign n13624 = n13623 ^ n13551 ^ n1283 ;
  assign n13625 = n11045 ^ n6259 ^ n2706 ;
  assign n13626 = n10997 ^ n1116 ^ 1'b0 ;
  assign n13627 = ~n4776 & n13626 ;
  assign n13628 = n13627 ^ n6038 ^ n5732 ;
  assign n13629 = ( n569 & n13625 ) | ( n569 & n13628 ) | ( n13625 & n13628 ) ;
  assign n13630 = n11710 ^ n8697 ^ n1299 ;
  assign n13631 = n9070 ^ n7387 ^ n1578 ;
  assign n13635 = n854 | n8521 ;
  assign n13634 = n2786 ^ n2033 ^ n1076 ;
  assign n13636 = n13635 ^ n13634 ^ n7506 ;
  assign n13637 = n6591 & ~n13636 ;
  assign n13632 = ( n747 & n791 ) | ( n747 & ~n1022 ) | ( n791 & ~n1022 ) ;
  assign n13633 = ~n10357 & n13632 ;
  assign n13638 = n13637 ^ n13633 ^ 1'b0 ;
  assign n13639 = ( ~n904 & n8986 ) | ( ~n904 & n12015 ) | ( n8986 & n12015 ) ;
  assign n13640 = n13639 ^ n7027 ^ n933 ;
  assign n13641 = ( ~n13631 & n13638 ) | ( ~n13631 & n13640 ) | ( n13638 & n13640 ) ;
  assign n13642 = ( n11714 & n13630 ) | ( n11714 & n13641 ) | ( n13630 & n13641 ) ;
  assign n13643 = ( n2719 & ~n6536 ) | ( n2719 & n10740 ) | ( ~n6536 & n10740 ) ;
  assign n13644 = ( n2146 & ~n3325 ) | ( n2146 & n5289 ) | ( ~n3325 & n5289 ) ;
  assign n13645 = n13644 ^ n5519 ^ n4430 ;
  assign n13646 = n5755 | n13645 ;
  assign n13647 = n10167 & ~n13646 ;
  assign n13648 = n13647 ^ n7430 ^ n4440 ;
  assign n13649 = n13648 ^ n10222 ^ n7372 ;
  assign n13650 = ( n12530 & ~n13643 ) | ( n12530 & n13649 ) | ( ~n13643 & n13649 ) ;
  assign n13651 = ( n1102 & n1315 ) | ( n1102 & n4819 ) | ( n1315 & n4819 ) ;
  assign n13652 = n13651 ^ n6871 ^ n1056 ;
  assign n13653 = ( n2426 & n7253 ) | ( n2426 & ~n11993 ) | ( n7253 & ~n11993 ) ;
  assign n13654 = n8053 ^ n4275 ^ n386 ;
  assign n13655 = ( n4578 & ~n13124 ) | ( n4578 & n13654 ) | ( ~n13124 & n13654 ) ;
  assign n13656 = n13655 ^ n10136 ^ n5091 ;
  assign n13657 = n6660 ^ n6427 ^ 1'b0 ;
  assign n13658 = n9557 ^ n6809 ^ 1'b0 ;
  assign n13659 = n13657 & ~n13658 ;
  assign n13660 = ( n1153 & ~n6313 ) | ( n1153 & n9888 ) | ( ~n6313 & n9888 ) ;
  assign n13662 = n2399 ^ x244 ^ x200 ;
  assign n13663 = n12505 & n13662 ;
  assign n13661 = ( ~n953 & n3257 ) | ( ~n953 & n4178 ) | ( n3257 & n4178 ) ;
  assign n13664 = n13663 ^ n13661 ^ n4501 ;
  assign n13665 = n11497 ^ n9381 ^ n3764 ;
  assign n13666 = ( n13660 & n13664 ) | ( n13660 & ~n13665 ) | ( n13664 & ~n13665 ) ;
  assign n13667 = ( n11612 & ~n13659 ) | ( n11612 & n13666 ) | ( ~n13659 & n13666 ) ;
  assign n13668 = x86 & n996 ;
  assign n13669 = ( n4480 & n4533 ) | ( n4480 & n9368 ) | ( n4533 & n9368 ) ;
  assign n13670 = ( ~n2937 & n5576 ) | ( ~n2937 & n13669 ) | ( n5576 & n13669 ) ;
  assign n13671 = n13670 ^ n13118 ^ n3081 ;
  assign n13672 = n13671 ^ n10318 ^ n265 ;
  assign n13673 = n13672 ^ n8597 ^ n5196 ;
  assign n13674 = ( ~n7785 & n13668 ) | ( ~n7785 & n13673 ) | ( n13668 & n13673 ) ;
  assign n13675 = n1864 | n8632 ;
  assign n13676 = n13675 ^ n2658 ^ 1'b0 ;
  assign n13677 = n9389 ^ n2469 ^ 1'b0 ;
  assign n13678 = n13677 ^ n1165 ^ x24 ;
  assign n13684 = n7509 ^ n5094 ^ 1'b0 ;
  assign n13685 = n12662 ^ x93 ^ 1'b0 ;
  assign n13686 = n13684 & ~n13685 ;
  assign n13683 = ( n7809 & n8513 ) | ( n7809 & ~n13082 ) | ( n8513 & ~n13082 ) ;
  assign n13681 = n8434 ^ n2589 ^ 1'b0 ;
  assign n13679 = n7044 ^ n3895 ^ n2564 ;
  assign n13680 = n13679 ^ n13212 ^ n11081 ;
  assign n13682 = n13681 ^ n13680 ^ x244 ;
  assign n13687 = n13686 ^ n13683 ^ n13682 ;
  assign n13688 = ( ~n5008 & n13678 ) | ( ~n5008 & n13687 ) | ( n13678 & n13687 ) ;
  assign n13689 = ( n1668 & n3320 ) | ( n1668 & n12621 ) | ( n3320 & n12621 ) ;
  assign n13690 = n13689 ^ n13385 ^ n1502 ;
  assign n13691 = n10994 ^ n2551 ^ 1'b0 ;
  assign n13692 = ~n10902 & n13691 ;
  assign n13693 = n10558 ^ n646 ^ 1'b0 ;
  assign n13694 = n13693 ^ n10065 ^ n688 ;
  assign n13695 = n13692 & ~n13694 ;
  assign n13696 = x130 & ~n12493 ;
  assign n13697 = ( n2252 & ~n10993 ) | ( n2252 & n13696 ) | ( ~n10993 & n13696 ) ;
  assign n13698 = n13697 ^ n12333 ^ 1'b0 ;
  assign n13699 = n13695 & ~n13698 ;
  assign n13700 = n1992 | n6638 ;
  assign n13701 = ( ~n6795 & n8303 ) | ( ~n6795 & n13700 ) | ( n8303 & n13700 ) ;
  assign n13702 = ( n4187 & ~n7770 ) | ( n4187 & n9605 ) | ( ~n7770 & n9605 ) ;
  assign n13703 = ( ~n5166 & n9481 ) | ( ~n5166 & n11016 ) | ( n9481 & n11016 ) ;
  assign n13704 = n13703 ^ n5399 ^ n3900 ;
  assign n13705 = x177 ^ x44 ^ x40 ;
  assign n13706 = n7602 ^ n782 ^ n293 ;
  assign n13707 = n13706 ^ n1836 ^ n442 ;
  assign n13708 = n10547 ^ n4727 ^ n3032 ;
  assign n13709 = ( n5219 & n13707 ) | ( n5219 & ~n13708 ) | ( n13707 & ~n13708 ) ;
  assign n13710 = ( n2722 & ~n12235 ) | ( n2722 & n13709 ) | ( ~n12235 & n13709 ) ;
  assign n13711 = ( n13537 & n13705 ) | ( n13537 & ~n13710 ) | ( n13705 & ~n13710 ) ;
  assign n13712 = ( n1650 & ~n13704 ) | ( n1650 & n13711 ) | ( ~n13704 & n13711 ) ;
  assign n13719 = n9379 ^ n5578 ^ 1'b0 ;
  assign n13717 = n9059 ^ n1996 ^ n283 ;
  assign n13713 = n4382 ^ n4238 ^ n2422 ;
  assign n13714 = ( ~n497 & n5480 ) | ( ~n497 & n13713 ) | ( n5480 & n13713 ) ;
  assign n13715 = n13714 ^ n7218 ^ x247 ;
  assign n13716 = n4662 & n13715 ;
  assign n13718 = n13717 ^ n13716 ^ n6798 ;
  assign n13720 = n13719 ^ n13718 ^ n2701 ;
  assign n13721 = ( ~n4682 & n5949 ) | ( ~n4682 & n13720 ) | ( n5949 & n13720 ) ;
  assign n13722 = n5107 ^ n2296 ^ 1'b0 ;
  assign n13723 = ( n5885 & ~n10822 ) | ( n5885 & n13722 ) | ( ~n10822 & n13722 ) ;
  assign n13724 = n3670 ^ n1356 ^ 1'b0 ;
  assign n13725 = ( n3032 & n12862 ) | ( n3032 & ~n13724 ) | ( n12862 & ~n13724 ) ;
  assign n13726 = ( n5299 & n9867 ) | ( n5299 & ~n13725 ) | ( n9867 & ~n13725 ) ;
  assign n13729 = n13670 ^ n1892 ^ 1'b0 ;
  assign n13727 = n8271 ^ n6917 ^ n1208 ;
  assign n13728 = ( n1368 & ~n11103 ) | ( n1368 & n13727 ) | ( ~n11103 & n13727 ) ;
  assign n13730 = n13729 ^ n13728 ^ n2499 ;
  assign n13731 = ( n1843 & n2981 ) | ( n1843 & n9269 ) | ( n2981 & n9269 ) ;
  assign n13732 = ( n13726 & n13730 ) | ( n13726 & ~n13731 ) | ( n13730 & ~n13731 ) ;
  assign n13733 = ~n538 & n3652 ;
  assign n13734 = n13733 ^ n10720 ^ n4201 ;
  assign n13736 = n4301 ^ n2611 ^ n580 ;
  assign n13737 = n13736 ^ n10035 ^ n2600 ;
  assign n13735 = n8592 ^ n6325 ^ n2058 ;
  assign n13738 = n13737 ^ n13735 ^ n6586 ;
  assign n13739 = n13738 ^ n3740 ^ n2381 ;
  assign n13751 = ( n3761 & n4018 ) | ( n3761 & ~n4189 ) | ( n4018 & ~n4189 ) ;
  assign n13749 = ( ~n481 & n4993 ) | ( ~n481 & n11016 ) | ( n4993 & n11016 ) ;
  assign n13750 = n13749 ^ n12056 ^ n4216 ;
  assign n13742 = n3658 ^ n1755 ^ n347 ;
  assign n13741 = n7540 ^ n3403 ^ n1448 ;
  assign n13740 = n5149 ^ n4538 ^ n1931 ;
  assign n13743 = n13742 ^ n13741 ^ n13740 ;
  assign n13744 = ( n2824 & ~n6384 ) | ( n2824 & n7725 ) | ( ~n6384 & n7725 ) ;
  assign n13745 = n13744 ^ n4370 ^ 1'b0 ;
  assign n13746 = n3082 | n13745 ;
  assign n13747 = n13743 | n13746 ;
  assign n13748 = n13747 ^ n1775 ^ 1'b0 ;
  assign n13752 = n13751 ^ n13750 ^ n13748 ;
  assign n13753 = n6832 & n7244 ;
  assign n13754 = n9218 ^ n5187 ^ 1'b0 ;
  assign n13755 = ~n9682 & n13754 ;
  assign n13756 = ( n2807 & ~n13753 ) | ( n2807 & n13755 ) | ( ~n13753 & n13755 ) ;
  assign n13757 = n11364 ^ n10436 ^ n2601 ;
  assign n13758 = ( n277 & n10285 ) | ( n277 & n13757 ) | ( n10285 & n13757 ) ;
  assign n13759 = ( n2870 & n6208 ) | ( n2870 & n9513 ) | ( n6208 & n9513 ) ;
  assign n13764 = ( n3788 & n5890 ) | ( n3788 & n7219 ) | ( n5890 & n7219 ) ;
  assign n13765 = n13764 ^ n4223 ^ n1101 ;
  assign n13763 = ( n2104 & ~n5719 ) | ( n2104 & n6147 ) | ( ~n5719 & n6147 ) ;
  assign n13760 = ( n1257 & n3954 ) | ( n1257 & n11781 ) | ( n3954 & n11781 ) ;
  assign n13761 = n13760 ^ n8464 ^ n4955 ;
  assign n13762 = ( ~n1270 & n11720 ) | ( ~n1270 & n13761 ) | ( n11720 & n13761 ) ;
  assign n13766 = n13765 ^ n13763 ^ n13762 ;
  assign n13767 = ( ~n331 & n9783 ) | ( ~n331 & n13766 ) | ( n9783 & n13766 ) ;
  assign n13768 = n8454 ^ n6804 ^ n6095 ;
  assign n13770 = ( ~x11 & n1595 ) | ( ~x11 & n4793 ) | ( n1595 & n4793 ) ;
  assign n13769 = ( n1160 & n4335 ) | ( n1160 & n5247 ) | ( n4335 & n5247 ) ;
  assign n13771 = n13770 ^ n13769 ^ n9375 ;
  assign n13772 = ( n3109 & n8734 ) | ( n3109 & n13771 ) | ( n8734 & n13771 ) ;
  assign n13773 = ( ~n13601 & n13768 ) | ( ~n13601 & n13772 ) | ( n13768 & n13772 ) ;
  assign n13774 = n13773 ^ n13592 ^ n1888 ;
  assign n13780 = n2152 ^ n1696 ^ n1195 ;
  assign n13777 = n9266 ^ n4102 ^ n3790 ;
  assign n13778 = ~n7054 & n13777 ;
  assign n13779 = n13778 ^ n9163 ^ 1'b0 ;
  assign n13775 = n9346 ^ n7455 ^ n2222 ;
  assign n13776 = n13775 ^ n8353 ^ n3396 ;
  assign n13781 = n13780 ^ n13779 ^ n13776 ;
  assign n13782 = n6360 ^ n3255 ^ n556 ;
  assign n13783 = n5848 ^ n3827 ^ n2842 ;
  assign n13784 = n13783 ^ n856 ^ 1'b0 ;
  assign n13785 = ~n1503 & n13784 ;
  assign n13786 = ( n1303 & n13782 ) | ( n1303 & n13785 ) | ( n13782 & n13785 ) ;
  assign n13787 = n4686 ^ n3451 ^ n1335 ;
  assign n13788 = ( x179 & ~x237 ) | ( x179 & n2510 ) | ( ~x237 & n2510 ) ;
  assign n13789 = ( n2960 & ~n4704 ) | ( n2960 & n13788 ) | ( ~n4704 & n13788 ) ;
  assign n13790 = n13789 ^ n6064 ^ n702 ;
  assign n13791 = n13790 ^ n11878 ^ n6604 ;
  assign n13792 = n3133 ^ n3069 ^ n2717 ;
  assign n13793 = n3076 ^ n2615 ^ n502 ;
  assign n13794 = ( ~n317 & n887 ) | ( ~n317 & n2679 ) | ( n887 & n2679 ) ;
  assign n13795 = n13794 ^ n6875 ^ n350 ;
  assign n13796 = ~n5106 & n13795 ;
  assign n13797 = n13796 ^ n4356 ^ 1'b0 ;
  assign n13798 = ( n13792 & ~n13793 ) | ( n13792 & n13797 ) | ( ~n13793 & n13797 ) ;
  assign n13799 = n13798 ^ n12427 ^ n3278 ;
  assign n13800 = n13799 ^ n12516 ^ 1'b0 ;
  assign n13801 = n13791 | n13800 ;
  assign n13821 = ~n2271 & n4233 ;
  assign n13822 = ~n1461 & n13821 ;
  assign n13823 = n13822 ^ n2386 ^ 1'b0 ;
  assign n13824 = n5841 & ~n13823 ;
  assign n13820 = ( n1850 & n5796 ) | ( n1850 & n6400 ) | ( n5796 & n6400 ) ;
  assign n13809 = ( n581 & n812 ) | ( n581 & ~n3873 ) | ( n812 & ~n3873 ) ;
  assign n13810 = n12781 ^ n3581 ^ n533 ;
  assign n13811 = n5308 | n13810 ;
  assign n13812 = n6228 | n13811 ;
  assign n13813 = n8065 ^ n4468 ^ n751 ;
  assign n13814 = n13813 ^ n1405 ^ x156 ;
  assign n13815 = n13814 ^ n11529 ^ n4321 ;
  assign n13816 = n13815 ^ n5087 ^ x150 ;
  assign n13817 = n13816 ^ n8572 ^ n4969 ;
  assign n13818 = ( ~n13809 & n13812 ) | ( ~n13809 & n13817 ) | ( n13812 & n13817 ) ;
  assign n13807 = n4298 | n10891 ;
  assign n13808 = ( ~n7094 & n10995 ) | ( ~n7094 & n13807 ) | ( n10995 & n13807 ) ;
  assign n13819 = n13818 ^ n13808 ^ n4342 ;
  assign n13825 = n13824 ^ n13820 ^ n13819 ;
  assign n13826 = n7552 | n13825 ;
  assign n13827 = n8712 & ~n13826 ;
  assign n13806 = n499 | n5685 ;
  assign n13803 = n10009 ^ n3184 ^ 1'b0 ;
  assign n13804 = ( x243 & n1204 ) | ( x243 & n13803 ) | ( n1204 & n13803 ) ;
  assign n13802 = n9627 ^ n7419 ^ n6307 ;
  assign n13805 = n13804 ^ n13802 ^ n11292 ;
  assign n13828 = n13827 ^ n13806 ^ n13805 ;
  assign n13829 = n12828 ^ n7071 ^ n2629 ;
  assign n13830 = ~n11567 & n13829 ;
  assign n13831 = n13830 ^ n9153 ^ n8818 ;
  assign n13832 = n1228 & n13052 ;
  assign n13833 = n13832 ^ n7335 ^ 1'b0 ;
  assign n13834 = ( ~n1585 & n2994 ) | ( ~n1585 & n13833 ) | ( n2994 & n13833 ) ;
  assign n13835 = n13834 ^ n11342 ^ n5248 ;
  assign n13836 = ( n11748 & n13831 ) | ( n11748 & n13835 ) | ( n13831 & n13835 ) ;
  assign n13854 = n1612 & ~n6260 ;
  assign n13855 = n13541 & n13854 ;
  assign n13856 = n5047 ^ n4445 ^ n3417 ;
  assign n13857 = ( n11943 & n13855 ) | ( n11943 & ~n13856 ) | ( n13855 & ~n13856 ) ;
  assign n13837 = ( n3101 & n5704 ) | ( n3101 & n7565 ) | ( n5704 & n7565 ) ;
  assign n13849 = n7441 ^ n4777 ^ 1'b0 ;
  assign n13850 = n13763 | n13849 ;
  assign n13844 = ( n3229 & n7259 ) | ( n3229 & n7964 ) | ( n7259 & n7964 ) ;
  assign n13845 = n4128 | n11438 ;
  assign n13846 = n11566 ^ n6950 ^ n1528 ;
  assign n13847 = ( n9182 & n13845 ) | ( n9182 & n13846 ) | ( n13845 & n13846 ) ;
  assign n13848 = ( n10011 & n13844 ) | ( n10011 & n13847 ) | ( n13844 & n13847 ) ;
  assign n13838 = n3353 ^ n2570 ^ x26 ;
  assign n13840 = ( n1957 & n1961 ) | ( n1957 & ~n5366 ) | ( n1961 & ~n5366 ) ;
  assign n13839 = ( n2063 & n4252 ) | ( n2063 & ~n7289 ) | ( n4252 & ~n7289 ) ;
  assign n13841 = n13840 ^ n13839 ^ n3391 ;
  assign n13842 = n13841 ^ n13245 ^ n4570 ;
  assign n13843 = ( ~n883 & n13838 ) | ( ~n883 & n13842 ) | ( n13838 & n13842 ) ;
  assign n13851 = n13850 ^ n13848 ^ n13843 ;
  assign n13852 = ( n12388 & ~n13837 ) | ( n12388 & n13851 ) | ( ~n13837 & n13851 ) ;
  assign n13853 = n13852 ^ n8381 ^ n5167 ;
  assign n13858 = n13857 ^ n13853 ^ n6120 ;
  assign n13870 = ( n2690 & n4506 ) | ( n2690 & ~n6316 ) | ( n4506 & ~n6316 ) ;
  assign n13871 = ( n1278 & n7248 ) | ( n1278 & ~n12736 ) | ( n7248 & ~n12736 ) ;
  assign n13872 = ( n8276 & n13870 ) | ( n8276 & ~n13871 ) | ( n13870 & ~n13871 ) ;
  assign n13860 = n521 & n12342 ;
  assign n13861 = n13860 ^ n7583 ^ 1'b0 ;
  assign n13859 = ( ~n9334 & n9622 ) | ( ~n9334 & n9843 ) | ( n9622 & n9843 ) ;
  assign n13862 = n13861 ^ n13859 ^ n3236 ;
  assign n13863 = ( n434 & n3184 ) | ( n434 & n4580 ) | ( n3184 & n4580 ) ;
  assign n13864 = ( ~n10948 & n12041 ) | ( ~n10948 & n13863 ) | ( n12041 & n13863 ) ;
  assign n13865 = n12257 ^ n8790 ^ n5096 ;
  assign n13866 = n8673 | n13865 ;
  assign n13867 = n13866 ^ n9213 ^ 1'b0 ;
  assign n13868 = ( n13862 & n13864 ) | ( n13862 & ~n13867 ) | ( n13864 & ~n13867 ) ;
  assign n13869 = ( n5880 & n7344 ) | ( n5880 & n13868 ) | ( n7344 & n13868 ) ;
  assign n13873 = n13872 ^ n13869 ^ n12762 ;
  assign n13874 = n3733 ^ n1781 ^ n1408 ;
  assign n13875 = n5191 & n13874 ;
  assign n13876 = n5621 & n13875 ;
  assign n13877 = n5411 | n13876 ;
  assign n13878 = n13877 ^ n2842 ^ 1'b0 ;
  assign n13879 = ( ~n8546 & n12746 ) | ( ~n8546 & n13878 ) | ( n12746 & n13878 ) ;
  assign n13880 = n12467 ^ n4476 ^ 1'b0 ;
  assign n13881 = ~n3292 & n13880 ;
  assign n13882 = ( ~n1556 & n4156 ) | ( ~n1556 & n6685 ) | ( n4156 & n6685 ) ;
  assign n13883 = n11557 ^ n5240 ^ n1356 ;
  assign n13884 = n6621 | n9193 ;
  assign n13885 = ( n2907 & n2945 ) | ( n2907 & ~n4063 ) | ( n2945 & ~n4063 ) ;
  assign n13886 = ( ~n13883 & n13884 ) | ( ~n13883 & n13885 ) | ( n13884 & n13885 ) ;
  assign n13887 = n13882 & ~n13886 ;
  assign n13888 = n3667 ^ n2999 ^ 1'b0 ;
  assign n13889 = n13888 ^ n8043 ^ 1'b0 ;
  assign n13890 = n13887 & ~n13889 ;
  assign n13891 = ( n6850 & ~n13881 ) | ( n6850 & n13890 ) | ( ~n13881 & n13890 ) ;
  assign n13892 = ( n1839 & n8364 ) | ( n1839 & ~n11562 ) | ( n8364 & ~n11562 ) ;
  assign n13893 = n13892 ^ n3956 ^ n2850 ;
  assign n13894 = ( n1668 & n3921 ) | ( n1668 & n5301 ) | ( n3921 & n5301 ) ;
  assign n13895 = ( n7653 & ~n11810 ) | ( n7653 & n13894 ) | ( ~n11810 & n13894 ) ;
  assign n13897 = n6251 ^ n4619 ^ n3710 ;
  assign n13896 = ( n4885 & ~n8593 ) | ( n4885 & n11858 ) | ( ~n8593 & n11858 ) ;
  assign n13898 = n13897 ^ n13896 ^ n4015 ;
  assign n13899 = n13898 ^ n7164 ^ 1'b0 ;
  assign n13900 = ( n13893 & n13895 ) | ( n13893 & ~n13899 ) | ( n13895 & ~n13899 ) ;
  assign n13901 = n11968 ^ n4319 ^ n1804 ;
  assign n13902 = n2778 ^ n997 ^ n619 ;
  assign n13903 = ( n974 & n1243 ) | ( n974 & ~n5490 ) | ( n1243 & ~n5490 ) ;
  assign n13904 = ( n1899 & n8170 ) | ( n1899 & ~n13903 ) | ( n8170 & ~n13903 ) ;
  assign n13905 = n13904 ^ n11357 ^ n4097 ;
  assign n13906 = n9262 & ~n13905 ;
  assign n13907 = ( ~n1835 & n13902 ) | ( ~n1835 & n13906 ) | ( n13902 & n13906 ) ;
  assign n13908 = ( n5908 & n6283 ) | ( n5908 & ~n13907 ) | ( n6283 & ~n13907 ) ;
  assign n13909 = n13908 ^ n12714 ^ n6563 ;
  assign n13910 = ( n13900 & n13901 ) | ( n13900 & n13909 ) | ( n13901 & n13909 ) ;
  assign n13911 = n11437 ^ n7903 ^ n7052 ;
  assign n13913 = n12162 ^ n7907 ^ n3917 ;
  assign n13912 = n5282 ^ n5047 ^ n2738 ;
  assign n13914 = n13913 ^ n13912 ^ n6643 ;
  assign n13915 = n13914 ^ n12082 ^ n884 ;
  assign n13916 = n6665 ^ n4988 ^ n4331 ;
  assign n13917 = ( n8768 & n12639 ) | ( n8768 & ~n13916 ) | ( n12639 & ~n13916 ) ;
  assign n13918 = n8523 ^ n5382 ^ n5269 ;
  assign n13919 = ( x113 & ~x199 ) | ( x113 & n13918 ) | ( ~x199 & n13918 ) ;
  assign n13920 = n6239 & ~n13919 ;
  assign n13921 = n13920 ^ n3565 ^ 1'b0 ;
  assign n13922 = n13921 ^ n8458 ^ n6905 ;
  assign n13923 = n10155 ^ n6661 ^ 1'b0 ;
  assign n13924 = ~n13259 & n13923 ;
  assign n13925 = n921 | n4335 ;
  assign n13926 = n4538 | n13925 ;
  assign n13927 = n13926 ^ n3509 ^ n3250 ;
  assign n13928 = n13927 ^ n4523 ^ 1'b0 ;
  assign n13929 = n6425 & n6691 ;
  assign n13930 = n12156 & n12917 ;
  assign n13931 = n8060 & n13930 ;
  assign n13936 = ( ~n739 & n4191 ) | ( ~n739 & n10527 ) | ( n4191 & n10527 ) ;
  assign n13937 = ( ~n6275 & n7780 ) | ( ~n6275 & n13936 ) | ( n7780 & n13936 ) ;
  assign n13935 = n9042 ^ n5581 ^ n4650 ;
  assign n13932 = n6326 ^ n3643 ^ n2980 ;
  assign n13933 = n13932 ^ n13449 ^ n9723 ;
  assign n13934 = n13933 ^ n3852 ^ n899 ;
  assign n13938 = n13937 ^ n13935 ^ n13934 ;
  assign n13939 = ( ~n450 & n1159 ) | ( ~n450 & n10603 ) | ( n1159 & n10603 ) ;
  assign n13940 = n13939 ^ n2493 ^ 1'b0 ;
  assign n13941 = ( n4950 & n8129 ) | ( n4950 & ~n13940 ) | ( n8129 & ~n13940 ) ;
  assign n13942 = n13941 ^ n8755 ^ x92 ;
  assign n13943 = n8319 ^ n2089 ^ n1766 ;
  assign n13944 = n13943 ^ n5946 ^ 1'b0 ;
  assign n13945 = n13942 & ~n13944 ;
  assign n13947 = ( n1687 & ~n1724 ) | ( n1687 & n4890 ) | ( ~n1724 & n4890 ) ;
  assign n13946 = n2181 | n10011 ;
  assign n13948 = n13947 ^ n13946 ^ 1'b0 ;
  assign n13949 = n13948 ^ n6117 ^ 1'b0 ;
  assign n13959 = n744 & n5545 ;
  assign n13960 = ~n1224 & n13959 ;
  assign n13957 = n10389 ^ n5688 ^ n1445 ;
  assign n13955 = ( ~n750 & n6010 ) | ( ~n750 & n9596 ) | ( n6010 & n9596 ) ;
  assign n13956 = n13955 ^ n1981 ^ n1199 ;
  assign n13958 = n13957 ^ n13956 ^ x41 ;
  assign n13961 = n13960 ^ n13958 ^ n6496 ;
  assign n13962 = ( n6000 & ~n8475 ) | ( n6000 & n13961 ) | ( ~n8475 & n13961 ) ;
  assign n13952 = ( n1670 & n7653 ) | ( n1670 & n8615 ) | ( n7653 & n8615 ) ;
  assign n13950 = n11826 ^ n5072 ^ n3696 ;
  assign n13951 = ~n6244 & n13950 ;
  assign n13953 = n13952 ^ n13951 ^ 1'b0 ;
  assign n13954 = ( n6161 & ~n8514 ) | ( n6161 & n13953 ) | ( ~n8514 & n13953 ) ;
  assign n13963 = n13962 ^ n13954 ^ n4637 ;
  assign n13964 = n11966 ^ n7914 ^ n4018 ;
  assign n13966 = n8489 ^ x235 ^ x18 ;
  assign n13965 = n1092 | n8454 ;
  assign n13967 = n13966 ^ n13965 ^ 1'b0 ;
  assign n13968 = n13967 ^ n10810 ^ n9434 ;
  assign n13970 = ( ~n357 & n751 ) | ( ~n357 & n3412 ) | ( n751 & n3412 ) ;
  assign n13971 = n13970 ^ n1786 ^ n903 ;
  assign n13969 = n2941 | n5643 ;
  assign n13972 = n13971 ^ n13969 ^ 1'b0 ;
  assign n13975 = ( x52 & n9825 ) | ( x52 & ~n10177 ) | ( n9825 & ~n10177 ) ;
  assign n13973 = n13713 ^ n5310 ^ n1709 ;
  assign n13974 = ( n3433 & n11430 ) | ( n3433 & ~n13973 ) | ( n11430 & ~n13973 ) ;
  assign n13976 = n13975 ^ n13974 ^ n12684 ;
  assign n13977 = n13976 ^ n2371 ^ 1'b0 ;
  assign n13978 = n13972 & n13977 ;
  assign n13979 = n13978 ^ n13729 ^ 1'b0 ;
  assign n13982 = ( n3009 & n4533 ) | ( n3009 & ~n5802 ) | ( n4533 & ~n5802 ) ;
  assign n13983 = ( ~n2174 & n7747 ) | ( ~n2174 & n13982 ) | ( n7747 & n13982 ) ;
  assign n13984 = n13983 ^ n9892 ^ n8636 ;
  assign n13985 = ( n1200 & n4819 ) | ( n1200 & ~n13984 ) | ( n4819 & ~n13984 ) ;
  assign n13980 = n8990 ^ n8240 ^ n4941 ;
  assign n13981 = n13980 ^ n11991 ^ n9004 ;
  assign n13986 = n13985 ^ n13981 ^ n10711 ;
  assign n13987 = ( n4263 & n5565 ) | ( n4263 & ~n11337 ) | ( n5565 & ~n11337 ) ;
  assign n13988 = n12510 & n13987 ;
  assign n13989 = ~n13986 & n13988 ;
  assign n13990 = ~n7542 & n9817 ;
  assign n13991 = n8365 & n13990 ;
  assign n13992 = n12505 ^ n5525 ^ n4257 ;
  assign n13993 = ( n1298 & n2661 ) | ( n1298 & n13992 ) | ( n2661 & n13992 ) ;
  assign n13995 = ( n3300 & n7552 ) | ( n3300 & ~n11468 ) | ( n7552 & ~n11468 ) ;
  assign n13994 = n5179 ^ n4801 ^ n4399 ;
  assign n13996 = n13995 ^ n13994 ^ n5888 ;
  assign n13997 = ( n11037 & n12230 ) | ( n11037 & ~n13996 ) | ( n12230 & ~n13996 ) ;
  assign n13998 = n7752 ^ n5576 ^ n2892 ;
  assign n13999 = n13998 ^ n7592 ^ n1448 ;
  assign n14000 = ( n3756 & n5502 ) | ( n3756 & n6138 ) | ( n5502 & n6138 ) ;
  assign n14001 = n14000 ^ n3404 ^ n1368 ;
  assign n14002 = ( ~n1803 & n8843 ) | ( ~n1803 & n14001 ) | ( n8843 & n14001 ) ;
  assign n14003 = ( n13749 & ~n13999 ) | ( n13749 & n14002 ) | ( ~n13999 & n14002 ) ;
  assign n14004 = ( n1540 & ~n8504 ) | ( n1540 & n10078 ) | ( ~n8504 & n10078 ) ;
  assign n14005 = ( n3104 & n14003 ) | ( n3104 & ~n14004 ) | ( n14003 & ~n14004 ) ;
  assign n14006 = n13045 ^ n7139 ^ n6514 ;
  assign n14007 = n14006 ^ n5658 ^ n1639 ;
  assign n14021 = n13742 ^ n6896 ^ 1'b0 ;
  assign n14022 = n7399 & n14021 ;
  assign n14015 = n1349 & n4576 ;
  assign n14013 = n8707 ^ n1029 ^ 1'b0 ;
  assign n14014 = n14013 ^ n2471 ^ x46 ;
  assign n14012 = ( n2537 & n4958 ) | ( n2537 & ~n7214 ) | ( n4958 & ~n7214 ) ;
  assign n14016 = n14015 ^ n14014 ^ n14012 ;
  assign n14017 = ( n7911 & n8546 ) | ( n7911 & n14016 ) | ( n8546 & n14016 ) ;
  assign n14011 = n1935 & n6506 ;
  assign n14018 = n14017 ^ n14011 ^ 1'b0 ;
  assign n14019 = ( n11382 & n13595 ) | ( n11382 & ~n14018 ) | ( n13595 & ~n14018 ) ;
  assign n14008 = n3487 | n3566 ;
  assign n14009 = n14008 ^ n7682 ^ n1095 ;
  assign n14010 = ( n1961 & n13902 ) | ( n1961 & ~n14009 ) | ( n13902 & ~n14009 ) ;
  assign n14020 = n14019 ^ n14010 ^ n1437 ;
  assign n14023 = n14022 ^ n14020 ^ n8489 ;
  assign n14026 = ( ~n1004 & n9448 ) | ( ~n1004 & n12876 ) | ( n9448 & n12876 ) ;
  assign n14024 = n9777 ^ n6354 ^ 1'b0 ;
  assign n14025 = n3475 & n14024 ;
  assign n14027 = n14026 ^ n14025 ^ n12966 ;
  assign n14028 = n14027 ^ n5386 ^ n3495 ;
  assign n14029 = n5907 ^ n4792 ^ n362 ;
  assign n14030 = ( n286 & n6799 ) | ( n286 & ~n14029 ) | ( n6799 & ~n14029 ) ;
  assign n14031 = n14030 ^ n4455 ^ 1'b0 ;
  assign n14032 = n3384 & n6903 ;
  assign n14033 = n14032 ^ n598 ^ 1'b0 ;
  assign n14034 = ( n13817 & n14031 ) | ( n13817 & n14033 ) | ( n14031 & n14033 ) ;
  assign n14035 = ( n7644 & ~n8636 ) | ( n7644 & n14034 ) | ( ~n8636 & n14034 ) ;
  assign n14036 = ( n4649 & ~n9030 ) | ( n4649 & n11162 ) | ( ~n9030 & n11162 ) ;
  assign n14037 = ( ~n1279 & n7234 ) | ( ~n1279 & n8060 ) | ( n7234 & n8060 ) ;
  assign n14038 = ( n5660 & n14036 ) | ( n5660 & n14037 ) | ( n14036 & n14037 ) ;
  assign n14044 = n9069 ^ n6263 ^ 1'b0 ;
  assign n14040 = n2605 ^ n548 ^ n291 ;
  assign n14041 = ( ~n2977 & n6929 ) | ( ~n2977 & n14040 ) | ( n6929 & n14040 ) ;
  assign n14042 = n14041 ^ n8324 ^ n5539 ;
  assign n14043 = ( n5379 & n8464 ) | ( n5379 & ~n14042 ) | ( n8464 & ~n14042 ) ;
  assign n14039 = n12486 ^ n4049 ^ n1484 ;
  assign n14045 = n14044 ^ n14043 ^ n14039 ;
  assign n14046 = n2563 ^ n2394 ^ x213 ;
  assign n14047 = ( ~n3501 & n6715 ) | ( ~n3501 & n14046 ) | ( n6715 & n14046 ) ;
  assign n14048 = n9601 ^ n1317 ^ n269 ;
  assign n14049 = n14048 ^ n5065 ^ n4299 ;
  assign n14050 = ( ~n873 & n7978 ) | ( ~n873 & n14049 ) | ( n7978 & n14049 ) ;
  assign n14051 = ( n7892 & ~n12840 ) | ( n7892 & n14050 ) | ( ~n12840 & n14050 ) ;
  assign n14052 = ( n3698 & n5705 ) | ( n3698 & n14051 ) | ( n5705 & n14051 ) ;
  assign n14053 = ( n2911 & ~n6166 ) | ( n2911 & n14052 ) | ( ~n6166 & n14052 ) ;
  assign n14054 = ( n6913 & n14047 ) | ( n6913 & ~n14053 ) | ( n14047 & ~n14053 ) ;
  assign n14055 = n8518 & n12372 ;
  assign n14056 = n10735 & n14055 ;
  assign n14057 = ~n2738 & n11097 ;
  assign n14059 = ( n439 & n1580 ) | ( n439 & n3264 ) | ( n1580 & n3264 ) ;
  assign n14058 = n319 | n4741 ;
  assign n14060 = n14059 ^ n14058 ^ 1'b0 ;
  assign n14061 = n13364 ^ n3941 ^ n2914 ;
  assign n14066 = x213 & ~n2317 ;
  assign n14067 = n3260 & n14066 ;
  assign n14068 = ( n3333 & ~n11672 ) | ( n3333 & n14067 ) | ( ~n11672 & n14067 ) ;
  assign n14062 = n4331 | n8042 ;
  assign n14063 = n14062 ^ n8484 ^ 1'b0 ;
  assign n14064 = ( n8428 & n10107 ) | ( n8428 & ~n14063 ) | ( n10107 & ~n14063 ) ;
  assign n14065 = ( ~n5867 & n9298 ) | ( ~n5867 & n14064 ) | ( n9298 & n14064 ) ;
  assign n14069 = n14068 ^ n14065 ^ n506 ;
  assign n14070 = ( ~n14060 & n14061 ) | ( ~n14060 & n14069 ) | ( n14061 & n14069 ) ;
  assign n14071 = ( n8430 & ~n9420 ) | ( n8430 & n10806 ) | ( ~n9420 & n10806 ) ;
  assign n14072 = n10862 ^ n10737 ^ n5946 ;
  assign n14073 = n14072 ^ n8345 ^ n3109 ;
  assign n14074 = ( n12116 & ~n14071 ) | ( n12116 & n14073 ) | ( ~n14071 & n14073 ) ;
  assign n14075 = n2741 & n3623 ;
  assign n14076 = ~n14074 & n14075 ;
  assign n14077 = ( n4352 & n8113 ) | ( n4352 & n8573 ) | ( n8113 & n8573 ) ;
  assign n14078 = ( n1513 & n5438 ) | ( n1513 & n14077 ) | ( n5438 & n14077 ) ;
  assign n14079 = ( n1487 & n1897 ) | ( n1487 & ~n3759 ) | ( n1897 & ~n3759 ) ;
  assign n14080 = ( n5245 & ~n7516 ) | ( n5245 & n14079 ) | ( ~n7516 & n14079 ) ;
  assign n14081 = n14080 ^ n9419 ^ n1424 ;
  assign n14082 = n8475 ^ n1102 ^ n1097 ;
  assign n14083 = ( ~n7251 & n10437 ) | ( ~n7251 & n11619 ) | ( n10437 & n11619 ) ;
  assign n14084 = ( n1620 & n3922 ) | ( n1620 & n13705 ) | ( n3922 & n13705 ) ;
  assign n14085 = n7553 ^ n6044 ^ n5268 ;
  assign n14086 = ( n1877 & n11392 ) | ( n1877 & ~n14085 ) | ( n11392 & ~n14085 ) ;
  assign n14087 = n14086 ^ n3087 ^ n291 ;
  assign n14088 = n632 & ~n758 ;
  assign n14089 = n14088 ^ n13995 ^ 1'b0 ;
  assign n14090 = ( ~n7306 & n12884 ) | ( ~n7306 & n14089 ) | ( n12884 & n14089 ) ;
  assign n14091 = ( n11980 & n14087 ) | ( n11980 & ~n14090 ) | ( n14087 & ~n14090 ) ;
  assign n14092 = n14091 ^ n4262 ^ 1'b0 ;
  assign n14093 = n14084 & ~n14092 ;
  assign n14094 = n12321 ^ n9654 ^ 1'b0 ;
  assign n14095 = ( n6013 & n6467 ) | ( n6013 & n14094 ) | ( n6467 & n14094 ) ;
  assign n14104 = ( n4278 & n4505 ) | ( n4278 & n4599 ) | ( n4505 & n4599 ) ;
  assign n14105 = n7110 & ~n10452 ;
  assign n14106 = ~n14104 & n14105 ;
  assign n14101 = n4460 ^ n1046 ^ n867 ;
  assign n14102 = ( n746 & n4040 ) | ( n746 & n14101 ) | ( n4040 & n14101 ) ;
  assign n14098 = ( n9446 & n10711 ) | ( n9446 & ~n13788 ) | ( n10711 & ~n13788 ) ;
  assign n14099 = n8973 ^ n2533 ^ 1'b0 ;
  assign n14100 = n14098 & n14099 ;
  assign n14103 = n14102 ^ n14100 ^ n11554 ;
  assign n14096 = n9189 ^ n5422 ^ n838 ;
  assign n14097 = n5298 & n14096 ;
  assign n14107 = n14106 ^ n14103 ^ n14097 ;
  assign n14108 = n14107 ^ n3783 ^ 1'b0 ;
  assign n14109 = ( n3869 & ~n4357 ) | ( n3869 & n4500 ) | ( ~n4357 & n4500 ) ;
  assign n14110 = n2767 | n14109 ;
  assign n14111 = n14108 | n14110 ;
  assign n14114 = n1619 ^ x220 ^ 1'b0 ;
  assign n14115 = n14114 ^ n13898 ^ n7255 ;
  assign n14112 = n6391 ^ n2555 ^ x50 ;
  assign n14113 = n14112 ^ n13845 ^ 1'b0 ;
  assign n14116 = n14115 ^ n14113 ^ n8346 ;
  assign n14117 = ( n979 & n9812 ) | ( n979 & ~n14116 ) | ( n9812 & ~n14116 ) ;
  assign n14118 = ( n584 & n1657 ) | ( n584 & ~n14117 ) | ( n1657 & ~n14117 ) ;
  assign n14119 = n895 & n14118 ;
  assign n14120 = n14119 ^ n12937 ^ 1'b0 ;
  assign n14121 = ( ~n4228 & n7110 ) | ( ~n4228 & n11135 ) | ( n7110 & n11135 ) ;
  assign n14122 = ( n1111 & ~n8098 ) | ( n1111 & n12814 ) | ( ~n8098 & n12814 ) ;
  assign n14123 = n2353 & ~n14122 ;
  assign n14124 = ~x203 & n14123 ;
  assign n14126 = n9492 ^ n4698 ^ n732 ;
  assign n14125 = n2929 & ~n8359 ;
  assign n14127 = n14126 ^ n14125 ^ n4737 ;
  assign n14128 = ( ~n12130 & n14124 ) | ( ~n12130 & n14127 ) | ( n14124 & n14127 ) ;
  assign n14131 = n1488 & n3335 ;
  assign n14132 = n3571 & n14131 ;
  assign n14129 = ( n2731 & n2869 ) | ( n2731 & n5612 ) | ( n2869 & n5612 ) ;
  assign n14130 = n3356 & ~n14129 ;
  assign n14133 = n14132 ^ n14130 ^ n3742 ;
  assign n14135 = n4850 ^ n4215 ^ x36 ;
  assign n14136 = n14135 ^ n6233 ^ 1'b0 ;
  assign n14134 = n8014 ^ n2627 ^ n485 ;
  assign n14137 = n14136 ^ n14134 ^ n2257 ;
  assign n14138 = ( n2398 & ~n4988 ) | ( n2398 & n14137 ) | ( ~n4988 & n14137 ) ;
  assign n14139 = n5492 | n9628 ;
  assign n14140 = n12632 ^ n8256 ^ n7377 ;
  assign n14141 = n14140 ^ n7155 ^ n2699 ;
  assign n14142 = ( n5302 & n14139 ) | ( n5302 & n14141 ) | ( n14139 & n14141 ) ;
  assign n14143 = ( ~n7774 & n8344 ) | ( ~n7774 & n11194 ) | ( n8344 & n11194 ) ;
  assign n14144 = ( n272 & n1362 ) | ( n272 & n8095 ) | ( n1362 & n8095 ) ;
  assign n14145 = n14144 ^ n10183 ^ n5106 ;
  assign n14146 = ( n14142 & n14143 ) | ( n14142 & n14145 ) | ( n14143 & n14145 ) ;
  assign n14147 = ~n6727 & n9040 ;
  assign n14148 = ( n3706 & n12641 ) | ( n3706 & ~n14147 ) | ( n12641 & ~n14147 ) ;
  assign n14149 = n2902 & n4839 ;
  assign n14150 = n14149 ^ n14029 ^ n6806 ;
  assign n14151 = ( n6587 & n9379 ) | ( n6587 & n14150 ) | ( n9379 & n14150 ) ;
  assign n14152 = ( ~n1571 & n3658 ) | ( ~n1571 & n5984 ) | ( n3658 & n5984 ) ;
  assign n14153 = n3983 & n14152 ;
  assign n14154 = n14153 ^ n12036 ^ 1'b0 ;
  assign n14155 = n11622 ^ n4029 ^ n660 ;
  assign n14156 = ( n8074 & n12561 ) | ( n8074 & n14155 ) | ( n12561 & n14155 ) ;
  assign n14157 = n14156 ^ n11002 ^ n1708 ;
  assign n14161 = n5808 | n8653 ;
  assign n14162 = n14161 ^ n7590 ^ n2618 ;
  assign n14158 = n13874 ^ n11692 ^ n2508 ;
  assign n14159 = n9960 ^ n7418 ^ n3356 ;
  assign n14160 = ( n4219 & ~n14158 ) | ( n4219 & n14159 ) | ( ~n14158 & n14159 ) ;
  assign n14163 = n14162 ^ n14160 ^ n3763 ;
  assign n14164 = n14163 ^ n8682 ^ n7338 ;
  assign n14165 = ( ~n3690 & n7192 ) | ( ~n3690 & n11994 ) | ( n7192 & n11994 ) ;
  assign n14166 = ( n1624 & n2913 ) | ( n1624 & ~n7640 ) | ( n2913 & ~n7640 ) ;
  assign n14167 = ( n940 & n10219 ) | ( n940 & n11009 ) | ( n10219 & n11009 ) ;
  assign n14168 = ( n9884 & n14166 ) | ( n9884 & ~n14167 ) | ( n14166 & ~n14167 ) ;
  assign n14169 = n14168 ^ n7395 ^ n4156 ;
  assign n14174 = ( n6281 & n7308 ) | ( n6281 & ~n8430 ) | ( n7308 & ~n8430 ) ;
  assign n14170 = n11443 ^ n7979 ^ n6812 ;
  assign n14171 = n6649 ^ n5850 ^ n3699 ;
  assign n14172 = ( ~n2168 & n6256 ) | ( ~n2168 & n14171 ) | ( n6256 & n14171 ) ;
  assign n14173 = n14170 & ~n14172 ;
  assign n14175 = n14174 ^ n14173 ^ 1'b0 ;
  assign n14176 = ( n14165 & n14169 ) | ( n14165 & n14175 ) | ( n14169 & n14175 ) ;
  assign n14178 = ( n962 & n1121 ) | ( n962 & ~n11169 ) | ( n1121 & ~n11169 ) ;
  assign n14177 = ( ~n6235 & n6478 ) | ( ~n6235 & n7395 ) | ( n6478 & n7395 ) ;
  assign n14179 = n14178 ^ n14177 ^ n487 ;
  assign n14180 = ( ~n1156 & n2153 ) | ( ~n1156 & n4361 ) | ( n2153 & n4361 ) ;
  assign n14181 = n14180 ^ n10256 ^ n3802 ;
  assign n14182 = n907 | n8216 ;
  assign n14183 = ( n1610 & n2015 ) | ( n1610 & ~n14182 ) | ( n2015 & ~n14182 ) ;
  assign n14184 = ( n3276 & n14181 ) | ( n3276 & n14183 ) | ( n14181 & n14183 ) ;
  assign n14185 = ( n2327 & n6527 ) | ( n2327 & ~n14184 ) | ( n6527 & ~n14184 ) ;
  assign n14186 = n11659 ^ n2254 ^ 1'b0 ;
  assign n14187 = n14185 & ~n14186 ;
  assign n14188 = ( n7714 & ~n10815 ) | ( n7714 & n14187 ) | ( ~n10815 & n14187 ) ;
  assign n14204 = n5706 ^ n2727 ^ n1162 ;
  assign n14198 = n8549 ^ n4565 ^ n2978 ;
  assign n14199 = n2759 | n4831 ;
  assign n14200 = n14199 ^ n738 ^ 1'b0 ;
  assign n14201 = ~n2618 & n14200 ;
  assign n14202 = ( n5924 & ~n6328 ) | ( n5924 & n14201 ) | ( ~n6328 & n14201 ) ;
  assign n14203 = ( ~n868 & n14198 ) | ( ~n868 & n14202 ) | ( n14198 & n14202 ) ;
  assign n14196 = ( n597 & n6205 ) | ( n597 & ~n8948 ) | ( n6205 & ~n8948 ) ;
  assign n14194 = n2787 & ~n10399 ;
  assign n14189 = n874 ^ n544 ^ x17 ;
  assign n14190 = n4354 ^ n3889 ^ n1402 ;
  assign n14191 = ( n4297 & ~n14189 ) | ( n4297 & n14190 ) | ( ~n14189 & n14190 ) ;
  assign n14192 = ( n3632 & ~n11153 ) | ( n3632 & n14191 ) | ( ~n11153 & n14191 ) ;
  assign n14193 = n14192 ^ n5577 ^ n3481 ;
  assign n14195 = n14194 ^ n14193 ^ 1'b0 ;
  assign n14197 = n14196 ^ n14195 ^ n11770 ;
  assign n14205 = n14204 ^ n14203 ^ n14197 ;
  assign n14206 = n14205 ^ n1378 ^ n880 ;
  assign n14207 = n9466 ^ n2127 ^ n375 ;
  assign n14208 = n14207 ^ n8902 ^ n8808 ;
  assign n14209 = n7685 ^ n3422 ^ n1933 ;
  assign n14210 = n14209 ^ n12343 ^ n10549 ;
  assign n14211 = n940 & n1294 ;
  assign n14212 = n14211 ^ n7416 ^ 1'b0 ;
  assign n14213 = ( n4498 & ~n11008 ) | ( n4498 & n14212 ) | ( ~n11008 & n14212 ) ;
  assign n14214 = n14213 ^ n6952 ^ n4990 ;
  assign n14215 = n6892 ^ n1482 ^ n1325 ;
  assign n14216 = ( ~n4115 & n8718 ) | ( ~n4115 & n14215 ) | ( n8718 & n14215 ) ;
  assign n14217 = ( ~n4689 & n14214 ) | ( ~n4689 & n14216 ) | ( n14214 & n14216 ) ;
  assign n14218 = n13084 ^ n1502 ^ n787 ;
  assign n14219 = ( n6392 & ~n13307 ) | ( n6392 & n14218 ) | ( ~n13307 & n14218 ) ;
  assign n14220 = ( ~n2200 & n9178 ) | ( ~n2200 & n14219 ) | ( n9178 & n14219 ) ;
  assign n14221 = n6967 & n7183 ;
  assign n14222 = ~n3502 & n14221 ;
  assign n14223 = n14222 ^ n2642 ^ 1'b0 ;
  assign n14224 = ~n4008 & n14223 ;
  assign n14225 = ( ~n977 & n5836 ) | ( ~n977 & n7786 ) | ( n5836 & n7786 ) ;
  assign n14226 = n14225 ^ n13616 ^ 1'b0 ;
  assign n14227 = ~n11005 & n14226 ;
  assign n14228 = ( n2705 & n9083 ) | ( n2705 & ~n14227 ) | ( n9083 & ~n14227 ) ;
  assign n14229 = ( n335 & n817 ) | ( n335 & n901 ) | ( n817 & n901 ) ;
  assign n14230 = n14229 ^ n11912 ^ n8943 ;
  assign n14231 = ( n7182 & n14228 ) | ( n7182 & ~n14230 ) | ( n14228 & ~n14230 ) ;
  assign n14232 = ( n14220 & n14224 ) | ( n14220 & ~n14231 ) | ( n14224 & ~n14231 ) ;
  assign n14233 = ( n760 & n2440 ) | ( n760 & n2857 ) | ( n2440 & n2857 ) ;
  assign n14234 = ( n1072 & ~n2578 ) | ( n1072 & n4087 ) | ( ~n2578 & n4087 ) ;
  assign n14235 = ( ~n2462 & n14233 ) | ( ~n2462 & n14234 ) | ( n14233 & n14234 ) ;
  assign n14236 = ( ~n8970 & n13657 ) | ( ~n8970 & n14235 ) | ( n13657 & n14235 ) ;
  assign n14237 = n9465 ^ n9022 ^ n544 ;
  assign n14238 = n9327 ^ n7343 ^ 1'b0 ;
  assign n14239 = ( n8162 & n10990 ) | ( n8162 & ~n14238 ) | ( n10990 & ~n14238 ) ;
  assign n14244 = n10322 ^ n7829 ^ n5359 ;
  assign n14245 = ( ~n3535 & n9777 ) | ( ~n3535 & n14244 ) | ( n9777 & n14244 ) ;
  assign n14240 = ( ~n2225 & n9507 ) | ( ~n2225 & n10130 ) | ( n9507 & n10130 ) ;
  assign n14241 = n9094 | n12390 ;
  assign n14242 = n14240 & ~n14241 ;
  assign n14243 = ( n3150 & n7276 ) | ( n3150 & n14242 ) | ( n7276 & n14242 ) ;
  assign n14246 = n14245 ^ n14243 ^ n6851 ;
  assign n14247 = ( n14237 & ~n14239 ) | ( n14237 & n14246 ) | ( ~n14239 & n14246 ) ;
  assign n14259 = n13363 ^ n5276 ^ 1'b0 ;
  assign n14253 = n7505 ^ n4364 ^ x108 ;
  assign n14254 = ( ~x133 & n589 ) | ( ~x133 & n10782 ) | ( n589 & n10782 ) ;
  assign n14255 = n14254 ^ n1586 ^ 1'b0 ;
  assign n14256 = n10523 & n14255 ;
  assign n14257 = ( n858 & n14253 ) | ( n858 & n14256 ) | ( n14253 & n14256 ) ;
  assign n14248 = n12261 ^ n4611 ^ n3860 ;
  assign n14249 = ( n1036 & ~n2267 ) | ( n1036 & n2445 ) | ( ~n2267 & n2445 ) ;
  assign n14250 = ( ~n838 & n1809 ) | ( ~n838 & n14249 ) | ( n1809 & n14249 ) ;
  assign n14251 = ( n5705 & n10368 ) | ( n5705 & n11650 ) | ( n10368 & n11650 ) ;
  assign n14252 = ( n14248 & n14250 ) | ( n14248 & ~n14251 ) | ( n14250 & ~n14251 ) ;
  assign n14258 = n14257 ^ n14252 ^ n4013 ;
  assign n14260 = n14259 ^ n14258 ^ n12172 ;
  assign n14262 = ( n309 & n1696 ) | ( n309 & n1906 ) | ( n1696 & n1906 ) ;
  assign n14261 = ( ~n1523 & n2566 ) | ( ~n1523 & n4314 ) | ( n2566 & n4314 ) ;
  assign n14263 = n14262 ^ n14261 ^ n5161 ;
  assign n14264 = n14040 ^ n9164 ^ n400 ;
  assign n14265 = n14264 ^ n3071 ^ n1989 ;
  assign n14266 = ( ~n875 & n14263 ) | ( ~n875 & n14265 ) | ( n14263 & n14265 ) ;
  assign n14267 = ( n3580 & ~n4625 ) | ( n3580 & n11438 ) | ( ~n4625 & n11438 ) ;
  assign n14268 = n10557 ^ n9841 ^ n2360 ;
  assign n14269 = n8291 & ~n13560 ;
  assign n14270 = ( n4925 & ~n14268 ) | ( n4925 & n14269 ) | ( ~n14268 & n14269 ) ;
  assign n14271 = n14270 ^ n8246 ^ n5808 ;
  assign n14272 = ( n12431 & ~n14267 ) | ( n12431 & n14271 ) | ( ~n14267 & n14271 ) ;
  assign n14276 = n6198 & ~n8968 ;
  assign n14273 = n1114 & ~n1116 ;
  assign n14274 = n14273 ^ n10889 ^ n807 ;
  assign n14275 = ( n659 & n8319 ) | ( n659 & n14274 ) | ( n8319 & n14274 ) ;
  assign n14277 = n14276 ^ n14275 ^ n11847 ;
  assign n14278 = ( n900 & ~n1452 ) | ( n900 & n4464 ) | ( ~n1452 & n4464 ) ;
  assign n14280 = n11249 ^ n9958 ^ n3525 ;
  assign n14279 = ~n3910 & n8485 ;
  assign n14281 = n14280 ^ n14279 ^ 1'b0 ;
  assign n14282 = ( n6652 & n14278 ) | ( n6652 & ~n14281 ) | ( n14278 & ~n14281 ) ;
  assign n14283 = n5548 ^ n448 ^ 1'b0 ;
  assign n14284 = ( n8666 & n10772 ) | ( n8666 & ~n14283 ) | ( n10772 & ~n14283 ) ;
  assign n14285 = n3406 ^ x180 ^ x85 ;
  assign n14286 = ( n3844 & ~n3864 ) | ( n3844 & n14285 ) | ( ~n3864 & n14285 ) ;
  assign n14287 = ( ~n487 & n5248 ) | ( ~n487 & n7476 ) | ( n5248 & n7476 ) ;
  assign n14288 = ( n3924 & n11557 ) | ( n3924 & ~n14287 ) | ( n11557 & ~n14287 ) ;
  assign n14289 = n9602 | n14288 ;
  assign n14290 = ( n1276 & ~n14286 ) | ( n1276 & n14289 ) | ( ~n14286 & n14289 ) ;
  assign n14293 = ( n3871 & n4237 ) | ( n3871 & ~n6906 ) | ( n4237 & ~n6906 ) ;
  assign n14291 = n6064 & ~n12120 ;
  assign n14292 = n14291 ^ n7563 ^ 1'b0 ;
  assign n14294 = n14293 ^ n14292 ^ n8703 ;
  assign n14295 = ( n5231 & n9905 ) | ( n5231 & ~n14294 ) | ( n9905 & ~n14294 ) ;
  assign n14296 = ( n469 & n9576 ) | ( n469 & n9773 ) | ( n9576 & n9773 ) ;
  assign n14297 = n2888 & n4140 ;
  assign n14298 = n14297 ^ n5322 ^ 1'b0 ;
  assign n14299 = n5637 | n14298 ;
  assign n14300 = ( ~n9267 & n14296 ) | ( ~n9267 & n14299 ) | ( n14296 & n14299 ) ;
  assign n14301 = ( n6099 & n8589 ) | ( n6099 & n13792 ) | ( n8589 & n13792 ) ;
  assign n14304 = n12142 ^ n5007 ^ n4963 ;
  assign n14305 = ~n6959 & n14304 ;
  assign n14306 = n14305 ^ n10422 ^ 1'b0 ;
  assign n14302 = ( n4074 & ~n8944 ) | ( n4074 & n9016 ) | ( ~n8944 & n9016 ) ;
  assign n14303 = ( n1104 & ~n11604 ) | ( n1104 & n14302 ) | ( ~n11604 & n14302 ) ;
  assign n14307 = n14306 ^ n14303 ^ 1'b0 ;
  assign n14308 = n12399 & ~n14307 ;
  assign n14309 = n7729 & ~n12582 ;
  assign n14310 = n8099 & n14309 ;
  assign n14311 = ( ~n3084 & n7178 ) | ( ~n3084 & n14310 ) | ( n7178 & n14310 ) ;
  assign n14312 = ~n3836 & n8045 ;
  assign n14313 = n14312 ^ n5131 ^ 1'b0 ;
  assign n14314 = ( n1756 & n3417 ) | ( n1756 & n14313 ) | ( n3417 & n14313 ) ;
  assign n14315 = n10977 ^ n9651 ^ 1'b0 ;
  assign n14316 = n772 & n1693 ;
  assign n14317 = n14316 ^ n6185 ^ n5721 ;
  assign n14318 = n14317 ^ n3302 ^ n1835 ;
  assign n14321 = n3432 ^ n1925 ^ n789 ;
  assign n14322 = n14321 ^ n8632 ^ n2639 ;
  assign n14323 = ( n346 & ~n1934 ) | ( n346 & n14322 ) | ( ~n1934 & n14322 ) ;
  assign n14324 = ( ~n7887 & n11322 ) | ( ~n7887 & n14323 ) | ( n11322 & n14323 ) ;
  assign n14319 = n1447 | n3237 ;
  assign n14320 = n10867 | n14319 ;
  assign n14325 = n14324 ^ n14320 ^ 1'b0 ;
  assign n14326 = n14325 ^ n12530 ^ n9020 ;
  assign n14327 = ( n2556 & ~n2751 ) | ( n2556 & n7466 ) | ( ~n2751 & n7466 ) ;
  assign n14328 = ( x0 & n8569 ) | ( x0 & n14327 ) | ( n8569 & n14327 ) ;
  assign n14329 = n14328 ^ n5870 ^ n3695 ;
  assign n14339 = ~x147 & n1767 ;
  assign n14330 = n3250 ^ n2091 ^ n896 ;
  assign n14331 = n14330 ^ n4787 ^ n1277 ;
  assign n14332 = n8766 ^ n4389 ^ n956 ;
  assign n14333 = n8983 | n14332 ;
  assign n14334 = ( n7441 & n14331 ) | ( n7441 & n14333 ) | ( n14331 & n14333 ) ;
  assign n14336 = ( ~n561 & n2934 ) | ( ~n561 & n7621 ) | ( n2934 & n7621 ) ;
  assign n14335 = n12257 ^ n7972 ^ n2320 ;
  assign n14337 = n14336 ^ n14335 ^ n1016 ;
  assign n14338 = ( x238 & n14334 ) | ( x238 & n14337 ) | ( n14334 & n14337 ) ;
  assign n14340 = n14339 ^ n14338 ^ 1'b0 ;
  assign n14341 = n4644 & n5189 ;
  assign n14342 = n2322 & n14341 ;
  assign n14343 = n3713 & n11274 ;
  assign n14344 = ~n9357 & n14343 ;
  assign n14345 = ( n4882 & n8297 ) | ( n4882 & n14344 ) | ( n8297 & n14344 ) ;
  assign n14346 = n9042 ^ n4794 ^ n1136 ;
  assign n14347 = ( n562 & n1694 ) | ( n562 & n14346 ) | ( n1694 & n14346 ) ;
  assign n14348 = ( n335 & n14345 ) | ( n335 & ~n14347 ) | ( n14345 & ~n14347 ) ;
  assign n14349 = n10734 ^ n9291 ^ x42 ;
  assign n14350 = ( x196 & ~n6216 ) | ( x196 & n14349 ) | ( ~n6216 & n14349 ) ;
  assign n14351 = n14350 ^ n12831 ^ n6737 ;
  assign n14356 = ( n1763 & n3282 ) | ( n1763 & n5188 ) | ( n3282 & n5188 ) ;
  assign n14357 = ( n6962 & n10162 ) | ( n6962 & ~n14356 ) | ( n10162 & ~n14356 ) ;
  assign n14358 = n14357 ^ n3214 ^ n2174 ;
  assign n14354 = ( ~n1879 & n3085 ) | ( ~n1879 & n9420 ) | ( n3085 & n9420 ) ;
  assign n14355 = n14354 ^ n9050 ^ n8525 ;
  assign n14352 = n917 & ~n2777 ;
  assign n14353 = n14352 ^ n13443 ^ n7471 ;
  assign n14359 = n14358 ^ n14355 ^ n14353 ;
  assign n14365 = ( ~n1398 & n5951 ) | ( ~n1398 & n6824 ) | ( n5951 & n6824 ) ;
  assign n14366 = ( n11214 & ~n11338 ) | ( n11214 & n14365 ) | ( ~n11338 & n14365 ) ;
  assign n14360 = ( n2588 & ~n4516 ) | ( n2588 & n11352 ) | ( ~n4516 & n11352 ) ;
  assign n14361 = n3461 ^ n3310 ^ 1'b0 ;
  assign n14362 = n14360 & n14361 ;
  assign n14363 = n14362 ^ n11487 ^ n1395 ;
  assign n14364 = n14363 ^ n7645 ^ n829 ;
  assign n14367 = n14366 ^ n14364 ^ n2265 ;
  assign n14368 = ( ~n1849 & n8279 ) | ( ~n1849 & n14367 ) | ( n8279 & n14367 ) ;
  assign n14369 = n11069 & n14368 ;
  assign n14370 = n14359 & n14369 ;
  assign n14371 = ( n1367 & n2871 ) | ( n1367 & ~n7064 ) | ( n2871 & ~n7064 ) ;
  assign n14372 = n5574 ^ n1594 ^ 1'b0 ;
  assign n14373 = ( n1298 & n14371 ) | ( n1298 & n14372 ) | ( n14371 & n14372 ) ;
  assign n14374 = n7338 ^ n3141 ^ 1'b0 ;
  assign n14375 = n14374 ^ n9079 ^ 1'b0 ;
  assign n14376 = n3093 & n10782 ;
  assign n14377 = n12338 & n14376 ;
  assign n14378 = n7015 & n14377 ;
  assign n14379 = n14378 ^ n8265 ^ n6310 ;
  assign n14380 = ( ~n2287 & n5432 ) | ( ~n2287 & n8615 ) | ( n5432 & n8615 ) ;
  assign n14381 = ( ~n5628 & n7919 ) | ( ~n5628 & n9602 ) | ( n7919 & n9602 ) ;
  assign n14382 = ( x233 & n14380 ) | ( x233 & ~n14381 ) | ( n14380 & ~n14381 ) ;
  assign n14383 = n7734 ^ n5796 ^ n5165 ;
  assign n14384 = ( ~n6172 & n6493 ) | ( ~n6172 & n12900 ) | ( n6493 & n12900 ) ;
  assign n14385 = n14384 ^ n8165 ^ 1'b0 ;
  assign n14386 = n2827 & n14385 ;
  assign n14387 = ( ~n10605 & n10969 ) | ( ~n10605 & n14386 ) | ( n10969 & n14386 ) ;
  assign n14388 = ( n14382 & n14383 ) | ( n14382 & ~n14387 ) | ( n14383 & ~n14387 ) ;
  assign n14389 = ( n475 & n14379 ) | ( n475 & n14388 ) | ( n14379 & n14388 ) ;
  assign n14390 = ( ~n5458 & n9211 ) | ( ~n5458 & n10792 ) | ( n9211 & n10792 ) ;
  assign n14392 = n10452 ^ n1182 ^ 1'b0 ;
  assign n14391 = n858 | n13446 ;
  assign n14393 = n14392 ^ n14391 ^ 1'b0 ;
  assign n14397 = n9924 ^ n4633 ^ n1552 ;
  assign n14395 = n8876 ^ n8627 ^ 1'b0 ;
  assign n14396 = ~n11671 & n14395 ;
  assign n14398 = n14397 ^ n14396 ^ n9081 ;
  assign n14394 = ( n4627 & n10367 ) | ( n4627 & n12122 ) | ( n10367 & n12122 ) ;
  assign n14399 = n14398 ^ n14394 ^ n6322 ;
  assign n14400 = n11764 ^ n9105 ^ n7665 ;
  assign n14401 = n6900 | n7412 ;
  assign n14402 = n9619 & n14401 ;
  assign n14403 = n14400 & n14402 ;
  assign n14404 = n14403 ^ n9458 ^ n8001 ;
  assign n14405 = n14227 ^ n10437 ^ n4694 ;
  assign n14406 = ( n7882 & n10807 ) | ( n7882 & n14405 ) | ( n10807 & n14405 ) ;
  assign n14407 = n14406 ^ n11115 ^ n4498 ;
  assign n14408 = n14407 ^ n12109 ^ n10171 ;
  assign n14411 = n3478 ^ n1837 ^ x66 ;
  assign n14409 = ( n732 & n3547 ) | ( n732 & ~n8301 ) | ( n3547 & ~n8301 ) ;
  assign n14410 = n14409 ^ n2437 ^ n1565 ;
  assign n14412 = n14411 ^ n14410 ^ x69 ;
  assign n14413 = ( x222 & n11039 ) | ( x222 & ~n14412 ) | ( n11039 & ~n14412 ) ;
  assign n14414 = n14413 ^ n5156 ^ n1371 ;
  assign n14415 = n14414 ^ n9918 ^ n8658 ;
  assign n14417 = ( n2651 & n3446 ) | ( n2651 & ~n3938 ) | ( n3446 & ~n3938 ) ;
  assign n14418 = ( n2821 & ~n13463 ) | ( n2821 & n14417 ) | ( ~n13463 & n14417 ) ;
  assign n14416 = n3084 | n4533 ;
  assign n14419 = n14418 ^ n14416 ^ 1'b0 ;
  assign n14422 = ( n9038 & n9086 ) | ( n9038 & n11928 ) | ( n9086 & n11928 ) ;
  assign n14423 = ( ~n2447 & n6258 ) | ( ~n2447 & n14422 ) | ( n6258 & n14422 ) ;
  assign n14424 = n14423 ^ n11514 ^ n10453 ;
  assign n14420 = n3734 ^ n1417 ^ 1'b0 ;
  assign n14421 = ( n6877 & n8379 ) | ( n6877 & ~n14420 ) | ( n8379 & ~n14420 ) ;
  assign n14425 = n14424 ^ n14421 ^ n8588 ;
  assign n14431 = ( n3731 & n3914 ) | ( n3731 & n4160 ) | ( n3914 & n4160 ) ;
  assign n14428 = ( x122 & n823 ) | ( x122 & ~n5548 ) | ( n823 & ~n5548 ) ;
  assign n14429 = ( ~n800 & n6951 ) | ( ~n800 & n14428 ) | ( n6951 & n14428 ) ;
  assign n14430 = n14429 ^ n12819 ^ n10753 ;
  assign n14426 = n8971 | n9052 ;
  assign n14427 = n14426 ^ n2521 ^ 1'b0 ;
  assign n14432 = n14431 ^ n14430 ^ n14427 ;
  assign n14433 = n14293 ^ n9364 ^ n2498 ;
  assign n14434 = n14433 ^ n13561 ^ n739 ;
  assign n14440 = n8119 ^ n5622 ^ n566 ;
  assign n14441 = ( ~n1805 & n6033 ) | ( ~n1805 & n12754 ) | ( n6033 & n12754 ) ;
  assign n14442 = n14441 ^ n13448 ^ n5263 ;
  assign n14443 = n14442 ^ n5314 ^ n659 ;
  assign n14444 = n967 & ~n3687 ;
  assign n14445 = ( ~n3558 & n6622 ) | ( ~n3558 & n14444 ) | ( n6622 & n14444 ) ;
  assign n14446 = n14445 ^ n11106 ^ n5094 ;
  assign n14447 = ( n14440 & n14443 ) | ( n14440 & n14446 ) | ( n14443 & n14446 ) ;
  assign n14435 = n8009 ^ n2512 ^ n2102 ;
  assign n14436 = ( ~n750 & n6255 ) | ( ~n750 & n11871 ) | ( n6255 & n11871 ) ;
  assign n14437 = ( n7665 & ~n10492 ) | ( n7665 & n14436 ) | ( ~n10492 & n14436 ) ;
  assign n14438 = n14437 ^ n10197 ^ x89 ;
  assign n14439 = ( n9483 & n14435 ) | ( n9483 & ~n14438 ) | ( n14435 & ~n14438 ) ;
  assign n14448 = n14447 ^ n14439 ^ n13610 ;
  assign n14452 = n1268 | n6589 ;
  assign n14449 = n7443 ^ n4811 ^ n3290 ;
  assign n14450 = n14449 ^ n6223 ^ n1790 ;
  assign n14451 = n14450 ^ n9386 ^ n8381 ;
  assign n14453 = n14452 ^ n14451 ^ n7809 ;
  assign n14454 = n4082 | n6763 ;
  assign n14455 = n14454 ^ n1243 ^ 1'b0 ;
  assign n14456 = n14455 ^ n9591 ^ n4683 ;
  assign n14457 = n6515 ^ n3515 ^ n649 ;
  assign n14458 = n7076 | n10198 ;
  assign n14459 = n3456 | n14458 ;
  assign n14460 = n14457 & n14459 ;
  assign n14461 = ( n6878 & n14456 ) | ( n6878 & ~n14460 ) | ( n14456 & ~n14460 ) ;
  assign n14462 = ( x195 & n4079 ) | ( x195 & ~n8099 ) | ( n4079 & ~n8099 ) ;
  assign n14463 = n14462 ^ n14332 ^ n13757 ;
  assign n14464 = n14463 ^ n13103 ^ n5625 ;
  assign n14465 = n14464 ^ n9454 ^ n751 ;
  assign n14466 = n4307 ^ n2743 ^ n2563 ;
  assign n14467 = n14466 ^ n13907 ^ n2244 ;
  assign n14468 = n1540 & ~n14467 ;
  assign n14469 = n13513 & n14468 ;
  assign n14470 = ( n2249 & ~n2652 ) | ( n2249 & n12269 ) | ( ~n2652 & n12269 ) ;
  assign n14471 = n13760 ^ n11812 ^ x79 ;
  assign n14472 = ( n9717 & ~n14470 ) | ( n9717 & n14471 ) | ( ~n14470 & n14471 ) ;
  assign n14473 = ( n2291 & n5262 ) | ( n2291 & n12994 ) | ( n5262 & n12994 ) ;
  assign n14474 = n14473 ^ n11053 ^ n760 ;
  assign n14475 = n4170 & n14474 ;
  assign n14478 = n10164 ^ n6935 ^ n1560 ;
  assign n14476 = n3520 ^ n2935 ^ n1364 ;
  assign n14477 = n14476 ^ n3613 ^ n2464 ;
  assign n14479 = n14478 ^ n14477 ^ 1'b0 ;
  assign n14480 = ~n14201 & n14479 ;
  assign n14481 = n14480 ^ n11169 ^ x64 ;
  assign n14482 = ( n2509 & n6009 ) | ( n2509 & n14170 ) | ( n6009 & n14170 ) ;
  assign n14483 = ( n878 & n2791 ) | ( n878 & n9492 ) | ( n2791 & n9492 ) ;
  assign n14484 = n2638 & n7581 ;
  assign n14485 = ( n955 & ~n5304 ) | ( n955 & n6816 ) | ( ~n5304 & n6816 ) ;
  assign n14486 = ( n6914 & n14484 ) | ( n6914 & n14485 ) | ( n14484 & n14485 ) ;
  assign n14487 = ( ~n5103 & n10717 ) | ( ~n5103 & n14486 ) | ( n10717 & n14486 ) ;
  assign n14489 = n4487 ^ n2602 ^ n2112 ;
  assign n14490 = ~n5480 & n14489 ;
  assign n14491 = ~n4100 & n14490 ;
  assign n14488 = x236 & ~n4637 ;
  assign n14492 = n14491 ^ n14488 ^ 1'b0 ;
  assign n14493 = ( n14483 & n14487 ) | ( n14483 & n14492 ) | ( n14487 & n14492 ) ;
  assign n14494 = ( n2477 & ~n9870 ) | ( n2477 & n11820 ) | ( ~n9870 & n11820 ) ;
  assign n14495 = n2412 & n3349 ;
  assign n14496 = n14495 ^ n4055 ^ 1'b0 ;
  assign n14497 = n1702 & n5948 ;
  assign n14498 = n14497 ^ n10725 ^ n2398 ;
  assign n14499 = n13906 ^ n6263 ^ n4105 ;
  assign n14500 = ( n1537 & ~n9325 ) | ( n1537 & n14499 ) | ( ~n9325 & n14499 ) ;
  assign n14501 = n8969 ^ n5609 ^ n1435 ;
  assign n14502 = n14501 ^ n4267 ^ n3960 ;
  assign n14503 = n14502 ^ n4011 ^ n2962 ;
  assign n14504 = n12961 ^ n4237 ^ 1'b0 ;
  assign n14505 = x19 & n14504 ;
  assign n14506 = n14505 ^ n8166 ^ n1085 ;
  assign n14507 = ( n6076 & ~n10878 ) | ( n6076 & n14506 ) | ( ~n10878 & n14506 ) ;
  assign n14512 = ~n4426 & n12490 ;
  assign n14510 = n8248 ^ n5954 ^ n3112 ;
  assign n14511 = n14510 ^ n494 ^ 1'b0 ;
  assign n14508 = ( n965 & n2557 ) | ( n965 & ~n13401 ) | ( n2557 & ~n13401 ) ;
  assign n14509 = ( n10053 & ~n10814 ) | ( n10053 & n14508 ) | ( ~n10814 & n14508 ) ;
  assign n14513 = n14512 ^ n14511 ^ n14509 ;
  assign n14514 = ( ~n14503 & n14507 ) | ( ~n14503 & n14513 ) | ( n14507 & n14513 ) ;
  assign n14515 = n10629 ^ n1345 ^ x125 ;
  assign n14516 = ( ~n1755 & n2106 ) | ( ~n1755 & n5078 ) | ( n2106 & n5078 ) ;
  assign n14519 = ( n1605 & ~n1903 ) | ( n1605 & n2995 ) | ( ~n1903 & n2995 ) ;
  assign n14520 = ( n10781 & n13063 ) | ( n10781 & ~n14519 ) | ( n13063 & ~n14519 ) ;
  assign n14517 = n871 | n4435 ;
  assign n14518 = n14517 ^ n5287 ^ 1'b0 ;
  assign n14521 = n14520 ^ n14518 ^ n6728 ;
  assign n14522 = ( n2546 & ~n14516 ) | ( n2546 & n14521 ) | ( ~n14516 & n14521 ) ;
  assign n14526 = n868 | n1250 ;
  assign n14527 = x173 | n14526 ;
  assign n14528 = n14527 ^ n6774 ^ n5550 ;
  assign n14525 = n7635 ^ n4973 ^ n1383 ;
  assign n14523 = ( n828 & ~n2461 ) | ( n828 & n4941 ) | ( ~n2461 & n4941 ) ;
  assign n14524 = ( n6470 & ~n11413 ) | ( n6470 & n14523 ) | ( ~n11413 & n14523 ) ;
  assign n14529 = n14528 ^ n14525 ^ n14524 ;
  assign n14530 = ( n862 & ~n10189 ) | ( n862 & n13794 ) | ( ~n10189 & n13794 ) ;
  assign n14531 = n7124 ^ n5345 ^ 1'b0 ;
  assign n14532 = n2796 | n14531 ;
  assign n14533 = n11801 ^ n5719 ^ n1044 ;
  assign n14534 = ~n14532 & n14533 ;
  assign n14535 = n14530 & n14534 ;
  assign n14538 = n4863 ^ n1150 ^ x169 ;
  assign n14539 = ( n2993 & n3375 ) | ( n2993 & n8926 ) | ( n3375 & n8926 ) ;
  assign n14540 = n14539 ^ n5970 ^ n4767 ;
  assign n14541 = ( n686 & n14538 ) | ( n686 & ~n14540 ) | ( n14538 & ~n14540 ) ;
  assign n14542 = ( n2700 & ~n12881 ) | ( n2700 & n14541 ) | ( ~n12881 & n14541 ) ;
  assign n14536 = ( n1859 & ~n3534 ) | ( n1859 & n4658 ) | ( ~n3534 & n4658 ) ;
  assign n14537 = n14536 ^ n4663 ^ n2741 ;
  assign n14543 = n14542 ^ n14537 ^ 1'b0 ;
  assign n14544 = n12038 & ~n14543 ;
  assign n14545 = n14544 ^ n6599 ^ n5844 ;
  assign n14546 = n14545 ^ n10587 ^ n2817 ;
  assign n14547 = ( ~x38 & n1083 ) | ( ~x38 & n8321 ) | ( n1083 & n8321 ) ;
  assign n14548 = n14547 ^ n13837 ^ n971 ;
  assign n14549 = ( n914 & ~n1544 ) | ( n914 & n9035 ) | ( ~n1544 & n9035 ) ;
  assign n14550 = n12340 ^ n11270 ^ 1'b0 ;
  assign n14551 = n14549 | n14550 ;
  assign n14552 = n14551 ^ n7259 ^ 1'b0 ;
  assign n14553 = n5105 ^ n2126 ^ n369 ;
  assign n14554 = n14553 ^ n6463 ^ n5746 ;
  assign n14555 = ( n2967 & ~n4869 ) | ( n2967 & n14554 ) | ( ~n4869 & n14554 ) ;
  assign n14556 = ( ~n1088 & n10835 ) | ( ~n1088 & n14555 ) | ( n10835 & n14555 ) ;
  assign n14557 = n14556 ^ n10962 ^ n1903 ;
  assign n14558 = n11148 ^ n11110 ^ n6993 ;
  assign n14559 = n7545 ^ n5248 ^ 1'b0 ;
  assign n14560 = ( n12429 & ~n14558 ) | ( n12429 & n14559 ) | ( ~n14558 & n14559 ) ;
  assign n14561 = n14560 ^ n9042 ^ n2162 ;
  assign n14562 = n14561 ^ n9601 ^ n3175 ;
  assign n14563 = ( n1637 & n3069 ) | ( n1637 & n4611 ) | ( n3069 & n4611 ) ;
  assign n14564 = ( n648 & n13522 ) | ( n648 & ~n14563 ) | ( n13522 & ~n14563 ) ;
  assign n14565 = n3796 ^ n375 ^ n282 ;
  assign n14566 = ( n7101 & n8290 ) | ( n7101 & ~n14565 ) | ( n8290 & ~n14565 ) ;
  assign n14567 = ( n3737 & n4883 ) | ( n3737 & ~n14566 ) | ( n4883 & ~n14566 ) ;
  assign n14568 = ( ~n5798 & n14564 ) | ( ~n5798 & n14567 ) | ( n14564 & n14567 ) ;
  assign n14570 = ( n3786 & n4238 ) | ( n3786 & n7551 ) | ( n4238 & n7551 ) ;
  assign n14571 = ( n2389 & n3024 ) | ( n2389 & n14570 ) | ( n3024 & n14570 ) ;
  assign n14569 = n14554 ^ n3480 ^ n1771 ;
  assign n14572 = n14571 ^ n14569 ^ 1'b0 ;
  assign n14573 = ( n13774 & n14568 ) | ( n13774 & n14572 ) | ( n14568 & n14572 ) ;
  assign n14574 = n13736 ^ n3602 ^ n2785 ;
  assign n14575 = n11235 ^ n8226 ^ n2219 ;
  assign n14576 = ~n639 & n14575 ;
  assign n14577 = n11153 & n14576 ;
  assign n14578 = n7644 ^ n6798 ^ 1'b0 ;
  assign n14579 = n308 & n14578 ;
  assign n14580 = n14579 ^ n13353 ^ n5567 ;
  assign n14581 = n14352 ^ n14073 ^ n1476 ;
  assign n14582 = n12897 & ~n14581 ;
  assign n14583 = ~n11405 & n12788 ;
  assign n14593 = n11464 ^ n2054 ^ n266 ;
  assign n14592 = ( n5520 & n6663 ) | ( n5520 & ~n12295 ) | ( n6663 & ~n12295 ) ;
  assign n14589 = n3118 ^ n2761 ^ 1'b0 ;
  assign n14588 = n12184 ^ n7324 ^ n4217 ;
  assign n14584 = n5116 ^ n4227 ^ n2435 ;
  assign n14585 = n7274 & n14584 ;
  assign n14586 = n13830 & n14585 ;
  assign n14587 = n14586 ^ n7845 ^ 1'b0 ;
  assign n14590 = n14589 ^ n14588 ^ n14587 ;
  assign n14591 = ( ~n6584 & n13118 ) | ( ~n6584 & n14590 ) | ( n13118 & n14590 ) ;
  assign n14594 = n14593 ^ n14592 ^ n14591 ;
  assign n14595 = ( ~n11000 & n12822 ) | ( ~n11000 & n13210 ) | ( n12822 & n13210 ) ;
  assign n14596 = n14595 ^ n2363 ^ 1'b0 ;
  assign n14597 = ~n2164 & n14596 ;
  assign n14598 = ( x173 & n1321 ) | ( x173 & ~n4228 ) | ( n1321 & ~n4228 ) ;
  assign n14599 = ( n2439 & ~n4475 ) | ( n2439 & n14598 ) | ( ~n4475 & n14598 ) ;
  assign n14600 = n14599 ^ n7685 ^ 1'b0 ;
  assign n14601 = n14600 ^ n13538 ^ n2497 ;
  assign n14602 = n7476 ^ n6052 ^ n3632 ;
  assign n14603 = ( ~n683 & n5491 ) | ( ~n683 & n14602 ) | ( n5491 & n14602 ) ;
  assign n14604 = ( n1130 & n6172 ) | ( n1130 & ~n14178 ) | ( n6172 & ~n14178 ) ;
  assign n14605 = ( ~n4956 & n14603 ) | ( ~n4956 & n14604 ) | ( n14603 & n14604 ) ;
  assign n14606 = n2491 & n12139 ;
  assign n14607 = n2401 & n9632 ;
  assign n14608 = ( ~n562 & n2375 ) | ( ~n562 & n2815 ) | ( n2375 & n2815 ) ;
  assign n14609 = n10197 ^ n9304 ^ n4559 ;
  assign n14610 = n12516 & n14609 ;
  assign n14623 = n1672 | n5775 ;
  assign n14611 = n9593 ^ n9415 ^ n2801 ;
  assign n14617 = n9880 ^ n5545 ^ n2526 ;
  assign n14612 = n5739 ^ n3715 ^ n1476 ;
  assign n14613 = n14612 ^ n7182 ^ n1427 ;
  assign n14614 = n14613 ^ n8891 ^ n6941 ;
  assign n14615 = ( n1305 & n3716 ) | ( n1305 & ~n14614 ) | ( n3716 & ~n14614 ) ;
  assign n14616 = n14615 ^ n12465 ^ n7216 ;
  assign n14618 = n14617 ^ n14616 ^ n2703 ;
  assign n14619 = n12078 | n14618 ;
  assign n14620 = n14619 ^ n13803 ^ 1'b0 ;
  assign n14621 = n14620 ^ n1291 ^ 1'b0 ;
  assign n14622 = ~n14611 & n14621 ;
  assign n14624 = n14623 ^ n14622 ^ n6809 ;
  assign n14625 = ( ~n561 & n7045 ) | ( ~n561 & n11168 ) | ( n7045 & n11168 ) ;
  assign n14626 = n14625 ^ n13718 ^ n5393 ;
  assign n14627 = n13630 ^ n3014 ^ 1'b0 ;
  assign n14628 = n14627 ^ n7274 ^ n959 ;
  assign n14629 = n14628 ^ n13256 ^ n6588 ;
  assign n14630 = ~n2356 & n14094 ;
  assign n14631 = ( n965 & n14629 ) | ( n965 & n14630 ) | ( n14629 & n14630 ) ;
  assign n14632 = n10688 ^ n650 ^ n640 ;
  assign n14633 = n11027 ^ n6601 ^ n5784 ;
  assign n14634 = ( n10341 & n14632 ) | ( n10341 & ~n14633 ) | ( n14632 & ~n14633 ) ;
  assign n14635 = ( n3703 & ~n5005 ) | ( n3703 & n6906 ) | ( ~n5005 & n6906 ) ;
  assign n14636 = n14635 ^ n3518 ^ n2268 ;
  assign n14637 = n2458 & ~n11525 ;
  assign n14638 = ( n3894 & ~n5881 ) | ( n3894 & n7510 ) | ( ~n5881 & n7510 ) ;
  assign n14639 = ( ~n2620 & n8320 ) | ( ~n2620 & n14638 ) | ( n8320 & n14638 ) ;
  assign n14640 = n4520 ^ n1041 ^ 1'b0 ;
  assign n14641 = n4874 | n14640 ;
  assign n14642 = n5953 ^ n4670 ^ n562 ;
  assign n14643 = n13704 ^ n13477 ^ n13003 ;
  assign n14644 = ( n2148 & ~n12989 ) | ( n2148 & n14643 ) | ( ~n12989 & n14643 ) ;
  assign n14645 = n11308 ^ n457 ^ 1'b0 ;
  assign n14647 = ( n2609 & n3419 ) | ( n2609 & ~n7789 ) | ( n3419 & ~n7789 ) ;
  assign n14646 = n11211 ^ n3591 ^ n3272 ;
  assign n14648 = n14647 ^ n14646 ^ n14187 ;
  assign n14659 = ~n515 & n755 ;
  assign n14660 = n14659 ^ n7501 ^ n660 ;
  assign n14655 = n4487 | n7124 ;
  assign n14656 = n14655 ^ n6748 ^ 1'b0 ;
  assign n14649 = n7387 ^ n2776 ^ n428 ;
  assign n14650 = ( ~n3874 & n5619 ) | ( ~n3874 & n14649 ) | ( n5619 & n14649 ) ;
  assign n14651 = n8285 ^ n347 ^ 1'b0 ;
  assign n14652 = ( n3903 & n4968 ) | ( n3903 & n14651 ) | ( n4968 & n14651 ) ;
  assign n14653 = ( x29 & n8569 ) | ( x29 & n14652 ) | ( n8569 & n14652 ) ;
  assign n14654 = ( n1657 & n14650 ) | ( n1657 & n14653 ) | ( n14650 & n14653 ) ;
  assign n14657 = n14656 ^ n14654 ^ n7793 ;
  assign n14658 = n14657 ^ n9493 ^ n7536 ;
  assign n14661 = n14660 ^ n14658 ^ 1'b0 ;
  assign n14662 = ~n5237 & n9934 ;
  assign n14667 = n8900 ^ n5543 ^ 1'b0 ;
  assign n14668 = n13388 & n14667 ;
  assign n14666 = n8168 ^ n7927 ^ n4000 ;
  assign n14663 = n4377 ^ n1062 ^ 1'b0 ;
  assign n14664 = n6804 & ~n7558 ;
  assign n14665 = ( n1584 & ~n14663 ) | ( n1584 & n14664 ) | ( ~n14663 & n14664 ) ;
  assign n14669 = n14668 ^ n14666 ^ n14665 ;
  assign n14675 = ~n7936 & n8297 ;
  assign n14676 = n14675 ^ n9053 ^ n3737 ;
  assign n14673 = n9928 ^ n9052 ^ n7888 ;
  assign n14672 = ( ~n1919 & n6759 ) | ( ~n1919 & n8265 ) | ( n6759 & n8265 ) ;
  assign n14674 = n14673 ^ n14672 ^ x223 ;
  assign n14670 = n5259 ^ n5156 ^ n3373 ;
  assign n14671 = n14670 ^ n8994 ^ n5135 ;
  assign n14677 = n14676 ^ n14674 ^ n14671 ;
  assign n14678 = ( n14662 & n14669 ) | ( n14662 & n14677 ) | ( n14669 & n14677 ) ;
  assign n14681 = ~n900 & n4855 ;
  assign n14679 = n7680 ^ n5521 ^ n1254 ;
  assign n14680 = ( ~n6778 & n7459 ) | ( ~n6778 & n14679 ) | ( n7459 & n14679 ) ;
  assign n14682 = n14681 ^ n14680 ^ n2146 ;
  assign n14683 = n14682 ^ n14079 ^ n9425 ;
  assign n14684 = n12344 ^ n10190 ^ n476 ;
  assign n14685 = ( ~n4515 & n5105 ) | ( ~n4515 & n14684 ) | ( n5105 & n14684 ) ;
  assign n14686 = ( n11598 & n14683 ) | ( n11598 & n14685 ) | ( n14683 & n14685 ) ;
  assign n14688 = n2389 | n7473 ;
  assign n14689 = n5173 & ~n14688 ;
  assign n14690 = n9081 ^ n8767 ^ 1'b0 ;
  assign n14691 = n14689 | n14690 ;
  assign n14692 = n13186 & ~n14691 ;
  assign n14687 = ( x24 & n901 ) | ( x24 & ~n11800 ) | ( n901 & ~n11800 ) ;
  assign n14693 = n14692 ^ n14687 ^ n6035 ;
  assign n14694 = ( ~n5905 & n8681 ) | ( ~n5905 & n12888 ) | ( n8681 & n12888 ) ;
  assign n14695 = n7258 & ~n10209 ;
  assign n14696 = n14695 ^ n12517 ^ n4816 ;
  assign n14699 = n6133 ^ n2653 ^ n1561 ;
  assign n14697 = n12028 ^ n11200 ^ n5262 ;
  assign n14698 = n14697 ^ n3247 ^ n2217 ;
  assign n14700 = n14699 ^ n14698 ^ n6313 ;
  assign n14701 = n6459 & ~n14700 ;
  assign n14702 = ~n14544 & n14701 ;
  assign n14703 = n11487 ^ n10663 ^ n5964 ;
  assign n14707 = ( n521 & n2889 ) | ( n521 & n6957 ) | ( n2889 & n6957 ) ;
  assign n14704 = n7710 ^ n2222 ^ n1356 ;
  assign n14705 = ( n428 & n4888 ) | ( n428 & n14704 ) | ( n4888 & n14704 ) ;
  assign n14706 = n6561 & ~n14705 ;
  assign n14708 = n14707 ^ n14706 ^ n962 ;
  assign n14709 = n9924 ^ n9537 ^ 1'b0 ;
  assign n14710 = n14708 & ~n14709 ;
  assign n14711 = n13669 ^ n10907 ^ n1750 ;
  assign n14712 = ( ~n6326 & n10281 ) | ( ~n6326 & n14711 ) | ( n10281 & n14711 ) ;
  assign n14713 = ( n5218 & n5321 ) | ( n5218 & n14712 ) | ( n5321 & n14712 ) ;
  assign n14714 = n8596 ^ n1194 ^ 1'b0 ;
  assign n14717 = ( n1030 & ~n4593 ) | ( n1030 & n8222 ) | ( ~n4593 & n8222 ) ;
  assign n14715 = ( n1380 & n3186 ) | ( n1380 & ~n5089 ) | ( n3186 & ~n5089 ) ;
  assign n14716 = ( n5104 & n13904 ) | ( n5104 & n14715 ) | ( n13904 & n14715 ) ;
  assign n14718 = n14717 ^ n14716 ^ n13763 ;
  assign n14719 = ( n320 & n6502 ) | ( n320 & n14356 ) | ( n6502 & n14356 ) ;
  assign n14720 = n14719 ^ n8068 ^ n726 ;
  assign n14721 = n14720 ^ n7260 ^ n6312 ;
  assign n14722 = ( n2072 & n5681 ) | ( n2072 & ~n7392 ) | ( n5681 & ~n7392 ) ;
  assign n14723 = ( n518 & n705 ) | ( n518 & ~n2367 ) | ( n705 & ~n2367 ) ;
  assign n14724 = ( n5511 & ~n5636 ) | ( n5511 & n14723 ) | ( ~n5636 & n14723 ) ;
  assign n14725 = ( ~n271 & n5321 ) | ( ~n271 & n14724 ) | ( n5321 & n14724 ) ;
  assign n14726 = ( n2807 & n10378 ) | ( n2807 & n14725 ) | ( n10378 & n14725 ) ;
  assign n14730 = ( ~n4010 & n8676 ) | ( ~n4010 & n12812 ) | ( n8676 & n12812 ) ;
  assign n14731 = ( ~n411 & n4959 ) | ( ~n411 & n14730 ) | ( n4959 & n14730 ) ;
  assign n14732 = ( n2889 & n8593 ) | ( n2889 & ~n11254 ) | ( n8593 & ~n11254 ) ;
  assign n14733 = ( n9817 & n14431 ) | ( n9817 & n14732 ) | ( n14431 & n14732 ) ;
  assign n14734 = ( n9359 & n14731 ) | ( n9359 & n14733 ) | ( n14731 & n14733 ) ;
  assign n14727 = ( n3700 & n4350 ) | ( n3700 & ~n12717 ) | ( n4350 & ~n12717 ) ;
  assign n14728 = n14727 ^ n13282 ^ n305 ;
  assign n14729 = ( n3079 & n3806 ) | ( n3079 & n14728 ) | ( n3806 & n14728 ) ;
  assign n14735 = n14734 ^ n14729 ^ n9577 ;
  assign n14736 = ( ~n9544 & n14726 ) | ( ~n9544 & n14735 ) | ( n14726 & n14735 ) ;
  assign n14737 = ( n5893 & n14722 ) | ( n5893 & n14736 ) | ( n14722 & n14736 ) ;
  assign n14738 = ( n6121 & ~n7329 ) | ( n6121 & n8921 ) | ( ~n7329 & n8921 ) ;
  assign n14742 = n6237 ^ n3596 ^ n3224 ;
  assign n14739 = ( n1534 & n1799 ) | ( n1534 & n3329 ) | ( n1799 & n3329 ) ;
  assign n14740 = ( n6425 & n8574 ) | ( n6425 & n14739 ) | ( n8574 & n14739 ) ;
  assign n14741 = n14740 ^ n6087 ^ n2500 ;
  assign n14743 = n14742 ^ n14741 ^ n600 ;
  assign n14744 = ( n1790 & n9661 ) | ( n1790 & n14743 ) | ( n9661 & n14743 ) ;
  assign n14745 = ( n3247 & ~n9357 ) | ( n3247 & n14744 ) | ( ~n9357 & n14744 ) ;
  assign n14746 = ( n11636 & ~n14738 ) | ( n11636 & n14745 ) | ( ~n14738 & n14745 ) ;
  assign n14747 = ~n12896 & n14746 ;
  assign n14748 = n12274 ^ n10877 ^ n9847 ;
  assign n14749 = ( n1042 & ~n1806 ) | ( n1042 & n14748 ) | ( ~n1806 & n14748 ) ;
  assign n14750 = n14749 ^ n13127 ^ n5965 ;
  assign n14752 = ( ~n3345 & n6266 ) | ( ~n3345 & n12590 ) | ( n6266 & n12590 ) ;
  assign n14751 = n2905 ^ x125 ^ x49 ;
  assign n14753 = n14752 ^ n14751 ^ n1424 ;
  assign n14754 = ( ~x45 & n11449 ) | ( ~x45 & n14753 ) | ( n11449 & n14753 ) ;
  assign n14755 = ( ~n3148 & n4952 ) | ( ~n3148 & n9492 ) | ( n4952 & n9492 ) ;
  assign n14757 = n2681 & n7078 ;
  assign n14758 = n14757 ^ n6512 ^ 1'b0 ;
  assign n14756 = ( n4566 & ~n7609 ) | ( n4566 & n14302 ) | ( ~n7609 & n14302 ) ;
  assign n14759 = n14758 ^ n14756 ^ n1006 ;
  assign n14760 = ( n2667 & ~n9059 ) | ( n2667 & n10247 ) | ( ~n9059 & n10247 ) ;
  assign n14761 = ( n2289 & n13119 ) | ( n2289 & n14566 ) | ( n13119 & n14566 ) ;
  assign n14762 = n14761 ^ n13799 ^ n13116 ;
  assign n14766 = ( n338 & n722 ) | ( n338 & n2616 ) | ( n722 & n2616 ) ;
  assign n14767 = n8728 & n14766 ;
  assign n14763 = n900 | n14122 ;
  assign n14764 = n14763 ^ n11124 ^ n9958 ;
  assign n14765 = n14764 ^ n14763 ^ n14278 ;
  assign n14768 = n14767 ^ n14765 ^ 1'b0 ;
  assign n14769 = ( n2221 & n6804 ) | ( n2221 & n11557 ) | ( n6804 & n11557 ) ;
  assign n14770 = n14769 ^ n7865 ^ n1939 ;
  assign n14771 = ( x182 & n1327 ) | ( x182 & ~n14770 ) | ( n1327 & ~n14770 ) ;
  assign n14772 = ( ~n9270 & n14768 ) | ( ~n9270 & n14771 ) | ( n14768 & n14771 ) ;
  assign n14773 = n3608 & n8407 ;
  assign n14774 = n14773 ^ n1288 ^ 1'b0 ;
  assign n14775 = n14774 ^ n11963 ^ n5738 ;
  assign n14778 = n1716 ^ n304 ^ 1'b0 ;
  assign n14779 = n7906 ^ n3554 ^ n1612 ;
  assign n14780 = ( n12834 & n14778 ) | ( n12834 & n14779 ) | ( n14778 & n14779 ) ;
  assign n14776 = n2509 & n4654 ;
  assign n14777 = ~n14127 & n14776 ;
  assign n14781 = n14780 ^ n14777 ^ 1'b0 ;
  assign n14782 = n478 & ~n2492 ;
  assign n14783 = n6482 & n14782 ;
  assign n14784 = n13888 ^ n389 ^ 1'b0 ;
  assign n14785 = ( n9690 & n14783 ) | ( n9690 & ~n14784 ) | ( n14783 & ~n14784 ) ;
  assign n14786 = n14785 ^ n14332 ^ n8747 ;
  assign n14787 = n1946 ^ n1392 ^ n889 ;
  assign n14788 = ( n3932 & n7214 ) | ( n3932 & n14787 ) | ( n7214 & n14787 ) ;
  assign n14789 = n10428 ^ n4319 ^ 1'b0 ;
  assign n14790 = n6091 | n14789 ;
  assign n14791 = ( n2136 & ~n10629 ) | ( n2136 & n14790 ) | ( ~n10629 & n14790 ) ;
  assign n14792 = ( n9608 & n14788 ) | ( n9608 & ~n14791 ) | ( n14788 & ~n14791 ) ;
  assign n14793 = ( ~n3976 & n8385 ) | ( ~n3976 & n12245 ) | ( n8385 & n12245 ) ;
  assign n14794 = ( n1599 & n6127 ) | ( n1599 & n9277 ) | ( n6127 & n9277 ) ;
  assign n14795 = n14793 & ~n14794 ;
  assign n14796 = ~n3538 & n14795 ;
  assign n14797 = n14796 ^ n272 ^ 1'b0 ;
  assign n14798 = ( n5903 & n7610 ) | ( n5903 & ~n14797 ) | ( n7610 & ~n14797 ) ;
  assign n14799 = n5686 ^ n1419 ^ n523 ;
  assign n14800 = n10554 ^ n3100 ^ 1'b0 ;
  assign n14801 = n14799 & n14800 ;
  assign n14807 = n4873 ^ n2657 ^ x239 ;
  assign n14808 = ~n6240 & n14807 ;
  assign n14802 = ( n1011 & ~n1926 ) | ( n1011 & n3000 ) | ( ~n1926 & n3000 ) ;
  assign n14803 = n4851 & ~n7784 ;
  assign n14804 = n7072 ^ n5567 ^ n3648 ;
  assign n14805 = ( n4047 & ~n14803 ) | ( n4047 & n14804 ) | ( ~n14803 & n14804 ) ;
  assign n14806 = ( n14322 & ~n14802 ) | ( n14322 & n14805 ) | ( ~n14802 & n14805 ) ;
  assign n14809 = n14808 ^ n14806 ^ n14102 ;
  assign n14810 = ( ~n327 & n2976 ) | ( ~n327 & n4320 ) | ( n2976 & n4320 ) ;
  assign n14811 = n11614 ^ n3503 ^ n2699 ;
  assign n14813 = ( n4606 & n6686 ) | ( n4606 & ~n7051 ) | ( n6686 & ~n7051 ) ;
  assign n14812 = n258 & n8053 ;
  assign n14814 = n14813 ^ n14812 ^ 1'b0 ;
  assign n14815 = n1422 & n10377 ;
  assign n14816 = ~n7442 & n14815 ;
  assign n14817 = ( n4147 & n14787 ) | ( n4147 & n14816 ) | ( n14787 & n14816 ) ;
  assign n14818 = n5082 ^ n4935 ^ n3260 ;
  assign n14819 = ~n11714 & n14818 ;
  assign n14820 = ( n5964 & n7100 ) | ( n5964 & ~n14819 ) | ( n7100 & ~n14819 ) ;
  assign n14821 = ( n14814 & n14817 ) | ( n14814 & n14820 ) | ( n14817 & n14820 ) ;
  assign n14822 = ( n11099 & n14811 ) | ( n11099 & n14821 ) | ( n14811 & n14821 ) ;
  assign n14823 = n14822 ^ n9716 ^ n3268 ;
  assign n14824 = n8666 ^ n5047 ^ n3120 ;
  assign n14825 = n7749 ^ n2498 ^ n2100 ;
  assign n14826 = n14824 & n14825 ;
  assign n14827 = ~n1470 & n12868 ;
  assign n14828 = n14826 & n14827 ;
  assign n14829 = n738 & ~n10158 ;
  assign n14830 = ( n917 & n3302 ) | ( n917 & ~n14829 ) | ( n3302 & ~n14829 ) ;
  assign n14831 = ( n3980 & n5575 ) | ( n3980 & n6315 ) | ( n5575 & n6315 ) ;
  assign n14832 = n4446 | n10528 ;
  assign n14833 = n10262 | n14832 ;
  assign n14834 = ( n1963 & n5689 ) | ( n1963 & n14833 ) | ( n5689 & n14833 ) ;
  assign n14835 = n14834 ^ n13545 ^ n9008 ;
  assign n14836 = n13384 ^ n2822 ^ n916 ;
  assign n14837 = n14836 ^ n8598 ^ n7557 ;
  assign n14838 = ( n7649 & ~n14835 ) | ( n7649 & n14837 ) | ( ~n14835 & n14837 ) ;
  assign n14839 = n4034 ^ x193 ^ 1'b0 ;
  assign n14840 = n14839 ^ n7540 ^ n396 ;
  assign n14841 = n14840 ^ n13903 ^ n4964 ;
  assign n14842 = n4120 ^ n3260 ^ 1'b0 ;
  assign n14843 = n14842 ^ n5223 ^ n4557 ;
  assign n14844 = ( ~n4931 & n10217 ) | ( ~n4931 & n14843 ) | ( n10217 & n14843 ) ;
  assign n14845 = n14844 ^ n12306 ^ x26 ;
  assign n14853 = n9266 ^ n7825 ^ n1644 ;
  assign n14854 = ( ~n5226 & n10720 ) | ( ~n5226 & n14853 ) | ( n10720 & n14853 ) ;
  assign n14850 = n14155 ^ n4018 ^ 1'b0 ;
  assign n14851 = ~n14233 & n14850 ;
  assign n14848 = n5115 ^ n2138 ^ n1740 ;
  assign n14846 = n7633 ^ n3051 ^ n578 ;
  assign n14847 = n8783 & ~n14846 ;
  assign n14849 = n14848 ^ n14847 ^ n1498 ;
  assign n14852 = n14851 ^ n14849 ^ n13733 ;
  assign n14855 = n14854 ^ n14852 ^ n1207 ;
  assign n14859 = ( n5973 & n8742 ) | ( n5973 & n11673 ) | ( n8742 & n11673 ) ;
  assign n14856 = n8772 & n13526 ;
  assign n14857 = ~n4890 & n9897 ;
  assign n14858 = ( n14730 & ~n14856 ) | ( n14730 & n14857 ) | ( ~n14856 & n14857 ) ;
  assign n14860 = n14859 ^ n14858 ^ n6912 ;
  assign n14861 = ( n1655 & ~n2963 ) | ( n1655 & n12042 ) | ( ~n2963 & n12042 ) ;
  assign n14862 = ( n4656 & n7025 ) | ( n4656 & ~n14861 ) | ( n7025 & ~n14861 ) ;
  assign n14863 = ( ~n9775 & n10142 ) | ( ~n9775 & n14862 ) | ( n10142 & n14862 ) ;
  assign n14864 = n6135 ^ n3118 ^ n2127 ;
  assign n14865 = n14864 ^ n520 ^ x41 ;
  assign n14866 = n5370 ^ n1012 ^ 1'b0 ;
  assign n14867 = n470 & n4316 ;
  assign n14868 = n14867 ^ n11928 ^ n4206 ;
  assign n14869 = n14868 ^ n3720 ^ 1'b0 ;
  assign n14870 = ~n11365 & n14869 ;
  assign n14871 = ~n321 & n14870 ;
  assign n14872 = ( n5416 & n14866 ) | ( n5416 & ~n14871 ) | ( n14866 & ~n14871 ) ;
  assign n14873 = ( ~n7288 & n9278 ) | ( ~n7288 & n11605 ) | ( n9278 & n11605 ) ;
  assign n14874 = n14873 ^ n4090 ^ n369 ;
  assign n14875 = ( n2754 & ~n2932 ) | ( n2754 & n14874 ) | ( ~n2932 & n14874 ) ;
  assign n14876 = ( n8474 & n13314 ) | ( n8474 & n14875 ) | ( n13314 & n14875 ) ;
  assign n14877 = n14876 ^ n11615 ^ 1'b0 ;
  assign n14878 = ( ~n2832 & n5535 ) | ( ~n2832 & n12342 ) | ( n5535 & n12342 ) ;
  assign n14879 = ( n2871 & ~n4663 ) | ( n2871 & n14878 ) | ( ~n4663 & n14878 ) ;
  assign n14880 = n14879 ^ n14560 ^ 1'b0 ;
  assign n14882 = n6318 ^ n2417 ^ n2416 ;
  assign n14883 = n14882 ^ n6905 ^ n6028 ;
  assign n14881 = n3729 & n5763 ;
  assign n14884 = n14883 ^ n14881 ^ 1'b0 ;
  assign n14885 = ( n1915 & n5594 ) | ( n1915 & n10807 ) | ( n5594 & n10807 ) ;
  assign n14886 = ( n3462 & n5528 ) | ( n3462 & n14885 ) | ( n5528 & n14885 ) ;
  assign n14887 = ( n6713 & ~n14884 ) | ( n6713 & n14886 ) | ( ~n14884 & n14886 ) ;
  assign n14888 = n14887 ^ n11546 ^ n3934 ;
  assign n14889 = n13300 ^ n4511 ^ n3862 ;
  assign n14890 = ( ~n4389 & n6155 ) | ( ~n4389 & n11853 ) | ( n6155 & n11853 ) ;
  assign n14891 = ( n2792 & n7857 ) | ( n2792 & n12652 ) | ( n7857 & n12652 ) ;
  assign n14892 = n14891 ^ n6255 ^ n3928 ;
  assign n14893 = ( n14889 & n14890 ) | ( n14889 & ~n14892 ) | ( n14890 & ~n14892 ) ;
  assign n14895 = ( n4751 & ~n8109 ) | ( n4751 & n13186 ) | ( ~n8109 & n13186 ) ;
  assign n14894 = x249 & n13567 ;
  assign n14896 = n14895 ^ n14894 ^ n1939 ;
  assign n14897 = n8323 & ~n14896 ;
  assign n14898 = ( n12489 & ~n13619 ) | ( n12489 & n14897 ) | ( ~n13619 & n14897 ) ;
  assign n14900 = ( ~n2456 & n4439 ) | ( ~n2456 & n7319 ) | ( n4439 & n7319 ) ;
  assign n14899 = n13422 ^ n12946 ^ n3600 ;
  assign n14901 = n14900 ^ n14899 ^ n7414 ;
  assign n14902 = n2004 | n14901 ;
  assign n14903 = n2379 ^ n1591 ^ n774 ;
  assign n14905 = n13152 ^ n7959 ^ n2694 ;
  assign n14904 = n10396 ^ n6726 ^ 1'b0 ;
  assign n14906 = n14905 ^ n14904 ^ 1'b0 ;
  assign n14907 = n14903 & n14906 ;
  assign n14908 = n14907 ^ n9779 ^ 1'b0 ;
  assign n14909 = n14902 | n14908 ;
  assign n14910 = n14909 ^ n13892 ^ n7459 ;
  assign n14912 = n3092 & n8188 ;
  assign n14913 = n14912 ^ n6301 ^ 1'b0 ;
  assign n14914 = n14913 ^ n12766 ^ n1033 ;
  assign n14911 = n4462 & n6849 ;
  assign n14915 = n14914 ^ n14911 ^ 1'b0 ;
  assign n14916 = n6057 & n12984 ;
  assign n14917 = n14916 ^ n10925 ^ 1'b0 ;
  assign n14918 = ( ~n4814 & n9471 ) | ( ~n4814 & n14917 ) | ( n9471 & n14917 ) ;
  assign n14919 = ( ~n2705 & n7294 ) | ( ~n2705 & n9880 ) | ( n7294 & n9880 ) ;
  assign n14926 = ( n2608 & ~n5419 ) | ( n2608 & n7518 ) | ( ~n5419 & n7518 ) ;
  assign n14923 = n4662 & ~n7080 ;
  assign n14924 = n14923 ^ n2539 ^ 1'b0 ;
  assign n14925 = n14924 ^ n5356 ^ x242 ;
  assign n14920 = ( n1727 & ~n2148 ) | ( n1727 & n6362 ) | ( ~n2148 & n6362 ) ;
  assign n14921 = n14920 ^ n7444 ^ n468 ;
  assign n14922 = ( n4478 & n7908 ) | ( n4478 & n14921 ) | ( n7908 & n14921 ) ;
  assign n14927 = n14926 ^ n14925 ^ n14922 ;
  assign n14928 = ( n12944 & ~n14919 ) | ( n12944 & n14927 ) | ( ~n14919 & n14927 ) ;
  assign n14929 = n10621 ^ n1869 ^ 1'b0 ;
  assign n14930 = n5442 & n14929 ;
  assign n14931 = n14930 ^ n6704 ^ 1'b0 ;
  assign n14932 = n3100 ^ n2747 ^ x172 ;
  assign n14933 = n333 & n9635 ;
  assign n14934 = ( n10583 & n13192 ) | ( n10583 & n14933 ) | ( n13192 & n14933 ) ;
  assign n14937 = ~n2945 & n5272 ;
  assign n14936 = n14174 ^ n9384 ^ n6565 ;
  assign n14935 = n11094 ^ n11018 ^ n1155 ;
  assign n14938 = n14937 ^ n14936 ^ n14935 ;
  assign n14954 = ( n310 & n3607 ) | ( n310 & ~n6628 ) | ( n3607 & ~n6628 ) ;
  assign n14955 = n14954 ^ n2681 ^ n1714 ;
  assign n14950 = n3621 ^ n2616 ^ x123 ;
  assign n14951 = n2186 & ~n2290 ;
  assign n14952 = ~n4234 & n14951 ;
  assign n14953 = ( ~n3495 & n14950 ) | ( ~n3495 & n14952 ) | ( n14950 & n14952 ) ;
  assign n14939 = ~n3841 & n4943 ;
  assign n14940 = ( x229 & n1018 ) | ( x229 & n2065 ) | ( n1018 & n2065 ) ;
  assign n14941 = ( n738 & ~n1446 ) | ( n738 & n6352 ) | ( ~n1446 & n6352 ) ;
  assign n14942 = ( n3723 & ~n14317 ) | ( n3723 & n14941 ) | ( ~n14317 & n14941 ) ;
  assign n14943 = ( n14939 & n14940 ) | ( n14939 & ~n14942 ) | ( n14940 & ~n14942 ) ;
  assign n14944 = ( n6044 & n9569 ) | ( n6044 & ~n14943 ) | ( n9569 & ~n14943 ) ;
  assign n14945 = n11178 ^ n3935 ^ 1'b0 ;
  assign n14946 = n14945 ^ n7990 ^ n7112 ;
  assign n14947 = n10568 ^ n8592 ^ n1078 ;
  assign n14948 = ( ~n4774 & n14946 ) | ( ~n4774 & n14947 ) | ( n14946 & n14947 ) ;
  assign n14949 = ( n6158 & ~n14944 ) | ( n6158 & n14948 ) | ( ~n14944 & n14948 ) ;
  assign n14956 = n14955 ^ n14953 ^ n14949 ;
  assign n14957 = ( n868 & ~n1861 ) | ( n868 & n9511 ) | ( ~n1861 & n9511 ) ;
  assign n14958 = n14957 ^ n8398 ^ 1'b0 ;
  assign n14960 = n6050 ^ n3757 ^ n804 ;
  assign n14961 = n14960 ^ n6138 ^ n3243 ;
  assign n14959 = n1994 & n7461 ;
  assign n14962 = n14961 ^ n14959 ^ 1'b0 ;
  assign n14984 = n2787 & ~n8620 ;
  assign n14985 = ( n2364 & n3672 ) | ( n2364 & n14984 ) | ( n3672 & n14984 ) ;
  assign n14983 = n5894 ^ n4903 ^ n4467 ;
  assign n14963 = n11915 ^ n2485 ^ 1'b0 ;
  assign n14964 = n12219 & n14963 ;
  assign n14965 = n475 | n2257 ;
  assign n14966 = ( n622 & n3173 ) | ( n622 & n14965 ) | ( n3173 & n14965 ) ;
  assign n14970 = ( n709 & ~n6200 ) | ( n709 & n8335 ) | ( ~n6200 & n8335 ) ;
  assign n14971 = n2820 | n14970 ;
  assign n14972 = n14971 ^ n5911 ^ 1'b0 ;
  assign n14973 = n14972 ^ n6589 ^ n719 ;
  assign n14974 = ( n4366 & n5774 ) | ( n4366 & ~n7188 ) | ( n5774 & ~n7188 ) ;
  assign n14975 = ( n7390 & ~n14973 ) | ( n7390 & n14974 ) | ( ~n14973 & n14974 ) ;
  assign n14976 = n14975 ^ n5804 ^ n931 ;
  assign n14967 = n5474 ^ n3151 ^ n2459 ;
  assign n14968 = ( n1505 & n7077 ) | ( n1505 & ~n14967 ) | ( n7077 & ~n14967 ) ;
  assign n14969 = n5042 | n14968 ;
  assign n14977 = n14976 ^ n14969 ^ 1'b0 ;
  assign n14978 = ~n4522 & n12555 ;
  assign n14979 = ( ~n14966 & n14977 ) | ( ~n14966 & n14978 ) | ( n14977 & n14978 ) ;
  assign n14980 = n14979 ^ n12528 ^ n682 ;
  assign n14981 = n14980 ^ n11504 ^ 1'b0 ;
  assign n14982 = n14964 & ~n14981 ;
  assign n14986 = n14985 ^ n14983 ^ n14982 ;
  assign n14987 = n11070 ^ n7367 ^ 1'b0 ;
  assign n14988 = n14987 ^ n9790 ^ n7667 ;
  assign n14989 = n9060 | n12476 ;
  assign n14990 = n4729 & n14989 ;
  assign n14991 = n14990 ^ n2168 ^ 1'b0 ;
  assign n14992 = n14991 ^ n12510 ^ n4643 ;
  assign n14993 = n13084 ^ n9803 ^ n4097 ;
  assign n14994 = n14993 ^ n11555 ^ n7699 ;
  assign n14995 = n5803 | n14994 ;
  assign n14996 = n14995 ^ n9292 ^ 1'b0 ;
  assign n14997 = n12781 ^ n6994 ^ n306 ;
  assign n14998 = ( ~n4102 & n12512 ) | ( ~n4102 & n14262 ) | ( n12512 & n14262 ) ;
  assign n14999 = ( n7319 & ~n14997 ) | ( n7319 & n14998 ) | ( ~n14997 & n14998 ) ;
  assign n15004 = ~n532 & n2224 ;
  assign n15001 = ( n1108 & n2179 ) | ( n1108 & n5175 ) | ( n2179 & n5175 ) ;
  assign n15002 = n15001 ^ n8431 ^ n5521 ;
  assign n15003 = ( n720 & n6633 ) | ( n720 & n15002 ) | ( n6633 & n15002 ) ;
  assign n15000 = n12673 ^ n10094 ^ n1357 ;
  assign n15005 = n15004 ^ n15003 ^ n15000 ;
  assign n15006 = n2506 ^ n2115 ^ n1781 ;
  assign n15007 = ( n713 & n7982 ) | ( n713 & ~n15006 ) | ( n7982 & ~n15006 ) ;
  assign n15008 = ~n1658 & n15007 ;
  assign n15009 = n12913 ^ n9459 ^ n8265 ;
  assign n15010 = n13293 ^ n8818 ^ n5343 ;
  assign n15011 = n10401 ^ n10312 ^ 1'b0 ;
  assign n15012 = ( n3134 & n15010 ) | ( n3134 & ~n15011 ) | ( n15010 & ~n15011 ) ;
  assign n15013 = n11110 ^ n8935 ^ n4367 ;
  assign n15014 = ( ~n277 & n3069 ) | ( ~n277 & n6010 ) | ( n3069 & n6010 ) ;
  assign n15015 = n15014 ^ n4959 ^ n3813 ;
  assign n15016 = ( n8761 & n13512 ) | ( n8761 & ~n14883 ) | ( n13512 & ~n14883 ) ;
  assign n15017 = n15016 ^ n2815 ^ 1'b0 ;
  assign n15018 = ~n15015 & n15017 ;
  assign n15019 = n15013 & n15018 ;
  assign n15020 = ( n3713 & n5727 ) | ( n3713 & n13288 ) | ( n5727 & n13288 ) ;
  assign n15021 = ( ~n2781 & n7565 ) | ( ~n2781 & n15020 ) | ( n7565 & n15020 ) ;
  assign n15022 = n8031 ^ n4944 ^ n4136 ;
  assign n15023 = ( n7912 & n13529 ) | ( n7912 & ~n15022 ) | ( n13529 & ~n15022 ) ;
  assign n15024 = n12973 ^ n8536 ^ n595 ;
  assign n15025 = n3793 | n9270 ;
  assign n15026 = n5932 | n15025 ;
  assign n15027 = ( ~n6745 & n15024 ) | ( ~n6745 & n15026 ) | ( n15024 & n15026 ) ;
  assign n15028 = n8858 ^ n5802 ^ n3206 ;
  assign n15029 = ( n4448 & n11500 ) | ( n4448 & n15028 ) | ( n11500 & n15028 ) ;
  assign n15036 = ( x48 & n5864 ) | ( x48 & ~n7423 ) | ( n5864 & ~n7423 ) ;
  assign n15033 = n3627 & ~n3872 ;
  assign n15034 = n15033 ^ n2682 ^ 1'b0 ;
  assign n15030 = ( n914 & n1425 ) | ( n914 & ~n12611 ) | ( n1425 & ~n12611 ) ;
  assign n15031 = ( n1983 & n2463 ) | ( n1983 & n15030 ) | ( n2463 & n15030 ) ;
  assign n15032 = n15031 ^ n1813 ^ n693 ;
  assign n15035 = n15034 ^ n15032 ^ x229 ;
  assign n15037 = n15036 ^ n15035 ^ n9987 ;
  assign n15038 = n15037 ^ n13765 ^ n13727 ;
  assign n15039 = n15038 ^ n1396 ^ 1'b0 ;
  assign n15040 = n15029 & n15039 ;
  assign n15041 = ( ~n4141 & n6884 ) | ( ~n4141 & n15040 ) | ( n6884 & n15040 ) ;
  assign n15042 = n15041 ^ n12261 ^ 1'b0 ;
  assign n15043 = n788 | n15042 ;
  assign n15044 = n14018 ^ n12279 ^ n646 ;
  assign n15045 = ( ~n7411 & n10560 ) | ( ~n7411 & n15044 ) | ( n10560 & n15044 ) ;
  assign n15050 = n1392 ^ n869 ^ 1'b0 ;
  assign n15048 = ( ~n480 & n1089 ) | ( ~n480 & n8842 ) | ( n1089 & n8842 ) ;
  assign n15049 = ( n1960 & ~n12520 ) | ( n1960 & n15048 ) | ( ~n12520 & n15048 ) ;
  assign n15051 = n15050 ^ n15049 ^ n7399 ;
  assign n15046 = n4981 ^ n4788 ^ n312 ;
  assign n15047 = n3376 & ~n15046 ;
  assign n15052 = n15051 ^ n15047 ^ n14594 ;
  assign n15057 = n2185 ^ n1619 ^ x159 ;
  assign n15058 = n15057 ^ n5944 ^ n2367 ;
  assign n15059 = ( n4668 & ~n7817 ) | ( n4668 & n15058 ) | ( ~n7817 & n15058 ) ;
  assign n15060 = n15059 ^ n2821 ^ n2052 ;
  assign n15056 = n13992 ^ n2601 ^ n1439 ;
  assign n15053 = ( n368 & n2984 ) | ( n368 & ~n3036 ) | ( n2984 & ~n3036 ) ;
  assign n15054 = ~n8018 & n15053 ;
  assign n15055 = n15054 ^ n3125 ^ 1'b0 ;
  assign n15061 = n15060 ^ n15056 ^ n15055 ;
  assign n15062 = n4772 ^ n3561 ^ n2700 ;
  assign n15063 = n15062 ^ n8214 ^ n1631 ;
  assign n15064 = n3352 & n4273 ;
  assign n15065 = n15064 ^ n10454 ^ n4266 ;
  assign n15066 = n15065 ^ n6497 ^ 1'b0 ;
  assign n15067 = ~n1533 & n15066 ;
  assign n15068 = ( ~n1838 & n7688 ) | ( ~n1838 & n15067 ) | ( n7688 & n15067 ) ;
  assign n15069 = ( ~n601 & n15063 ) | ( ~n601 & n15068 ) | ( n15063 & n15068 ) ;
  assign n15070 = ( n2082 & n9958 ) | ( n2082 & n12202 ) | ( n9958 & n12202 ) ;
  assign n15071 = ( n10707 & n15069 ) | ( n10707 & n15070 ) | ( n15069 & n15070 ) ;
  assign n15073 = n12120 ^ n5918 ^ n407 ;
  assign n15072 = n6320 & ~n8145 ;
  assign n15074 = n15073 ^ n15072 ^ n5004 ;
  assign n15075 = n5393 ^ n5295 ^ n2688 ;
  assign n15076 = n15075 ^ n7978 ^ n4295 ;
  assign n15077 = ( n519 & n13856 ) | ( n519 & n15076 ) | ( n13856 & n15076 ) ;
  assign n15078 = n7106 ^ n5601 ^ n1499 ;
  assign n15079 = n15078 ^ n7930 ^ n3575 ;
  assign n15080 = n15079 ^ n10459 ^ n565 ;
  assign n15081 = ( n13048 & ~n13378 ) | ( n13048 & n15080 ) | ( ~n13378 & n15080 ) ;
  assign n15082 = n6378 ^ n5383 ^ n3804 ;
  assign n15083 = ( n1437 & ~n4708 ) | ( n1437 & n15082 ) | ( ~n4708 & n15082 ) ;
  assign n15084 = ( n3988 & ~n4354 ) | ( n3988 & n11128 ) | ( ~n4354 & n11128 ) ;
  assign n15085 = ( n14717 & n15083 ) | ( n14717 & ~n15084 ) | ( n15083 & ~n15084 ) ;
  assign n15086 = ( n1009 & n5822 ) | ( n1009 & n15085 ) | ( n5822 & n15085 ) ;
  assign n15087 = ( n3223 & n4747 ) | ( n3223 & n5056 ) | ( n4747 & n5056 ) ;
  assign n15088 = n15087 ^ n2254 ^ n643 ;
  assign n15089 = n9677 & n15088 ;
  assign n15090 = n12311 | n15089 ;
  assign n15092 = n10955 ^ n359 ^ n335 ;
  assign n15091 = n10202 ^ n9106 ^ n8885 ;
  assign n15093 = n15092 ^ n15091 ^ n2962 ;
  assign n15094 = ( ~n625 & n5850 ) | ( ~n625 & n15093 ) | ( n5850 & n15093 ) ;
  assign n15095 = ( ~x81 & n1492 ) | ( ~x81 & n3243 ) | ( n1492 & n3243 ) ;
  assign n15096 = n10488 ^ n9772 ^ n2624 ;
  assign n15097 = ( n1223 & ~n9004 ) | ( n1223 & n15096 ) | ( ~n9004 & n15096 ) ;
  assign n15098 = ( n10216 & n15095 ) | ( n10216 & ~n15097 ) | ( n15095 & ~n15097 ) ;
  assign n15099 = ( n2143 & n9879 ) | ( n2143 & n14905 ) | ( n9879 & n14905 ) ;
  assign n15104 = n7770 | n11937 ;
  assign n15100 = n11688 ^ n10081 ^ n4292 ;
  assign n15101 = ( n2492 & n9605 ) | ( n2492 & n15100 ) | ( n9605 & n15100 ) ;
  assign n15102 = ( n905 & ~n12867 ) | ( n905 & n15101 ) | ( ~n12867 & n15101 ) ;
  assign n15103 = ( ~n5908 & n8541 ) | ( ~n5908 & n15102 ) | ( n8541 & n15102 ) ;
  assign n15105 = n15104 ^ n15103 ^ n12533 ;
  assign n15106 = n2476 | n5412 ;
  assign n15107 = n15106 ^ n9143 ^ 1'b0 ;
  assign n15109 = ( n916 & n1010 ) | ( n916 & ~n8740 ) | ( n1010 & ~n8740 ) ;
  assign n15108 = n14925 ^ n11844 ^ n1559 ;
  assign n15110 = n15109 ^ n15108 ^ 1'b0 ;
  assign n15111 = n7565 ^ n3840 ^ n3699 ;
  assign n15112 = ( n1851 & ~n13822 ) | ( n1851 & n15111 ) | ( ~n13822 & n15111 ) ;
  assign n15117 = ( n1336 & ~n3102 ) | ( n1336 & n8138 ) | ( ~n3102 & n8138 ) ;
  assign n15118 = ( n1706 & n6192 ) | ( n1706 & n6832 ) | ( n6192 & n6832 ) ;
  assign n15119 = ( n7082 & ~n11160 ) | ( n7082 & n14048 ) | ( ~n11160 & n14048 ) ;
  assign n15120 = n15119 ^ n4768 ^ 1'b0 ;
  assign n15121 = n15118 & ~n15120 ;
  assign n15122 = ~n15117 & n15121 ;
  assign n15113 = n12249 ^ n533 ^ 1'b0 ;
  assign n15114 = ( ~n8188 & n12264 ) | ( ~n8188 & n15113 ) | ( n12264 & n15113 ) ;
  assign n15115 = ( n3367 & n12623 ) | ( n3367 & ~n15114 ) | ( n12623 & ~n15114 ) ;
  assign n15116 = ( n2485 & n10513 ) | ( n2485 & ~n15115 ) | ( n10513 & ~n15115 ) ;
  assign n15123 = n15122 ^ n15116 ^ n8212 ;
  assign n15129 = n3886 | n7182 ;
  assign n15124 = n11703 ^ n9867 ^ 1'b0 ;
  assign n15125 = n535 & n15124 ;
  assign n15126 = n10075 ^ n4696 ^ x102 ;
  assign n15127 = n15126 ^ n4888 ^ n2900 ;
  assign n15128 = ( n2371 & n15125 ) | ( n2371 & n15127 ) | ( n15125 & n15127 ) ;
  assign n15130 = n15129 ^ n15128 ^ n6003 ;
  assign n15131 = n11292 ^ n10686 ^ n851 ;
  assign n15135 = ( n1176 & ~n5277 ) | ( n1176 & n7128 ) | ( ~n5277 & n7128 ) ;
  assign n15136 = ( n745 & ~n2063 ) | ( n745 & n15135 ) | ( ~n2063 & n15135 ) ;
  assign n15137 = n15136 ^ n6910 ^ n2229 ;
  assign n15138 = n15137 ^ n8288 ^ n8163 ;
  assign n15132 = ( ~n854 & n5286 ) | ( ~n854 & n9175 ) | ( n5286 & n9175 ) ;
  assign n15133 = ( n4236 & n8067 ) | ( n4236 & n15132 ) | ( n8067 & n15132 ) ;
  assign n15134 = n15133 ^ n11678 ^ n4199 ;
  assign n15139 = n15138 ^ n15134 ^ n9566 ;
  assign n15140 = ( n2425 & ~n5624 ) | ( n2425 & n6148 ) | ( ~n5624 & n6148 ) ;
  assign n15141 = n5702 ^ n4798 ^ n1696 ;
  assign n15142 = ( n4659 & ~n15140 ) | ( n4659 & n15141 ) | ( ~n15140 & n15141 ) ;
  assign n15143 = n15142 ^ n5377 ^ n4441 ;
  assign n15162 = n6993 ^ n2494 ^ 1'b0 ;
  assign n15144 = ~n1794 & n6169 ;
  assign n15146 = n3348 & n4195 ;
  assign n15147 = ~n5075 & n15146 ;
  assign n15145 = n7134 ^ n3403 ^ n1966 ;
  assign n15148 = n15147 ^ n15145 ^ n1193 ;
  assign n15149 = ( n2438 & n4504 ) | ( n2438 & n15148 ) | ( n4504 & n15148 ) ;
  assign n15154 = ( n3804 & n3899 ) | ( n3804 & ~n8279 ) | ( n3899 & ~n8279 ) ;
  assign n15150 = n6761 ^ n671 ^ n623 ;
  assign n15151 = n15150 ^ n10808 ^ n8048 ;
  assign n15152 = n2480 | n11587 ;
  assign n15153 = ( n2824 & ~n15151 ) | ( n2824 & n15152 ) | ( ~n15151 & n15152 ) ;
  assign n15155 = n15154 ^ n15153 ^ 1'b0 ;
  assign n15156 = n6433 ^ n6051 ^ 1'b0 ;
  assign n15157 = n15156 ^ n11468 ^ n4957 ;
  assign n15158 = n5355 | n15157 ;
  assign n15159 = n15158 ^ n1328 ^ x243 ;
  assign n15160 = n15155 | n15159 ;
  assign n15161 = ( n15144 & n15149 ) | ( n15144 & ~n15160 ) | ( n15149 & ~n15160 ) ;
  assign n15163 = n15162 ^ n15161 ^ 1'b0 ;
  assign n15164 = ~n1777 & n15163 ;
  assign n15165 = n9042 | n10127 ;
  assign n15166 = n15165 ^ n2324 ^ 1'b0 ;
  assign n15167 = n8980 | n10073 ;
  assign n15168 = n9067 ^ n5989 ^ n5324 ;
  assign n15172 = ( n1249 & n2264 ) | ( n1249 & n13850 ) | ( n2264 & n13850 ) ;
  assign n15173 = ( n1636 & ~n13015 ) | ( n1636 & n15172 ) | ( ~n13015 & n15172 ) ;
  assign n15169 = ( ~n1952 & n4173 ) | ( ~n1952 & n6446 ) | ( n4173 & n6446 ) ;
  assign n15170 = ( n3903 & n5790 ) | ( n3903 & n15169 ) | ( n5790 & n15169 ) ;
  assign n15171 = ( n4379 & n14656 ) | ( n4379 & ~n15170 ) | ( n14656 & ~n15170 ) ;
  assign n15174 = n15173 ^ n15171 ^ n1656 ;
  assign n15175 = n4285 & ~n15174 ;
  assign n15176 = ( n940 & n1629 ) | ( n940 & ~n4850 ) | ( n1629 & ~n4850 ) ;
  assign n15177 = ~n2378 & n15176 ;
  assign n15178 = n15177 ^ n10163 ^ n3519 ;
  assign n15179 = ( n482 & ~n992 ) | ( n482 & n4597 ) | ( ~n992 & n4597 ) ;
  assign n15180 = ( n2163 & n7433 ) | ( n2163 & ~n15179 ) | ( n7433 & ~n15179 ) ;
  assign n15183 = ( n1531 & ~n10682 ) | ( n1531 & n12489 ) | ( ~n10682 & n12489 ) ;
  assign n15181 = n10281 ^ n499 ^ x233 ;
  assign n15182 = n878 | n15181 ;
  assign n15184 = n15183 ^ n15182 ^ 1'b0 ;
  assign n15185 = ( n15178 & n15180 ) | ( n15178 & n15184 ) | ( n15180 & n15184 ) ;
  assign n15186 = ( n5285 & n6092 ) | ( n5285 & n8841 ) | ( n6092 & n8841 ) ;
  assign n15197 = ( ~n3346 & n5711 ) | ( ~n3346 & n5954 ) | ( n5711 & n5954 ) ;
  assign n15187 = n7979 ^ n7510 ^ n1052 ;
  assign n15188 = ( ~n4469 & n6334 ) | ( ~n4469 & n15187 ) | ( n6334 & n15187 ) ;
  assign n15189 = ( n2951 & n7579 ) | ( n2951 & n15188 ) | ( n7579 & n15188 ) ;
  assign n15190 = n15189 ^ n5152 ^ n2710 ;
  assign n15191 = n1863 & ~n9946 ;
  assign n15192 = n15191 ^ n477 ^ 1'b0 ;
  assign n15193 = ( ~n8048 & n11014 ) | ( ~n8048 & n15192 ) | ( n11014 & n15192 ) ;
  assign n15194 = n1172 | n15193 ;
  assign n15195 = n15190 & ~n15194 ;
  assign n15196 = n15195 ^ n13424 ^ n9918 ;
  assign n15198 = n15197 ^ n15196 ^ n6887 ;
  assign n15199 = n12462 ^ n1460 ^ x2 ;
  assign n15200 = n15199 ^ n13855 ^ 1'b0 ;
  assign n15201 = ( n272 & n8030 ) | ( n272 & n15200 ) | ( n8030 & n15200 ) ;
  assign n15202 = n8513 | n15201 ;
  assign n15207 = x192 & n8860 ;
  assign n15208 = n15207 ^ n3766 ^ 1'b0 ;
  assign n15203 = ( n5785 & n6636 ) | ( n5785 & n9803 ) | ( n6636 & n9803 ) ;
  assign n15204 = n6312 & n15203 ;
  assign n15205 = n7064 & n15204 ;
  assign n15206 = n13518 & ~n15205 ;
  assign n15209 = n15208 ^ n15206 ^ 1'b0 ;
  assign n15210 = n2481 & ~n11824 ;
  assign n15211 = n15210 ^ n6798 ^ 1'b0 ;
  assign n15212 = n15211 ^ n12036 ^ n10740 ;
  assign n15213 = ( n1998 & ~n3881 ) | ( n1998 & n5053 ) | ( ~n3881 & n5053 ) ;
  assign n15214 = n6334 ^ n2651 ^ 1'b0 ;
  assign n15215 = n15213 & n15214 ;
  assign n15216 = ~n8850 & n15215 ;
  assign n15217 = ~n6952 & n15216 ;
  assign n15219 = n8138 ^ n2919 ^ 1'b0 ;
  assign n15218 = ( n1638 & n6066 ) | ( n1638 & ~n11400 ) | ( n6066 & ~n11400 ) ;
  assign n15220 = n15219 ^ n15218 ^ n4001 ;
  assign n15221 = ( n15212 & n15217 ) | ( n15212 & ~n15220 ) | ( n15217 & ~n15220 ) ;
  assign n15225 = n2886 ^ n532 ^ 1'b0 ;
  assign n15226 = n3185 & ~n15225 ;
  assign n15222 = ( ~n354 & n5828 ) | ( ~n354 & n8437 ) | ( n5828 & n8437 ) ;
  assign n15223 = ( n7407 & ~n10811 ) | ( n7407 & n15222 ) | ( ~n10811 & n15222 ) ;
  assign n15224 = n15223 ^ n8925 ^ n993 ;
  assign n15227 = n15226 ^ n15224 ^ n921 ;
  assign n15234 = n7500 ^ n4923 ^ n2774 ;
  assign n15228 = n4474 ^ n766 ^ 1'b0 ;
  assign n15229 = ~n8071 & n15228 ;
  assign n15230 = n3192 ^ n1772 ^ n1556 ;
  assign n15231 = ~n6022 & n15230 ;
  assign n15232 = n15231 ^ n4926 ^ 1'b0 ;
  assign n15233 = ( n5002 & n15229 ) | ( n5002 & ~n15232 ) | ( n15229 & ~n15232 ) ;
  assign n15235 = n15234 ^ n15233 ^ n4223 ;
  assign n15236 = n10042 ^ n9996 ^ 1'b0 ;
  assign n15237 = n5045 ^ n1889 ^ 1'b0 ;
  assign n15238 = ( ~n13304 & n14512 ) | ( ~n13304 & n15237 ) | ( n14512 & n15237 ) ;
  assign n15239 = n14330 ^ n11538 ^ x101 ;
  assign n15240 = ( n15236 & n15238 ) | ( n15236 & n15239 ) | ( n15238 & n15239 ) ;
  assign n15241 = ( n13143 & n15235 ) | ( n13143 & ~n15240 ) | ( n15235 & ~n15240 ) ;
  assign n15242 = n15241 ^ n14743 ^ n13575 ;
  assign n15247 = n7560 | n11051 ;
  assign n15243 = ( n5309 & n7977 ) | ( n5309 & ~n8045 ) | ( n7977 & ~n8045 ) ;
  assign n15244 = n10891 ^ n10357 ^ n2016 ;
  assign n15245 = n5990 ^ n2066 ^ 1'b0 ;
  assign n15246 = ( ~n15243 & n15244 ) | ( ~n15243 & n15245 ) | ( n15244 & n15245 ) ;
  assign n15248 = n15247 ^ n15246 ^ 1'b0 ;
  assign n15249 = ~n15242 & n15248 ;
  assign n15250 = n11468 ^ n3336 ^ n1007 ;
  assign n15251 = n1682 & n15250 ;
  assign n15252 = ~n8913 & n15251 ;
  assign n15253 = n15252 ^ n7934 ^ n6464 ;
  assign n15254 = n13051 ^ n7146 ^ n3531 ;
  assign n15259 = ( n7855 & n13469 ) | ( n7855 & n14233 ) | ( n13469 & n14233 ) ;
  assign n15260 = n15259 ^ n4519 ^ n3261 ;
  assign n15257 = n11557 ^ n2028 ^ n1515 ;
  assign n15255 = n685 ^ n582 ^ 1'b0 ;
  assign n15256 = ( ~n1312 & n5768 ) | ( ~n1312 & n15255 ) | ( n5768 & n15255 ) ;
  assign n15258 = n15257 ^ n15256 ^ n4543 ;
  assign n15261 = n15260 ^ n15258 ^ 1'b0 ;
  assign n15262 = ( n3605 & n7071 ) | ( n3605 & ~n13686 ) | ( n7071 & ~n13686 ) ;
  assign n15263 = ( ~x150 & n12613 ) | ( ~x150 & n15262 ) | ( n12613 & n15262 ) ;
  assign n15275 = n11818 ^ n4667 ^ 1'b0 ;
  assign n15276 = ( n3937 & n9353 ) | ( n3937 & n15275 ) | ( n9353 & n15275 ) ;
  assign n15269 = ( n623 & n4922 ) | ( n623 & ~n12952 ) | ( n4922 & ~n12952 ) ;
  assign n15270 = n5772 ^ n3631 ^ n1137 ;
  assign n15271 = ( ~n2796 & n4288 ) | ( ~n2796 & n15270 ) | ( n4288 & n15270 ) ;
  assign n15272 = ( n4223 & n15269 ) | ( n4223 & ~n15271 ) | ( n15269 & ~n15271 ) ;
  assign n15273 = n15272 ^ n13436 ^ n523 ;
  assign n15274 = n15273 ^ n9596 ^ n1095 ;
  assign n15264 = n3076 & n3549 ;
  assign n15265 = n8483 ^ n7211 ^ 1'b0 ;
  assign n15266 = n11006 ^ n2920 ^ 1'b0 ;
  assign n15267 = ~n15265 & n15266 ;
  assign n15268 = ( n14344 & ~n15264 ) | ( n14344 & n15267 ) | ( ~n15264 & n15267 ) ;
  assign n15277 = n15276 ^ n15274 ^ n15268 ;
  assign n15278 = n2346 & n11194 ;
  assign n15279 = ~n1194 & n15278 ;
  assign n15282 = n11078 ^ n10738 ^ n4237 ;
  assign n15280 = n2189 | n10584 ;
  assign n15281 = n15280 ^ n13785 ^ n1889 ;
  assign n15283 = n15282 ^ n15281 ^ n12313 ;
  assign n15284 = n13545 ^ n6620 ^ n4637 ;
  assign n15290 = n14849 ^ n12652 ^ n4103 ;
  assign n15285 = n7414 & n13852 ;
  assign n15286 = n7480 & n15285 ;
  assign n15287 = ( ~n13535 & n15199 ) | ( ~n13535 & n15286 ) | ( n15199 & n15286 ) ;
  assign n15288 = n10642 ^ n9525 ^ n8467 ;
  assign n15289 = ( n12002 & ~n15287 ) | ( n12002 & n15288 ) | ( ~n15287 & n15288 ) ;
  assign n15291 = n15290 ^ n15289 ^ n3964 ;
  assign n15294 = n2112 | n3518 ;
  assign n15295 = n15294 ^ n6819 ^ 1'b0 ;
  assign n15293 = ( n2494 & ~n7880 ) | ( n2494 & n11230 ) | ( ~n7880 & n11230 ) ;
  assign n15292 = n14008 ^ n9930 ^ 1'b0 ;
  assign n15296 = n15295 ^ n15293 ^ n15292 ;
  assign n15297 = ~n2384 & n6782 ;
  assign n15298 = n15296 & n15297 ;
  assign n15299 = ( n5864 & ~n10154 ) | ( n5864 & n13662 ) | ( ~n10154 & n13662 ) ;
  assign n15300 = ( n1751 & ~n4872 ) | ( n1751 & n15299 ) | ( ~n4872 & n15299 ) ;
  assign n15301 = n13240 ^ n737 ^ n537 ;
  assign n15303 = n732 | n10820 ;
  assign n15304 = n15303 ^ n1328 ^ 1'b0 ;
  assign n15302 = ( ~x36 & n722 ) | ( ~x36 & n5650 ) | ( n722 & n5650 ) ;
  assign n15305 = n15304 ^ n15302 ^ n13994 ;
  assign n15306 = ( n8853 & ~n15301 ) | ( n8853 & n15305 ) | ( ~n15301 & n15305 ) ;
  assign n15307 = ( n7590 & n10430 ) | ( n7590 & ~n11987 ) | ( n10430 & ~n11987 ) ;
  assign n15308 = n15307 ^ n9412 ^ n8119 ;
  assign n15309 = ( n5981 & ~n15306 ) | ( n5981 & n15308 ) | ( ~n15306 & n15308 ) ;
  assign n15310 = n9105 ^ n8805 ^ 1'b0 ;
  assign n15311 = ( ~n12593 & n15307 ) | ( ~n12593 & n15310 ) | ( n15307 & n15310 ) ;
  assign n15317 = ( x224 & n2561 ) | ( x224 & ~n5605 ) | ( n2561 & ~n5605 ) ;
  assign n15316 = n12753 ^ n5068 ^ n1971 ;
  assign n15312 = ( n1557 & n3056 ) | ( n1557 & n3104 ) | ( n3056 & n3104 ) ;
  assign n15313 = n15312 ^ n15113 ^ 1'b0 ;
  assign n15314 = ( n3088 & ~n9634 ) | ( n3088 & n15313 ) | ( ~n9634 & n15313 ) ;
  assign n15315 = n15314 ^ n6335 ^ n6240 ;
  assign n15318 = n15317 ^ n15316 ^ n15315 ;
  assign n15319 = n1779 & n14484 ;
  assign n15320 = n15319 ^ n13567 ^ n2902 ;
  assign n15321 = n5816 ^ n4939 ^ n2511 ;
  assign n15322 = ( n1491 & ~n14989 ) | ( n1491 & n15321 ) | ( ~n14989 & n15321 ) ;
  assign n15328 = ( n896 & n2602 ) | ( n896 & n2703 ) | ( n2602 & n2703 ) ;
  assign n15329 = n15328 ^ n14774 ^ x198 ;
  assign n15330 = n15329 ^ n1587 ^ n1492 ;
  assign n15325 = n13282 & ~n14049 ;
  assign n15326 = n13644 & n15325 ;
  assign n15323 = n8054 | n12446 ;
  assign n15324 = n15323 ^ n3555 ^ 1'b0 ;
  assign n15327 = n15326 ^ n15324 ^ n13570 ;
  assign n15331 = n15330 ^ n15327 ^ n12517 ;
  assign n15333 = ( x213 & n1452 ) | ( x213 & n5874 ) | ( n1452 & n5874 ) ;
  assign n15332 = ( n419 & ~n3492 ) | ( n419 & n3578 ) | ( ~n3492 & n3578 ) ;
  assign n15334 = n15333 ^ n15332 ^ n1342 ;
  assign n15335 = n15334 ^ n5101 ^ n1588 ;
  assign n15336 = n12639 ^ n8035 ^ 1'b0 ;
  assign n15337 = n13513 ^ n6864 ^ n2085 ;
  assign n15338 = n15336 & n15337 ;
  assign n15339 = ( n1971 & n3568 ) | ( n1971 & ~n9410 ) | ( n3568 & ~n9410 ) ;
  assign n15340 = n15339 ^ n7102 ^ n4847 ;
  assign n15342 = n2526 | n5817 ;
  assign n15343 = n6999 & ~n15342 ;
  assign n15344 = ( ~n3750 & n5540 ) | ( ~n3750 & n15102 ) | ( n5540 & n15102 ) ;
  assign n15345 = ( ~n12403 & n15343 ) | ( ~n12403 & n15344 ) | ( n15343 & n15344 ) ;
  assign n15341 = ( n1664 & ~n11136 ) | ( n1664 & n13689 ) | ( ~n11136 & n13689 ) ;
  assign n15346 = n15345 ^ n15341 ^ n3005 ;
  assign n15347 = n15346 ^ n4284 ^ 1'b0 ;
  assign n15348 = n15340 | n15347 ;
  assign n15351 = ( n4910 & ~n9498 ) | ( n4910 & n9847 ) | ( ~n9498 & n9847 ) ;
  assign n15349 = n8082 ^ n3622 ^ n2894 ;
  assign n15350 = ( n12818 & ~n14554 ) | ( n12818 & n15349 ) | ( ~n14554 & n15349 ) ;
  assign n15352 = n15351 ^ n15350 ^ n6102 ;
  assign n15353 = ( n2449 & ~n2521 ) | ( n2449 & n7609 ) | ( ~n2521 & n7609 ) ;
  assign n15354 = n15353 ^ n842 ^ 1'b0 ;
  assign n15355 = n7088 ^ n5941 ^ 1'b0 ;
  assign n15356 = ~n14790 & n15355 ;
  assign n15357 = ( n7212 & n7706 ) | ( n7212 & n15356 ) | ( n7706 & n15356 ) ;
  assign n15358 = ( n10941 & n11274 ) | ( n10941 & ~n15357 ) | ( n11274 & ~n15357 ) ;
  assign n15359 = n6892 & n12476 ;
  assign n15360 = n15359 ^ n1674 ^ 1'b0 ;
  assign n15361 = n15360 ^ n15178 ^ n575 ;
  assign n15362 = n4571 ^ n1731 ^ 1'b0 ;
  assign n15363 = ( n3813 & n4522 ) | ( n3813 & ~n6400 ) | ( n4522 & ~n6400 ) ;
  assign n15364 = n2623 & n15363 ;
  assign n15365 = n14558 & ~n15192 ;
  assign n15366 = n15365 ^ n725 ^ 1'b0 ;
  assign n15367 = n15366 ^ n1941 ^ 1'b0 ;
  assign n15368 = ( n4283 & ~n4922 ) | ( n4283 & n12380 ) | ( ~n4922 & n12380 ) ;
  assign n15369 = n15368 ^ n867 ^ n262 ;
  assign n15370 = ~n10403 & n15369 ;
  assign n15371 = n10965 & ~n15370 ;
  assign n15372 = n15367 & n15371 ;
  assign n15373 = n6638 ^ n6417 ^ n2698 ;
  assign n15374 = ~n3608 & n15373 ;
  assign n15375 = ( ~n1829 & n2047 ) | ( ~n1829 & n13481 ) | ( n2047 & n13481 ) ;
  assign n15376 = ( ~n989 & n2818 ) | ( ~n989 & n8335 ) | ( n2818 & n8335 ) ;
  assign n15377 = n15376 ^ n5966 ^ n1894 ;
  assign n15378 = ( n5714 & ~n11053 ) | ( n5714 & n15377 ) | ( ~n11053 & n15377 ) ;
  assign n15379 = n15378 ^ n4197 ^ n1621 ;
  assign n15380 = ( n2039 & ~n6099 ) | ( n2039 & n14286 ) | ( ~n6099 & n14286 ) ;
  assign n15381 = ~n839 & n14873 ;
  assign n15382 = ~n15380 & n15381 ;
  assign n15383 = ~n10423 & n14040 ;
  assign n15384 = ( ~n477 & n7423 ) | ( ~n477 & n10079 ) | ( n7423 & n10079 ) ;
  assign n15390 = ( n2548 & ~n2602 ) | ( n2548 & n3917 ) | ( ~n2602 & n3917 ) ;
  assign n15385 = n6693 ^ n4760 ^ n3047 ;
  assign n15386 = n2494 ^ n2096 ^ 1'b0 ;
  assign n15387 = n3820 | n15386 ;
  assign n15388 = ( x20 & ~n7088 ) | ( x20 & n15387 ) | ( ~n7088 & n15387 ) ;
  assign n15389 = ( n13078 & n15385 ) | ( n13078 & ~n15388 ) | ( n15385 & ~n15388 ) ;
  assign n15391 = n15390 ^ n15389 ^ n1114 ;
  assign n15392 = ( n956 & n8153 ) | ( n956 & n15391 ) | ( n8153 & n15391 ) ;
  assign n15393 = ( ~n2747 & n6790 ) | ( ~n2747 & n13245 ) | ( n6790 & n13245 ) ;
  assign n15394 = n15393 ^ n8763 ^ n1843 ;
  assign n15395 = n15394 ^ n8047 ^ x174 ;
  assign n15396 = ( n6192 & n7459 ) | ( n6192 & ~n15395 ) | ( n7459 & ~n15395 ) ;
  assign n15403 = ( n1434 & n10129 ) | ( n1434 & ~n11401 ) | ( n10129 & ~n11401 ) ;
  assign n15404 = n15403 ^ n5111 ^ n3042 ;
  assign n15397 = n9812 ^ n5514 ^ n1547 ;
  assign n15398 = ( n1404 & n7760 ) | ( n1404 & n9607 ) | ( n7760 & n9607 ) ;
  assign n15399 = n14967 ^ n3171 ^ 1'b0 ;
  assign n15400 = ( n1359 & ~n5269 ) | ( n1359 & n15399 ) | ( ~n5269 & n15399 ) ;
  assign n15401 = ( n744 & n15398 ) | ( n744 & ~n15400 ) | ( n15398 & ~n15400 ) ;
  assign n15402 = ( n5733 & n15397 ) | ( n5733 & n15401 ) | ( n15397 & n15401 ) ;
  assign n15405 = n15404 ^ n15402 ^ n11908 ;
  assign n15406 = n9803 ^ n5456 ^ n2127 ;
  assign n15407 = n6819 ^ n5376 ^ n1077 ;
  assign n15408 = n15407 ^ n5940 ^ 1'b0 ;
  assign n15409 = n15406 & n15408 ;
  assign n15410 = n11272 ^ n5196 ^ x52 ;
  assign n15411 = n15410 ^ n8996 ^ n3719 ;
  assign n15412 = n15411 ^ n6217 ^ n3749 ;
  assign n15413 = n15109 ^ n3228 ^ n894 ;
  assign n15415 = ( n1810 & ~n3385 ) | ( n1810 & n6192 ) | ( ~n3385 & n6192 ) ;
  assign n15414 = n3091 | n10572 ;
  assign n15416 = n15415 ^ n15414 ^ 1'b0 ;
  assign n15417 = ( n2438 & n15413 ) | ( n2438 & n15416 ) | ( n15413 & n15416 ) ;
  assign n15418 = n15417 ^ n3416 ^ 1'b0 ;
  assign n15419 = ~n15412 & n15418 ;
  assign n15420 = n11748 ^ n5338 ^ 1'b0 ;
  assign n15421 = ( n5880 & n8887 ) | ( n5880 & ~n12712 ) | ( n8887 & ~n12712 ) ;
  assign n15422 = ( n12695 & ~n14322 ) | ( n12695 & n15421 ) | ( ~n14322 & n15421 ) ;
  assign n15423 = n15422 ^ n9679 ^ n8924 ;
  assign n15424 = ( n1667 & n15420 ) | ( n1667 & ~n15423 ) | ( n15420 & ~n15423 ) ;
  assign n15429 = ( n2235 & n2504 ) | ( n2235 & n4293 ) | ( n2504 & n4293 ) ;
  assign n15430 = n15429 ^ n13025 ^ n9865 ;
  assign n15431 = ( n1535 & n12739 ) | ( n1535 & ~n15430 ) | ( n12739 & ~n15430 ) ;
  assign n15425 = ( n389 & ~n990 ) | ( n389 & n5564 ) | ( ~n990 & n5564 ) ;
  assign n15426 = n11782 ^ n2980 ^ n2411 ;
  assign n15427 = ( n1182 & ~n15425 ) | ( n1182 & n15426 ) | ( ~n15425 & n15426 ) ;
  assign n15428 = n15427 ^ n14803 ^ n14756 ;
  assign n15432 = n15431 ^ n15428 ^ n15272 ;
  assign n15433 = n6608 ^ n5012 ^ n955 ;
  assign n15434 = ( n12991 & n14383 ) | ( n12991 & n15433 ) | ( n14383 & n15433 ) ;
  assign n15435 = ( n10669 & n13312 ) | ( n10669 & n13619 ) | ( n13312 & n13619 ) ;
  assign n15436 = ( n6886 & n11169 ) | ( n6886 & ~n13936 ) | ( n11169 & ~n13936 ) ;
  assign n15437 = ( x75 & ~n6347 ) | ( x75 & n9854 ) | ( ~n6347 & n9854 ) ;
  assign n15438 = n6164 & ~n15437 ;
  assign n15439 = ( n4198 & ~n12684 ) | ( n4198 & n15438 ) | ( ~n12684 & n15438 ) ;
  assign n15440 = ( n6947 & n7675 ) | ( n6947 & ~n15439 ) | ( n7675 & ~n15439 ) ;
  assign n15441 = ( n15435 & ~n15436 ) | ( n15435 & n15440 ) | ( ~n15436 & n15440 ) ;
  assign n15442 = n15441 ^ n5103 ^ n1673 ;
  assign n15443 = n1135 & ~n1247 ;
  assign n15444 = n15443 ^ n11091 ^ 1'b0 ;
  assign n15445 = n15444 ^ n11581 ^ n4458 ;
  assign n15446 = n10381 ^ n10107 ^ n6694 ;
  assign n15447 = n4354 ^ n4011 ^ n3832 ;
  assign n15448 = n15447 ^ n6214 ^ x222 ;
  assign n15449 = ( n3302 & n5339 ) | ( n3302 & n6950 ) | ( n5339 & n6950 ) ;
  assign n15450 = ( ~n1526 & n6982 ) | ( ~n1526 & n15449 ) | ( n6982 & n15449 ) ;
  assign n15451 = ~n625 & n6975 ;
  assign n15452 = ~n15450 & n15451 ;
  assign n15453 = n15452 ^ n2974 ^ n2303 ;
  assign n15454 = ( n1686 & n9816 ) | ( n1686 & ~n15453 ) | ( n9816 & ~n15453 ) ;
  assign n15455 = n15454 ^ n9707 ^ n5179 ;
  assign n15456 = ( n1175 & ~n9627 ) | ( n1175 & n10203 ) | ( ~n9627 & n10203 ) ;
  assign n15457 = ( ~n3865 & n4648 ) | ( ~n3865 & n15456 ) | ( n4648 & n15456 ) ;
  assign n15458 = n15457 ^ n8041 ^ n3949 ;
  assign n15459 = n12902 ^ n1983 ^ 1'b0 ;
  assign n15460 = ( ~n1132 & n1522 ) | ( ~n1132 & n9366 ) | ( n1522 & n9366 ) ;
  assign n15461 = ( n3634 & n12242 ) | ( n3634 & ~n15460 ) | ( n12242 & ~n15460 ) ;
  assign n15462 = n561 & ~n14920 ;
  assign n15463 = n15462 ^ n12357 ^ 1'b0 ;
  assign n15464 = n15463 ^ n5595 ^ n504 ;
  assign n15465 = n15464 ^ n3899 ^ 1'b0 ;
  assign n15466 = n12496 & ~n15465 ;
  assign n15471 = n8862 ^ n4472 ^ n2112 ;
  assign n15467 = n10774 & ~n11005 ;
  assign n15468 = n2943 & n15467 ;
  assign n15469 = ( n9918 & n12218 ) | ( n9918 & ~n15468 ) | ( n12218 & ~n15468 ) ;
  assign n15470 = n15469 ^ n5758 ^ n3323 ;
  assign n15472 = n15471 ^ n15470 ^ n13231 ;
  assign n15473 = n15472 ^ n6576 ^ 1'b0 ;
  assign n15474 = ( n1171 & n9931 ) | ( n1171 & n10570 ) | ( n9931 & n10570 ) ;
  assign n15475 = n13596 ^ n1870 ^ 1'b0 ;
  assign n15476 = n15474 & ~n15475 ;
  assign n15477 = n10156 ^ n9433 ^ n4385 ;
  assign n15478 = ( ~n10729 & n11991 ) | ( ~n10729 & n15477 ) | ( n11991 & n15477 ) ;
  assign n15479 = ( n7973 & ~n11182 ) | ( n7973 & n15478 ) | ( ~n11182 & n15478 ) ;
  assign n15480 = ( n11438 & ~n13700 ) | ( n11438 & n15479 ) | ( ~n13700 & n15479 ) ;
  assign n15481 = n11989 ^ n8521 ^ n3567 ;
  assign n15482 = n11396 ^ n4343 ^ 1'b0 ;
  assign n15483 = ~n1636 & n15482 ;
  assign n15484 = ( n4412 & n6413 ) | ( n4412 & n15483 ) | ( n6413 & n15483 ) ;
  assign n15486 = n11304 ^ n10395 ^ n4635 ;
  assign n15487 = ( n4226 & ~n6991 ) | ( n4226 & n8727 ) | ( ~n6991 & n8727 ) ;
  assign n15488 = ( n3866 & n15486 ) | ( n3866 & n15487 ) | ( n15486 & n15487 ) ;
  assign n15485 = n9414 ^ n2013 ^ n1949 ;
  assign n15489 = n15488 ^ n15485 ^ n8414 ;
  assign n15490 = ( n6219 & n13073 ) | ( n6219 & n15489 ) | ( n13073 & n15489 ) ;
  assign n15491 = n15484 & ~n15490 ;
  assign n15492 = ( n1324 & n4403 ) | ( n1324 & ~n8736 ) | ( n4403 & ~n8736 ) ;
  assign n15493 = ( n782 & n8238 ) | ( n782 & n15492 ) | ( n8238 & n15492 ) ;
  assign n15494 = ( n3511 & ~n13967 ) | ( n3511 & n15493 ) | ( ~n13967 & n15493 ) ;
  assign n15495 = n11705 ^ n10059 ^ n951 ;
  assign n15497 = ( n3141 & n6859 ) | ( n3141 & ~n13340 ) | ( n6859 & ~n13340 ) ;
  assign n15496 = n9585 ^ n7178 ^ n4978 ;
  assign n15498 = n15497 ^ n15496 ^ n2484 ;
  assign n15500 = n9932 ^ n1656 ^ 1'b0 ;
  assign n15501 = n15500 ^ n4529 ^ 1'b0 ;
  assign n15499 = n2493 & ~n5141 ;
  assign n15502 = n15501 ^ n15499 ^ 1'b0 ;
  assign n15503 = n15502 ^ n7384 ^ n1998 ;
  assign n15507 = n14040 ^ n6296 ^ 1'b0 ;
  assign n15508 = ~n7926 & n15507 ;
  assign n15509 = ( n4646 & n5161 ) | ( n4646 & ~n15508 ) | ( n5161 & ~n15508 ) ;
  assign n15506 = ( ~n3449 & n4278 ) | ( ~n3449 & n13705 ) | ( n4278 & n13705 ) ;
  assign n15505 = n3135 ^ n2843 ^ n2462 ;
  assign n15510 = n15509 ^ n15506 ^ n15505 ;
  assign n15504 = ( n5310 & n12389 ) | ( n5310 & ~n13335 ) | ( n12389 & ~n13335 ) ;
  assign n15511 = n15510 ^ n15504 ^ n1971 ;
  assign n15512 = n15511 ^ n11428 ^ n518 ;
  assign n15513 = n11659 ^ n10241 ^ n3784 ;
  assign n15514 = ( x252 & n10060 ) | ( x252 & ~n15513 ) | ( n10060 & ~n15513 ) ;
  assign n15515 = n4317 ^ n2838 ^ n1109 ;
  assign n15516 = n15515 ^ n14212 ^ n13103 ;
  assign n15517 = n10372 ^ n6560 ^ n4177 ;
  assign n15518 = n10556 ^ n3845 ^ n884 ;
  assign n15519 = ( n15516 & ~n15517 ) | ( n15516 & n15518 ) | ( ~n15517 & n15518 ) ;
  assign n15521 = n6792 & ~n9088 ;
  assign n15522 = ( n2240 & n4015 ) | ( n2240 & ~n4645 ) | ( n4015 & ~n4645 ) ;
  assign n15523 = n15522 ^ n2240 ^ 1'b0 ;
  assign n15524 = n3199 & n15523 ;
  assign n15525 = ( n13822 & n15521 ) | ( n13822 & ~n15524 ) | ( n15521 & ~n15524 ) ;
  assign n15526 = n15525 ^ n11175 ^ n5557 ;
  assign n15520 = n14748 ^ n12359 ^ n2799 ;
  assign n15527 = n15526 ^ n15520 ^ 1'b0 ;
  assign n15528 = n15519 & n15527 ;
  assign n15529 = ( n1310 & n5099 ) | ( n1310 & n14839 ) | ( n5099 & n14839 ) ;
  assign n15530 = n7449 & ~n15529 ;
  assign n15531 = ( n3065 & n12556 ) | ( n3065 & ~n15530 ) | ( n12556 & ~n15530 ) ;
  assign n15532 = ( n1564 & ~n3984 ) | ( n1564 & n11214 ) | ( ~n3984 & n11214 ) ;
  assign n15533 = ( ~n5935 & n6496 ) | ( ~n5935 & n15532 ) | ( n6496 & n15532 ) ;
  assign n15534 = n4250 & ~n11413 ;
  assign n15535 = ~n3576 & n15534 ;
  assign n15536 = ( n2171 & n15533 ) | ( n2171 & n15535 ) | ( n15533 & n15535 ) ;
  assign n15537 = n12460 ^ n2412 ^ 1'b0 ;
  assign n15538 = n15537 ^ n12795 ^ n3132 ;
  assign n15539 = n13364 ^ n8279 ^ n5149 ;
  assign n15540 = n15539 ^ n2669 ^ n2332 ;
  assign n15541 = ( n10832 & n15176 ) | ( n10832 & n15540 ) | ( n15176 & n15540 ) ;
  assign n15542 = n15541 ^ n14591 ^ n6655 ;
  assign n15543 = n7925 ^ n3296 ^ n1390 ;
  assign n15544 = n15543 ^ n3378 ^ 1'b0 ;
  assign n15545 = ( n5981 & ~n8804 ) | ( n5981 & n15544 ) | ( ~n8804 & n15544 ) ;
  assign n15546 = n9848 ^ n7731 ^ 1'b0 ;
  assign n15547 = n15546 ^ n11107 ^ n6060 ;
  assign n15548 = ( n1357 & n6160 ) | ( n1357 & n9010 ) | ( n6160 & n9010 ) ;
  assign n15549 = n15548 ^ n6250 ^ 1'b0 ;
  assign n15550 = ( ~n1152 & n6540 ) | ( ~n1152 & n15549 ) | ( n6540 & n15549 ) ;
  assign n15551 = n14715 & ~n15550 ;
  assign n15552 = n6491 ^ n4077 ^ x88 ;
  assign n15553 = ( n3495 & n12871 ) | ( n3495 & ~n15552 ) | ( n12871 & ~n15552 ) ;
  assign n15554 = ( n1799 & n6809 ) | ( n1799 & n10523 ) | ( n6809 & n10523 ) ;
  assign n15555 = ( n9892 & n15553 ) | ( n9892 & n15554 ) | ( n15553 & n15554 ) ;
  assign n15556 = ( ~n2805 & n14658 ) | ( ~n2805 & n15555 ) | ( n14658 & n15555 ) ;
  assign n15557 = ( x220 & n1203 ) | ( x220 & ~n8448 ) | ( n1203 & ~n8448 ) ;
  assign n15558 = ( ~n4275 & n7214 ) | ( ~n4275 & n15557 ) | ( n7214 & n15557 ) ;
  assign n15559 = n15558 ^ n5637 ^ n987 ;
  assign n15560 = ~n1300 & n1560 ;
  assign n15561 = n15560 ^ n1702 ^ 1'b0 ;
  assign n15562 = n15561 ^ n3513 ^ n1759 ;
  assign n15563 = n15562 ^ n11037 ^ 1'b0 ;
  assign n15565 = n4903 ^ n2799 ^ 1'b0 ;
  assign n15566 = ~n12929 & n15565 ;
  assign n15564 = n5942 ^ n2607 ^ x51 ;
  assign n15567 = n15566 ^ n15564 ^ n2628 ;
  assign n15568 = n345 & n15567 ;
  assign n15569 = n5078 & n15568 ;
  assign n15570 = ( n8286 & ~n10144 ) | ( n8286 & n15569 ) | ( ~n10144 & n15569 ) ;
  assign n15571 = ( n15559 & n15563 ) | ( n15559 & ~n15570 ) | ( n15563 & ~n15570 ) ;
  assign n15580 = ~n1914 & n2064 ;
  assign n15581 = ~n4154 & n15580 ;
  assign n15582 = ( ~n1388 & n6729 ) | ( ~n1388 & n15581 ) | ( n6729 & n15581 ) ;
  assign n15576 = ( n8260 & n10690 ) | ( n8260 & n12797 ) | ( n10690 & n12797 ) ;
  assign n15577 = n15576 ^ n15272 ^ n2516 ;
  assign n15578 = n15577 ^ n1103 ^ 1'b0 ;
  assign n15579 = ~n1334 & n15578 ;
  assign n15572 = n8668 ^ n3437 ^ 1'b0 ;
  assign n15573 = n15572 ^ n9251 ^ n5310 ;
  assign n15574 = n9143 ^ n3701 ^ n3146 ;
  assign n15575 = ( n13607 & n15573 ) | ( n13607 & ~n15574 ) | ( n15573 & ~n15574 ) ;
  assign n15583 = n15582 ^ n15579 ^ n15575 ;
  assign n15585 = ( x103 & n1368 ) | ( x103 & n7764 ) | ( n1368 & n7764 ) ;
  assign n15586 = n15585 ^ n9917 ^ 1'b0 ;
  assign n15584 = n5157 & n12473 ;
  assign n15587 = n15586 ^ n15584 ^ 1'b0 ;
  assign n15588 = ( n7162 & ~n12704 ) | ( n7162 & n15587 ) | ( ~n12704 & n15587 ) ;
  assign n15589 = n8484 ^ n1990 ^ n657 ;
  assign n15590 = ~n4269 & n15053 ;
  assign n15591 = n15590 ^ n11319 ^ 1'b0 ;
  assign n15593 = n10678 ^ n4911 ^ n2837 ;
  assign n15592 = n12162 ^ n8257 ^ 1'b0 ;
  assign n15594 = n15593 ^ n15592 ^ n1332 ;
  assign n15595 = ( ~n15589 & n15591 ) | ( ~n15589 & n15594 ) | ( n15591 & n15594 ) ;
  assign n15596 = n10842 ^ n9190 ^ n8653 ;
  assign n15597 = ( n1795 & n8639 ) | ( n1795 & n10599 ) | ( n8639 & n10599 ) ;
  assign n15598 = ( n12977 & n15596 ) | ( n12977 & n15597 ) | ( n15596 & n15597 ) ;
  assign n15599 = n4304 & n8829 ;
  assign n15600 = n15599 ^ n13530 ^ 1'b0 ;
  assign n15601 = n8157 ^ n2546 ^ 1'b0 ;
  assign n15602 = ( n3298 & n8131 ) | ( n3298 & ~n15601 ) | ( n8131 & ~n15601 ) ;
  assign n15603 = ~n7766 & n15602 ;
  assign n15604 = ( n15598 & n15600 ) | ( n15598 & ~n15603 ) | ( n15600 & ~n15603 ) ;
  assign n15605 = n11529 ^ n7183 ^ 1'b0 ;
  assign n15606 = n12425 & n15605 ;
  assign n15607 = ( ~n3034 & n12457 ) | ( ~n3034 & n14512 ) | ( n12457 & n14512 ) ;
  assign n15608 = n10697 ^ n6803 ^ n4403 ;
  assign n15609 = n15608 ^ n4115 ^ 1'b0 ;
  assign n15610 = n3183 | n15609 ;
  assign n15611 = ( n10727 & n15521 ) | ( n10727 & n15610 ) | ( n15521 & n15610 ) ;
  assign n15612 = n6205 ^ n5816 ^ n547 ;
  assign n15613 = n15612 ^ n9569 ^ n1217 ;
  assign n15614 = n15613 ^ n3464 ^ n1873 ;
  assign n15615 = ( ~n2573 & n4128 ) | ( ~n2573 & n14769 ) | ( n4128 & n14769 ) ;
  assign n15616 = ( n13132 & ~n15614 ) | ( n13132 & n15615 ) | ( ~n15614 & n15615 ) ;
  assign n15618 = n7723 ^ n4858 ^ n1067 ;
  assign n15619 = n987 & ~n15618 ;
  assign n15620 = ~n3949 & n15619 ;
  assign n15621 = n15620 ^ n2655 ^ n839 ;
  assign n15617 = n5496 ^ n5251 ^ n2042 ;
  assign n15622 = n15621 ^ n15617 ^ 1'b0 ;
  assign n15624 = n12854 ^ n8522 ^ x195 ;
  assign n15623 = n6319 & ~n9427 ;
  assign n15625 = n15624 ^ n15623 ^ 1'b0 ;
  assign n15626 = ( n3048 & n11824 ) | ( n3048 & ~n15625 ) | ( n11824 & ~n15625 ) ;
  assign n15627 = n15626 ^ n10684 ^ 1'b0 ;
  assign n15628 = n2796 ^ n1655 ^ n752 ;
  assign n15629 = ( n11556 & ~n14079 ) | ( n11556 & n15628 ) | ( ~n14079 & n15628 ) ;
  assign n15630 = ( ~n1950 & n7451 ) | ( ~n1950 & n14059 ) | ( n7451 & n14059 ) ;
  assign n15631 = ( n493 & ~n2328 ) | ( n493 & n5084 ) | ( ~n2328 & n5084 ) ;
  assign n15632 = ~n627 & n15631 ;
  assign n15633 = n11954 & n14729 ;
  assign n15634 = n15632 & n15633 ;
  assign n15635 = x154 & ~n15634 ;
  assign n15636 = n15630 & n15635 ;
  assign n15637 = ( n12030 & n13842 ) | ( n12030 & ~n15169 ) | ( n13842 & ~n15169 ) ;
  assign n15638 = ( n1314 & ~n8246 ) | ( n1314 & n11546 ) | ( ~n8246 & n11546 ) ;
  assign n15639 = n1120 ^ n830 ^ 1'b0 ;
  assign n15640 = ~n15638 & n15639 ;
  assign n15641 = ( n2658 & n6653 ) | ( n2658 & ~n9493 ) | ( n6653 & ~n9493 ) ;
  assign n15642 = n12462 & ~n15641 ;
  assign n15643 = ~n15640 & n15642 ;
  assign n15644 = ( ~n4786 & n15637 ) | ( ~n4786 & n15643 ) | ( n15637 & n15643 ) ;
  assign n15645 = ~n3580 & n7724 ;
  assign n15646 = ( n5900 & n10510 ) | ( n5900 & n12702 ) | ( n10510 & n12702 ) ;
  assign n15648 = ( n2228 & ~n4665 ) | ( n2228 & n8146 ) | ( ~n4665 & n8146 ) ;
  assign n15649 = ( ~n2471 & n10070 ) | ( ~n2471 & n15648 ) | ( n10070 & n15648 ) ;
  assign n15647 = ( n3273 & ~n12052 ) | ( n3273 & n12378 ) | ( ~n12052 & n12378 ) ;
  assign n15650 = n15649 ^ n15647 ^ n14034 ;
  assign n15651 = x99 & ~n4930 ;
  assign n15652 = x185 & n15651 ;
  assign n15653 = n15652 ^ n11255 ^ 1'b0 ;
  assign n15655 = n3721 ^ x237 ^ 1'b0 ;
  assign n15654 = n8668 | n12607 ;
  assign n15656 = n15655 ^ n15654 ^ n10897 ;
  assign n15657 = ( n11945 & ~n15653 ) | ( n11945 & n15656 ) | ( ~n15653 & n15656 ) ;
  assign n15658 = n11005 ^ n7312 ^ n1495 ;
  assign n15659 = ( n9918 & n15100 ) | ( n9918 & n15658 ) | ( n15100 & n15658 ) ;
  assign n15660 = ( n698 & n1540 ) | ( n698 & n15659 ) | ( n1540 & n15659 ) ;
  assign n15661 = n15660 ^ n11579 ^ n2385 ;
  assign n15662 = ( ~n9466 & n9720 ) | ( ~n9466 & n15661 ) | ( n9720 & n15661 ) ;
  assign n15663 = ( n716 & n2678 ) | ( n716 & n7196 ) | ( n2678 & n7196 ) ;
  assign n15664 = ( n1906 & n3598 ) | ( n1906 & n7509 ) | ( n3598 & n7509 ) ;
  assign n15665 = n15664 ^ n13803 ^ n5474 ;
  assign n15666 = ( ~n1929 & n15663 ) | ( ~n1929 & n15665 ) | ( n15663 & n15665 ) ;
  assign n15667 = n15666 ^ n2435 ^ n2359 ;
  assign n15668 = n13874 ^ n3984 ^ n954 ;
  assign n15669 = ( n3718 & ~n14790 ) | ( n3718 & n15668 ) | ( ~n14790 & n15668 ) ;
  assign n15671 = n345 & ~n2122 ;
  assign n15672 = ( ~n2817 & n8862 ) | ( ~n2817 & n15671 ) | ( n8862 & n15671 ) ;
  assign n15670 = ~n3363 & n7313 ;
  assign n15673 = n15672 ^ n15670 ^ 1'b0 ;
  assign n15678 = ( n4671 & n14478 ) | ( n4671 & ~n14503 ) | ( n14478 & ~n14503 ) ;
  assign n15677 = ( n3826 & ~n8274 ) | ( n3826 & n11858 ) | ( ~n8274 & n11858 ) ;
  assign n15674 = n9042 ^ n3395 ^ n1592 ;
  assign n15675 = ( ~n4646 & n14955 ) | ( ~n4646 & n15674 ) | ( n14955 & n15674 ) ;
  assign n15676 = n15675 ^ n4606 ^ 1'b0 ;
  assign n15679 = n15678 ^ n15677 ^ n15676 ;
  assign n15680 = ( n15669 & n15673 ) | ( n15669 & n15679 ) | ( n15673 & n15679 ) ;
  assign n15681 = ~n1272 & n11314 ;
  assign n15686 = n11211 ^ n4538 ^ 1'b0 ;
  assign n15682 = n12812 ^ n10095 ^ n3956 ;
  assign n15683 = ~n4521 & n15682 ;
  assign n15684 = n15683 ^ n4611 ^ 1'b0 ;
  assign n15685 = ( ~n11948 & n12603 ) | ( ~n11948 & n15684 ) | ( n12603 & n15684 ) ;
  assign n15687 = n15686 ^ n15685 ^ n7094 ;
  assign n15688 = n15687 ^ n3737 ^ n3146 ;
  assign n15690 = ( n5463 & n6198 ) | ( n5463 & ~n10907 ) | ( n6198 & ~n10907 ) ;
  assign n15691 = ( n1624 & n10775 ) | ( n1624 & n15690 ) | ( n10775 & n15690 ) ;
  assign n15692 = ( n4423 & n6361 ) | ( n4423 & n15691 ) | ( n6361 & n15691 ) ;
  assign n15693 = n15692 ^ n4289 ^ 1'b0 ;
  assign n15689 = ~n2434 & n14418 ;
  assign n15694 = n15693 ^ n15689 ^ 1'b0 ;
  assign n15695 = n13419 | n15694 ;
  assign n15696 = ( n865 & ~n9627 ) | ( n865 & n11374 ) | ( ~n9627 & n11374 ) ;
  assign n15697 = n15696 ^ n8067 ^ n3692 ;
  assign n15698 = n10490 ^ n10467 ^ n8398 ;
  assign n15699 = ( n2218 & n2716 ) | ( n2218 & n14189 ) | ( n2716 & n14189 ) ;
  assign n15700 = ( ~n5800 & n13645 ) | ( ~n5800 & n15699 ) | ( n13645 & n15699 ) ;
  assign n15701 = ( n15697 & n15698 ) | ( n15697 & n15700 ) | ( n15698 & n15700 ) ;
  assign n15702 = ( n8113 & ~n9605 ) | ( n8113 & n12356 ) | ( ~n9605 & n12356 ) ;
  assign n15703 = n15702 ^ n5827 ^ 1'b0 ;
  assign n15704 = n14310 ^ n4191 ^ n1578 ;
  assign n15714 = n8720 ^ n5892 ^ n5396 ;
  assign n15711 = n8664 ^ n6038 ^ n5442 ;
  assign n15712 = ( n5439 & n7244 ) | ( n5439 & n15711 ) | ( n7244 & n15711 ) ;
  assign n15713 = n15712 ^ n5491 ^ 1'b0 ;
  assign n15705 = n3819 ^ n2689 ^ n523 ;
  assign n15706 = n7165 ^ n1490 ^ 1'b0 ;
  assign n15707 = ~n15705 & n15706 ;
  assign n15708 = n7308 ^ n5983 ^ 1'b0 ;
  assign n15709 = ( ~x40 & n7731 ) | ( ~x40 & n15708 ) | ( n7731 & n15708 ) ;
  assign n15710 = ( n13896 & n15707 ) | ( n13896 & n15709 ) | ( n15707 & n15709 ) ;
  assign n15715 = n15714 ^ n15713 ^ n15710 ;
  assign n15716 = n15704 | n15715 ;
  assign n15717 = n8068 ^ n7368 ^ n5803 ;
  assign n15718 = ( ~n7289 & n12056 ) | ( ~n7289 & n15717 ) | ( n12056 & n15717 ) ;
  assign n15719 = n10072 ^ n9858 ^ n5950 ;
  assign n15720 = n7956 ^ n7931 ^ n6861 ;
  assign n15721 = ( n11481 & ~n15719 ) | ( n11481 & n15720 ) | ( ~n15719 & n15720 ) ;
  assign n15722 = ( n2905 & ~n4984 ) | ( n2905 & n5295 ) | ( ~n4984 & n5295 ) ;
  assign n15723 = n12747 ^ n8374 ^ n4858 ;
  assign n15724 = ( n2443 & ~n4844 ) | ( n2443 & n13196 ) | ( ~n4844 & n13196 ) ;
  assign n15725 = n2259 & ~n15724 ;
  assign n15726 = n15723 & n15725 ;
  assign n15727 = ( n1712 & n7576 ) | ( n1712 & ~n14748 ) | ( n7576 & ~n14748 ) ;
  assign n15728 = n11356 ^ n3312 ^ n688 ;
  assign n15729 = n15728 ^ n2919 ^ n2455 ;
  assign n15730 = n15729 ^ n7669 ^ n1997 ;
  assign n15731 = ( ~n4027 & n15727 ) | ( ~n4027 & n15730 ) | ( n15727 & n15730 ) ;
  assign n15732 = n819 & n1337 ;
  assign n15733 = n15732 ^ n10979 ^ n1531 ;
  assign n15734 = ( n2391 & n7101 ) | ( n2391 & ~n8970 ) | ( n7101 & ~n8970 ) ;
  assign n15735 = n7247 ^ n5715 ^ n5360 ;
  assign n15736 = n14063 ^ n13717 ^ n13530 ;
  assign n15737 = n1362 & n15736 ;
  assign n15738 = ( ~n6686 & n15735 ) | ( ~n6686 & n15737 ) | ( n15735 & n15737 ) ;
  assign n15739 = ( n7192 & ~n15734 ) | ( n7192 & n15738 ) | ( ~n15734 & n15738 ) ;
  assign n15740 = n8042 ^ n8007 ^ 1'b0 ;
  assign n15741 = ~n2603 & n15740 ;
  assign n15742 = n15741 ^ n3746 ^ n2727 ;
  assign n15749 = n5649 ^ n4455 ^ n2431 ;
  assign n15748 = n13760 ^ n10746 ^ n8859 ;
  assign n15743 = n9514 ^ n3917 ^ 1'b0 ;
  assign n15744 = n8668 | n15743 ;
  assign n15745 = n4103 & ~n11235 ;
  assign n15746 = n15745 ^ n1841 ^ 1'b0 ;
  assign n15747 = ( ~n12895 & n15744 ) | ( ~n12895 & n15746 ) | ( n15744 & n15746 ) ;
  assign n15750 = n15749 ^ n15748 ^ n15747 ;
  assign n15751 = n9852 ^ n2587 ^ 1'b0 ;
  assign n15752 = ~n5853 & n15751 ;
  assign n15753 = ( n415 & n2139 ) | ( n415 & ~n15752 ) | ( n2139 & ~n15752 ) ;
  assign n15754 = n15753 ^ n15064 ^ 1'b0 ;
  assign n15755 = n14536 ^ n12967 ^ n9591 ;
  assign n15756 = n13423 ^ n9716 ^ n5765 ;
  assign n15757 = n8060 ^ n290 ^ 1'b0 ;
  assign n15758 = ( ~n1173 & n3612 ) | ( ~n1173 & n8929 ) | ( n3612 & n8929 ) ;
  assign n15759 = ( ~n8758 & n9361 ) | ( ~n8758 & n15758 ) | ( n9361 & n15758 ) ;
  assign n15760 = ( n5485 & n6746 ) | ( n5485 & n15150 ) | ( n6746 & n15150 ) ;
  assign n15761 = ~n4954 & n13283 ;
  assign n15762 = n12192 & n15761 ;
  assign n15763 = ( ~n11982 & n15760 ) | ( ~n11982 & n15762 ) | ( n15760 & n15762 ) ;
  assign n15764 = n14155 ^ n8022 ^ n1615 ;
  assign n15765 = n4559 & ~n15764 ;
  assign n15766 = ~n341 & n15765 ;
  assign n15767 = n8645 ^ x130 ^ 1'b0 ;
  assign n15768 = n15767 ^ n7350 ^ n6581 ;
  assign n15769 = ( ~n4021 & n7634 ) | ( ~n4021 & n10636 ) | ( n7634 & n10636 ) ;
  assign n15770 = n15769 ^ n9173 ^ n827 ;
  assign n15771 = ( n11731 & n13354 ) | ( n11731 & n15770 ) | ( n13354 & n15770 ) ;
  assign n15782 = n5831 ^ n5490 ^ n3304 ;
  assign n15779 = n13814 ^ n12047 ^ n6319 ;
  assign n15780 = n15779 ^ n4820 ^ 1'b0 ;
  assign n15781 = ~n9570 & n15780 ;
  assign n15775 = ( n450 & n4549 ) | ( n450 & n5834 ) | ( n4549 & n5834 ) ;
  assign n15773 = n1893 & n8524 ;
  assign n15774 = n7335 | n15773 ;
  assign n15776 = n15775 ^ n15774 ^ 1'b0 ;
  assign n15777 = ( n2335 & ~n7276 ) | ( n2335 & n15776 ) | ( ~n7276 & n15776 ) ;
  assign n15772 = n3661 & ~n5064 ;
  assign n15778 = n15777 ^ n15772 ^ 1'b0 ;
  assign n15783 = n15782 ^ n15781 ^ n15778 ;
  assign n15784 = x151 | n1704 ;
  assign n15785 = ( n11478 & n11810 ) | ( n11478 & ~n15784 ) | ( n11810 & ~n15784 ) ;
  assign n15786 = n12700 ^ n9575 ^ 1'b0 ;
  assign n15787 = n1421 & ~n1427 ;
  assign n15788 = n15787 ^ n1512 ^ 1'b0 ;
  assign n15789 = n368 & n15788 ;
  assign n15790 = n15789 ^ n6183 ^ 1'b0 ;
  assign n15791 = n1559 & ~n5053 ;
  assign n15792 = ( n4095 & ~n15790 ) | ( n4095 & n15791 ) | ( ~n15790 & n15791 ) ;
  assign n15793 = ( n2386 & ~n5465 ) | ( n2386 & n13219 ) | ( ~n5465 & n13219 ) ;
  assign n15794 = n15793 ^ n2097 ^ x192 ;
  assign n15795 = ( ~x247 & n15792 ) | ( ~x247 & n15794 ) | ( n15792 & n15794 ) ;
  assign n15796 = ~n1559 & n12381 ;
  assign n15797 = n15498 ^ x185 ^ 1'b0 ;
  assign n15798 = n602 & n15797 ;
  assign n15799 = n4303 ^ n2580 ^ n1031 ;
  assign n15800 = n7383 ^ n4262 ^ 1'b0 ;
  assign n15801 = n15800 ^ n10133 ^ n7467 ;
  assign n15802 = ( ~n4493 & n11057 ) | ( ~n4493 & n15801 ) | ( n11057 & n15801 ) ;
  assign n15804 = n2235 | n4636 ;
  assign n15805 = n8241 | n15804 ;
  assign n15803 = n9236 ^ n8752 ^ 1'b0 ;
  assign n15806 = n15805 ^ n15803 ^ n12793 ;
  assign n15807 = ( x177 & ~n4954 ) | ( x177 & n5501 ) | ( ~n4954 & n5501 ) ;
  assign n15808 = n15807 ^ n7919 ^ n1709 ;
  assign n15809 = ( n7134 & ~n15806 ) | ( n7134 & n15808 ) | ( ~n15806 & n15808 ) ;
  assign n15811 = n4540 ^ n2492 ^ n2377 ;
  assign n15810 = n2035 ^ n1342 ^ n1189 ;
  assign n15812 = n15811 ^ n15810 ^ n11337 ;
  assign n15813 = ~n13357 & n15812 ;
  assign n15814 = n10338 & n15813 ;
  assign n15815 = ( x190 & n3267 ) | ( x190 & n9991 ) | ( n3267 & n9991 ) ;
  assign n15816 = ( n555 & n3724 ) | ( n555 & ~n9414 ) | ( n3724 & ~n9414 ) ;
  assign n15817 = ( ~n6357 & n11049 ) | ( ~n6357 & n15816 ) | ( n11049 & n15816 ) ;
  assign n15818 = ( n7087 & n15815 ) | ( n7087 & n15817 ) | ( n15815 & n15817 ) ;
  assign n15819 = ( n3047 & ~n4243 ) | ( n3047 & n6816 ) | ( ~n4243 & n6816 ) ;
  assign n15820 = ( n8249 & n14155 ) | ( n8249 & n15819 ) | ( n14155 & n15819 ) ;
  assign n15821 = n15820 ^ n14192 ^ x161 ;
  assign n15822 = ( n6070 & n15818 ) | ( n6070 & n15821 ) | ( n15818 & n15821 ) ;
  assign n15823 = n10086 & ~n13976 ;
  assign n15824 = n15823 ^ n491 ^ 1'b0 ;
  assign n15825 = n15230 & n15824 ;
  assign n15826 = ( n2742 & n4873 ) | ( n2742 & ~n8827 ) | ( n4873 & ~n8827 ) ;
  assign n15827 = n15826 ^ n10751 ^ 1'b0 ;
  assign n15828 = ( ~n1717 & n7706 ) | ( ~n1717 & n11792 ) | ( n7706 & n11792 ) ;
  assign n15829 = n5500 | n15828 ;
  assign n15830 = n15829 ^ n9900 ^ 1'b0 ;
  assign n15831 = ( n11647 & n15807 ) | ( n11647 & ~n15830 ) | ( n15807 & ~n15830 ) ;
  assign n15832 = n12045 ^ n8429 ^ 1'b0 ;
  assign n15833 = n12867 | n15832 ;
  assign n15834 = n11699 ^ n10643 ^ n3515 ;
  assign n15835 = n15834 ^ n14512 ^ n5884 ;
  assign n15836 = ( ~n5449 & n6874 ) | ( ~n5449 & n9931 ) | ( n6874 & n9931 ) ;
  assign n15837 = n15836 ^ n9119 ^ 1'b0 ;
  assign n15840 = n4094 ^ n2585 ^ n304 ;
  assign n15838 = ( n3022 & n5448 ) | ( n3022 & ~n5502 ) | ( n5448 & ~n5502 ) ;
  assign n15839 = x193 & ~n15838 ;
  assign n15841 = n15840 ^ n15839 ^ 1'b0 ;
  assign n15842 = ( n2964 & n13861 ) | ( n2964 & ~n15841 ) | ( n13861 & ~n15841 ) ;
  assign n15843 = ~n1347 & n15842 ;
  assign n15844 = ~n15837 & n15843 ;
  assign n15845 = ( n6608 & n15835 ) | ( n6608 & n15844 ) | ( n15835 & n15844 ) ;
  assign n15849 = n9006 ^ n6010 ^ n2217 ;
  assign n15846 = n4658 & n4748 ;
  assign n15847 = ( ~n4962 & n11814 ) | ( ~n4962 & n12490 ) | ( n11814 & n12490 ) ;
  assign n15848 = ( ~n7811 & n15846 ) | ( ~n7811 & n15847 ) | ( n15846 & n15847 ) ;
  assign n15850 = n15849 ^ n15848 ^ n9865 ;
  assign n15851 = ( ~n15833 & n15845 ) | ( ~n15833 & n15850 ) | ( n15845 & n15850 ) ;
  assign n15852 = n7807 ^ n5450 ^ 1'b0 ;
  assign n15853 = n12815 ^ n7545 ^ 1'b0 ;
  assign n15854 = n15852 & ~n15853 ;
  assign n15855 = n15854 ^ n2795 ^ n2738 ;
  assign n15856 = n7657 ^ n7350 ^ n1461 ;
  assign n15857 = n15856 ^ n3037 ^ n2913 ;
  assign n15858 = ( n7518 & n15855 ) | ( n7518 & n15857 ) | ( n15855 & n15857 ) ;
  assign n15863 = n2479 ^ n1137 ^ x217 ;
  assign n15861 = n848 & ~n5343 ;
  assign n15859 = n7260 ^ n2723 ^ 1'b0 ;
  assign n15860 = ~n12246 & n15859 ;
  assign n15862 = n15861 ^ n15860 ^ n5650 ;
  assign n15864 = n15863 ^ n15862 ^ n7838 ;
  assign n15865 = ( n2279 & n4605 ) | ( n2279 & n15864 ) | ( n4605 & n15864 ) ;
  assign n15866 = ( n6332 & ~n6378 ) | ( n6332 & n8894 ) | ( ~n6378 & n8894 ) ;
  assign n15867 = n15866 ^ n10548 ^ n5155 ;
  assign n15868 = n15867 ^ n5324 ^ x4 ;
  assign n15869 = n5659 & n15868 ;
  assign n15870 = n8501 ^ n7196 ^ n4498 ;
  assign n15871 = ( n3605 & n9498 ) | ( n3605 & n15870 ) | ( n9498 & n15870 ) ;
  assign n15872 = ( ~n14002 & n15746 ) | ( ~n14002 & n15871 ) | ( n15746 & n15871 ) ;
  assign n15873 = n1189 & ~n15872 ;
  assign n15874 = n15873 ^ n13208 ^ n11172 ;
  assign n15878 = n13803 ^ n6366 ^ n3296 ;
  assign n15879 = n15878 ^ n4605 ^ n3526 ;
  assign n15880 = n2716 ^ n491 ^ x79 ;
  assign n15881 = n15880 ^ n10760 ^ n5576 ;
  assign n15882 = ( n11286 & n15879 ) | ( n11286 & n15881 ) | ( n15879 & n15881 ) ;
  assign n15875 = n2274 & n4627 ;
  assign n15876 = n15875 ^ n6640 ^ n486 ;
  assign n15877 = n15876 ^ n8852 ^ n7020 ;
  assign n15883 = n15882 ^ n15877 ^ n6346 ;
  assign n15884 = ( ~n1199 & n4916 ) | ( ~n1199 & n8621 ) | ( n4916 & n8621 ) ;
  assign n15885 = n3691 & n9155 ;
  assign n15886 = ~n4437 & n15885 ;
  assign n15887 = ( n3015 & n4047 ) | ( n3015 & n15886 ) | ( n4047 & n15886 ) ;
  assign n15888 = ( ~n1255 & n15884 ) | ( ~n1255 & n15887 ) | ( n15884 & n15887 ) ;
  assign n15889 = ( x69 & n15319 ) | ( x69 & n15888 ) | ( n15319 & n15888 ) ;
  assign n15890 = ~n10263 & n15889 ;
  assign n15891 = n4788 & n15890 ;
  assign n15892 = ( n4343 & n6234 ) | ( n4343 & n14715 ) | ( n6234 & n14715 ) ;
  assign n15893 = ~n4648 & n15892 ;
  assign n15894 = ( n585 & n1259 ) | ( n585 & ~n5433 ) | ( n1259 & ~n5433 ) ;
  assign n15895 = n15894 ^ n6486 ^ n3803 ;
  assign n15902 = n2860 & n3615 ;
  assign n15903 = n15902 ^ n6420 ^ 1'b0 ;
  assign n15896 = n15544 ^ n1099 ^ 1'b0 ;
  assign n15897 = n4843 & ~n15896 ;
  assign n15898 = ( ~n6073 & n6596 ) | ( ~n6073 & n8385 ) | ( n6596 & n8385 ) ;
  assign n15899 = n13216 & ~n15898 ;
  assign n15900 = n15899 ^ n843 ^ 1'b0 ;
  assign n15901 = ( n7353 & n15897 ) | ( n7353 & ~n15900 ) | ( n15897 & ~n15900 ) ;
  assign n15904 = n15903 ^ n15901 ^ n6531 ;
  assign n15905 = n11557 ^ n9182 ^ n2777 ;
  assign n15906 = n15905 ^ n8951 ^ n6398 ;
  assign n15907 = ( ~n15895 & n15904 ) | ( ~n15895 & n15906 ) | ( n15904 & n15906 ) ;
  assign n15908 = n13494 ^ n2288 ^ n1934 ;
  assign n15909 = ( n268 & n7597 ) | ( n268 & n15908 ) | ( n7597 & n15908 ) ;
  assign n15910 = n9841 & ~n15909 ;
  assign n15911 = ( x76 & ~n1846 ) | ( x76 & n3682 ) | ( ~n1846 & n3682 ) ;
  assign n15912 = n15911 ^ n10111 ^ n6709 ;
  assign n15913 = ( n4698 & ~n7666 ) | ( n4698 & n10680 ) | ( ~n7666 & n10680 ) ;
  assign n15914 = n15913 ^ n4060 ^ 1'b0 ;
  assign n15915 = n11205 ^ n5195 ^ n3632 ;
  assign n15916 = n15915 ^ n2094 ^ 1'b0 ;
  assign n15917 = n4042 & n15916 ;
  assign n15918 = n15917 ^ n10818 ^ n1954 ;
  assign n15925 = n4504 ^ n1430 ^ x166 ;
  assign n15926 = n15925 ^ n7789 ^ n3006 ;
  assign n15927 = ( n2456 & ~n8216 ) | ( n2456 & n15926 ) | ( ~n8216 & n15926 ) ;
  assign n15920 = n1896 & ~n5244 ;
  assign n15921 = ~n4283 & n15920 ;
  assign n15922 = n15921 ^ n5563 ^ n1379 ;
  assign n15923 = n15922 ^ n13266 ^ n8911 ;
  assign n15924 = n15923 ^ n8853 ^ n7975 ;
  assign n15919 = ( n4070 & n8573 ) | ( n4070 & ~n13202 ) | ( n8573 & ~n13202 ) ;
  assign n15928 = n15927 ^ n15924 ^ n15919 ;
  assign n15929 = ( ~x171 & n10118 ) | ( ~x171 & n13485 ) | ( n10118 & n13485 ) ;
  assign n15930 = n1598 & n13727 ;
  assign n15934 = n3942 ^ n2538 ^ n2141 ;
  assign n15935 = n15934 ^ n965 ^ 1'b0 ;
  assign n15931 = n4935 & ~n8872 ;
  assign n15932 = n15931 ^ n7253 ^ 1'b0 ;
  assign n15933 = ~x10 & n15932 ;
  assign n15936 = n15935 ^ n15933 ^ n13509 ;
  assign n15939 = n7643 ^ n4718 ^ n3627 ;
  assign n15940 = n15939 ^ n5424 ^ n3971 ;
  assign n15937 = ( n3211 & n6587 ) | ( n3211 & ~n6717 ) | ( n6587 & ~n6717 ) ;
  assign n15938 = n15937 ^ n14973 ^ 1'b0 ;
  assign n15941 = n15940 ^ n15938 ^ n2530 ;
  assign n15942 = n12771 & n15941 ;
  assign n15943 = n10773 ^ n3865 ^ 1'b0 ;
  assign n15944 = n10740 ^ n3483 ^ n1072 ;
  assign n15945 = n3652 | n15944 ;
  assign n15946 = n13703 ^ n1799 ^ 1'b0 ;
  assign n15947 = n9739 & ~n15946 ;
  assign n15948 = ( n15943 & ~n15945 ) | ( n15943 & n15947 ) | ( ~n15945 & n15947 ) ;
  assign n15949 = n15948 ^ n6403 ^ 1'b0 ;
  assign n15950 = n15942 & ~n15949 ;
  assign n15951 = n7844 ^ n6638 ^ n3872 ;
  assign n15952 = ( x185 & n6286 ) | ( x185 & ~n15951 ) | ( n6286 & ~n15951 ) ;
  assign n15953 = ( n971 & n4675 ) | ( n971 & n8301 ) | ( n4675 & n8301 ) ;
  assign n15954 = n2782 & ~n15953 ;
  assign n15955 = ~n15952 & n15954 ;
  assign n15956 = ~n11770 & n15955 ;
  assign n15957 = n6426 ^ n2925 ^ 1'b0 ;
  assign n15958 = x204 & n15957 ;
  assign n15959 = n15958 ^ n3202 ^ n801 ;
  assign n15960 = n5463 ^ n1395 ^ 1'b0 ;
  assign n15961 = ( n6640 & n10164 ) | ( n6640 & ~n15960 ) | ( n10164 & ~n15960 ) ;
  assign n15962 = ( n8283 & n15959 ) | ( n8283 & ~n15961 ) | ( n15959 & ~n15961 ) ;
  assign n15964 = n1220 & ~n1281 ;
  assign n15965 = n2608 & n15964 ;
  assign n15966 = n2651 | n15965 ;
  assign n15967 = n15966 ^ n382 ^ 1'b0 ;
  assign n15963 = ( n6908 & n8737 ) | ( n6908 & n14048 ) | ( n8737 & n14048 ) ;
  assign n15968 = n15967 ^ n15963 ^ n8548 ;
  assign n15969 = n8793 ^ n8297 ^ n901 ;
  assign n15970 = ( n2613 & n8970 ) | ( n2613 & ~n15969 ) | ( n8970 & ~n15969 ) ;
  assign n15971 = ( n6013 & n8710 ) | ( n6013 & ~n15970 ) | ( n8710 & ~n15970 ) ;
  assign n15972 = n9151 ^ n4228 ^ n1093 ;
  assign n15973 = ( n3926 & ~n5872 ) | ( n3926 & n15972 ) | ( ~n5872 & n15972 ) ;
  assign n15974 = n10167 ^ n10022 ^ n4000 ;
  assign n15975 = ( ~n9844 & n15973 ) | ( ~n9844 & n15974 ) | ( n15973 & n15974 ) ;
  assign n15976 = n12324 ^ n12237 ^ n9819 ;
  assign n15977 = n6819 & ~n15976 ;
  assign n15978 = n7739 ^ n1638 ^ 1'b0 ;
  assign n15979 = n9483 & ~n10650 ;
  assign n15980 = n13841 & n15979 ;
  assign n15981 = n6483 | n15980 ;
  assign n15982 = n15981 ^ n14339 ^ 1'b0 ;
  assign n15983 = ( ~n7846 & n11477 ) | ( ~n7846 & n15982 ) | ( n11477 & n15982 ) ;
  assign n15984 = ( x69 & n14384 ) | ( x69 & ~n15983 ) | ( n14384 & ~n15983 ) ;
  assign n15985 = ~n15816 & n15984 ;
  assign n15986 = ( n9541 & n15978 ) | ( n9541 & n15985 ) | ( n15978 & n15985 ) ;
  assign n15987 = ( n12246 & n15977 ) | ( n12246 & ~n15986 ) | ( n15977 & ~n15986 ) ;
  assign n15990 = n8429 ^ n1009 ^ n665 ;
  assign n15991 = ( n3748 & n9147 ) | ( n3748 & n15990 ) | ( n9147 & n15990 ) ;
  assign n15988 = n13831 ^ n4582 ^ n1077 ;
  assign n15989 = n15988 ^ n15169 ^ n5798 ;
  assign n15992 = n15991 ^ n15989 ^ 1'b0 ;
  assign n15993 = ( n5437 & ~n5956 ) | ( n5437 & n12964 ) | ( ~n5956 & n12964 ) ;
  assign n15994 = n15846 ^ n402 ^ 1'b0 ;
  assign n15995 = n2129 & ~n15994 ;
  assign n15996 = ( n3206 & n4218 ) | ( n3206 & n8071 ) | ( n4218 & n8071 ) ;
  assign n15997 = n15996 ^ n8412 ^ n7183 ;
  assign n15998 = n15997 ^ n1510 ^ 1'b0 ;
  assign n15999 = n2235 | n15998 ;
  assign n16000 = x59 & n2425 ;
  assign n16001 = ~x221 & n16000 ;
  assign n16007 = n12027 ^ n1754 ^ n796 ;
  assign n16008 = ~n7909 & n16007 ;
  assign n16004 = ( n818 & n1327 ) | ( n818 & n1684 ) | ( n1327 & n1684 ) ;
  assign n16002 = n10583 ^ n5341 ^ n3331 ;
  assign n16003 = n16002 ^ n14840 ^ n4214 ;
  assign n16005 = n16004 ^ n16003 ^ n6106 ;
  assign n16006 = ( n1413 & n8442 ) | ( n1413 & ~n16005 ) | ( n8442 & ~n16005 ) ;
  assign n16009 = n16008 ^ n16006 ^ n3924 ;
  assign n16010 = n7295 ^ n6281 ^ n5742 ;
  assign n16011 = n16010 ^ n15637 ^ n3380 ;
  assign n16012 = n16011 ^ n8121 ^ n1849 ;
  assign n16013 = ( ~n16001 & n16009 ) | ( ~n16001 & n16012 ) | ( n16009 & n16012 ) ;
  assign n16030 = ( n1533 & ~n1707 ) | ( n1533 & n3204 ) | ( ~n1707 & n3204 ) ;
  assign n16031 = ( n1158 & n2347 ) | ( n1158 & ~n16030 ) | ( n2347 & ~n16030 ) ;
  assign n16028 = ( n522 & n1745 ) | ( n522 & n4412 ) | ( n1745 & n4412 ) ;
  assign n16029 = n16028 ^ n9435 ^ n8158 ;
  assign n16032 = n16031 ^ n16029 ^ n12731 ;
  assign n16022 = ( n426 & n5659 ) | ( n426 & ~n7886 ) | ( n5659 & ~n7886 ) ;
  assign n16023 = n16022 ^ n9891 ^ n3042 ;
  assign n16021 = n10162 ^ n8627 ^ n3602 ;
  assign n16024 = n16023 ^ n16021 ^ n8986 ;
  assign n16025 = n15497 ^ n11463 ^ n9162 ;
  assign n16026 = ~n341 & n16025 ;
  assign n16027 = n16024 & n16026 ;
  assign n16019 = n5499 | n12150 ;
  assign n16017 = n11962 ^ n9741 ^ n2063 ;
  assign n16014 = n902 | n4917 ;
  assign n16015 = n16014 ^ n9970 ^ 1'b0 ;
  assign n16016 = n16015 ^ n2626 ^ 1'b0 ;
  assign n16018 = n16017 ^ n16016 ^ n4407 ;
  assign n16020 = n16019 ^ n16018 ^ n14149 ;
  assign n16033 = n16032 ^ n16027 ^ n16020 ;
  assign n16034 = n5072 ^ n4159 ^ n2311 ;
  assign n16035 = ( ~n8522 & n15471 ) | ( ~n8522 & n16034 ) | ( n15471 & n16034 ) ;
  assign n16036 = ( ~n3773 & n11234 ) | ( ~n3773 & n16035 ) | ( n11234 & n16035 ) ;
  assign n16038 = ( n2049 & n2744 ) | ( n2049 & n2781 ) | ( n2744 & n2781 ) ;
  assign n16039 = ( x190 & ~n5376 ) | ( x190 & n16038 ) | ( ~n5376 & n16038 ) ;
  assign n16037 = ( n10538 & ~n11528 ) | ( n10538 & n14428 ) | ( ~n11528 & n14428 ) ;
  assign n16040 = n16039 ^ n16037 ^ n8212 ;
  assign n16041 = n16040 ^ n6903 ^ 1'b0 ;
  assign n16042 = ( n1004 & ~n5251 ) | ( n1004 & n5400 ) | ( ~n5251 & n5400 ) ;
  assign n16043 = ( ~n6506 & n11507 ) | ( ~n6506 & n16042 ) | ( n11507 & n16042 ) ;
  assign n16044 = n16043 ^ n10949 ^ n8598 ;
  assign n16045 = ( n1321 & n2279 ) | ( n1321 & ~n4557 ) | ( n2279 & ~n4557 ) ;
  assign n16061 = n4525 ^ n793 ^ n404 ;
  assign n16057 = n9856 ^ n4599 ^ 1'b0 ;
  assign n16058 = n5024 | n16057 ;
  assign n16059 = ( n13498 & n13768 ) | ( n13498 & n16058 ) | ( n13768 & n16058 ) ;
  assign n16060 = ( ~n3072 & n7988 ) | ( ~n3072 & n16059 ) | ( n7988 & n16059 ) ;
  assign n16054 = n1596 & ~n3907 ;
  assign n16055 = n16054 ^ n3520 ^ n1795 ;
  assign n16052 = n6369 & n10197 ;
  assign n16053 = n8739 & n16052 ;
  assign n16056 = n16055 ^ n16053 ^ n656 ;
  assign n16062 = n16061 ^ n16060 ^ n16056 ;
  assign n16046 = n2314 ^ n884 ^ 1'b0 ;
  assign n16047 = n13030 | n16046 ;
  assign n16048 = n8170 ^ n3282 ^ 1'b0 ;
  assign n16049 = ~n16047 & n16048 ;
  assign n16050 = n16049 ^ n2735 ^ n2427 ;
  assign n16051 = ( n11153 & n11315 ) | ( n11153 & ~n16050 ) | ( n11315 & ~n16050 ) ;
  assign n16063 = n16062 ^ n16051 ^ n12517 ;
  assign n16064 = ( n4319 & n16045 ) | ( n4319 & ~n16063 ) | ( n16045 & ~n16063 ) ;
  assign n16066 = ( n1142 & n3525 ) | ( n1142 & ~n9928 ) | ( n3525 & ~n9928 ) ;
  assign n16067 = n16066 ^ n15317 ^ n2112 ;
  assign n16068 = n8978 ^ n1781 ^ n1706 ;
  assign n16069 = n16068 ^ n11646 ^ n9278 ;
  assign n16070 = ( n1639 & n13512 ) | ( n1639 & n16069 ) | ( n13512 & n16069 ) ;
  assign n16071 = ( n855 & ~n2640 ) | ( n855 & n16070 ) | ( ~n2640 & n16070 ) ;
  assign n16072 = ( n1475 & n3687 ) | ( n1475 & n16071 ) | ( n3687 & n16071 ) ;
  assign n16073 = ( n13112 & ~n16067 ) | ( n13112 & n16072 ) | ( ~n16067 & n16072 ) ;
  assign n16065 = n8751 & n15202 ;
  assign n16074 = n16073 ^ n16065 ^ 1'b0 ;
  assign n16075 = ( ~n3858 & n5321 ) | ( ~n3858 & n8422 ) | ( n5321 & n8422 ) ;
  assign n16076 = ( n2719 & ~n10225 ) | ( n2719 & n10295 ) | ( ~n10225 & n10295 ) ;
  assign n16077 = n16075 & n16076 ;
  assign n16078 = n12989 & n16077 ;
  assign n16079 = n12441 ^ n3290 ^ n3242 ;
  assign n16080 = n12005 | n16079 ;
  assign n16081 = n13567 ^ n4586 ^ n3110 ;
  assign n16082 = n16081 ^ n9280 ^ n3274 ;
  assign n16083 = ( ~x244 & n14524 ) | ( ~x244 & n16082 ) | ( n14524 & n16082 ) ;
  assign n16084 = ( ~n4770 & n6432 ) | ( ~n4770 & n7169 ) | ( n6432 & n7169 ) ;
  assign n16085 = ( n6168 & n7590 ) | ( n6168 & ~n16084 ) | ( n7590 & ~n16084 ) ;
  assign n16086 = n9037 ^ n6361 ^ n1698 ;
  assign n16087 = n7660 ^ n824 ^ x201 ;
  assign n16088 = ( n9095 & n16086 ) | ( n9095 & n16087 ) | ( n16086 & n16087 ) ;
  assign n16089 = n10492 ^ n2491 ^ n884 ;
  assign n16105 = ( n430 & n710 ) | ( n430 & n9682 ) | ( n710 & n9682 ) ;
  assign n16106 = ( n7527 & n8203 ) | ( n7527 & ~n16105 ) | ( n8203 & ~n16105 ) ;
  assign n16102 = n15879 ^ n11013 ^ n2578 ;
  assign n16103 = n16102 ^ n7518 ^ n6766 ;
  assign n16104 = ~n11364 & n16103 ;
  assign n16090 = ( n1813 & n4267 ) | ( n1813 & n11272 ) | ( n4267 & n11272 ) ;
  assign n16091 = ( n1563 & n5977 ) | ( n1563 & ~n16090 ) | ( n5977 & ~n16090 ) ;
  assign n16092 = n14067 ^ n9433 ^ n1164 ;
  assign n16093 = n16092 ^ n12662 ^ 1'b0 ;
  assign n16094 = ~n12067 & n16093 ;
  assign n16095 = n8924 ^ n430 ^ 1'b0 ;
  assign n16096 = n16095 ^ n6440 ^ n3592 ;
  assign n16097 = ( x150 & n4581 ) | ( x150 & n5835 ) | ( n4581 & n5835 ) ;
  assign n16098 = n16097 ^ n15826 ^ 1'b0 ;
  assign n16099 = n2841 | n16098 ;
  assign n16100 = ( n6189 & ~n16096 ) | ( n6189 & n16099 ) | ( ~n16096 & n16099 ) ;
  assign n16101 = ( n16091 & ~n16094 ) | ( n16091 & n16100 ) | ( ~n16094 & n16100 ) ;
  assign n16107 = n16106 ^ n16104 ^ n16101 ;
  assign n16108 = ( n2113 & n8340 ) | ( n2113 & ~n13716 ) | ( n8340 & ~n13716 ) ;
  assign n16109 = n14816 ^ n11296 ^ n5416 ;
  assign n16110 = ( n8987 & n9232 ) | ( n8987 & n16109 ) | ( n9232 & n16109 ) ;
  assign n16111 = n2711 & ~n9212 ;
  assign n16112 = n16111 ^ n3373 ^ 1'b0 ;
  assign n16113 = n16110 | n16112 ;
  assign n16114 = ( n437 & ~n1911 ) | ( n437 & n3164 ) | ( ~n1911 & n3164 ) ;
  assign n16115 = n16114 ^ n3224 ^ n2602 ;
  assign n16116 = ( n799 & n8785 ) | ( n799 & ~n16115 ) | ( n8785 & ~n16115 ) ;
  assign n16117 = n3773 ^ n3058 ^ n1694 ;
  assign n16118 = n16117 ^ n7214 ^ x75 ;
  assign n16119 = ( n669 & n16116 ) | ( n669 & n16118 ) | ( n16116 & n16118 ) ;
  assign n16120 = n11233 & n16119 ;
  assign n16121 = ( ~n9500 & n12841 ) | ( ~n9500 & n16120 ) | ( n12841 & n16120 ) ;
  assign n16123 = n10477 ^ n8508 ^ 1'b0 ;
  assign n16124 = n4496 & ~n16123 ;
  assign n16122 = ( x82 & x232 ) | ( x82 & n9555 ) | ( x232 & n9555 ) ;
  assign n16125 = n16124 ^ n16122 ^ n8464 ;
  assign n16126 = n16125 ^ n9645 ^ 1'b0 ;
  assign n16127 = ( n5993 & n10230 ) | ( n5993 & ~n16126 ) | ( n10230 & ~n16126 ) ;
  assign n16129 = ( n1489 & n5135 ) | ( n1489 & ~n12743 ) | ( n5135 & ~n12743 ) ;
  assign n16130 = n13175 ^ n4744 ^ n3832 ;
  assign n16131 = ( n3857 & n16129 ) | ( n3857 & n16130 ) | ( n16129 & n16130 ) ;
  assign n16128 = n15317 ^ n5973 ^ n3101 ;
  assign n16132 = n16131 ^ n16128 ^ n14449 ;
  assign n16133 = ( n1556 & n5332 ) | ( n1556 & ~n6691 ) | ( n5332 & ~n6691 ) ;
  assign n16134 = n16133 ^ n6346 ^ n1284 ;
  assign n16135 = n16134 ^ n12161 ^ n4585 ;
  assign n16136 = ( n14612 & n14895 ) | ( n14612 & n16135 ) | ( n14895 & n16135 ) ;
  assign n16137 = ( n981 & n2697 ) | ( n981 & ~n16136 ) | ( n2697 & ~n16136 ) ;
  assign n16138 = n16137 ^ n14758 ^ n3980 ;
  assign n16139 = ( n2344 & n13726 ) | ( n2344 & ~n16138 ) | ( n13726 & ~n16138 ) ;
  assign n16140 = n9159 ^ n6137 ^ n4578 ;
  assign n16141 = n16140 ^ n6275 ^ n3522 ;
  assign n16142 = ( x146 & ~x249 ) | ( x146 & n6654 ) | ( ~x249 & n6654 ) ;
  assign n16143 = n16141 & n16142 ;
  assign n16144 = ~n15660 & n16143 ;
  assign n16145 = n16139 | n16144 ;
  assign n16146 = n16145 ^ n11167 ^ 1'b0 ;
  assign n16147 = n16146 ^ n8457 ^ n1795 ;
  assign n16148 = n12627 ^ n4952 ^ n2959 ;
  assign n16149 = x196 & ~n2014 ;
  assign n16150 = ~n16148 & n16149 ;
  assign n16151 = n16150 ^ n13601 ^ n2623 ;
  assign n16152 = n7238 ^ n6741 ^ n3842 ;
  assign n16153 = n16152 ^ n11800 ^ n11473 ;
  assign n16154 = n16153 ^ n728 ^ 1'b0 ;
  assign n16155 = n16151 & ~n16154 ;
  assign n16160 = ( n5679 & ~n10580 ) | ( n5679 & n10892 ) | ( ~n10580 & n10892 ) ;
  assign n16161 = n16160 ^ n13895 ^ n470 ;
  assign n16156 = ( n5716 & n8025 ) | ( n5716 & n8668 ) | ( n8025 & n8668 ) ;
  assign n16157 = n11876 ^ n3720 ^ n2230 ;
  assign n16158 = ~n1056 & n16157 ;
  assign n16159 = ( n4072 & n16156 ) | ( n4072 & n16158 ) | ( n16156 & n16158 ) ;
  assign n16162 = n16161 ^ n16159 ^ n11945 ;
  assign n16163 = n16162 ^ n14195 ^ n2975 ;
  assign n16164 = n10304 ^ n7094 ^ n2299 ;
  assign n16165 = n16164 ^ n15240 ^ n3601 ;
  assign n16166 = ( ~n4390 & n15159 ) | ( ~n4390 & n16165 ) | ( n15159 & n16165 ) ;
  assign n16171 = n4094 ^ n3878 ^ 1'b0 ;
  assign n16172 = ~n1115 & n16171 ;
  assign n16173 = ~n12277 & n16172 ;
  assign n16169 = n12812 ^ n1652 ^ 1'b0 ;
  assign n16170 = ( n3283 & n8698 ) | ( n3283 & n16169 ) | ( n8698 & n16169 ) ;
  assign n16167 = ( ~x140 & n6296 ) | ( ~x140 & n7113 ) | ( n6296 & n7113 ) ;
  assign n16168 = n16167 ^ n15838 ^ 1'b0 ;
  assign n16174 = n16173 ^ n16170 ^ n16168 ;
  assign n16175 = n6543 & n15974 ;
  assign n16176 = ( n2953 & n11660 ) | ( n2953 & n16175 ) | ( n11660 & n16175 ) ;
  assign n16179 = n12465 ^ n5140 ^ n4234 ;
  assign n16180 = n16179 ^ n15525 ^ n3784 ;
  assign n16177 = n3110 & ~n7157 ;
  assign n16178 = n13895 & n16177 ;
  assign n16181 = n16180 ^ n16178 ^ 1'b0 ;
  assign n16182 = n10077 & n16181 ;
  assign n16183 = ( n1899 & n10280 ) | ( n1899 & ~n10654 ) | ( n10280 & ~n10654 ) ;
  assign n16184 = ( ~n6363 & n13634 ) | ( ~n6363 & n16183 ) | ( n13634 & n16183 ) ;
  assign n16185 = ( n1764 & n9673 ) | ( n1764 & ~n16184 ) | ( n9673 & ~n16184 ) ;
  assign n16196 = ( ~n1740 & n4182 ) | ( ~n1740 & n11126 ) | ( n4182 & n11126 ) ;
  assign n16197 = ( n991 & n5989 ) | ( n991 & n16196 ) | ( n5989 & n16196 ) ;
  assign n16198 = ( n14321 & n14818 ) | ( n14321 & n16197 ) | ( n14818 & n16197 ) ;
  assign n16199 = n16198 ^ n9346 ^ n1164 ;
  assign n16186 = n1578 | n5281 ;
  assign n16187 = n14867 | n16186 ;
  assign n16188 = n9578 ^ n3761 ^ n3554 ;
  assign n16189 = ( n4702 & n16187 ) | ( n4702 & n16188 ) | ( n16187 & n16188 ) ;
  assign n16190 = n16189 ^ n7578 ^ n1311 ;
  assign n16191 = n10461 ^ n5682 ^ 1'b0 ;
  assign n16192 = n10697 & ~n16191 ;
  assign n16193 = n7037 & n16192 ;
  assign n16194 = n16193 ^ n6578 ^ 1'b0 ;
  assign n16195 = n16190 & ~n16194 ;
  assign n16200 = n16199 ^ n16195 ^ 1'b0 ;
  assign n16204 = n1696 & ~n2210 ;
  assign n16202 = n15925 ^ n7735 ^ n3848 ;
  assign n16201 = n10921 ^ n7888 ^ n2216 ;
  assign n16203 = n16202 ^ n16201 ^ 1'b0 ;
  assign n16205 = n16204 ^ n16203 ^ n11973 ;
  assign n16206 = n7001 ^ n6913 ^ n530 ;
  assign n16208 = ( x121 & ~n923 ) | ( x121 & n7822 ) | ( ~n923 & n7822 ) ;
  assign n16207 = n14218 ^ n13112 ^ n7810 ;
  assign n16209 = n16208 ^ n16207 ^ 1'b0 ;
  assign n16210 = n2716 & n16209 ;
  assign n16211 = n5407 ^ n5094 ^ 1'b0 ;
  assign n16212 = n14193 ^ n6472 ^ x201 ;
  assign n16213 = ( x246 & n6281 ) | ( x246 & n15007 ) | ( n6281 & n15007 ) ;
  assign n16214 = ( n16211 & ~n16212 ) | ( n16211 & n16213 ) | ( ~n16212 & n16213 ) ;
  assign n16215 = ( ~n4630 & n7414 ) | ( ~n4630 & n8636 ) | ( n7414 & n8636 ) ;
  assign n16216 = n16215 ^ n369 ^ 1'b0 ;
  assign n16217 = n16216 ^ n6994 ^ x3 ;
  assign n16218 = n16217 ^ n11933 ^ n10786 ;
  assign n16227 = n13507 ^ n13443 ^ x89 ;
  assign n16228 = n16227 ^ n1677 ^ n1319 ;
  assign n16224 = ~n6254 & n9447 ;
  assign n16225 = n7306 & n16224 ;
  assign n16221 = n15664 ^ n14730 ^ n1534 ;
  assign n16219 = ( n2990 & ~n7930 ) | ( n2990 & n13980 ) | ( ~n7930 & n13980 ) ;
  assign n16220 = n16219 ^ n11232 ^ n3572 ;
  assign n16222 = n16221 ^ n16220 ^ 1'b0 ;
  assign n16223 = n16222 ^ n13829 ^ x144 ;
  assign n16226 = n16225 ^ n16223 ^ n12375 ;
  assign n16229 = n16228 ^ n16226 ^ n13006 ;
  assign n16230 = n15233 ^ n8144 ^ n578 ;
  assign n16231 = n2854 & ~n16230 ;
  assign n16232 = n16231 ^ n4885 ^ 1'b0 ;
  assign n16234 = n7009 ^ n2237 ^ 1'b0 ;
  assign n16235 = ~n1149 & n16234 ;
  assign n16236 = n16235 ^ n2275 ^ n1874 ;
  assign n16237 = ( n3555 & n16079 ) | ( n3555 & ~n16236 ) | ( n16079 & ~n16236 ) ;
  assign n16233 = n6193 ^ n1785 ^ n799 ;
  assign n16238 = n16237 ^ n16233 ^ n6908 ;
  assign n16239 = n13631 ^ n7534 ^ n453 ;
  assign n16240 = ( n5570 & ~n9911 ) | ( n5570 & n16239 ) | ( ~n9911 & n16239 ) ;
  assign n16241 = ( n7873 & n8921 ) | ( n7873 & n15570 ) | ( n8921 & n15570 ) ;
  assign n16242 = n9242 ^ n4312 ^ 1'b0 ;
  assign n16243 = n16242 ^ n12122 ^ 1'b0 ;
  assign n16244 = n11078 ^ n10152 ^ n6539 ;
  assign n16245 = n16244 ^ n6914 ^ n5177 ;
  assign n16246 = ( n4361 & n16243 ) | ( n4361 & n16245 ) | ( n16243 & n16245 ) ;
  assign n16247 = n16246 ^ n15675 ^ n4665 ;
  assign n16250 = ( n2318 & ~n5390 ) | ( n2318 & n6493 ) | ( ~n5390 & n6493 ) ;
  assign n16251 = n12611 ^ n8376 ^ n997 ;
  assign n16252 = ( ~n7656 & n16250 ) | ( ~n7656 & n16251 ) | ( n16250 & n16251 ) ;
  assign n16249 = n5733 ^ n5552 ^ n916 ;
  assign n16248 = n13943 ^ n10266 ^ 1'b0 ;
  assign n16253 = n16252 ^ n16249 ^ n16248 ;
  assign n16254 = n13381 ^ n5040 ^ 1'b0 ;
  assign n16255 = ~n16253 & n16254 ;
  assign n16263 = n5177 & n6617 ;
  assign n16264 = ( ~n6805 & n8879 ) | ( ~n6805 & n16263 ) | ( n8879 & n16263 ) ;
  assign n16256 = ( n1645 & n4343 ) | ( n1645 & ~n11718 ) | ( n4343 & ~n11718 ) ;
  assign n16257 = n1819 ^ n1088 ^ n264 ;
  assign n16258 = ( x105 & ~n5171 ) | ( x105 & n8655 ) | ( ~n5171 & n8655 ) ;
  assign n16259 = ( n2128 & n3071 ) | ( n2128 & n6432 ) | ( n3071 & n6432 ) ;
  assign n16260 = n16259 ^ x241 ^ x12 ;
  assign n16261 = ( n16257 & ~n16258 ) | ( n16257 & n16260 ) | ( ~n16258 & n16260 ) ;
  assign n16262 = ( ~n16125 & n16256 ) | ( ~n16125 & n16261 ) | ( n16256 & n16261 ) ;
  assign n16265 = n16264 ^ n16262 ^ n15056 ;
  assign n16266 = n15548 ^ n12559 ^ n1117 ;
  assign n16267 = n15183 ^ n450 ^ 1'b0 ;
  assign n16274 = n1624 & n3960 ;
  assign n16275 = n16274 ^ n13566 ^ 1'b0 ;
  assign n16271 = n8166 ^ n1198 ^ n982 ;
  assign n16272 = n16271 ^ n15861 ^ n1213 ;
  assign n16268 = n2081 ^ n1974 ^ x103 ;
  assign n16269 = ( ~n1351 & n3149 ) | ( ~n1351 & n5022 ) | ( n3149 & n5022 ) ;
  assign n16270 = ( n11928 & n16268 ) | ( n11928 & ~n16269 ) | ( n16268 & ~n16269 ) ;
  assign n16273 = n16272 ^ n16270 ^ n7222 ;
  assign n16276 = n16275 ^ n16273 ^ n10141 ;
  assign n16277 = ~n4617 & n4702 ;
  assign n16278 = n8745 & n16277 ;
  assign n16279 = n11009 ^ n2521 ^ 1'b0 ;
  assign n16280 = ( x108 & n2412 ) | ( x108 & ~n7313 ) | ( n2412 & ~n7313 ) ;
  assign n16281 = n16280 ^ n2178 ^ 1'b0 ;
  assign n16293 = n5191 ^ n3840 ^ x91 ;
  assign n16287 = n3630 ^ n574 ^ 1'b0 ;
  assign n16288 = n1793 | n16287 ;
  assign n16289 = ( ~n5340 & n7506 ) | ( ~n5340 & n16288 ) | ( n7506 & n16288 ) ;
  assign n16290 = ( n4032 & ~n4439 ) | ( n4032 & n7609 ) | ( ~n4439 & n7609 ) ;
  assign n16291 = ( n5899 & ~n16289 ) | ( n5899 & n16290 ) | ( ~n16289 & n16290 ) ;
  assign n16286 = ( n2309 & n4852 ) | ( n2309 & ~n14135 ) | ( n4852 & ~n14135 ) ;
  assign n16282 = ( ~n3426 & n3759 ) | ( ~n3426 & n5242 ) | ( n3759 & n5242 ) ;
  assign n16283 = n16282 ^ n15004 ^ n2874 ;
  assign n16284 = ( n5646 & ~n11015 ) | ( n5646 & n16283 ) | ( ~n11015 & n16283 ) ;
  assign n16285 = ( ~n5319 & n13718 ) | ( ~n5319 & n16284 ) | ( n13718 & n16284 ) ;
  assign n16292 = n16291 ^ n16286 ^ n16285 ;
  assign n16294 = n16293 ^ n16292 ^ n8959 ;
  assign n16295 = ( ~n512 & n1800 ) | ( ~n512 & n5213 ) | ( n1800 & n5213 ) ;
  assign n16296 = ( n5479 & ~n6826 ) | ( n5479 & n16295 ) | ( ~n6826 & n16295 ) ;
  assign n16308 = ( ~n3347 & n4729 ) | ( ~n3347 & n9337 ) | ( n4729 & n9337 ) ;
  assign n16309 = n16308 ^ n13624 ^ n1993 ;
  assign n16304 = ( n2037 & ~n7216 ) | ( n2037 & n9609 ) | ( ~n7216 & n9609 ) ;
  assign n16302 = ( n2287 & n5869 ) | ( n2287 & ~n7295 ) | ( n5869 & ~n7295 ) ;
  assign n16301 = ( ~n3492 & n4720 ) | ( ~n3492 & n5468 ) | ( n4720 & n5468 ) ;
  assign n16298 = ( n7444 & ~n8064 ) | ( n7444 & n9565 ) | ( ~n8064 & n9565 ) ;
  assign n16299 = ( n4501 & ~n8146 ) | ( n4501 & n16298 ) | ( ~n8146 & n16298 ) ;
  assign n16300 = n6998 & ~n16299 ;
  assign n16303 = n16302 ^ n16301 ^ n16300 ;
  assign n16305 = n16304 ^ n16303 ^ 1'b0 ;
  assign n16297 = n13113 ^ n2693 ^ 1'b0 ;
  assign n16306 = n16305 ^ n16297 ^ n14544 ;
  assign n16307 = n8931 | n16306 ;
  assign n16310 = n16309 ^ n16307 ^ 1'b0 ;
  assign n16311 = ( n1461 & n6584 ) | ( n1461 & ~n15815 ) | ( n6584 & ~n15815 ) ;
  assign n16312 = n16311 ^ n8161 ^ n5021 ;
  assign n16313 = n1709 | n9555 ;
  assign n16314 = ( n10687 & n11573 ) | ( n10687 & ~n16313 ) | ( n11573 & ~n16313 ) ;
  assign n16315 = n10824 ^ n1169 ^ 1'b0 ;
  assign n16316 = ( n16312 & ~n16314 ) | ( n16312 & n16315 ) | ( ~n16314 & n16315 ) ;
  assign n16317 = ( ~n5806 & n16310 ) | ( ~n5806 & n16316 ) | ( n16310 & n16316 ) ;
  assign n16325 = ( n9089 & n10329 ) | ( n9089 & n16038 ) | ( n10329 & n16038 ) ;
  assign n16326 = n16325 ^ n15935 ^ n8593 ;
  assign n16327 = n16326 ^ n10395 ^ n7627 ;
  assign n16319 = n12744 ^ n10554 ^ n4191 ;
  assign n16320 = ( n2259 & n4068 ) | ( n2259 & n11710 ) | ( n4068 & n11710 ) ;
  assign n16321 = n14485 & n16320 ;
  assign n16322 = n3013 & ~n16321 ;
  assign n16323 = ( n3331 & n6844 ) | ( n3331 & ~n15356 ) | ( n6844 & ~n15356 ) ;
  assign n16324 = ( n16319 & n16322 ) | ( n16319 & ~n16323 ) | ( n16322 & ~n16323 ) ;
  assign n16318 = ( n1160 & n7913 ) | ( n1160 & n12175 ) | ( n7913 & n12175 ) ;
  assign n16328 = n16327 ^ n16324 ^ n16318 ;
  assign n16330 = ( n3513 & ~n7136 ) | ( n3513 & n11891 ) | ( ~n7136 & n11891 ) ;
  assign n16329 = ( n2085 & ~n11767 ) | ( n2085 & n12821 ) | ( ~n11767 & n12821 ) ;
  assign n16331 = n16330 ^ n16329 ^ 1'b0 ;
  assign n16332 = ( ~n1162 & n2418 ) | ( ~n1162 & n3078 ) | ( n2418 & n3078 ) ;
  assign n16333 = ( n1507 & n8105 ) | ( n1507 & n16332 ) | ( n8105 & n16332 ) ;
  assign n16334 = n10673 ^ n2823 ^ x95 ;
  assign n16335 = n10118 ^ n6296 ^ n2031 ;
  assign n16336 = ( n3012 & ~n9125 ) | ( n3012 & n16335 ) | ( ~n9125 & n16335 ) ;
  assign n16337 = n12873 ^ n4455 ^ n3115 ;
  assign n16338 = n16337 ^ n11731 ^ n8966 ;
  assign n16339 = ~n16336 & n16338 ;
  assign n16340 = n15505 & n16339 ;
  assign n16345 = ( ~n4151 & n4775 ) | ( ~n4151 & n9372 ) | ( n4775 & n9372 ) ;
  assign n16343 = n2399 | n7952 ;
  assign n16344 = n16343 ^ n3856 ^ 1'b0 ;
  assign n16341 = n4860 ^ n3904 ^ n3090 ;
  assign n16342 = n5608 & n16341 ;
  assign n16346 = n16345 ^ n16344 ^ n16342 ;
  assign n16347 = ( n6327 & n13395 ) | ( n6327 & ~n16346 ) | ( n13395 & ~n16346 ) ;
  assign n16348 = n16340 | n16347 ;
  assign n16349 = n16334 & ~n16348 ;
  assign n16363 = n6096 & ~n11483 ;
  assign n16364 = n16363 ^ n3400 ^ 1'b0 ;
  assign n16355 = n10914 ^ n3669 ^ n2540 ;
  assign n16356 = n16355 ^ n14145 ^ n8144 ;
  assign n16357 = n3679 & ~n15468 ;
  assign n16358 = ~n6428 & n16357 ;
  assign n16359 = ( ~n4180 & n15212 ) | ( ~n4180 & n16358 ) | ( n15212 & n16358 ) ;
  assign n16360 = ( n5365 & ~n15653 ) | ( n5365 & n16359 ) | ( ~n15653 & n16359 ) ;
  assign n16361 = n3630 | n16360 ;
  assign n16362 = n16356 & ~n16361 ;
  assign n16365 = n16364 ^ n16362 ^ n12604 ;
  assign n16350 = n8294 ^ n4714 ^ 1'b0 ;
  assign n16351 = n14256 ^ n5722 ^ n3976 ;
  assign n16352 = n16351 ^ n5577 ^ 1'b0 ;
  assign n16353 = ~n16350 & n16352 ;
  assign n16354 = n16353 ^ n14417 ^ n11376 ;
  assign n16366 = n16365 ^ n16354 ^ n8718 ;
  assign n16367 = n7028 ^ n4115 ^ 1'b0 ;
  assign n16368 = n1448 & ~n16367 ;
  assign n16369 = n11891 ^ n8605 ^ n1051 ;
  assign n16370 = n16369 ^ n13602 ^ n10621 ;
  assign n16371 = ( ~n477 & n8348 ) | ( ~n477 & n16370 ) | ( n8348 & n16370 ) ;
  assign n16372 = n16371 ^ n13537 ^ n3465 ;
  assign n16373 = ( n3628 & n16368 ) | ( n3628 & n16372 ) | ( n16368 & n16372 ) ;
  assign n16374 = n4467 ^ n945 ^ 1'b0 ;
  assign n16375 = ( n2938 & n11162 ) | ( n2938 & ~n16374 ) | ( n11162 & ~n16374 ) ;
  assign n16376 = n16375 ^ n6808 ^ n2921 ;
  assign n16377 = n16376 ^ n9169 ^ 1'b0 ;
  assign n16378 = n6854 & n16377 ;
  assign n16382 = ( n5082 & n9311 ) | ( n5082 & n15501 ) | ( n9311 & n15501 ) ;
  assign n16379 = ( n981 & ~n2091 ) | ( n981 & n11095 ) | ( ~n2091 & n11095 ) ;
  assign n16380 = n16379 ^ n8833 ^ n1691 ;
  assign n16381 = n16380 ^ n10171 ^ n6891 ;
  assign n16383 = n16382 ^ n16381 ^ n10753 ;
  assign n16384 = n16383 ^ n16160 ^ n2497 ;
  assign n16385 = n13245 ^ n1536 ^ n1148 ;
  assign n16386 = ( n331 & ~n5629 ) | ( n331 & n6473 ) | ( ~n5629 & n6473 ) ;
  assign n16387 = n16386 ^ n5470 ^ n4429 ;
  assign n16388 = n10922 ^ n9098 ^ n7290 ;
  assign n16389 = ( n5725 & n5923 ) | ( n5725 & ~n15376 ) | ( n5923 & ~n15376 ) ;
  assign n16390 = ( n371 & ~n16388 ) | ( n371 & n16389 ) | ( ~n16388 & n16389 ) ;
  assign n16391 = ~n489 & n11335 ;
  assign n16392 = n16391 ^ n3413 ^ 1'b0 ;
  assign n16393 = ( n2478 & n12125 ) | ( n2478 & n16392 ) | ( n12125 & n16392 ) ;
  assign n16394 = ( ~n3079 & n8569 ) | ( ~n3079 & n16393 ) | ( n8569 & n16393 ) ;
  assign n16395 = n563 | n10519 ;
  assign n16396 = n5394 | n16395 ;
  assign n16397 = n12863 ^ n3205 ^ n1988 ;
  assign n16398 = ( n6379 & ~n6977 ) | ( n6379 & n16397 ) | ( ~n6977 & n16397 ) ;
  assign n16399 = ( n4478 & n15275 ) | ( n4478 & ~n16398 ) | ( n15275 & ~n16398 ) ;
  assign n16400 = n6089 ^ n3423 ^ n1936 ;
  assign n16401 = n7102 & ~n16400 ;
  assign n16402 = n16401 ^ n3138 ^ 1'b0 ;
  assign n16403 = n3910 ^ n1105 ^ 1'b0 ;
  assign n16404 = n14668 & n16403 ;
  assign n16405 = n16404 ^ n7543 ^ n5675 ;
  assign n16406 = n6550 ^ x229 ^ 1'b0 ;
  assign n16407 = n7341 | n16406 ;
  assign n16411 = n13285 ^ n11854 ^ n6312 ;
  assign n16412 = ( n806 & n4275 ) | ( n806 & n16068 ) | ( n4275 & n16068 ) ;
  assign n16413 = ( n1998 & ~n5086 ) | ( n1998 & n16412 ) | ( ~n5086 & n16412 ) ;
  assign n16414 = ( ~n13855 & n16411 ) | ( ~n13855 & n16413 ) | ( n16411 & n16413 ) ;
  assign n16408 = n8494 ^ n1688 ^ x242 ;
  assign n16409 = n6423 | n16408 ;
  assign n16410 = n16409 ^ n1806 ^ 1'b0 ;
  assign n16415 = n16414 ^ n16410 ^ 1'b0 ;
  assign n16416 = ( ~n2245 & n6970 ) | ( ~n2245 & n16415 ) | ( n6970 & n16415 ) ;
  assign n16417 = n16416 ^ n7276 ^ n5044 ;
  assign n16419 = n8747 ^ n5944 ^ n5894 ;
  assign n16418 = ( n2587 & n5437 ) | ( n2587 & n10478 ) | ( n5437 & n10478 ) ;
  assign n16420 = n16419 ^ n16418 ^ n8669 ;
  assign n16421 = n12313 & ~n16420 ;
  assign n16422 = n14719 & n16421 ;
  assign n16423 = ( n5451 & ~n10326 ) | ( n5451 & n12834 ) | ( ~n10326 & n12834 ) ;
  assign n16424 = n16423 ^ n2749 ^ 1'b0 ;
  assign n16425 = n13483 | n16424 ;
  assign n16426 = ( n11215 & n16197 ) | ( n11215 & n16425 ) | ( n16197 & n16425 ) ;
  assign n16427 = n8533 ^ n4465 ^ n4063 ;
  assign n16428 = n8331 ^ n6276 ^ n5987 ;
  assign n16429 = n16428 ^ n15240 ^ n1311 ;
  assign n16430 = n16429 ^ n3652 ^ 1'b0 ;
  assign n16431 = n16430 ^ n8766 ^ n1566 ;
  assign n16432 = n15097 ^ n6247 ^ n4877 ;
  assign n16435 = ( ~x192 & n2389 ) | ( ~x192 & n6690 ) | ( n2389 & n6690 ) ;
  assign n16436 = n16435 ^ n4704 ^ n3999 ;
  assign n16433 = ~n445 & n2653 ;
  assign n16434 = ~n11497 & n16433 ;
  assign n16437 = n16436 ^ n16434 ^ n8267 ;
  assign n16438 = n10519 ^ n5495 ^ n339 ;
  assign n16439 = ( n8134 & n14732 ) | ( n8134 & ~n16438 ) | ( n14732 & ~n16438 ) ;
  assign n16440 = ( n1781 & ~n6297 ) | ( n1781 & n15775 ) | ( ~n6297 & n15775 ) ;
  assign n16441 = n7841 ^ n5884 ^ n3748 ;
  assign n16442 = ( ~n14491 & n16440 ) | ( ~n14491 & n16441 ) | ( n16440 & n16441 ) ;
  assign n16443 = n16442 ^ n12481 ^ 1'b0 ;
  assign n16444 = n16443 ^ n1705 ^ x82 ;
  assign n16451 = n14466 ^ n13724 ^ n4647 ;
  assign n16452 = ( n5911 & n9420 ) | ( n5911 & ~n16451 ) | ( n9420 & ~n16451 ) ;
  assign n16447 = ( n11103 & n14864 ) | ( n11103 & ~n15840 ) | ( n14864 & ~n15840 ) ;
  assign n16448 = ( ~n3930 & n8826 ) | ( ~n3930 & n16447 ) | ( n8826 & n16447 ) ;
  assign n16449 = ( ~n4617 & n12757 ) | ( ~n4617 & n16448 ) | ( n12757 & n16448 ) ;
  assign n16445 = ( n2910 & n3260 ) | ( n2910 & ~n3308 ) | ( n3260 & ~n3308 ) ;
  assign n16446 = ( ~n2243 & n8074 ) | ( ~n2243 & n16445 ) | ( n8074 & n16445 ) ;
  assign n16450 = n16449 ^ n16446 ^ n14346 ;
  assign n16453 = n16452 ^ n16450 ^ n11321 ;
  assign n16454 = n8534 ^ n831 ^ 1'b0 ;
  assign n16455 = n16454 ^ n16312 ^ n10293 ;
  assign n16456 = n16455 ^ n6976 ^ 1'b0 ;
  assign n16457 = ( n3207 & n4631 ) | ( n3207 & ~n9316 ) | ( n4631 & ~n9316 ) ;
  assign n16458 = n16457 ^ n7553 ^ n1161 ;
  assign n16460 = n8964 ^ n7717 ^ n5053 ;
  assign n16461 = ( ~n7784 & n8586 ) | ( ~n7784 & n12321 ) | ( n8586 & n12321 ) ;
  assign n16462 = ( n11783 & n13376 ) | ( n11783 & ~n16461 ) | ( n13376 & ~n16461 ) ;
  assign n16463 = ( ~n5851 & n16460 ) | ( ~n5851 & n16462 ) | ( n16460 & n16462 ) ;
  assign n16459 = n13503 ^ n11916 ^ n1266 ;
  assign n16464 = n16463 ^ n16459 ^ 1'b0 ;
  assign n16465 = n6414 & ~n16464 ;
  assign n16472 = x248 & ~n12031 ;
  assign n16473 = n16472 ^ n14122 ^ 1'b0 ;
  assign n16470 = n10538 ^ n4930 ^ 1'b0 ;
  assign n16466 = ( n3288 & ~n8670 ) | ( n3288 & n12295 ) | ( ~n8670 & n12295 ) ;
  assign n16467 = n11617 ^ n6857 ^ n3439 ;
  assign n16468 = ( ~n1063 & n8347 ) | ( ~n1063 & n16467 ) | ( n8347 & n16467 ) ;
  assign n16469 = ( n16376 & n16466 ) | ( n16376 & n16468 ) | ( n16466 & n16468 ) ;
  assign n16471 = n16470 ^ n16469 ^ n1521 ;
  assign n16474 = n16473 ^ n16471 ^ n301 ;
  assign n16475 = n12283 ^ n3431 ^ n3355 ;
  assign n16476 = n6379 ^ n4350 ^ 1'b0 ;
  assign n16477 = n6846 | n16476 ;
  assign n16478 = ( ~n2483 & n10308 ) | ( ~n2483 & n16477 ) | ( n10308 & n16477 ) ;
  assign n16484 = n12457 ^ n7816 ^ x76 ;
  assign n16479 = x106 & n6161 ;
  assign n16480 = n16479 ^ n6906 ^ 1'b0 ;
  assign n16481 = n16480 ^ n8125 ^ n5748 ;
  assign n16482 = n16481 ^ n13376 ^ 1'b0 ;
  assign n16483 = n7118 & ~n16482 ;
  assign n16485 = n16484 ^ n16483 ^ n15553 ;
  assign n16486 = ( ~n16475 & n16478 ) | ( ~n16475 & n16485 ) | ( n16478 & n16485 ) ;
  assign n16487 = n2190 & n15185 ;
  assign n16496 = ( n1018 & n7409 ) | ( n1018 & n14589 ) | ( n7409 & n14589 ) ;
  assign n16499 = ~x113 & n574 ;
  assign n16497 = n14298 ^ n13330 ^ n3139 ;
  assign n16498 = n14049 | n16497 ;
  assign n16500 = n16499 ^ n16498 ^ 1'b0 ;
  assign n16501 = ( n1656 & n16496 ) | ( n1656 & n16500 ) | ( n16496 & n16500 ) ;
  assign n16490 = n2702 & n5795 ;
  assign n16491 = ~n2473 & n16490 ;
  assign n16489 = n16114 ^ n8153 ^ n4812 ;
  assign n16488 = ( n2110 & ~n6316 ) | ( n2110 & n13844 ) | ( ~n6316 & n13844 ) ;
  assign n16492 = n16491 ^ n16489 ^ n16488 ;
  assign n16493 = n16492 ^ n10997 ^ 1'b0 ;
  assign n16494 = n4854 & ~n16493 ;
  assign n16495 = ( n5161 & n15390 ) | ( n5161 & n16494 ) | ( n15390 & n16494 ) ;
  assign n16502 = n16501 ^ n16495 ^ n12641 ;
  assign n16503 = n292 & n5808 ;
  assign n16504 = n16503 ^ n1174 ^ 1'b0 ;
  assign n16505 = ( n2544 & n6867 ) | ( n2544 & ~n16504 ) | ( n6867 & ~n16504 ) ;
  assign n16506 = n14274 | n16499 ;
  assign n16507 = n16506 ^ n10712 ^ 1'b0 ;
  assign n16508 = ( n3449 & ~n12783 ) | ( n3449 & n16507 ) | ( ~n12783 & n16507 ) ;
  assign n16509 = ( n282 & n16505 ) | ( n282 & n16508 ) | ( n16505 & n16508 ) ;
  assign n16519 = n6334 | n6643 ;
  assign n16520 = n16519 ^ n12588 ^ 1'b0 ;
  assign n16510 = n9628 ^ n8690 ^ 1'b0 ;
  assign n16511 = n16510 ^ n7780 ^ 1'b0 ;
  assign n16512 = ( n2171 & n5782 ) | ( n2171 & ~n8225 ) | ( n5782 & ~n8225 ) ;
  assign n16513 = n1605 & ~n12583 ;
  assign n16514 = n16513 ^ n2865 ^ 1'b0 ;
  assign n16515 = n2692 | n16514 ;
  assign n16516 = n16512 & n16515 ;
  assign n16517 = n16516 ^ n4424 ^ n3731 ;
  assign n16518 = ( n14191 & n16511 ) | ( n14191 & ~n16517 ) | ( n16511 & ~n16517 ) ;
  assign n16521 = n16520 ^ n16518 ^ n9900 ;
  assign n16526 = n7040 ^ n4708 ^ n1113 ;
  assign n16524 = n14357 ^ n10304 ^ n8065 ;
  assign n16522 = n14527 ^ n6147 ^ 1'b0 ;
  assign n16523 = n16522 ^ n2256 ^ 1'b0 ;
  assign n16525 = n16524 ^ n16523 ^ n10175 ;
  assign n16527 = n16526 ^ n16525 ^ n6037 ;
  assign n16531 = x201 & n14349 ;
  assign n16528 = n7925 ^ n5576 ^ n1937 ;
  assign n16529 = n16528 ^ n3451 ^ n479 ;
  assign n16530 = n9166 & ~n16529 ;
  assign n16532 = n16531 ^ n16530 ^ n6660 ;
  assign n16535 = n15154 ^ n2594 ^ n881 ;
  assign n16536 = n16535 ^ n12146 ^ 1'b0 ;
  assign n16533 = n15566 ^ n7510 ^ n1196 ;
  assign n16534 = ( n6898 & n9078 ) | ( n6898 & n16533 ) | ( n9078 & n16533 ) ;
  assign n16537 = n16536 ^ n16534 ^ n4515 ;
  assign n16538 = n6347 ^ n3383 ^ n1325 ;
  assign n16539 = ( ~n10978 & n13077 ) | ( ~n10978 & n16538 ) | ( n13077 & n16538 ) ;
  assign n16540 = n10179 ^ n9870 ^ n2649 ;
  assign n16541 = n7112 & n8134 ;
  assign n16542 = n8222 & n16541 ;
  assign n16543 = n3650 ^ n3451 ^ n315 ;
  assign n16544 = ( n1680 & ~n8473 ) | ( n1680 & n16543 ) | ( ~n8473 & n16543 ) ;
  assign n16545 = ( n1535 & n16542 ) | ( n1535 & ~n16544 ) | ( n16542 & ~n16544 ) ;
  assign n16546 = n16545 ^ n6323 ^ 1'b0 ;
  assign n16547 = n5824 & ~n16546 ;
  assign n16548 = n3188 & n16547 ;
  assign n16549 = n16548 ^ n7860 ^ n4314 ;
  assign n16550 = n2898 & ~n16549 ;
  assign n16551 = ~n10262 & n16550 ;
  assign n16552 = ( n6541 & n7073 ) | ( n6541 & n9277 ) | ( n7073 & n9277 ) ;
  assign n16553 = n11223 | n15760 ;
  assign n16556 = ( ~n5417 & n7576 ) | ( ~n5417 & n11803 ) | ( n7576 & n11803 ) ;
  assign n16554 = ( n5785 & n7513 ) | ( n5785 & ~n9864 ) | ( n7513 & ~n9864 ) ;
  assign n16555 = n16554 ^ n3164 ^ 1'b0 ;
  assign n16557 = n16556 ^ n16555 ^ n5558 ;
  assign n16558 = n14379 ^ n11021 ^ n8822 ;
  assign n16559 = n16558 ^ n16471 ^ n15268 ;
  assign n16565 = ( n2097 & n2679 ) | ( n2097 & ~n8412 ) | ( n2679 & ~n8412 ) ;
  assign n16560 = n2253 ^ x97 ^ 1'b0 ;
  assign n16561 = n1571 & n16560 ;
  assign n16562 = ( n2333 & n5530 ) | ( n2333 & ~n16561 ) | ( n5530 & ~n16561 ) ;
  assign n16563 = ( x249 & n6595 ) | ( x249 & ~n16562 ) | ( n6595 & ~n16562 ) ;
  assign n16564 = ( n8001 & ~n9952 ) | ( n8001 & n16563 ) | ( ~n9952 & n16563 ) ;
  assign n16566 = n16565 ^ n16564 ^ 1'b0 ;
  assign n16567 = n13814 ^ n11262 ^ n3805 ;
  assign n16570 = n4715 ^ n1705 ^ 1'b0 ;
  assign n16571 = ( n1282 & n11781 ) | ( n1282 & ~n16570 ) | ( n11781 & ~n16570 ) ;
  assign n16568 = ( n1319 & n2019 ) | ( n1319 & ~n14724 ) | ( n2019 & ~n14724 ) ;
  assign n16569 = n16568 ^ n13043 ^ n4497 ;
  assign n16572 = n16571 ^ n16569 ^ n664 ;
  assign n16573 = ( n8640 & ~n16567 ) | ( n8640 & n16572 ) | ( ~n16567 & n16572 ) ;
  assign n16574 = ( n750 & n2085 ) | ( n750 & n3025 ) | ( n2085 & n3025 ) ;
  assign n16575 = ( n9852 & ~n12485 ) | ( n9852 & n16574 ) | ( ~n12485 & n16574 ) ;
  assign n16576 = n13318 ^ n11698 ^ n7055 ;
  assign n16577 = n2836 | n14939 ;
  assign n16578 = n16577 ^ n9378 ^ n2572 ;
  assign n16579 = n16578 ^ n3309 ^ 1'b0 ;
  assign n16580 = n8464 & n16579 ;
  assign n16581 = ( n1071 & n16576 ) | ( n1071 & n16580 ) | ( n16576 & n16580 ) ;
  assign n16582 = n3825 & n7857 ;
  assign n16583 = ~n7982 & n16582 ;
  assign n16584 = ( n6760 & n11695 ) | ( n6760 & n16583 ) | ( n11695 & n16583 ) ;
  assign n16585 = ( ~n10815 & n13025 ) | ( ~n10815 & n16584 ) | ( n13025 & n16584 ) ;
  assign n16586 = n2131 & ~n4750 ;
  assign n16587 = n16585 & n16586 ;
  assign n16588 = ( n16350 & n16581 ) | ( n16350 & n16587 ) | ( n16581 & n16587 ) ;
  assign n16589 = ( n2349 & n5932 ) | ( n2349 & n14598 ) | ( n5932 & n14598 ) ;
  assign n16590 = ( ~x57 & n6115 ) | ( ~x57 & n16589 ) | ( n6115 & n16589 ) ;
  assign n16592 = n7321 ^ n922 ^ n818 ;
  assign n16593 = ~n9786 & n16592 ;
  assign n16591 = n12541 ^ n1293 ^ 1'b0 ;
  assign n16594 = n16593 ^ n16591 ^ n3854 ;
  assign n16595 = n1644 ^ n1153 ^ n985 ;
  assign n16596 = ( ~n12407 & n12555 ) | ( ~n12407 & n16595 ) | ( n12555 & n16595 ) ;
  assign n16597 = ( n5905 & n6144 ) | ( n5905 & n15429 ) | ( n6144 & n15429 ) ;
  assign n16598 = n9704 ^ n3830 ^ n1633 ;
  assign n16599 = ( n2631 & ~n4005 ) | ( n2631 & n16598 ) | ( ~n4005 & n16598 ) ;
  assign n16600 = ( n7568 & ~n15053 ) | ( n7568 & n16599 ) | ( ~n15053 & n16599 ) ;
  assign n16601 = n4189 | n9128 ;
  assign n16602 = n16601 ^ n14049 ^ 1'b0 ;
  assign n16603 = n16602 ^ n5618 ^ 1'b0 ;
  assign n16604 = ~n11358 & n16603 ;
  assign n16605 = ~n4791 & n9448 ;
  assign n16606 = ~n16604 & n16605 ;
  assign n16610 = ( ~n1213 & n2550 ) | ( ~n1213 & n2584 ) | ( n2550 & n2584 ) ;
  assign n16607 = n16466 ^ n9296 ^ n5234 ;
  assign n16608 = n7746 ^ n6165 ^ x95 ;
  assign n16609 = ( n1541 & ~n16607 ) | ( n1541 & n16608 ) | ( ~n16607 & n16608 ) ;
  assign n16611 = n16610 ^ n16609 ^ n15403 ;
  assign n16612 = n16611 ^ n7993 ^ n3834 ;
  assign n16613 = ( n3792 & ~n16606 ) | ( n3792 & n16612 ) | ( ~n16606 & n16612 ) ;
  assign n16614 = n8345 ^ n901 ^ n256 ;
  assign n16615 = n286 & ~n2487 ;
  assign n16616 = n4109 & n16615 ;
  assign n16617 = n16616 ^ n4521 ^ n3989 ;
  assign n16618 = n16617 ^ n14682 ^ n4710 ;
  assign n16619 = n7715 ^ n6549 ^ n2144 ;
  assign n16620 = n2895 & n16619 ;
  assign n16621 = n16620 ^ n8629 ^ 1'b0 ;
  assign n16622 = n16621 ^ n15543 ^ n12869 ;
  assign n16623 = ( n2912 & n9940 ) | ( n2912 & ~n12667 ) | ( n9940 & ~n12667 ) ;
  assign n16624 = ( n2041 & n6728 ) | ( n2041 & ~n8944 ) | ( n6728 & ~n8944 ) ;
  assign n16625 = ( ~n10567 & n16623 ) | ( ~n10567 & n16624 ) | ( n16623 & n16624 ) ;
  assign n16626 = ( n12156 & n12418 ) | ( n12156 & n16625 ) | ( n12418 & n16625 ) ;
  assign n16627 = n16626 ^ n10495 ^ 1'b0 ;
  assign n16628 = n16622 | n16627 ;
  assign n16629 = n16628 ^ n15233 ^ n883 ;
  assign n16630 = ( n16614 & n16618 ) | ( n16614 & ~n16629 ) | ( n16618 & ~n16629 ) ;
  assign n16631 = n5675 ^ n3451 ^ n590 ;
  assign n16632 = ( n4704 & n6458 ) | ( n4704 & n16631 ) | ( n6458 & n16631 ) ;
  assign n16633 = ( n3200 & ~n3835 ) | ( n3200 & n16632 ) | ( ~n3835 & n16632 ) ;
  assign n16634 = n15224 ^ n2369 ^ n1561 ;
  assign n16635 = n5235 ^ n2309 ^ n993 ;
  assign n16636 = ( n2986 & n10934 ) | ( n2986 & n16635 ) | ( n10934 & n16635 ) ;
  assign n16637 = n16636 ^ n10727 ^ n7921 ;
  assign n16638 = ~n5396 & n13995 ;
  assign n16639 = n16638 ^ n5178 ^ n5116 ;
  assign n16640 = ( n4824 & n5374 ) | ( n4824 & ~n14997 ) | ( n5374 & ~n14997 ) ;
  assign n16641 = n16640 ^ n16460 ^ n9486 ;
  assign n16642 = n16641 ^ n14749 ^ n11524 ;
  assign n16643 = n2470 ^ n1109 ^ 1'b0 ;
  assign n16644 = ( n1139 & n10230 ) | ( n1139 & n16643 ) | ( n10230 & n16643 ) ;
  assign n16645 = n16644 ^ n10239 ^ 1'b0 ;
  assign n16646 = n14352 | n16645 ;
  assign n16647 = n11363 ^ n7832 ^ n4264 ;
  assign n16648 = n16647 ^ n2268 ^ 1'b0 ;
  assign n16649 = n16648 ^ n10447 ^ n3390 ;
  assign n16659 = ( n2195 & n5302 ) | ( n2195 & n8592 ) | ( n5302 & n8592 ) ;
  assign n16652 = n6021 ^ n2484 ^ n930 ;
  assign n16653 = n2211 ^ n1732 ^ n1709 ;
  assign n16654 = n16653 ^ n4338 ^ n1359 ;
  assign n16655 = n12102 ^ n524 ^ 1'b0 ;
  assign n16656 = n16654 & ~n16655 ;
  assign n16657 = n16656 ^ n9972 ^ 1'b0 ;
  assign n16658 = n16652 & ~n16657 ;
  assign n16660 = n16659 ^ n16658 ^ n2960 ;
  assign n16661 = n11912 & ~n16660 ;
  assign n16662 = n16661 ^ n7968 ^ 1'b0 ;
  assign n16650 = n7643 ^ n4401 ^ n652 ;
  assign n16651 = n16650 ^ n9963 ^ n5751 ;
  assign n16663 = n16662 ^ n16651 ^ n11795 ;
  assign n16664 = ( n371 & n13923 ) | ( n371 & n16059 ) | ( n13923 & n16059 ) ;
  assign n16665 = x10 & ~n13519 ;
  assign n16666 = n16665 ^ n9498 ^ 1'b0 ;
  assign n16667 = n3863 ^ n3499 ^ n1396 ;
  assign n16668 = ( n1203 & ~n4131 ) | ( n1203 & n9407 ) | ( ~n4131 & n9407 ) ;
  assign n16669 = ( ~n7739 & n8399 ) | ( ~n7739 & n16668 ) | ( n8399 & n16668 ) ;
  assign n16670 = n6283 ^ n2576 ^ n1195 ;
  assign n16671 = ( n5160 & n8665 ) | ( n5160 & n16670 ) | ( n8665 & n16670 ) ;
  assign n16672 = n11451 ^ n7223 ^ 1'b0 ;
  assign n16673 = n13652 ^ n4132 ^ 1'b0 ;
  assign n16674 = ~n16672 & n16673 ;
  assign n16675 = n11827 ^ n7473 ^ n6918 ;
  assign n16676 = n16675 ^ n9501 ^ 1'b0 ;
  assign n16677 = n16676 ^ n5347 ^ 1'b0 ;
  assign n16678 = n12463 ^ n7919 ^ n6947 ;
  assign n16679 = n5689 | n15222 ;
  assign n16680 = n16679 ^ n589 ^ 1'b0 ;
  assign n16681 = ( n4091 & n8768 ) | ( n4091 & ~n16680 ) | ( n8768 & ~n16680 ) ;
  assign n16682 = n6080 & ~n16681 ;
  assign n16683 = ~n16678 & n16682 ;
  assign n16685 = n5688 ^ n4611 ^ n3027 ;
  assign n16686 = n16685 ^ n6691 ^ n6631 ;
  assign n16684 = ~n446 & n8939 ;
  assign n16687 = n16686 ^ n16684 ^ 1'b0 ;
  assign n16688 = ( n3760 & n15958 ) | ( n3760 & n16687 ) | ( n15958 & n16687 ) ;
  assign n16689 = ~n2186 & n8323 ;
  assign n16690 = n16689 ^ n16525 ^ n8087 ;
  assign n16691 = n16690 ^ n16222 ^ n3879 ;
  assign n16693 = ( ~n1851 & n5775 ) | ( ~n1851 & n8500 ) | ( n5775 & n8500 ) ;
  assign n16694 = n16693 ^ n4988 ^ n1348 ;
  assign n16692 = n8708 ^ n5696 ^ 1'b0 ;
  assign n16695 = n16694 ^ n16692 ^ n9397 ;
  assign n16696 = n14263 ^ n9846 ^ n5577 ;
  assign n16697 = n16696 ^ n12084 ^ n4168 ;
  assign n16698 = ( ~n5264 & n5276 ) | ( ~n5264 & n5489 ) | ( n5276 & n5489 ) ;
  assign n16700 = n6995 ^ n6538 ^ n4618 ;
  assign n16699 = ~n2871 & n6079 ;
  assign n16701 = n16700 ^ n16699 ^ 1'b0 ;
  assign n16702 = n10069 ^ n6421 ^ n2471 ;
  assign n16703 = ( n1949 & n16235 ) | ( n1949 & n16702 ) | ( n16235 & n16702 ) ;
  assign n16704 = ( ~n16698 & n16701 ) | ( ~n16698 & n16703 ) | ( n16701 & n16703 ) ;
  assign n16705 = n13595 ^ n8654 ^ n7613 ;
  assign n16706 = n16705 ^ n14544 ^ n6510 ;
  assign n16714 = ( ~n3691 & n6200 ) | ( ~n3691 & n16068 ) | ( n6200 & n16068 ) ;
  assign n16709 = ( n298 & n2390 ) | ( n298 & n7752 ) | ( n2390 & n7752 ) ;
  assign n16707 = ( n2192 & n3664 ) | ( n2192 & ~n4448 ) | ( n3664 & ~n4448 ) ;
  assign n16708 = ( n1036 & n4080 ) | ( n1036 & n16707 ) | ( n4080 & n16707 ) ;
  assign n16710 = n16709 ^ n16708 ^ n3625 ;
  assign n16711 = n11740 | n16710 ;
  assign n16712 = n16364 & ~n16711 ;
  assign n16713 = n3442 & ~n16712 ;
  assign n16715 = n16714 ^ n16713 ^ 1'b0 ;
  assign n16717 = n2981 & n8833 ;
  assign n16718 = ( ~n2879 & n4116 ) | ( ~n2879 & n16717 ) | ( n4116 & n16717 ) ;
  assign n16716 = ~n842 & n15220 ;
  assign n16719 = n16718 ^ n16716 ^ 1'b0 ;
  assign n16725 = n2074 | n6776 ;
  assign n16726 = n16725 ^ n4290 ^ 1'b0 ;
  assign n16720 = n4621 & n6328 ;
  assign n16721 = n16720 ^ n14530 ^ 1'b0 ;
  assign n16722 = n13487 ^ n12315 ^ n5764 ;
  assign n16723 = ( n9233 & ~n16721 ) | ( n9233 & n16722 ) | ( ~n16721 & n16722 ) ;
  assign n16724 = ( n1906 & n3389 ) | ( n1906 & n16723 ) | ( n3389 & n16723 ) ;
  assign n16727 = n16726 ^ n16724 ^ n11000 ;
  assign n16728 = n16727 ^ n7674 ^ n6527 ;
  assign n16729 = x242 & n303 ;
  assign n16730 = n16729 ^ n510 ^ 1'b0 ;
  assign n16731 = n16730 ^ n9971 ^ n9922 ;
  assign n16732 = n12120 ^ n5359 ^ n5280 ;
  assign n16733 = n16732 ^ n11393 ^ n1928 ;
  assign n16734 = n12979 ^ n7153 ^ 1'b0 ;
  assign n16735 = n16733 & ~n16734 ;
  assign n16737 = n6557 & ~n16692 ;
  assign n16736 = ( n1211 & n1352 ) | ( n1211 & ~n7646 ) | ( n1352 & ~n7646 ) ;
  assign n16738 = n16737 ^ n16736 ^ n9528 ;
  assign n16739 = ( x43 & n6780 ) | ( x43 & n16738 ) | ( n6780 & n16738 ) ;
  assign n16740 = ~n449 & n7303 ;
  assign n16741 = n16740 ^ n7206 ^ 1'b0 ;
  assign n16742 = ( n1514 & ~n16016 ) | ( n1514 & n16741 ) | ( ~n16016 & n16741 ) ;
  assign n16743 = n10263 ^ n3826 ^ n2099 ;
  assign n16744 = n16743 ^ n12657 ^ n4218 ;
  assign n16745 = n16744 ^ n16158 ^ n2432 ;
  assign n16751 = n7706 & ~n15444 ;
  assign n16746 = n7239 ^ n2548 ^ 1'b0 ;
  assign n16747 = n11786 & n16746 ;
  assign n16748 = ~n2351 & n16747 ;
  assign n16749 = n16748 ^ n15319 ^ n4721 ;
  assign n16750 = n10857 & n16749 ;
  assign n16752 = n16751 ^ n16750 ^ 1'b0 ;
  assign n16758 = ( x101 & n10442 ) | ( x101 & ~n15450 ) | ( n10442 & ~n15450 ) ;
  assign n16757 = n12161 ^ n7345 ^ n5007 ;
  assign n16753 = ( n1803 & n2282 ) | ( n1803 & ~n13599 ) | ( n2282 & ~n13599 ) ;
  assign n16754 = n16753 ^ n15177 ^ n11450 ;
  assign n16755 = ( x200 & n4265 ) | ( x200 & ~n16754 ) | ( n4265 & ~n16754 ) ;
  assign n16756 = ( n11068 & n15003 ) | ( n11068 & n16755 ) | ( n15003 & n16755 ) ;
  assign n16759 = n16758 ^ n16757 ^ n16756 ;
  assign n16775 = ( ~n3861 & n7565 ) | ( ~n3861 & n11922 ) | ( n7565 & n11922 ) ;
  assign n16760 = ~n1784 & n6330 ;
  assign n16761 = n16760 ^ n6510 ^ n5748 ;
  assign n16762 = ( x140 & n1696 ) | ( x140 & ~n12840 ) | ( n1696 & ~n12840 ) ;
  assign n16763 = n5321 ^ n1374 ^ n1312 ;
  assign n16764 = ~n699 & n5255 ;
  assign n16765 = ( n2993 & n3858 ) | ( n2993 & ~n16764 ) | ( n3858 & ~n16764 ) ;
  assign n16766 = n4615 | n7456 ;
  assign n16767 = ( n1349 & ~n2360 ) | ( n1349 & n14356 ) | ( ~n2360 & n14356 ) ;
  assign n16768 = ( ~n15848 & n16766 ) | ( ~n15848 & n16767 ) | ( n16766 & n16767 ) ;
  assign n16769 = ( ~n1656 & n16765 ) | ( ~n1656 & n16768 ) | ( n16765 & n16768 ) ;
  assign n16770 = n16769 ^ n7654 ^ n5125 ;
  assign n16771 = ( n6264 & ~n16763 ) | ( n6264 & n16770 ) | ( ~n16763 & n16770 ) ;
  assign n16772 = n16771 ^ n13614 ^ n721 ;
  assign n16773 = ( n10692 & n16762 ) | ( n10692 & ~n16772 ) | ( n16762 & ~n16772 ) ;
  assign n16774 = n16761 | n16773 ;
  assign n16776 = n16775 ^ n16774 ^ 1'b0 ;
  assign n16777 = n13805 ^ n9600 ^ n3345 ;
  assign n16778 = n16499 ^ n6921 ^ 1'b0 ;
  assign n16779 = n2136 ^ n614 ^ x4 ;
  assign n16780 = ( n2480 & n10933 ) | ( n2480 & ~n16779 ) | ( n10933 & ~n16779 ) ;
  assign n16781 = n1418 & ~n9537 ;
  assign n16782 = n12374 ^ n2487 ^ 1'b0 ;
  assign n16783 = n3547 & n16782 ;
  assign n16784 = ( n1794 & n3864 ) | ( n1794 & n16783 ) | ( n3864 & n16783 ) ;
  assign n16790 = n12729 ^ n8452 ^ n2935 ;
  assign n16791 = n16790 ^ n1722 ^ n601 ;
  assign n16785 = ( n657 & n748 ) | ( n657 & ~n3487 ) | ( n748 & ~n3487 ) ;
  assign n16786 = n16785 ^ n7640 ^ x84 ;
  assign n16787 = n16786 ^ n6038 ^ 1'b0 ;
  assign n16788 = n10848 & ~n16787 ;
  assign n16789 = ( n10035 & n12716 ) | ( n10035 & ~n16788 ) | ( n12716 & ~n16788 ) ;
  assign n16792 = n16791 ^ n16789 ^ n2174 ;
  assign n16793 = n16784 & ~n16792 ;
  assign n16794 = n12439 & n12665 ;
  assign n16795 = ~n16793 & n16794 ;
  assign n16797 = n2864 ^ n2818 ^ n1469 ;
  assign n16796 = ( n2738 & n5146 ) | ( n2738 & n9070 ) | ( n5146 & n9070 ) ;
  assign n16798 = n16797 ^ n16796 ^ n11005 ;
  assign n16802 = n9457 ^ n5401 ^ x214 ;
  assign n16803 = ( n2133 & ~n4984 ) | ( n2133 & n16802 ) | ( ~n4984 & n16802 ) ;
  assign n16799 = ( n3591 & n5370 ) | ( n3591 & ~n6462 ) | ( n5370 & ~n6462 ) ;
  assign n16800 = n16799 ^ n9254 ^ n1557 ;
  assign n16801 = ( ~n8817 & n16369 ) | ( ~n8817 & n16800 ) | ( n16369 & n16800 ) ;
  assign n16804 = n16803 ^ n16801 ^ n2486 ;
  assign n16806 = n9730 ^ n6716 ^ x34 ;
  assign n16805 = n14234 ^ n5229 ^ n2929 ;
  assign n16807 = n16806 ^ n16805 ^ n7965 ;
  assign n16808 = ( n973 & n9681 ) | ( n973 & n10099 ) | ( n9681 & n10099 ) ;
  assign n16809 = ( n4693 & n6094 ) | ( n4693 & ~n16808 ) | ( n6094 & ~n16808 ) ;
  assign n16810 = ( n312 & n3000 ) | ( n312 & ~n16802 ) | ( n3000 & ~n16802 ) ;
  assign n16811 = ( ~n2371 & n13850 ) | ( ~n2371 & n13957 ) | ( n13850 & n13957 ) ;
  assign n16812 = n16811 ^ n3306 ^ n974 ;
  assign n16813 = ( ~n965 & n16810 ) | ( ~n965 & n16812 ) | ( n16810 & n16812 ) ;
  assign n16814 = ( n766 & ~n4556 ) | ( n766 & n5681 ) | ( ~n4556 & n5681 ) ;
  assign n16815 = ( ~n1167 & n8853 ) | ( ~n1167 & n16814 ) | ( n8853 & n16814 ) ;
  assign n16816 = n16815 ^ n9287 ^ x57 ;
  assign n16817 = n12663 | n13635 ;
  assign n16818 = n16816 & ~n16817 ;
  assign n16819 = ( n711 & n721 ) | ( n711 & n8698 ) | ( n721 & n8698 ) ;
  assign n16826 = n14625 ^ n9606 ^ n5591 ;
  assign n16827 = n6366 ^ n3109 ^ n2777 ;
  assign n16828 = n16826 | n16827 ;
  assign n16829 = ( n4505 & n10338 ) | ( n4505 & ~n16828 ) | ( n10338 & ~n16828 ) ;
  assign n16820 = ( n491 & n2185 ) | ( n491 & ~n2711 ) | ( n2185 & ~n2711 ) ;
  assign n16821 = ( n3403 & n12042 ) | ( n3403 & ~n16820 ) | ( n12042 & ~n16820 ) ;
  assign n16822 = ( n1601 & n5426 ) | ( n1601 & n16821 ) | ( n5426 & n16821 ) ;
  assign n16823 = n16803 ^ n3634 ^ 1'b0 ;
  assign n16824 = n16822 & n16823 ;
  assign n16825 = n16824 ^ n13483 ^ n2571 ;
  assign n16830 = n16829 ^ n16825 ^ n3186 ;
  assign n16831 = ( n2175 & n16819 ) | ( n2175 & n16830 ) | ( n16819 & n16830 ) ;
  assign n16832 = n16236 ^ n5456 ^ n4563 ;
  assign n16833 = n16832 ^ n4600 ^ n2692 ;
  assign n16834 = n11076 ^ n7201 ^ n4400 ;
  assign n16835 = n16834 ^ n2038 ^ x200 ;
  assign n16836 = n13102 ^ n3593 ^ n1095 ;
  assign n16837 = ( ~n16332 & n16835 ) | ( ~n16332 & n16836 ) | ( n16835 & n16836 ) ;
  assign n16838 = n3815 & ~n4563 ;
  assign n16839 = n12781 ^ n10013 ^ 1'b0 ;
  assign n16840 = n8279 & n16839 ;
  assign n16841 = ( n1210 & ~n6301 ) | ( n1210 & n16840 ) | ( ~n6301 & n16840 ) ;
  assign n16842 = n10605 ^ n7185 ^ 1'b0 ;
  assign n16843 = n13043 ^ n8494 ^ n1335 ;
  assign n16844 = n16842 & n16843 ;
  assign n16845 = ~n16841 & n16844 ;
  assign n16846 = n16838 & ~n16845 ;
  assign n16847 = ( n7552 & n15330 ) | ( n7552 & ~n16846 ) | ( n15330 & ~n16846 ) ;
  assign n16848 = n16847 ^ n14403 ^ n12646 ;
  assign n16849 = ~n10717 & n14366 ;
  assign n16850 = n16849 ^ n16504 ^ n14957 ;
  assign n16851 = ( n2754 & n11124 ) | ( n2754 & ~n16850 ) | ( n11124 & ~n16850 ) ;
  assign n16852 = ( n10592 & ~n10689 ) | ( n10592 & n16851 ) | ( ~n10689 & n16851 ) ;
  assign n16854 = ( n5417 & n8737 ) | ( n5417 & ~n14365 ) | ( n8737 & ~n14365 ) ;
  assign n16855 = n16854 ^ n12528 ^ n5462 ;
  assign n16856 = n16855 ^ n9278 ^ 1'b0 ;
  assign n16857 = ~n15985 & n16856 ;
  assign n16853 = ~n14398 & n16346 ;
  assign n16858 = n16857 ^ n16853 ^ n11937 ;
  assign n16859 = n16858 ^ n15989 ^ n2127 ;
  assign n16860 = n1199 ^ n314 ^ 1'b0 ;
  assign n16861 = n11683 & n16860 ;
  assign n16862 = n16861 ^ n4337 ^ 1'b0 ;
  assign n16863 = n2386 & n4701 ;
  assign n16864 = n1339 & ~n15585 ;
  assign n16865 = ( n5519 & n8671 ) | ( n5519 & ~n16864 ) | ( n8671 & ~n16864 ) ;
  assign n16866 = ( n1288 & n1379 ) | ( n1288 & ~n1755 ) | ( n1379 & ~n1755 ) ;
  assign n16867 = ( n5268 & ~n9280 ) | ( n5268 & n16866 ) | ( ~n9280 & n16866 ) ;
  assign n16868 = ( n2749 & ~n8225 ) | ( n2749 & n16867 ) | ( ~n8225 & n16867 ) ;
  assign n16869 = n16868 ^ n8707 ^ 1'b0 ;
  assign n16870 = ( n16863 & ~n16865 ) | ( n16863 & n16869 ) | ( ~n16865 & n16869 ) ;
  assign n16871 = ( n3723 & n5619 ) | ( n3723 & n8640 ) | ( n5619 & n8640 ) ;
  assign n16872 = ~x216 & n1080 ;
  assign n16873 = n16872 ^ n15255 ^ n12714 ;
  assign n16875 = n8556 ^ n5860 ^ n5113 ;
  assign n16876 = ( ~n5090 & n10726 ) | ( ~n5090 & n16875 ) | ( n10726 & n16875 ) ;
  assign n16874 = ( x187 & ~n9334 ) | ( x187 & n16286 ) | ( ~n9334 & n16286 ) ;
  assign n16877 = n16876 ^ n16874 ^ 1'b0 ;
  assign n16878 = n16873 & n16877 ;
  assign n16879 = ~n4160 & n14882 ;
  assign n16880 = n8338 ^ n5322 ^ n2055 ;
  assign n16881 = n10488 ^ n3325 ^ 1'b0 ;
  assign n16882 = ( n9076 & n16880 ) | ( n9076 & n16881 ) | ( n16880 & n16881 ) ;
  assign n16883 = n10457 & ~n16882 ;
  assign n16884 = n13463 & n16883 ;
  assign n16885 = n8181 ^ n4041 ^ n3974 ;
  assign n16886 = n16885 ^ n11050 ^ n1905 ;
  assign n16887 = ( n16879 & ~n16884 ) | ( n16879 & n16886 ) | ( ~n16884 & n16886 ) ;
  assign n16888 = ( ~n5265 & n8993 ) | ( ~n5265 & n16887 ) | ( n8993 & n16887 ) ;
  assign n16889 = ( n2470 & n10307 ) | ( n2470 & ~n16888 ) | ( n10307 & ~n16888 ) ;
  assign n16890 = n1048 ^ n876 ^ 1'b0 ;
  assign n16891 = ( ~n13182 & n14424 ) | ( ~n13182 & n16890 ) | ( n14424 & n16890 ) ;
  assign n16895 = n5314 ^ n4048 ^ n364 ;
  assign n16892 = ( n734 & ~n1077 ) | ( n734 & n2485 ) | ( ~n1077 & n2485 ) ;
  assign n16893 = n16892 ^ n14016 ^ n13345 ;
  assign n16894 = n16893 ^ n8743 ^ n1563 ;
  assign n16896 = n16895 ^ n16894 ^ n13623 ;
  assign n16897 = n16896 ^ n15895 ^ n7844 ;
  assign n16898 = n13587 ^ n7836 ^ n5184 ;
  assign n16899 = n16898 ^ n10536 ^ n3681 ;
  assign n16900 = ( n957 & ~n3184 ) | ( n957 & n5883 ) | ( ~n3184 & n5883 ) ;
  assign n16901 = ( n2429 & ~n4518 ) | ( n2429 & n16900 ) | ( ~n4518 & n16900 ) ;
  assign n16902 = ( n6653 & ~n16899 ) | ( n6653 & n16901 ) | ( ~n16899 & n16901 ) ;
  assign n16903 = n11865 ^ n8365 ^ 1'b0 ;
  assign n16904 = ( ~n1473 & n7541 ) | ( ~n1473 & n12514 ) | ( n7541 & n12514 ) ;
  assign n16905 = n5990 & n6747 ;
  assign n16906 = n16905 ^ n2433 ^ 1'b0 ;
  assign n16907 = ( n1777 & n4429 ) | ( n1777 & n6545 ) | ( n4429 & n6545 ) ;
  assign n16908 = ( ~n2240 & n16906 ) | ( ~n2240 & n16907 ) | ( n16906 & n16907 ) ;
  assign n16909 = ( n1870 & ~n4725 ) | ( n1870 & n10809 ) | ( ~n4725 & n10809 ) ;
  assign n16910 = n16909 ^ n2432 ^ 1'b0 ;
  assign n16911 = ~n16908 & n16910 ;
  assign n16912 = ~n16904 & n16911 ;
  assign n16913 = n16912 ^ n11981 ^ 1'b0 ;
  assign n16914 = n11837 & n15700 ;
  assign n16915 = ~n16913 & n16914 ;
  assign n16916 = n8268 ^ n5799 ^ n5496 ;
  assign n16917 = ( ~n3168 & n5152 ) | ( ~n3168 & n5993 ) | ( n5152 & n5993 ) ;
  assign n16918 = ( n2840 & ~n5960 ) | ( n2840 & n16512 ) | ( ~n5960 & n16512 ) ;
  assign n16919 = ( ~n9534 & n16917 ) | ( ~n9534 & n16918 ) | ( n16917 & n16918 ) ;
  assign n16920 = ( n3319 & n16203 ) | ( n3319 & ~n16919 ) | ( n16203 & ~n16919 ) ;
  assign n16921 = n16916 & ~n16920 ;
  assign n16922 = n5601 ^ n5229 ^ 1'b0 ;
  assign n16923 = n8168 & ~n16922 ;
  assign n16927 = n378 | n2378 ;
  assign n16924 = x45 & n8568 ;
  assign n16925 = n16924 ^ n15574 ^ 1'b0 ;
  assign n16926 = ( n3922 & ~n8617 ) | ( n3922 & n16925 ) | ( ~n8617 & n16925 ) ;
  assign n16928 = n16927 ^ n16926 ^ n12654 ;
  assign n16929 = ( n1749 & n1762 ) | ( n1749 & ~n4517 ) | ( n1762 & ~n4517 ) ;
  assign n16930 = ( ~n2374 & n3015 ) | ( ~n2374 & n9282 ) | ( n3015 & n9282 ) ;
  assign n16931 = ( n4011 & n6299 ) | ( n4011 & ~n16930 ) | ( n6299 & ~n16930 ) ;
  assign n16932 = n9339 ^ n2429 ^ n1823 ;
  assign n16933 = n16932 ^ n6536 ^ n4373 ;
  assign n16934 = n5093 ^ n2945 ^ x188 ;
  assign n16935 = n11474 | n16934 ;
  assign n16936 = n5122 & n16935 ;
  assign n16937 = n16936 ^ n13833 ^ 1'b0 ;
  assign n16944 = n1547 | n10567 ;
  assign n16938 = n10192 ^ n1436 ^ x171 ;
  assign n16939 = ( n3461 & n3568 ) | ( n3461 & ~n10221 ) | ( n3568 & ~n10221 ) ;
  assign n16940 = n2937 & n16939 ;
  assign n16941 = n16940 ^ n15295 ^ n6784 ;
  assign n16942 = n16941 ^ n14287 ^ n4784 ;
  assign n16943 = ~n16938 & n16942 ;
  assign n16945 = n16944 ^ n16943 ^ 1'b0 ;
  assign n16946 = n16945 ^ n8841 ^ n2521 ;
  assign n16947 = n3539 ^ n2210 ^ n1260 ;
  assign n16948 = ~n792 & n16947 ;
  assign n16949 = ( ~n1947 & n8607 ) | ( ~n1947 & n16948 ) | ( n8607 & n16948 ) ;
  assign n16950 = ( n3645 & n4514 ) | ( n3645 & n6096 ) | ( n4514 & n6096 ) ;
  assign n16951 = n16950 ^ n5853 ^ n5779 ;
  assign n16952 = ( ~n2052 & n7690 ) | ( ~n2052 & n16951 ) | ( n7690 & n16951 ) ;
  assign n16953 = n4423 & n8901 ;
  assign n16954 = n7905 ^ n3219 ^ 1'b0 ;
  assign n16955 = ~n4599 & n5544 ;
  assign n16956 = n16954 & n16955 ;
  assign n16957 = n13443 ^ n9063 ^ n6124 ;
  assign n16958 = n16957 ^ n13684 ^ n12540 ;
  assign n16971 = ( x109 & n1810 ) | ( x109 & ~n16007 ) | ( n1810 & ~n16007 ) ;
  assign n16969 = n1777 ^ n1663 ^ n1156 ;
  assign n16968 = n3453 ^ n3082 ^ x23 ;
  assign n16970 = n16969 ^ n16968 ^ n6543 ;
  assign n16962 = ( n3165 & ~n5239 ) | ( n3165 & n15784 ) | ( ~n5239 & n15784 ) ;
  assign n16963 = n16962 ^ n4875 ^ n3790 ;
  assign n16964 = n5451 & n16963 ;
  assign n16965 = ~n6608 & n16964 ;
  assign n16966 = n16965 ^ n11407 ^ n7370 ;
  assign n16959 = n5650 ^ n1855 ^ n1142 ;
  assign n16960 = n16959 ^ n6610 ^ n513 ;
  assign n16961 = n16960 ^ n8502 ^ n4862 ;
  assign n16967 = n16966 ^ n16961 ^ n3181 ;
  assign n16972 = n16971 ^ n16970 ^ n16967 ;
  assign n16973 = ( n16956 & ~n16958 ) | ( n16956 & n16972 ) | ( ~n16958 & n16972 ) ;
  assign n16974 = n7906 & n12929 ;
  assign n16975 = n16974 ^ n10930 ^ n4374 ;
  assign n16976 = ( n8860 & n10182 ) | ( n8860 & n16975 ) | ( n10182 & n16975 ) ;
  assign n16977 = ~n4239 & n16055 ;
  assign n16978 = ( n7501 & ~n8158 ) | ( n7501 & n13709 ) | ( ~n8158 & n13709 ) ;
  assign n16979 = n16978 ^ n15951 ^ n2774 ;
  assign n16980 = ( n5520 & n7159 ) | ( n5520 & ~n16979 ) | ( n7159 & ~n16979 ) ;
  assign n16981 = ( n16976 & n16977 ) | ( n16976 & ~n16980 ) | ( n16977 & ~n16980 ) ;
  assign n16990 = ( x22 & n497 ) | ( x22 & ~n1790 ) | ( n497 & ~n1790 ) ;
  assign n16991 = ( n2732 & n6332 ) | ( n2732 & n16990 ) | ( n6332 & n16990 ) ;
  assign n16982 = n4880 ^ n1193 ^ n654 ;
  assign n16983 = x249 & ~n15811 ;
  assign n16984 = n3044 & n16983 ;
  assign n16985 = ( n327 & n770 ) | ( n327 & n4804 ) | ( n770 & n4804 ) ;
  assign n16986 = ( ~n16982 & n16984 ) | ( ~n16982 & n16985 ) | ( n16984 & n16985 ) ;
  assign n16987 = ( n1945 & ~n4289 ) | ( n1945 & n7183 ) | ( ~n4289 & n7183 ) ;
  assign n16988 = ( n666 & ~n9257 ) | ( n666 & n16987 ) | ( ~n9257 & n16987 ) ;
  assign n16989 = ( ~n8755 & n16986 ) | ( ~n8755 & n16988 ) | ( n16986 & n16988 ) ;
  assign n16992 = n16991 ^ n16989 ^ n8974 ;
  assign n16993 = ~n1861 & n16992 ;
  assign n16994 = ( ~n2251 & n12848 ) | ( ~n2251 & n16993 ) | ( n12848 & n16993 ) ;
  assign n16995 = ( x240 & n4428 ) | ( x240 & ~n5530 ) | ( n4428 & ~n5530 ) ;
  assign n16996 = ( n3342 & n7472 ) | ( n3342 & ~n16995 ) | ( n7472 & ~n16995 ) ;
  assign n16997 = ( n2369 & ~n5556 ) | ( n2369 & n9141 ) | ( ~n5556 & n9141 ) ;
  assign n16998 = n3930 ^ n1708 ^ n839 ;
  assign n16999 = ( n4820 & ~n15532 ) | ( n4820 & n16998 ) | ( ~n15532 & n16998 ) ;
  assign n17000 = ( n1154 & n11337 ) | ( n1154 & n16999 ) | ( n11337 & n16999 ) ;
  assign n17001 = ( n3031 & n16997 ) | ( n3031 & ~n17000 ) | ( n16997 & ~n17000 ) ;
  assign n17002 = n13304 ^ n4797 ^ n2804 ;
  assign n17003 = n17002 ^ n11080 ^ n2956 ;
  assign n17004 = ( n3262 & ~n3654 ) | ( n3262 & n14235 ) | ( ~n3654 & n14235 ) ;
  assign n17005 = n9983 ^ n788 ^ n313 ;
  assign n17006 = n17005 ^ n7412 ^ n6726 ;
  assign n17007 = n2647 & ~n17006 ;
  assign n17008 = n839 & n17007 ;
  assign n17009 = ~n4953 & n12007 ;
  assign n17010 = n17009 ^ n8929 ^ 1'b0 ;
  assign n17011 = n17010 ^ n14168 ^ n3846 ;
  assign n17012 = n17011 ^ n16993 ^ n11496 ;
  assign n17013 = n9057 ^ n8330 ^ n2875 ;
  assign n17019 = ( n663 & ~n2028 ) | ( n663 & n11199 ) | ( ~n2028 & n11199 ) ;
  assign n17020 = ( n1822 & n16524 ) | ( n1822 & ~n17019 ) | ( n16524 & ~n17019 ) ;
  assign n17014 = n1220 & n10817 ;
  assign n17015 = n17014 ^ n4022 ^ 1'b0 ;
  assign n17016 = n17015 ^ n2230 ^ n2100 ;
  assign n17017 = n12021 ^ n8134 ^ 1'b0 ;
  assign n17018 = n17016 & ~n17017 ;
  assign n17021 = n17020 ^ n17018 ^ 1'b0 ;
  assign n17022 = ( n4075 & ~n5993 ) | ( n4075 & n14155 ) | ( ~n5993 & n14155 ) ;
  assign n17023 = n17022 ^ n3202 ^ n3036 ;
  assign n17030 = n15195 ^ n10166 ^ n8254 ;
  assign n17024 = n5147 ^ n391 ^ 1'b0 ;
  assign n17025 = n12542 & ~n17024 ;
  assign n17026 = n17025 ^ n5711 ^ n3392 ;
  assign n17027 = n13143 | n17026 ;
  assign n17028 = n11120 & ~n17027 ;
  assign n17029 = ( n12360 & n13164 ) | ( n12360 & ~n17028 ) | ( n13164 & ~n17028 ) ;
  assign n17031 = n17030 ^ n17029 ^ 1'b0 ;
  assign n17032 = n17023 | n17031 ;
  assign n17033 = n11265 ^ n8198 ^ n5185 ;
  assign n17034 = ~n11427 & n17033 ;
  assign n17035 = n17034 ^ n10524 ^ 1'b0 ;
  assign n17036 = n10525 ^ n2421 ^ n1036 ;
  assign n17037 = ( n2644 & ~n4894 ) | ( n2644 & n12783 ) | ( ~n4894 & n12783 ) ;
  assign n17038 = ( n11469 & n12940 ) | ( n11469 & n17037 ) | ( n12940 & n17037 ) ;
  assign n17039 = n5394 ^ n2884 ^ 1'b0 ;
  assign n17040 = n5863 & n17039 ;
  assign n17041 = ( n6413 & ~n15717 ) | ( n6413 & n17040 ) | ( ~n15717 & n17040 ) ;
  assign n17043 = ( n4564 & n4643 ) | ( n4564 & n4879 ) | ( n4643 & n4879 ) ;
  assign n17042 = ( ~n1387 & n13578 ) | ( ~n1387 & n16169 ) | ( n13578 & n16169 ) ;
  assign n17044 = n17043 ^ n17042 ^ n7411 ;
  assign n17045 = n5553 ^ n5173 ^ n4217 ;
  assign n17046 = n17045 ^ n10820 ^ 1'b0 ;
  assign n17047 = n11936 | n17046 ;
  assign n17048 = ( ~n1016 & n4318 ) | ( ~n1016 & n9597 ) | ( n4318 & n9597 ) ;
  assign n17049 = ~n5751 & n17048 ;
  assign n17050 = n17049 ^ n2407 ^ 1'b0 ;
  assign n17051 = ( n7396 & ~n11726 ) | ( n7396 & n17050 ) | ( ~n11726 & n17050 ) ;
  assign n17061 = n11052 ^ n4129 ^ n710 ;
  assign n17060 = ( n3988 & n5113 ) | ( n3988 & n16570 ) | ( n5113 & n16570 ) ;
  assign n17062 = n17061 ^ n17060 ^ n1614 ;
  assign n17052 = ( ~n7049 & n7847 ) | ( ~n7049 & n11677 ) | ( n7847 & n11677 ) ;
  assign n17053 = ( n7618 & n10331 ) | ( n7618 & n16455 ) | ( n10331 & n16455 ) ;
  assign n17054 = ( n3725 & ~n17052 ) | ( n3725 & n17053 ) | ( ~n17052 & n17053 ) ;
  assign n17055 = ( n407 & n4341 ) | ( n407 & ~n5098 ) | ( n4341 & ~n5098 ) ;
  assign n17056 = ( ~n973 & n7653 ) | ( ~n973 & n17055 ) | ( n7653 & n17055 ) ;
  assign n17057 = ( ~n298 & n6487 ) | ( ~n298 & n17056 ) | ( n6487 & n17056 ) ;
  assign n17058 = ( x159 & n17054 ) | ( x159 & ~n17057 ) | ( n17054 & ~n17057 ) ;
  assign n17059 = ~n13536 & n17058 ;
  assign n17063 = n17062 ^ n17059 ^ 1'b0 ;
  assign n17064 = ( n17047 & n17051 ) | ( n17047 & n17063 ) | ( n17051 & n17063 ) ;
  assign n17066 = ~n9025 & n15944 ;
  assign n17065 = n3589 ^ n1856 ^ n743 ;
  assign n17067 = n17066 ^ n17065 ^ n8443 ;
  assign n17068 = ( n2481 & n3401 ) | ( n2481 & n9299 ) | ( n3401 & n9299 ) ;
  assign n17069 = ( ~n6309 & n17067 ) | ( ~n6309 & n17068 ) | ( n17067 & n17068 ) ;
  assign n17070 = n17069 ^ n13867 ^ n5530 ;
  assign n17071 = n4235 & ~n14360 ;
  assign n17072 = ( n3753 & ~n4422 ) | ( n3753 & n12961 ) | ( ~n4422 & n12961 ) ;
  assign n17073 = n17072 ^ n16070 ^ n5424 ;
  assign n17075 = n2280 | n13272 ;
  assign n17074 = ( ~n2765 & n3680 ) | ( ~n2765 & n5251 ) | ( n3680 & n5251 ) ;
  assign n17076 = n17075 ^ n17074 ^ n15530 ;
  assign n17077 = ( n1452 & n3601 ) | ( n1452 & n5767 ) | ( n3601 & n5767 ) ;
  assign n17078 = n12621 ^ n7529 ^ n3182 ;
  assign n17079 = n17078 ^ n4799 ^ n2800 ;
  assign n17080 = ( n12577 & n17077 ) | ( n12577 & n17079 ) | ( n17077 & n17079 ) ;
  assign n17081 = ( n17073 & n17076 ) | ( n17073 & n17080 ) | ( n17076 & n17080 ) ;
  assign n17082 = n16272 ^ n4940 ^ 1'b0 ;
  assign n17083 = n12834 | n17082 ;
  assign n17084 = n5843 ^ n4542 ^ n812 ;
  assign n17085 = n17084 ^ n16992 ^ 1'b0 ;
  assign n17086 = n17083 | n17085 ;
  assign n17087 = ( ~n9987 & n14354 ) | ( ~n9987 & n16962 ) | ( n14354 & n16962 ) ;
  assign n17088 = ( n3531 & n13664 ) | ( n3531 & ~n17087 ) | ( n13664 & ~n17087 ) ;
  assign n17089 = n2398 & ~n17088 ;
  assign n17090 = n9204 ^ n7898 ^ n3804 ;
  assign n17091 = n17090 ^ n11872 ^ n4141 ;
  assign n17092 = n13740 ^ n3510 ^ n2667 ;
  assign n17093 = ( n2564 & ~n3890 ) | ( n2564 & n17092 ) | ( ~n3890 & n17092 ) ;
  assign n17095 = n13025 ^ n4310 ^ n1898 ;
  assign n17094 = ( n5435 & ~n8500 ) | ( n5435 & n12790 ) | ( ~n8500 & n12790 ) ;
  assign n17096 = n17095 ^ n17094 ^ 1'b0 ;
  assign n17097 = n10985 ^ n10025 ^ n1813 ;
  assign n17098 = n13318 ^ n12161 ^ n11323 ;
  assign n17099 = n583 & n17098 ;
  assign n17100 = n17099 ^ n5276 ^ 1'b0 ;
  assign n17101 = ( n1178 & n17097 ) | ( n1178 & n17100 ) | ( n17097 & n17100 ) ;
  assign n17102 = n17101 ^ n8479 ^ n6717 ;
  assign n17103 = ( n3310 & n4381 ) | ( n3310 & n6553 ) | ( n4381 & n6553 ) ;
  assign n17104 = ( n8174 & ~n17098 ) | ( n8174 & n17103 ) | ( ~n17098 & n17103 ) ;
  assign n17105 = n10057 ^ n10010 ^ 1'b0 ;
  assign n17106 = n7771 & n17105 ;
  assign n17107 = n11785 ^ n1598 ^ x156 ;
  assign n17108 = n7239 ^ n6799 ^ n2432 ;
  assign n17109 = ~n5263 & n11211 ;
  assign n17110 = n17109 ^ n4564 ^ 1'b0 ;
  assign n17111 = ( n3992 & ~n17108 ) | ( n3992 & n17110 ) | ( ~n17108 & n17110 ) ;
  assign n17112 = n17107 | n17111 ;
  assign n17113 = n10813 ^ n2647 ^ n1740 ;
  assign n17114 = n14467 ^ n3974 ^ 1'b0 ;
  assign n17115 = n5259 & n17114 ;
  assign n17116 = ( ~n7138 & n13291 ) | ( ~n7138 & n17115 ) | ( n13291 & n17115 ) ;
  assign n17117 = n4545 ^ n1710 ^ 1'b0 ;
  assign n17118 = n6183 | n17117 ;
  assign n17119 = ( n4767 & ~n8807 ) | ( n4767 & n17118 ) | ( ~n8807 & n17118 ) ;
  assign n17120 = n12494 & n17119 ;
  assign n17121 = n8193 ^ n2797 ^ 1'b0 ;
  assign n17122 = n10941 ^ n534 ^ 1'b0 ;
  assign n17123 = n17122 ^ n16341 ^ n11429 ;
  assign n17124 = ~n2245 & n17123 ;
  assign n17125 = n17121 & n17124 ;
  assign n17126 = ( ~n8803 & n17120 ) | ( ~n8803 & n17125 ) | ( n17120 & n17125 ) ;
  assign n17127 = n2206 & n14729 ;
  assign n17128 = ~n4131 & n17127 ;
  assign n17132 = n7938 ^ n6875 ^ n5331 ;
  assign n17131 = n7514 ^ n2393 ^ 1'b0 ;
  assign n17129 = n10278 ^ n5554 ^ 1'b0 ;
  assign n17130 = n2274 & ~n17129 ;
  assign n17133 = n17132 ^ n17131 ^ n17130 ;
  assign n17134 = ( n6933 & ~n17128 ) | ( n6933 & n17133 ) | ( ~n17128 & n17133 ) ;
  assign n17135 = ( n846 & n3888 ) | ( n846 & ~n5008 ) | ( n3888 & ~n5008 ) ;
  assign n17136 = ( ~n2698 & n5835 ) | ( ~n2698 & n8104 ) | ( n5835 & n8104 ) ;
  assign n17137 = n17136 ^ n7832 ^ n2978 ;
  assign n17138 = ( ~n5897 & n8451 ) | ( ~n5897 & n17137 ) | ( n8451 & n17137 ) ;
  assign n17139 = n17135 & ~n17138 ;
  assign n17140 = n4170 & n6260 ;
  assign n17141 = n14177 ^ n7415 ^ 1'b0 ;
  assign n17142 = n8134 & n17141 ;
  assign n17143 = ( n10745 & ~n17140 ) | ( n10745 & n17142 ) | ( ~n17140 & n17142 ) ;
  assign n17144 = ( ~n3544 & n17139 ) | ( ~n3544 & n17143 ) | ( n17139 & n17143 ) ;
  assign n17146 = n10862 ^ n5961 ^ n3261 ;
  assign n17145 = n7581 ^ n1297 ^ 1'b0 ;
  assign n17147 = n17146 ^ n17145 ^ n9090 ;
  assign n17148 = n17147 ^ n10931 ^ n10088 ;
  assign n17149 = n7211 ^ n4873 ^ 1'b0 ;
  assign n17150 = n5189 & ~n17149 ;
  assign n17151 = ( n1289 & n9015 ) | ( n1289 & n10916 ) | ( n9015 & n10916 ) ;
  assign n17152 = ( n5707 & ~n17150 ) | ( n5707 & n17151 ) | ( ~n17150 & n17151 ) ;
  assign n17164 = n5916 ^ n4554 ^ 1'b0 ;
  assign n17165 = ( n2345 & ~n5427 ) | ( n2345 & n17164 ) | ( ~n5427 & n17164 ) ;
  assign n17166 = ( n6580 & n9998 ) | ( n6580 & n12647 ) | ( n9998 & n12647 ) ;
  assign n17167 = ( n14248 & ~n17165 ) | ( n14248 & n17166 ) | ( ~n17165 & n17166 ) ;
  assign n17154 = ( x199 & n3855 ) | ( x199 & ~n5921 ) | ( n3855 & ~n5921 ) ;
  assign n17153 = n4315 ^ n4229 ^ n2295 ;
  assign n17155 = n17154 ^ n17153 ^ n1008 ;
  assign n17156 = n8869 & n14484 ;
  assign n17157 = n17156 ^ n16685 ^ 1'b0 ;
  assign n17158 = ( n572 & n17155 ) | ( n572 & n17157 ) | ( n17155 & n17157 ) ;
  assign n17159 = n3805 ^ n1861 ^ 1'b0 ;
  assign n17160 = n15856 & ~n17159 ;
  assign n17161 = ~n2921 & n17160 ;
  assign n17162 = ( n3910 & ~n5726 ) | ( n3910 & n17161 ) | ( ~n5726 & n17161 ) ;
  assign n17163 = ( n10990 & n17158 ) | ( n10990 & ~n17162 ) | ( n17158 & ~n17162 ) ;
  assign n17168 = n17167 ^ n17163 ^ n12481 ;
  assign n17169 = n17168 ^ n5148 ^ 1'b0 ;
  assign n17170 = n2153 & n17169 ;
  assign n17174 = n11627 ^ n1439 ^ n473 ;
  assign n17175 = n17174 ^ n12753 ^ x239 ;
  assign n17172 = n2927 & ~n14091 ;
  assign n17171 = n1909 | n2389 ;
  assign n17173 = n17172 ^ n17171 ^ 1'b0 ;
  assign n17176 = n17175 ^ n17173 ^ n4390 ;
  assign n17177 = n14480 ^ n8163 ^ 1'b0 ;
  assign n17178 = n17177 ^ n8796 ^ 1'b0 ;
  assign n17185 = n17025 ^ x245 ^ 1'b0 ;
  assign n17179 = n4993 ^ n4750 ^ n4476 ;
  assign n17180 = n10504 ^ n8085 ^ n6345 ;
  assign n17181 = n17180 ^ n6530 ^ n1188 ;
  assign n17182 = n12028 ^ n2086 ^ 1'b0 ;
  assign n17183 = n17182 ^ n6472 ^ n5974 ;
  assign n17184 = ( ~n17179 & n17181 ) | ( ~n17179 & n17183 ) | ( n17181 & n17183 ) ;
  assign n17186 = n17185 ^ n17184 ^ n12288 ;
  assign n17187 = ( n7430 & ~n12405 ) | ( n7430 & n17186 ) | ( ~n12405 & n17186 ) ;
  assign n17188 = ~n17178 & n17187 ;
  assign n17189 = ~n13589 & n14253 ;
  assign n17190 = n17188 & n17189 ;
  assign n17191 = n8171 ^ n3622 ^ n692 ;
  assign n17192 = ~n7088 & n8124 ;
  assign n17193 = n17192 ^ n4888 ^ 1'b0 ;
  assign n17194 = ( n847 & ~n9323 ) | ( n847 & n17193 ) | ( ~n9323 & n17193 ) ;
  assign n17195 = ( ~n10277 & n14275 ) | ( ~n10277 & n17194 ) | ( n14275 & n17194 ) ;
  assign n17196 = n4007 & ~n6112 ;
  assign n17197 = n482 & n1393 ;
  assign n17198 = ( ~n556 & n6439 ) | ( ~n556 & n17197 ) | ( n6439 & n17197 ) ;
  assign n17199 = n17198 ^ n2987 ^ n2640 ;
  assign n17200 = n6334 | n17199 ;
  assign n17201 = n17200 ^ n3755 ^ 1'b0 ;
  assign n17202 = ( n4707 & n6981 ) | ( n4707 & n14811 ) | ( n6981 & n14811 ) ;
  assign n17203 = ( n578 & n6199 ) | ( n578 & n13660 ) | ( n6199 & n13660 ) ;
  assign n17204 = ( n5391 & ~n6464 ) | ( n5391 & n17203 ) | ( ~n6464 & n17203 ) ;
  assign n17205 = ( ~n17201 & n17202 ) | ( ~n17201 & n17204 ) | ( n17202 & n17204 ) ;
  assign n17206 = n11244 ^ n950 ^ 1'b0 ;
  assign n17207 = ( n2033 & n16030 ) | ( n2033 & n16211 ) | ( n16030 & n16211 ) ;
  assign n17208 = n4913 & ~n17207 ;
  assign n17209 = n17208 ^ n8273 ^ n5760 ;
  assign n17210 = n12697 ^ n1551 ^ 1'b0 ;
  assign n17211 = n6563 & ~n17210 ;
  assign n17212 = ( n2941 & ~n17209 ) | ( n2941 & n17211 ) | ( ~n17209 & n17211 ) ;
  assign n17219 = n635 | n1336 ;
  assign n17220 = n17219 ^ n3994 ^ 1'b0 ;
  assign n17221 = n3149 & ~n17220 ;
  assign n17214 = ( n521 & ~n3279 ) | ( n521 & n4922 ) | ( ~n3279 & n4922 ) ;
  assign n17215 = n17214 ^ n14096 ^ n3023 ;
  assign n17216 = ( n2327 & ~n12815 ) | ( n2327 & n17215 ) | ( ~n12815 & n17215 ) ;
  assign n17217 = n17216 ^ n7717 ^ 1'b0 ;
  assign n17218 = n8399 | n17217 ;
  assign n17222 = n17221 ^ n17218 ^ x241 ;
  assign n17213 = n2435 | n14803 ;
  assign n17223 = n17222 ^ n17213 ^ 1'b0 ;
  assign n17224 = n5587 & n17223 ;
  assign n17225 = ~n17212 & n17224 ;
  assign n17226 = ( n1697 & n2327 ) | ( n1697 & ~n5759 ) | ( n2327 & ~n5759 ) ;
  assign n17227 = n3227 & n17226 ;
  assign n17228 = n6452 & n17227 ;
  assign n17229 = ( n13285 & ~n15416 ) | ( n13285 & n17228 ) | ( ~n15416 & n17228 ) ;
  assign n17230 = n9211 ^ n6561 ^ 1'b0 ;
  assign n17231 = ( n582 & n969 ) | ( n582 & n2527 ) | ( n969 & n2527 ) ;
  assign n17232 = n17231 ^ n11731 ^ n8619 ;
  assign n17233 = ( n850 & n2884 ) | ( n850 & n6555 ) | ( n2884 & n6555 ) ;
  assign n17234 = ( n1937 & n2164 ) | ( n1937 & n17233 ) | ( n2164 & n17233 ) ;
  assign n17235 = ( n4562 & n17232 ) | ( n4562 & ~n17234 ) | ( n17232 & ~n17234 ) ;
  assign n17236 = ( ~n1041 & n5000 ) | ( ~n1041 & n6839 ) | ( n5000 & n6839 ) ;
  assign n17237 = n13106 ^ n3968 ^ n2291 ;
  assign n17238 = n16374 ^ n13002 ^ n4338 ;
  assign n17239 = ( n17236 & ~n17237 ) | ( n17236 & n17238 ) | ( ~n17237 & n17238 ) ;
  assign n17240 = n17172 ^ n16096 ^ 1'b0 ;
  assign n17241 = n12655 ^ n12340 ^ n1911 ;
  assign n17242 = n8665 ^ n3672 ^ n773 ;
  assign n17245 = ( x213 & ~n2836 ) | ( x213 & n5955 ) | ( ~n2836 & n5955 ) ;
  assign n17246 = n17245 ^ n15394 ^ n7609 ;
  assign n17243 = n11552 | n12929 ;
  assign n17244 = n2834 & ~n17243 ;
  assign n17247 = n17246 ^ n17244 ^ n11645 ;
  assign n17248 = ( ~n14944 & n17242 ) | ( ~n14944 & n17247 ) | ( n17242 & n17247 ) ;
  assign n17249 = ( n3742 & ~n17241 ) | ( n3742 & n17248 ) | ( ~n17241 & n17248 ) ;
  assign n17250 = n14165 ^ n8355 ^ n6387 ;
  assign n17251 = ( n2376 & n4875 ) | ( n2376 & ~n14997 ) | ( n4875 & ~n14997 ) ;
  assign n17252 = n8686 ^ n3134 ^ n2601 ;
  assign n17253 = ( ~n8129 & n17251 ) | ( ~n8129 & n17252 ) | ( n17251 & n17252 ) ;
  assign n17254 = x254 & ~n14364 ;
  assign n17255 = n336 & n17254 ;
  assign n17256 = ( n13887 & n17253 ) | ( n13887 & n17255 ) | ( n17253 & n17255 ) ;
  assign n17257 = n15679 ^ n14624 ^ n4580 ;
  assign n17258 = n8270 & ~n9601 ;
  assign n17259 = ( n6100 & n10470 ) | ( n6100 & ~n12729 ) | ( n10470 & ~n12729 ) ;
  assign n17260 = n11955 & ~n17259 ;
  assign n17261 = ( n7059 & n14975 ) | ( n7059 & ~n15035 ) | ( n14975 & ~n15035 ) ;
  assign n17262 = ( ~n1330 & n7902 ) | ( ~n1330 & n17261 ) | ( n7902 & n17261 ) ;
  assign n17266 = ( n5188 & n9268 ) | ( n5188 & n17061 ) | ( n9268 & n17061 ) ;
  assign n17263 = n4464 & n13664 ;
  assign n17264 = ~n6996 & n17263 ;
  assign n17265 = n17264 ^ n12784 ^ n2566 ;
  assign n17267 = n17266 ^ n17265 ^ n9352 ;
  assign n17268 = n17262 & ~n17267 ;
  assign n17271 = n12296 ^ n6005 ^ n4699 ;
  assign n17269 = ( ~n3654 & n6824 ) | ( ~n3654 & n8742 ) | ( n6824 & n8742 ) ;
  assign n17270 = ( n6088 & n12880 ) | ( n6088 & ~n17269 ) | ( n12880 & ~n17269 ) ;
  assign n17272 = n17271 ^ n17270 ^ n286 ;
  assign n17273 = ( n10237 & n11563 ) | ( n10237 & ~n13601 ) | ( n11563 & ~n13601 ) ;
  assign n17274 = n17273 ^ n11744 ^ x96 ;
  assign n17275 = n6291 ^ n4117 ^ n384 ;
  assign n17276 = ( x136 & ~n10709 ) | ( x136 & n17275 ) | ( ~n10709 & n17275 ) ;
  assign n17278 = n14659 ^ n3084 ^ n2267 ;
  assign n17277 = n10901 ^ n8946 ^ n2432 ;
  assign n17279 = n17278 ^ n17277 ^ n10930 ;
  assign n17280 = ( n922 & n17276 ) | ( n922 & n17279 ) | ( n17276 & n17279 ) ;
  assign n17281 = ( n1010 & n2902 ) | ( n1010 & n6664 ) | ( n2902 & n6664 ) ;
  assign n17282 = n368 & n17281 ;
  assign n17283 = n6676 & n17282 ;
  assign n17284 = ~n3958 & n17283 ;
  assign n17285 = n11194 & ~n17284 ;
  assign n17286 = n17285 ^ n2709 ^ 1'b0 ;
  assign n17287 = ( n4893 & n10719 ) | ( n4893 & ~n17286 ) | ( n10719 & ~n17286 ) ;
  assign n17288 = ( n13735 & ~n17280 ) | ( n13735 & n17287 ) | ( ~n17280 & n17287 ) ;
  assign n17294 = n8634 & n9010 ;
  assign n17292 = n9328 ^ n5477 ^ n513 ;
  assign n17289 = ( ~n1504 & n7593 ) | ( ~n1504 & n7618 ) | ( n7593 & n7618 ) ;
  assign n17290 = ( n8666 & n8983 ) | ( n8666 & ~n17289 ) | ( n8983 & ~n17289 ) ;
  assign n17291 = ( ~n984 & n16606 ) | ( ~n984 & n17290 ) | ( n16606 & n17290 ) ;
  assign n17293 = n17292 ^ n17291 ^ n7952 ;
  assign n17295 = n17294 ^ n17293 ^ 1'b0 ;
  assign n17296 = n17288 & n17295 ;
  assign n17297 = n2036 & ~n7165 ;
  assign n17298 = n7768 ^ n2761 ^ 1'b0 ;
  assign n17299 = n410 | n17298 ;
  assign n17300 = n17299 ^ n14976 ^ n13532 ;
  assign n17305 = n7747 ^ n7284 ^ n2241 ;
  assign n17303 = ( n3636 & n5457 ) | ( n3636 & n9299 ) | ( n5457 & n9299 ) ;
  assign n17302 = n10901 ^ n6747 ^ n5618 ;
  assign n17304 = n17303 ^ n17302 ^ n1793 ;
  assign n17301 = n15336 ^ n12977 ^ n1223 ;
  assign n17306 = n17305 ^ n17304 ^ n17301 ;
  assign n17307 = n6264 ^ n4289 ^ n1912 ;
  assign n17308 = n17307 ^ n5758 ^ n1717 ;
  assign n17309 = n17308 ^ n8458 ^ 1'b0 ;
  assign n17310 = n607 | n10439 ;
  assign n17311 = n17310 ^ n12510 ^ x36 ;
  assign n17312 = ( n11464 & n11569 ) | ( n11464 & n13532 ) | ( n11569 & n13532 ) ;
  assign n17313 = n17312 ^ n11315 ^ n10161 ;
  assign n17314 = ( ~n10658 & n11058 ) | ( ~n10658 & n17313 ) | ( n11058 & n17313 ) ;
  assign n17315 = ( n785 & n6234 ) | ( n785 & ~n17314 ) | ( n6234 & ~n17314 ) ;
  assign n17316 = ( n17309 & n17311 ) | ( n17309 & n17315 ) | ( n17311 & n17315 ) ;
  assign n17317 = n3089 ^ n1824 ^ n1600 ;
  assign n17318 = ( n1481 & ~n3780 ) | ( n1481 & n17317 ) | ( ~n3780 & n17317 ) ;
  assign n17319 = n5878 & n17318 ;
  assign n17320 = ~n5615 & n17319 ;
  assign n17321 = n556 & ~n6999 ;
  assign n17322 = n17321 ^ n3294 ^ 1'b0 ;
  assign n17323 = ( ~n3805 & n17320 ) | ( ~n3805 & n17322 ) | ( n17320 & n17322 ) ;
  assign n17324 = n12441 ^ n12262 ^ n9503 ;
  assign n17325 = ( ~n9140 & n17323 ) | ( ~n9140 & n17324 ) | ( n17323 & n17324 ) ;
  assign n17327 = n7361 ^ n4670 ^ n907 ;
  assign n17326 = n7576 & n12440 ;
  assign n17328 = n17327 ^ n17326 ^ 1'b0 ;
  assign n17329 = ( n4408 & ~n5450 ) | ( n4408 & n17328 ) | ( ~n5450 & n17328 ) ;
  assign n17330 = n4718 & n6226 ;
  assign n17331 = n13134 & n17330 ;
  assign n17332 = n17331 ^ n11210 ^ n6534 ;
  assign n17333 = n8220 ^ n6241 ^ 1'b0 ;
  assign n17334 = ( n689 & n16743 ) | ( n689 & n17333 ) | ( n16743 & n17333 ) ;
  assign n17335 = n17334 ^ n16631 ^ n10156 ;
  assign n17336 = n2532 ^ n2397 ^ 1'b0 ;
  assign n17337 = n17336 ^ n12007 ^ n9090 ;
  assign n17338 = ( n17332 & n17335 ) | ( n17332 & ~n17337 ) | ( n17335 & ~n17337 ) ;
  assign n17339 = n8943 ^ n7943 ^ 1'b0 ;
  assign n17340 = n17339 ^ n13987 ^ 1'b0 ;
  assign n17341 = ( ~n14227 & n17338 ) | ( ~n14227 & n17340 ) | ( n17338 & n17340 ) ;
  assign n17342 = ( ~n9627 & n11230 ) | ( ~n9627 & n15517 ) | ( n11230 & n15517 ) ;
  assign n17343 = n13259 ^ n11379 ^ n3602 ;
  assign n17344 = ( n2600 & n5891 ) | ( n2600 & n17343 ) | ( n5891 & n17343 ) ;
  assign n17348 = n5344 ^ n3655 ^ n3303 ;
  assign n17349 = ( ~n8842 & n11720 ) | ( ~n8842 & n17348 ) | ( n11720 & n17348 ) ;
  assign n17350 = n11563 & n17349 ;
  assign n17351 = n17350 ^ n10392 ^ n7650 ;
  assign n17345 = ( n1905 & n7509 ) | ( n1905 & ~n15197 ) | ( n7509 & ~n15197 ) ;
  assign n17346 = ( n2236 & n6057 ) | ( n2236 & n12779 ) | ( n6057 & n12779 ) ;
  assign n17347 = ( ~n9229 & n17345 ) | ( ~n9229 & n17346 ) | ( n17345 & n17346 ) ;
  assign n17352 = n17351 ^ n17347 ^ n11667 ;
  assign n17356 = ( n1002 & ~n2843 ) | ( n1002 & n10326 ) | ( ~n2843 & n10326 ) ;
  assign n17354 = ~n2943 & n3818 ;
  assign n17355 = ~n10227 & n17354 ;
  assign n17357 = n17356 ^ n17355 ^ n1186 ;
  assign n17353 = ( ~n320 & n9408 ) | ( ~n320 & n10476 ) | ( n9408 & n10476 ) ;
  assign n17358 = n17357 ^ n17353 ^ n15729 ;
  assign n17359 = n16034 ^ n11591 ^ 1'b0 ;
  assign n17360 = n11406 & n17359 ;
  assign n17361 = n17360 ^ n13662 ^ 1'b0 ;
  assign n17365 = n13589 ^ n4830 ^ n2175 ;
  assign n17366 = ( x97 & ~n3054 ) | ( x97 & n17365 ) | ( ~n3054 & n17365 ) ;
  assign n17362 = ( n1652 & n6696 ) | ( n1652 & ~n7233 ) | ( n6696 & ~n7233 ) ;
  assign n17363 = n17362 ^ n11877 ^ x180 ;
  assign n17364 = ( n5521 & n6684 ) | ( n5521 & ~n17363 ) | ( n6684 & ~n17363 ) ;
  assign n17367 = n17366 ^ n17364 ^ n6235 ;
  assign n17368 = n13294 ^ n3573 ^ n3152 ;
  assign n17369 = n16959 ^ n13994 ^ n8577 ;
  assign n17370 = n6574 ^ n4222 ^ n374 ;
  assign n17371 = ( n2331 & n17369 ) | ( n2331 & ~n17370 ) | ( n17369 & ~n17370 ) ;
  assign n17372 = n17371 ^ n15562 ^ n8200 ;
  assign n17373 = n8450 ^ n6216 ^ n1940 ;
  assign n17374 = ( x138 & n1309 ) | ( x138 & n17373 ) | ( n1309 & n17373 ) ;
  assign n17375 = ( n7499 & n9159 ) | ( n7499 & ~n10091 ) | ( n9159 & ~n10091 ) ;
  assign n17376 = n13138 ^ n9988 ^ n5835 ;
  assign n17377 = n17376 ^ n16624 ^ n12297 ;
  assign n17378 = n17377 ^ n12812 ^ n2514 ;
  assign n17379 = ( ~n2052 & n11222 ) | ( ~n2052 & n11671 ) | ( n11222 & n11671 ) ;
  assign n17380 = n17379 ^ n7333 ^ 1'b0 ;
  assign n17381 = n6898 | n17380 ;
  assign n17382 = ( ~n17375 & n17378 ) | ( ~n17375 & n17381 ) | ( n17378 & n17381 ) ;
  assign n17383 = n17374 | n17382 ;
  assign n17384 = ( ~n13584 & n16933 ) | ( ~n13584 & n17383 ) | ( n16933 & n17383 ) ;
  assign n17385 = n6269 | n7286 ;
  assign n17386 = ( n2752 & n5091 ) | ( n2752 & n8425 ) | ( n5091 & n8425 ) ;
  assign n17387 = n17386 ^ n10367 ^ n7881 ;
  assign n17388 = n4496 ^ n905 ^ n851 ;
  assign n17389 = n17388 ^ n1991 ^ 1'b0 ;
  assign n17390 = n17389 ^ n10440 ^ 1'b0 ;
  assign n17391 = ( n4627 & ~n17387 ) | ( n4627 & n17390 ) | ( ~n17387 & n17390 ) ;
  assign n17392 = n16890 ^ n12057 ^ n4223 ;
  assign n17393 = ( n625 & n3098 ) | ( n625 & n17392 ) | ( n3098 & n17392 ) ;
  assign n17394 = ( ~n1865 & n8268 ) | ( ~n1865 & n15133 ) | ( n8268 & n15133 ) ;
  assign n17395 = n5077 & n17394 ;
  assign n17396 = ~n2570 & n17395 ;
  assign n17397 = n7610 & ~n16640 ;
  assign n17398 = n17397 ^ n675 ^ 1'b0 ;
  assign n17399 = ( ~n3700 & n14994 ) | ( ~n3700 & n17398 ) | ( n14994 & n17398 ) ;
  assign n17400 = ( n3877 & n4837 ) | ( n3877 & n17311 ) | ( n4837 & n17311 ) ;
  assign n17401 = ( n1015 & n3473 ) | ( n1015 & ~n11897 ) | ( n3473 & ~n11897 ) ;
  assign n17402 = ( n4617 & n8699 ) | ( n4617 & n17401 ) | ( n8699 & n17401 ) ;
  assign n17403 = n17402 ^ n14735 ^ n10849 ;
  assign n17404 = ( ~n6079 & n10855 ) | ( ~n6079 & n17403 ) | ( n10855 & n17403 ) ;
  assign n17405 = ~n4916 & n10474 ;
  assign n17406 = ( n3448 & n4701 ) | ( n3448 & n16208 ) | ( n4701 & n16208 ) ;
  assign n17407 = ( n6585 & ~n9831 ) | ( n6585 & n17406 ) | ( ~n9831 & n17406 ) ;
  assign n17408 = n15312 ^ n8025 ^ n3098 ;
  assign n17410 = n3893 | n6705 ;
  assign n17411 = n17410 ^ n10345 ^ 1'b0 ;
  assign n17409 = n8789 & ~n9464 ;
  assign n17412 = n17411 ^ n17409 ^ n2122 ;
  assign n17413 = ( n17407 & ~n17408 ) | ( n17407 & n17412 ) | ( ~n17408 & n17412 ) ;
  assign n17414 = n7264 ^ n3540 ^ n1114 ;
  assign n17415 = n5980 ^ n5672 ^ n1104 ;
  assign n17416 = n4358 & ~n15353 ;
  assign n17417 = n1702 & n17416 ;
  assign n17418 = ( n4702 & ~n6160 ) | ( n4702 & n17417 ) | ( ~n6160 & n17417 ) ;
  assign n17419 = n2168 ^ x47 ^ 1'b0 ;
  assign n17420 = n6667 & n17419 ;
  assign n17421 = ( x107 & n6601 ) | ( x107 & n17420 ) | ( n6601 & n17420 ) ;
  assign n17422 = n17421 ^ n14739 ^ 1'b0 ;
  assign n17423 = ( n7175 & ~n17418 ) | ( n7175 & n17422 ) | ( ~n17418 & n17422 ) ;
  assign n17424 = ( ~n15752 & n17415 ) | ( ~n15752 & n17423 ) | ( n17415 & n17423 ) ;
  assign n17425 = n17378 ^ n15314 ^ 1'b0 ;
  assign n17426 = ( n4134 & ~n17424 ) | ( n4134 & n17425 ) | ( ~n17424 & n17425 ) ;
  assign n17427 = ( n13461 & ~n17414 ) | ( n13461 & n17426 ) | ( ~n17414 & n17426 ) ;
  assign n17428 = ( n17405 & n17413 ) | ( n17405 & n17427 ) | ( n17413 & n17427 ) ;
  assign n17429 = ( n13424 & ~n13500 ) | ( n13424 & n14671 ) | ( ~n13500 & n14671 ) ;
  assign n17430 = ~x144 & n3240 ;
  assign n17431 = ( n1468 & n12140 ) | ( n1468 & ~n17430 ) | ( n12140 & ~n17430 ) ;
  assign n17432 = ( n8788 & ~n17429 ) | ( n8788 & n17431 ) | ( ~n17429 & n17431 ) ;
  assign n17433 = n17432 ^ n14057 ^ n13584 ;
  assign n17434 = n2857 & n3768 ;
  assign n17435 = n3441 ^ n1146 ^ 1'b0 ;
  assign n17436 = n10193 & ~n17435 ;
  assign n17437 = ( n2080 & ~n17434 ) | ( n2080 & n17436 ) | ( ~n17434 & n17436 ) ;
  assign n17443 = n6652 ^ n4599 ^ x50 ;
  assign n17438 = n2672 ^ n2427 ^ n2393 ;
  assign n17439 = n7767 ^ n6498 ^ n4103 ;
  assign n17440 = n3949 & ~n17439 ;
  assign n17441 = ( n3734 & n17438 ) | ( n3734 & ~n17440 ) | ( n17438 & ~n17440 ) ;
  assign n17442 = n17441 ^ n12495 ^ x197 ;
  assign n17444 = n17443 ^ n17442 ^ n14924 ;
  assign n17445 = n10725 ^ n2061 ^ n882 ;
  assign n17446 = ( n10955 & n13631 ) | ( n10955 & ~n17445 ) | ( n13631 & ~n17445 ) ;
  assign n17447 = n8955 & n17446 ;
  assign n17448 = ~n11866 & n17447 ;
  assign n17449 = n9087 ^ n1373 ^ 1'b0 ;
  assign n17450 = ( n1279 & ~n17140 ) | ( n1279 & n17449 ) | ( ~n17140 & n17449 ) ;
  assign n17454 = n14724 ^ n4464 ^ n2869 ;
  assign n17452 = ( n762 & ~n4986 ) | ( n762 & n8928 ) | ( ~n4986 & n8928 ) ;
  assign n17451 = n7490 ^ n3730 ^ n2329 ;
  assign n17453 = n17452 ^ n17451 ^ n2464 ;
  assign n17455 = n17454 ^ n17453 ^ n3980 ;
  assign n17456 = n7554 ^ n7432 ^ n4092 ;
  assign n17457 = ( ~n2908 & n5599 ) | ( ~n2908 & n17456 ) | ( n5599 & n17456 ) ;
  assign n17458 = ( ~n1481 & n4093 ) | ( ~n1481 & n5677 ) | ( n4093 & n5677 ) ;
  assign n17459 = n17458 ^ n608 ^ 1'b0 ;
  assign n17460 = n5824 & ~n17459 ;
  assign n17461 = ( ~n7259 & n12113 ) | ( ~n7259 & n17460 ) | ( n12113 & n17460 ) ;
  assign n17462 = n17457 & n17461 ;
  assign n17463 = n7389 ^ n3496 ^ n1614 ;
  assign n17464 = n17463 ^ n10631 ^ n1974 ;
  assign n17465 = n13564 & ~n17464 ;
  assign n17466 = n17465 ^ n15324 ^ 1'b0 ;
  assign n17467 = ( n1649 & ~n1666 ) | ( n1649 & n16034 ) | ( ~n1666 & n16034 ) ;
  assign n17468 = ( n1822 & n5051 ) | ( n1822 & ~n7089 ) | ( n5051 & ~n7089 ) ;
  assign n17469 = n17468 ^ n4722 ^ n1485 ;
  assign n17470 = n17469 ^ n6004 ^ n4440 ;
  assign n17471 = ( ~n4355 & n11881 ) | ( ~n4355 & n17470 ) | ( n11881 & n17470 ) ;
  assign n17472 = ( ~n11318 & n17467 ) | ( ~n11318 & n17471 ) | ( n17467 & n17471 ) ;
  assign n17473 = ( n7270 & ~n14548 ) | ( n7270 & n17472 ) | ( ~n14548 & n17472 ) ;
  assign n17479 = ( n514 & ~n622 ) | ( n514 & n7324 ) | ( ~n622 & n7324 ) ;
  assign n17480 = n17479 ^ n1822 ^ 1'b0 ;
  assign n17477 = n7398 ^ n6971 ^ n3719 ;
  assign n17478 = ( n7656 & n10930 ) | ( n7656 & n17477 ) | ( n10930 & n17477 ) ;
  assign n17481 = n17480 ^ n17478 ^ n11566 ;
  assign n17474 = n7247 ^ n4244 ^ n1690 ;
  assign n17475 = n17474 ^ n3513 ^ n823 ;
  assign n17476 = n7264 & ~n17475 ;
  assign n17482 = n17481 ^ n17476 ^ 1'b0 ;
  assign n17483 = n17482 ^ n1065 ^ n510 ;
  assign n17484 = n8270 ^ n7509 ^ n2196 ;
  assign n17485 = n6929 & n10631 ;
  assign n17486 = n17485 ^ n8990 ^ 1'b0 ;
  assign n17487 = ( n2221 & n3495 ) | ( n2221 & ~n17486 ) | ( n3495 & ~n17486 ) ;
  assign n17488 = n17487 ^ n4614 ^ 1'b0 ;
  assign n17489 = n12502 & n17488 ;
  assign n17490 = ( ~n4659 & n9408 ) | ( ~n4659 & n13509 ) | ( n9408 & n13509 ) ;
  assign n17491 = ( n11308 & n17489 ) | ( n11308 & ~n17490 ) | ( n17489 & ~n17490 ) ;
  assign n17492 = n9164 ^ n7289 ^ n3718 ;
  assign n17493 = ( n10758 & n15773 ) | ( n10758 & ~n17492 ) | ( n15773 & ~n17492 ) ;
  assign n17494 = ( n17484 & ~n17491 ) | ( n17484 & n17493 ) | ( ~n17491 & n17493 ) ;
  assign n17495 = n3195 & ~n4292 ;
  assign n17496 = n17495 ^ n1825 ^ 1'b0 ;
  assign n17497 = n17496 ^ n2511 ^ n1239 ;
  assign n17498 = n12693 ^ n12235 ^ n1235 ;
  assign n17499 = n17199 ^ n11071 ^ n3989 ;
  assign n17500 = ( n17497 & n17498 ) | ( n17497 & ~n17499 ) | ( n17498 & ~n17499 ) ;
  assign n17501 = n2366 ^ n979 ^ 1'b0 ;
  assign n17502 = n17501 ^ n10841 ^ n9599 ;
  assign n17503 = n1611 | n16090 ;
  assign n17504 = n17503 ^ n2426 ^ n480 ;
  assign n17505 = n3541 & n17504 ;
  assign n17506 = n17505 ^ n824 ^ 1'b0 ;
  assign n17507 = ( n2935 & n13040 ) | ( n2935 & n15668 ) | ( n13040 & n15668 ) ;
  assign n17508 = n2957 | n5817 ;
  assign n17509 = n7554 & ~n17508 ;
  assign n17510 = ( n1184 & n14846 ) | ( n1184 & n17509 ) | ( n14846 & n17509 ) ;
  assign n17511 = n15777 | n17510 ;
  assign n17512 = n17090 | n17511 ;
  assign n17513 = n17512 ^ n5145 ^ n933 ;
  assign n17514 = ( n10822 & ~n17507 ) | ( n10822 & n17513 ) | ( ~n17507 & n17513 ) ;
  assign n17519 = n9950 ^ n1164 ^ n889 ;
  assign n17520 = n17519 ^ x34 ^ 1'b0 ;
  assign n17521 = n17520 ^ n13010 ^ 1'b0 ;
  assign n17522 = n6238 | n17521 ;
  assign n17515 = n5946 & ~n9063 ;
  assign n17516 = ~n972 & n5902 ;
  assign n17517 = n17516 ^ n7019 ^ 1'b0 ;
  assign n17518 = n17515 | n17517 ;
  assign n17523 = n17522 ^ n17518 ^ 1'b0 ;
  assign n17529 = ~n4805 & n5350 ;
  assign n17530 = ~n12988 & n17529 ;
  assign n17531 = ( n6560 & ~n11528 ) | ( n6560 & n17530 ) | ( ~n11528 & n17530 ) ;
  assign n17532 = ( ~n3749 & n4386 ) | ( ~n3749 & n10328 ) | ( n4386 & n10328 ) ;
  assign n17533 = n17532 ^ n13192 ^ n9103 ;
  assign n17534 = ( n10857 & ~n17531 ) | ( n10857 & n17533 ) | ( ~n17531 & n17533 ) ;
  assign n17535 = n10411 | n17534 ;
  assign n17526 = ( n1348 & ~n6849 ) | ( n1348 & n16786 ) | ( ~n6849 & n16786 ) ;
  assign n17524 = n6715 ^ x44 ^ 1'b0 ;
  assign n17525 = n17524 ^ n2240 ^ 1'b0 ;
  assign n17527 = n17526 ^ n17525 ^ 1'b0 ;
  assign n17528 = n17527 ^ n13357 ^ n1186 ;
  assign n17536 = n17535 ^ n17528 ^ 1'b0 ;
  assign n17537 = n9653 & n17536 ;
  assign n17538 = ( n3526 & n9645 ) | ( n3526 & ~n15171 ) | ( n9645 & ~n15171 ) ;
  assign n17542 = ( ~n1550 & n3267 ) | ( ~n1550 & n4565 ) | ( n3267 & n4565 ) ;
  assign n17540 = n6938 ^ x140 ^ 1'b0 ;
  assign n17539 = ( n4637 & n7134 ) | ( n4637 & n14285 ) | ( n7134 & n14285 ) ;
  assign n17541 = n17540 ^ n17539 ^ n513 ;
  assign n17543 = n17542 ^ n17541 ^ n17030 ;
  assign n17544 = ( ~x245 & n3874 ) | ( ~x245 & n7076 ) | ( n3874 & n7076 ) ;
  assign n17545 = ( n4707 & n6221 ) | ( n4707 & n17544 ) | ( n6221 & n17544 ) ;
  assign n17546 = n17545 ^ n13950 ^ n12869 ;
  assign n17547 = ( n3560 & n17074 ) | ( n3560 & n17546 ) | ( n17074 & n17546 ) ;
  assign n17548 = n17547 ^ n6362 ^ n298 ;
  assign n17549 = n17548 ^ n9134 ^ 1'b0 ;
  assign n17550 = ~n10191 & n17549 ;
  assign n17551 = n11100 ^ n9482 ^ x176 ;
  assign n17552 = n4909 & ~n9121 ;
  assign n17553 = ~n17551 & n17552 ;
  assign n17554 = n17553 ^ n15506 ^ n8371 ;
  assign n17555 = ( x178 & n3240 ) | ( x178 & n5295 ) | ( n3240 & n5295 ) ;
  assign n17556 = ( n9041 & n17554 ) | ( n9041 & n17555 ) | ( n17554 & n17555 ) ;
  assign n17557 = ( n7047 & n13833 ) | ( n7047 & n15010 ) | ( n13833 & n15010 ) ;
  assign n17561 = n5088 | n12121 ;
  assign n17558 = ( n2626 & ~n8758 ) | ( n2626 & n11829 ) | ( ~n8758 & n11829 ) ;
  assign n17559 = n17558 ^ n12512 ^ 1'b0 ;
  assign n17560 = ~n4945 & n17559 ;
  assign n17562 = n17561 ^ n17560 ^ n12272 ;
  assign n17563 = n15921 ^ n2097 ^ n1879 ;
  assign n17564 = ( n7060 & n15897 ) | ( n7060 & n17563 ) | ( n15897 & n17563 ) ;
  assign n17565 = n4931 & ~n17564 ;
  assign n17566 = ( n14149 & ~n17562 ) | ( n14149 & n17565 ) | ( ~n17562 & n17565 ) ;
  assign n17570 = ( n1150 & n5540 ) | ( n1150 & ~n7947 ) | ( n5540 & ~n7947 ) ;
  assign n17571 = ( ~n7274 & n7370 ) | ( ~n7274 & n17570 ) | ( n7370 & n17570 ) ;
  assign n17567 = ( n2171 & n9536 ) | ( n2171 & ~n10118 ) | ( n9536 & ~n10118 ) ;
  assign n17568 = n17567 ^ n11147 ^ 1'b0 ;
  assign n17569 = n17568 ^ n4968 ^ n3417 ;
  assign n17572 = n17571 ^ n17569 ^ n4238 ;
  assign n17573 = n17572 ^ n11856 ^ n2723 ;
  assign n17574 = ( ~n8919 & n11614 ) | ( ~n8919 & n13095 ) | ( n11614 & n13095 ) ;
  assign n17575 = n16430 & ~n17574 ;
  assign n17576 = ( x101 & n4714 ) | ( x101 & n17077 ) | ( n4714 & n17077 ) ;
  assign n17577 = n12047 ^ n5749 ^ 1'b0 ;
  assign n17578 = n9189 & n17577 ;
  assign n17579 = n17578 ^ n8578 ^ 1'b0 ;
  assign n17580 = ~n17576 & n17579 ;
  assign n17585 = ( n659 & n3927 ) | ( n659 & ~n4339 ) | ( n3927 & ~n4339 ) ;
  assign n17586 = ( ~n3822 & n8024 ) | ( ~n3822 & n17585 ) | ( n8024 & n17585 ) ;
  assign n17587 = ( n5877 & n10091 ) | ( n5877 & n17586 ) | ( n10091 & n17586 ) ;
  assign n17581 = ( n1298 & n7536 ) | ( n1298 & n7745 ) | ( n7536 & n7745 ) ;
  assign n17582 = ( ~n2947 & n8969 ) | ( ~n2947 & n10558 ) | ( n8969 & n10558 ) ;
  assign n17583 = ( n2505 & n17581 ) | ( n2505 & n17582 ) | ( n17581 & n17582 ) ;
  assign n17584 = ( n1841 & n9911 ) | ( n1841 & n17583 ) | ( n9911 & n17583 ) ;
  assign n17588 = n17587 ^ n17584 ^ n1181 ;
  assign n17589 = ( n3068 & ~n17580 ) | ( n3068 & n17588 ) | ( ~n17580 & n17588 ) ;
  assign n17590 = n13710 ^ n4326 ^ n3003 ;
  assign n17593 = n13788 ^ n10144 ^ n8968 ;
  assign n17592 = n10246 ^ n9420 ^ n6477 ;
  assign n17591 = ~n2907 & n3134 ;
  assign n17594 = n17593 ^ n17592 ^ n17591 ;
  assign n17595 = n15187 ^ n9347 ^ n4118 ;
  assign n17596 = n2180 & n17595 ;
  assign n17597 = n17596 ^ n15238 ^ 1'b0 ;
  assign n17598 = n17597 ^ x144 ^ 1'b0 ;
  assign n17599 = ~n17594 & n17598 ;
  assign n17600 = ( n11032 & n12124 ) | ( n11032 & n17599 ) | ( n12124 & n17599 ) ;
  assign n17601 = ( n966 & n17590 ) | ( n966 & ~n17600 ) | ( n17590 & ~n17600 ) ;
  assign n17606 = ( n8838 & n9980 ) | ( n8838 & ~n14726 ) | ( n9980 & ~n14726 ) ;
  assign n17604 = ( n1207 & ~n2264 ) | ( n1207 & n8430 ) | ( ~n2264 & n8430 ) ;
  assign n17602 = ( n1167 & ~n3579 ) | ( n1167 & n4935 ) | ( ~n3579 & n4935 ) ;
  assign n17603 = ( n10148 & n10541 ) | ( n10148 & ~n17602 ) | ( n10541 & ~n17602 ) ;
  assign n17605 = n17604 ^ n17603 ^ n1315 ;
  assign n17607 = n17606 ^ n17605 ^ 1'b0 ;
  assign n17612 = ( n1788 & n2026 ) | ( n1788 & n9868 ) | ( n2026 & n9868 ) ;
  assign n17611 = n10815 ^ n6141 ^ n4513 ;
  assign n17613 = n17612 ^ n17611 ^ n2020 ;
  assign n17614 = n17613 ^ n1342 ^ 1'b0 ;
  assign n17615 = ~n12260 & n17614 ;
  assign n17608 = n8458 ^ n4031 ^ n2006 ;
  assign n17609 = n17608 ^ n12960 ^ n1579 ;
  assign n17610 = ( n13354 & n14575 ) | ( n13354 & n17609 ) | ( n14575 & n17609 ) ;
  assign n17616 = n17615 ^ n17610 ^ n17471 ;
  assign n17617 = ( n5452 & n8880 ) | ( n5452 & n9949 ) | ( n8880 & n9949 ) ;
  assign n17618 = ( n4656 & n11549 ) | ( n4656 & ~n17617 ) | ( n11549 & ~n17617 ) ;
  assign n17619 = ( n7478 & ~n10637 ) | ( n7478 & n17618 ) | ( ~n10637 & n17618 ) ;
  assign n17620 = n15369 ^ n10592 ^ n2074 ;
  assign n17621 = ~n6625 & n6782 ;
  assign n17622 = n17621 ^ n888 ^ 1'b0 ;
  assign n17623 = n10527 ^ n9280 ^ n5969 ;
  assign n17624 = ( n13365 & n17622 ) | ( n13365 & ~n17623 ) | ( n17622 & ~n17623 ) ;
  assign n17625 = ( ~n1567 & n17620 ) | ( ~n1567 & n17624 ) | ( n17620 & n17624 ) ;
  assign n17626 = n9260 & ~n12386 ;
  assign n17627 = n17626 ^ n16243 ^ 1'b0 ;
  assign n17628 = n7099 | n17627 ;
  assign n17629 = n17628 ^ n6861 ^ 1'b0 ;
  assign n17630 = n17629 ^ n10848 ^ n2476 ;
  assign n17631 = n11497 ^ n10292 ^ x252 ;
  assign n17632 = ( n2298 & n2572 ) | ( n2298 & ~n7895 ) | ( n2572 & ~n7895 ) ;
  assign n17633 = ( ~n868 & n17631 ) | ( ~n868 & n17632 ) | ( n17631 & n17632 ) ;
  assign n17634 = n4387 ^ n1905 ^ n780 ;
  assign n17635 = ( n1201 & ~n4031 ) | ( n1201 & n11856 ) | ( ~n4031 & n11856 ) ;
  assign n17636 = ( n6490 & n17634 ) | ( n6490 & ~n17635 ) | ( n17634 & ~n17635 ) ;
  assign n17637 = x225 & ~n9937 ;
  assign n17638 = n17636 & n17637 ;
  assign n17640 = n7399 ^ n5347 ^ n824 ;
  assign n17639 = n14060 ^ n8347 ^ n597 ;
  assign n17641 = n17640 ^ n17639 ^ n6767 ;
  assign n17642 = n4584 & n17641 ;
  assign n17643 = ( ~n527 & n1239 ) | ( ~n527 & n17642 ) | ( n1239 & n17642 ) ;
  assign n17662 = n1716 ^ n1321 ^ x68 ;
  assign n17663 = ( ~n12485 & n13919 ) | ( ~n12485 & n17662 ) | ( n13919 & n17662 ) ;
  assign n17646 = n14339 ^ n3812 ^ n3471 ;
  assign n17644 = n1358 & n14538 ;
  assign n17645 = ( n13839 & ~n14101 ) | ( n13839 & n17644 ) | ( ~n14101 & n17644 ) ;
  assign n17647 = n17646 ^ n17645 ^ n10730 ;
  assign n17648 = n2751 | n17647 ;
  assign n17649 = n17648 ^ n8194 ^ 1'b0 ;
  assign n17657 = n972 | n7203 ;
  assign n17658 = n17657 ^ n6273 ^ n4571 ;
  assign n17659 = n7739 & n17658 ;
  assign n17650 = n10809 ^ n9421 ^ n8760 ;
  assign n17651 = n5593 ^ n4413 ^ n2664 ;
  assign n17652 = n17651 ^ n5527 ^ n890 ;
  assign n17653 = ( n502 & n9589 ) | ( n502 & ~n17652 ) | ( n9589 & ~n17652 ) ;
  assign n17654 = n17653 ^ n11588 ^ 1'b0 ;
  assign n17655 = ~n17650 & n17654 ;
  assign n17656 = ( n4928 & ~n5932 ) | ( n4928 & n17655 ) | ( ~n5932 & n17655 ) ;
  assign n17660 = n17659 ^ n17656 ^ n11523 ;
  assign n17661 = n17649 & ~n17660 ;
  assign n17664 = n17663 ^ n17661 ^ 1'b0 ;
  assign n17667 = n9125 ^ n605 ^ 1'b0 ;
  assign n17668 = ( ~n7574 & n9099 ) | ( ~n7574 & n17667 ) | ( n9099 & n17667 ) ;
  assign n17665 = ( n5176 & n12933 ) | ( n5176 & n15775 ) | ( n12933 & n15775 ) ;
  assign n17666 = n17665 ^ n7722 ^ n5800 ;
  assign n17669 = n17668 ^ n17666 ^ n8382 ;
  assign n17673 = n4010 & ~n13804 ;
  assign n17674 = n17673 ^ n5586 ^ 1'b0 ;
  assign n17670 = n7988 ^ n4463 ^ n1413 ;
  assign n17671 = n5473 & n12264 ;
  assign n17672 = ( n1928 & ~n17670 ) | ( n1928 & n17671 ) | ( ~n17670 & n17671 ) ;
  assign n17675 = n17674 ^ n17672 ^ n7064 ;
  assign n17678 = ( n806 & n3851 ) | ( n806 & n5827 ) | ( n3851 & n5827 ) ;
  assign n17676 = ( ~n1136 & n12971 ) | ( ~n1136 & n16954 ) | ( n12971 & n16954 ) ;
  assign n17677 = n17676 ^ n13936 ^ n1793 ;
  assign n17679 = n17678 ^ n17677 ^ n5263 ;
  assign n17680 = ( n1378 & n1921 ) | ( n1378 & ~n2869 ) | ( n1921 & ~n2869 ) ;
  assign n17681 = n17680 ^ n11595 ^ n6561 ;
  assign n17682 = ( ~n9747 & n12902 ) | ( ~n9747 & n17681 ) | ( n12902 & n17681 ) ;
  assign n17683 = n1891 | n2435 ;
  assign n17684 = n17683 ^ n7037 ^ n828 ;
  assign n17685 = ~n16227 & n17684 ;
  assign n17686 = n17682 & n17685 ;
  assign n17687 = ( n6084 & n7022 ) | ( n6084 & n11326 ) | ( n7022 & n11326 ) ;
  assign n17688 = n17687 ^ n15111 ^ n1517 ;
  assign n17689 = ( ~n10441 & n10525 ) | ( ~n10441 & n15082 ) | ( n10525 & n15082 ) ;
  assign n17690 = n5445 | n12722 ;
  assign n17691 = n17690 ^ n883 ^ 1'b0 ;
  assign n17692 = n17691 ^ n7346 ^ n3167 ;
  assign n17693 = n14847 ^ n13245 ^ n7680 ;
  assign n17694 = ( n2268 & n13708 ) | ( n2268 & n17693 ) | ( n13708 & n17693 ) ;
  assign n17699 = n11326 ^ n5175 ^ n4896 ;
  assign n17696 = n11046 ^ n4025 ^ 1'b0 ;
  assign n17697 = ( n5347 & n12198 ) | ( n5347 & n17696 ) | ( n12198 & n17696 ) ;
  assign n17698 = n17697 ^ n11597 ^ n10011 ;
  assign n17695 = ~n4820 & n6711 ;
  assign n17700 = n17699 ^ n17698 ^ n17695 ;
  assign n17701 = n14796 ^ n7743 ^ n4980 ;
  assign n17702 = n14213 & ~n17701 ;
  assign n17703 = n1593 & n17702 ;
  assign n17709 = n889 | n3237 ;
  assign n17710 = n17709 ^ n16115 ^ 1'b0 ;
  assign n17711 = ( n301 & ~n15304 ) | ( n301 & n17710 ) | ( ~n15304 & n17710 ) ;
  assign n17707 = n8926 | n8978 ;
  assign n17705 = ( n784 & n4159 ) | ( n784 & n15784 ) | ( n4159 & n15784 ) ;
  assign n17706 = n17705 ^ n13246 ^ 1'b0 ;
  assign n17704 = ( n506 & n6829 ) | ( n506 & ~n12590 ) | ( n6829 & ~n12590 ) ;
  assign n17708 = n17707 ^ n17706 ^ n17704 ;
  assign n17712 = n17711 ^ n17708 ^ n1176 ;
  assign n17713 = n3969 | n17712 ;
  assign n17721 = n9655 ^ n523 ^ 1'b0 ;
  assign n17722 = n5439 & n17721 ;
  assign n17723 = n17722 ^ n5920 ^ n5301 ;
  assign n17724 = n17723 ^ n7034 ^ n1286 ;
  assign n17715 = n11646 ^ n8191 ^ n7359 ;
  assign n17716 = n17715 ^ n14190 ^ 1'b0 ;
  assign n17717 = n14650 & n17716 ;
  assign n17718 = ( n2993 & n14899 ) | ( n2993 & n17717 ) | ( n14899 & n17717 ) ;
  assign n17719 = ~n13043 & n17718 ;
  assign n17720 = n17719 ^ n9918 ^ n8499 ;
  assign n17714 = n14231 ^ n6030 ^ n3371 ;
  assign n17725 = n17724 ^ n17720 ^ n17714 ;
  assign n17726 = ( n263 & ~n7624 ) | ( n263 & n9094 ) | ( ~n7624 & n9094 ) ;
  assign n17727 = n17726 ^ n9256 ^ n3373 ;
  assign n17728 = n10782 ^ n3923 ^ n2495 ;
  assign n17729 = ( ~n13206 & n17727 ) | ( ~n13206 & n17728 ) | ( n17727 & n17728 ) ;
  assign n17730 = ( ~n2355 & n3433 ) | ( ~n2355 & n6322 ) | ( n3433 & n6322 ) ;
  assign n17731 = n14276 ^ n1061 ^ x178 ;
  assign n17732 = n17731 ^ n5536 ^ n1539 ;
  assign n17733 = n17732 ^ n415 ^ x163 ;
  assign n17734 = n15145 ^ n4174 ^ n1976 ;
  assign n17735 = n17734 ^ n13064 ^ n11577 ;
  assign n17736 = n11141 & n17735 ;
  assign n17737 = ( ~n1214 & n5685 ) | ( ~n1214 & n12713 ) | ( n5685 & n12713 ) ;
  assign n17738 = n17737 ^ n14503 ^ n12716 ;
  assign n17739 = ( n5599 & ~n13051 ) | ( n5599 & n15815 ) | ( ~n13051 & n15815 ) ;
  assign n17740 = ( n4702 & n13096 ) | ( n4702 & n17739 ) | ( n13096 & n17739 ) ;
  assign n17741 = ( ~n12508 & n17738 ) | ( ~n12508 & n17740 ) | ( n17738 & n17740 ) ;
  assign n17742 = ( n1981 & ~n10280 ) | ( n1981 & n17741 ) | ( ~n10280 & n17741 ) ;
  assign n17743 = n5504 ^ n4236 ^ n899 ;
  assign n17744 = n10445 & ~n17743 ;
  assign n17745 = ( ~n1888 & n7147 ) | ( ~n1888 & n13961 ) | ( n7147 & n13961 ) ;
  assign n17746 = n14902 ^ n5790 ^ n4488 ;
  assign n17747 = ( ~n4952 & n15980 ) | ( ~n4952 & n17746 ) | ( n15980 & n17746 ) ;
  assign n17748 = ( ~n7922 & n17745 ) | ( ~n7922 & n17747 ) | ( n17745 & n17747 ) ;
  assign n17749 = n15504 ^ n8447 ^ n8041 ;
  assign n17750 = ( n1764 & ~n3650 ) | ( n1764 & n17749 ) | ( ~n3650 & n17749 ) ;
  assign n17751 = ( n2362 & ~n4602 ) | ( n2362 & n11553 ) | ( ~n4602 & n11553 ) ;
  assign n17752 = ( n5918 & ~n12809 ) | ( n5918 & n16140 ) | ( ~n12809 & n16140 ) ;
  assign n17753 = ( n2985 & ~n3074 ) | ( n2985 & n13321 ) | ( ~n3074 & n13321 ) ;
  assign n17754 = n17753 ^ n12576 ^ n11329 ;
  assign n17755 = n17754 ^ n7774 ^ n4555 ;
  assign n17756 = ( n1178 & ~n3040 ) | ( n1178 & n9138 ) | ( ~n3040 & n9138 ) ;
  assign n17757 = ( ~n452 & n3174 ) | ( ~n452 & n17756 ) | ( n3174 & n17756 ) ;
  assign n17758 = ~n468 & n2750 ;
  assign n17759 = ( n6981 & ~n16530 ) | ( n6981 & n17758 ) | ( ~n16530 & n17758 ) ;
  assign n17760 = ( n363 & n3389 ) | ( n363 & ~n10312 ) | ( n3389 & ~n10312 ) ;
  assign n17761 = ( n4061 & ~n4791 ) | ( n4061 & n17760 ) | ( ~n4791 & n17760 ) ;
  assign n17769 = n2454 & n3457 ;
  assign n17770 = n14181 & n17769 ;
  assign n17771 = ( n8678 & n10605 ) | ( n8678 & n17770 ) | ( n10605 & n17770 ) ;
  assign n17766 = n4932 & ~n8632 ;
  assign n17767 = n17766 ^ n15390 ^ 1'b0 ;
  assign n17768 = n6615 & n17767 ;
  assign n17763 = n10421 ^ n6000 ^ 1'b0 ;
  assign n17762 = ( n5635 & ~n5787 ) | ( n5635 & n16256 ) | ( ~n5787 & n16256 ) ;
  assign n17764 = n17763 ^ n17762 ^ n17644 ;
  assign n17765 = ( n758 & ~n4735 ) | ( n758 & n17764 ) | ( ~n4735 & n17764 ) ;
  assign n17772 = n17771 ^ n17768 ^ n17765 ;
  assign n17773 = n9626 & n10111 ;
  assign n17774 = ( n4686 & n5691 ) | ( n4686 & n10933 ) | ( n5691 & n10933 ) ;
  assign n17775 = ( ~n1255 & n16225 ) | ( ~n1255 & n17774 ) | ( n16225 & n17774 ) ;
  assign n17776 = ( n6169 & n7688 ) | ( n6169 & ~n17414 ) | ( n7688 & ~n17414 ) ;
  assign n17777 = ( n10291 & n11507 ) | ( n10291 & ~n17776 ) | ( n11507 & ~n17776 ) ;
  assign n17778 = n17777 ^ n11531 ^ 1'b0 ;
  assign n17780 = ( n349 & n11886 ) | ( n349 & n13096 ) | ( n11886 & n13096 ) ;
  assign n17779 = n1013 & ~n11848 ;
  assign n17781 = n17780 ^ n17779 ^ 1'b0 ;
  assign n17782 = ( n7093 & ~n13172 ) | ( n7093 & n17781 ) | ( ~n13172 & n17781 ) ;
  assign n17783 = n13881 ^ n8857 ^ n6267 ;
  assign n17784 = n17346 ^ n8953 ^ n2186 ;
  assign n17785 = ( n8099 & n8549 ) | ( n8099 & ~n17784 ) | ( n8549 & ~n17784 ) ;
  assign n17786 = ( n4404 & ~n8549 ) | ( n4404 & n17785 ) | ( ~n8549 & n17785 ) ;
  assign n17792 = n2696 | n16990 ;
  assign n17793 = n17792 ^ n10864 ^ n6108 ;
  assign n17794 = ( n4169 & n6368 ) | ( n4169 & n17793 ) | ( n6368 & n17793 ) ;
  assign n17795 = n17794 ^ n12440 ^ 1'b0 ;
  assign n17787 = n4615 | n12818 ;
  assign n17788 = ( n817 & n12609 ) | ( n817 & ~n16963 ) | ( n12609 & ~n16963 ) ;
  assign n17789 = n1609 ^ n1594 ^ n875 ;
  assign n17790 = n17789 ^ n6046 ^ 1'b0 ;
  assign n17791 = ( n17787 & n17788 ) | ( n17787 & ~n17790 ) | ( n17788 & ~n17790 ) ;
  assign n17796 = n17795 ^ n17791 ^ n10498 ;
  assign n17797 = ( n2046 & n12570 ) | ( n2046 & n13484 ) | ( n12570 & n13484 ) ;
  assign n17801 = ( n815 & ~n11613 ) | ( n815 & n12184 ) | ( ~n11613 & n12184 ) ;
  assign n17802 = n17801 ^ n11674 ^ n10083 ;
  assign n17803 = n17802 ^ n13082 ^ n1856 ;
  assign n17804 = n14649 ^ n1964 ^ 1'b0 ;
  assign n17805 = n6223 | n17804 ;
  assign n17806 = n17805 ^ n7431 ^ 1'b0 ;
  assign n17807 = n17042 | n17806 ;
  assign n17808 = n17807 ^ n5889 ^ n3386 ;
  assign n17809 = ( ~n7282 & n17803 ) | ( ~n7282 & n17808 ) | ( n17803 & n17808 ) ;
  assign n17798 = n7395 & ~n7684 ;
  assign n17799 = n17798 ^ n1256 ^ 1'b0 ;
  assign n17800 = n7640 & ~n17799 ;
  assign n17810 = n17809 ^ n17800 ^ 1'b0 ;
  assign n17811 = ( n17223 & n17797 ) | ( n17223 & ~n17810 ) | ( n17797 & ~n17810 ) ;
  assign n17812 = n16389 ^ n14104 ^ n13542 ;
  assign n17818 = n16280 ^ n7416 ^ n5150 ;
  assign n17813 = ( n429 & n4394 ) | ( n429 & n10711 ) | ( n4394 & n10711 ) ;
  assign n17814 = n8090 ^ n7527 ^ n1976 ;
  assign n17815 = n17814 ^ n3963 ^ x29 ;
  assign n17816 = ( n6208 & n12633 ) | ( n6208 & n17815 ) | ( n12633 & n17815 ) ;
  assign n17817 = ( n14367 & ~n17813 ) | ( n14367 & n17816 ) | ( ~n17813 & n17816 ) ;
  assign n17819 = n17818 ^ n17817 ^ n9020 ;
  assign n17825 = n9862 ^ n5754 ^ n3374 ;
  assign n17824 = ( n15369 & n16165 ) | ( n15369 & n16797 ) | ( n16165 & n16797 ) ;
  assign n17820 = ~n6834 & n17662 ;
  assign n17821 = ~n4018 & n17820 ;
  assign n17822 = n14313 ^ n10002 ^ n8042 ;
  assign n17823 = ( n2133 & n17821 ) | ( n2133 & n17822 ) | ( n17821 & n17822 ) ;
  assign n17826 = n17825 ^ n17824 ^ n17823 ;
  assign n17827 = ( ~n13561 & n17819 ) | ( ~n13561 & n17826 ) | ( n17819 & n17826 ) ;
  assign n17840 = n1910 ^ n1660 ^ n1242 ;
  assign n17834 = n5563 ^ n4850 ^ n922 ;
  assign n17835 = n7048 ^ n6732 ^ n3242 ;
  assign n17836 = n17835 ^ n4884 ^ 1'b0 ;
  assign n17837 = ( x120 & ~n1180 ) | ( x120 & n17836 ) | ( ~n1180 & n17836 ) ;
  assign n17838 = ( n837 & n1678 ) | ( n837 & n17837 ) | ( n1678 & n17837 ) ;
  assign n17839 = ( n13955 & n17834 ) | ( n13955 & n17838 ) | ( n17834 & n17838 ) ;
  assign n17841 = n17840 ^ n17839 ^ n14873 ;
  assign n17833 = n12374 ^ n11388 ^ n2826 ;
  assign n17830 = ( n2094 & n4967 ) | ( n2094 & ~n7117 ) | ( n4967 & ~n7117 ) ;
  assign n17828 = n16118 ^ n14354 ^ n10510 ;
  assign n17829 = n17828 ^ n13117 ^ n12781 ;
  assign n17831 = n17830 ^ n17829 ^ n7362 ;
  assign n17832 = ( n7259 & n10708 ) | ( n7259 & n17831 ) | ( n10708 & n17831 ) ;
  assign n17842 = n17841 ^ n17833 ^ n17832 ;
  assign n17843 = ( ~n9182 & n13420 ) | ( ~n9182 & n17603 ) | ( n13420 & n17603 ) ;
  assign n17848 = n3282 & ~n6625 ;
  assign n17847 = n1235 & ~n14741 ;
  assign n17849 = n17848 ^ n17847 ^ 1'b0 ;
  assign n17845 = n17305 ^ n1472 ^ n1457 ;
  assign n17846 = ( n1578 & n1986 ) | ( n1578 & ~n17845 ) | ( n1986 & ~n17845 ) ;
  assign n17844 = ( n1205 & ~n4321 ) | ( n1205 & n14763 ) | ( ~n4321 & n14763 ) ;
  assign n17850 = n17849 ^ n17846 ^ n17844 ;
  assign n17851 = ( n4088 & ~n17843 ) | ( n4088 & n17850 ) | ( ~n17843 & n17850 ) ;
  assign n17852 = n15508 ^ n5213 ^ n2731 ;
  assign n17853 = n863 | n2826 ;
  assign n17854 = ( ~n8568 & n8611 ) | ( ~n8568 & n17853 ) | ( n8611 & n17853 ) ;
  assign n17855 = n17854 ^ n3891 ^ n2506 ;
  assign n17856 = n11647 ^ n3279 ^ n3091 ;
  assign n17861 = ( n2807 & n5149 ) | ( n2807 & ~n11795 ) | ( n5149 & ~n11795 ) ;
  assign n17857 = ( n552 & ~n2256 ) | ( n552 & n2577 ) | ( ~n2256 & n2577 ) ;
  assign n17858 = ( n2060 & n3078 ) | ( n2060 & ~n4887 ) | ( n3078 & ~n4887 ) ;
  assign n17859 = n17858 ^ n4063 ^ n3369 ;
  assign n17860 = ( n1934 & ~n17857 ) | ( n1934 & n17859 ) | ( ~n17857 & n17859 ) ;
  assign n17862 = n17861 ^ n17860 ^ n17530 ;
  assign n17863 = n17862 ^ n13819 ^ n3630 ;
  assign n17864 = n13407 ^ n11320 ^ 1'b0 ;
  assign n17865 = n10126 ^ n7114 ^ n1593 ;
  assign n17866 = ( n3781 & n4073 ) | ( n3781 & n17865 ) | ( n4073 & n17865 ) ;
  assign n17867 = ( n1427 & ~n5946 ) | ( n1427 & n16659 ) | ( ~n5946 & n16659 ) ;
  assign n17868 = ( n11920 & n17866 ) | ( n11920 & ~n17867 ) | ( n17866 & ~n17867 ) ;
  assign n17869 = ( n1377 & n13697 ) | ( n1377 & n17868 ) | ( n13697 & n17868 ) ;
  assign n17870 = ( n10007 & n17864 ) | ( n10007 & n17869 ) | ( n17864 & n17869 ) ;
  assign n17874 = ~n2223 & n10477 ;
  assign n17871 = n8369 ^ n2378 ^ n1837 ;
  assign n17872 = ( n5019 & n5545 ) | ( n5019 & n17871 ) | ( n5545 & n17871 ) ;
  assign n17873 = n17872 ^ n9615 ^ n1946 ;
  assign n17875 = n17874 ^ n17873 ^ n3589 ;
  assign n17876 = ( n1947 & n5779 ) | ( n1947 & ~n17875 ) | ( n5779 & ~n17875 ) ;
  assign n17877 = ( n605 & ~n9163 ) | ( n605 & n13522 ) | ( ~n9163 & n13522 ) ;
  assign n17878 = ( n3733 & n4737 ) | ( n3733 & n17877 ) | ( n4737 & n17877 ) ;
  assign n17879 = n15088 ^ n12237 ^ n7494 ;
  assign n17882 = ( n4941 & n8429 ) | ( n4941 & ~n14940 ) | ( n8429 & ~n14940 ) ;
  assign n17880 = n4621 & n7595 ;
  assign n17881 = n693 & n17880 ;
  assign n17883 = n17882 ^ n17881 ^ n11493 ;
  assign n17884 = ( n462 & n7236 ) | ( n462 & ~n16998 ) | ( n7236 & ~n16998 ) ;
  assign n17885 = n17884 ^ n7085 ^ n6606 ;
  assign n17886 = n10316 ^ n10175 ^ n1269 ;
  assign n17888 = n3489 ^ n3405 ^ n1435 ;
  assign n17889 = n17888 ^ n13119 ^ n3560 ;
  assign n17887 = ~n15001 & n16256 ;
  assign n17890 = n17889 ^ n17887 ^ n14113 ;
  assign n17891 = n8821 | n17890 ;
  assign n17892 = n17886 | n17891 ;
  assign n17893 = n17334 ^ n4483 ^ n2089 ;
  assign n17894 = n8364 & ~n17893 ;
  assign n17895 = ( ~n2418 & n14965 ) | ( ~n2418 & n15150 ) | ( n14965 & n15150 ) ;
  assign n17896 = n17895 ^ n12281 ^ 1'b0 ;
  assign n17897 = n8676 & ~n17896 ;
  assign n17898 = ( ~n391 & n9386 ) | ( ~n391 & n17897 ) | ( n9386 & n17897 ) ;
  assign n17899 = ( ~n4463 & n16308 ) | ( ~n4463 & n16972 ) | ( n16308 & n16972 ) ;
  assign n17902 = n4170 | n6375 ;
  assign n17903 = n17902 ^ n6237 ^ 1'b0 ;
  assign n17900 = n14386 ^ n7528 ^ n2363 ;
  assign n17901 = n17900 ^ n16110 ^ n11312 ;
  assign n17904 = n17903 ^ n17901 ^ x6 ;
  assign n17905 = n13437 ^ n13240 ^ n5843 ;
  assign n17906 = ( n4448 & n8234 ) | ( n4448 & ~n14639 ) | ( n8234 & ~n14639 ) ;
  assign n17907 = n15007 ^ n13643 ^ n9089 ;
  assign n17908 = ( ~n2715 & n12146 ) | ( ~n2715 & n17907 ) | ( n12146 & n17907 ) ;
  assign n17909 = ( n4337 & n10927 ) | ( n4337 & n17441 ) | ( n10927 & n17441 ) ;
  assign n17910 = ~n11187 & n17909 ;
  assign n17913 = ( n2332 & ~n9180 ) | ( n2332 & n10096 ) | ( ~n9180 & n10096 ) ;
  assign n17911 = n17723 ^ n9213 ^ 1'b0 ;
  assign n17912 = n17911 ^ n17649 ^ n7084 ;
  assign n17914 = n17913 ^ n17912 ^ n8080 ;
  assign n17915 = n3270 & ~n14240 ;
  assign n17916 = n15980 ^ n10474 ^ n7909 ;
  assign n17917 = n17916 ^ n13617 ^ n9911 ;
  assign n17918 = ~n6160 & n17917 ;
  assign n17919 = n17918 ^ n12652 ^ 1'b0 ;
  assign n17920 = ~n10969 & n17919 ;
  assign n17921 = n17762 ^ n6001 ^ n2697 ;
  assign n17922 = ( ~x230 & n7334 ) | ( ~x230 & n12367 ) | ( n7334 & n12367 ) ;
  assign n17923 = ( n445 & n3842 ) | ( n445 & ~n6581 ) | ( n3842 & ~n6581 ) ;
  assign n17924 = ( n1720 & ~n10544 ) | ( n1720 & n17923 ) | ( ~n10544 & n17923 ) ;
  assign n17925 = n17924 ^ n15587 ^ n8146 ;
  assign n17926 = n17925 ^ n2562 ^ 1'b0 ;
  assign n17927 = n3408 & n17926 ;
  assign n17928 = ( n13771 & n17922 ) | ( n13771 & n17927 ) | ( n17922 & n17927 ) ;
  assign n17929 = ( n4852 & ~n12151 ) | ( n4852 & n13717 ) | ( ~n12151 & n13717 ) ;
  assign n17933 = n7100 ^ n2064 ^ 1'b0 ;
  assign n17934 = n17933 ^ n15069 ^ n851 ;
  assign n17930 = n2936 ^ n1377 ^ n284 ;
  assign n17931 = n17930 ^ n473 ^ x108 ;
  assign n17932 = n17931 ^ n10611 ^ n6214 ;
  assign n17935 = n17934 ^ n17932 ^ n2067 ;
  assign n17938 = n2167 & ~n4012 ;
  assign n17939 = ( n5138 & n9880 ) | ( n5138 & n17938 ) | ( n9880 & n17938 ) ;
  assign n17936 = n14613 ^ n9370 ^ 1'b0 ;
  assign n17937 = n8450 & n17936 ;
  assign n17940 = n17939 ^ n17937 ^ n14746 ;
  assign n17941 = ( ~n12855 & n13526 ) | ( ~n12855 & n17940 ) | ( n13526 & n17940 ) ;
  assign n17942 = ( n2134 & n2970 ) | ( n2134 & ~n4350 ) | ( n2970 & ~n4350 ) ;
  assign n17943 = n14869 ^ n13178 ^ n7730 ;
  assign n17944 = ( n12957 & n17942 ) | ( n12957 & n17943 ) | ( n17942 & n17943 ) ;
  assign n17945 = ( x192 & n2159 ) | ( x192 & n11307 ) | ( n2159 & n11307 ) ;
  assign n17946 = n6476 ^ n4724 ^ n256 ;
  assign n17947 = ( n1884 & ~n6217 ) | ( n1884 & n17946 ) | ( ~n6217 & n17946 ) ;
  assign n17948 = ~n10721 & n17418 ;
  assign n17949 = ( n6672 & n8653 ) | ( n6672 & ~n17948 ) | ( n8653 & ~n17948 ) ;
  assign n17950 = ( n922 & ~n17947 ) | ( n922 & n17949 ) | ( ~n17947 & n17949 ) ;
  assign n17953 = ( ~n6548 & n8994 ) | ( ~n6548 & n10474 ) | ( n8994 & n10474 ) ;
  assign n17951 = n10062 ^ n2701 ^ n2626 ;
  assign n17952 = n17951 ^ n10330 ^ n5147 ;
  assign n17954 = n17953 ^ n17952 ^ n1210 ;
  assign n17955 = ( n5343 & ~n6368 ) | ( n5343 & n17954 ) | ( ~n6368 & n17954 ) ;
  assign n17956 = n17955 ^ n14700 ^ n4779 ;
  assign n17957 = ( n6551 & n8374 ) | ( n6551 & n8904 ) | ( n8374 & n8904 ) ;
  assign n17958 = n17957 ^ n7137 ^ n5852 ;
  assign n17959 = n16332 ^ n14273 ^ n4749 ;
  assign n17960 = n10454 ^ n10431 ^ n7031 ;
  assign n17961 = n17959 & ~n17960 ;
  assign n17962 = n17961 ^ n6291 ^ 1'b0 ;
  assign n17965 = n17787 ^ n1700 ^ 1'b0 ;
  assign n17966 = n1741 & n17965 ;
  assign n17967 = ~x63 & n17966 ;
  assign n17963 = ( n313 & n946 ) | ( n313 & ~n7383 ) | ( n946 & ~n7383 ) ;
  assign n17964 = ( n6374 & n6681 ) | ( n6374 & n17963 ) | ( n6681 & n17963 ) ;
  assign n17968 = n17967 ^ n17964 ^ 1'b0 ;
  assign n17969 = ~n13964 & n17968 ;
  assign n17970 = n5833 & n11605 ;
  assign n17972 = n17683 ^ n10143 ^ n1160 ;
  assign n17971 = n290 & ~n6685 ;
  assign n17973 = n17972 ^ n17971 ^ 1'b0 ;
  assign n17974 = n17973 ^ n9547 ^ n3535 ;
  assign n17975 = n16799 ^ n12169 ^ n10473 ;
  assign n17976 = ( n8513 & n17882 ) | ( n8513 & n17975 ) | ( n17882 & n17975 ) ;
  assign n17977 = ( ~n10019 & n17974 ) | ( ~n10019 & n17976 ) | ( n17974 & n17976 ) ;
  assign n17978 = n10501 ^ n8673 ^ n6261 ;
  assign n17979 = ~n7107 & n17978 ;
  assign n17980 = n17977 & n17979 ;
  assign n17988 = n14000 ^ n4748 ^ 1'b0 ;
  assign n17989 = ~n10547 & n17988 ;
  assign n17990 = n9203 ^ n4494 ^ n2687 ;
  assign n17991 = ( n12580 & n17989 ) | ( n12580 & ~n17990 ) | ( n17989 & ~n17990 ) ;
  assign n17992 = ( n4283 & n17787 ) | ( n4283 & ~n17991 ) | ( n17787 & ~n17991 ) ;
  assign n17986 = n14848 ^ n1011 ^ x210 ;
  assign n17987 = n17986 ^ n10370 ^ n322 ;
  assign n17981 = n2396 & ~n6659 ;
  assign n17982 = n17981 ^ n10815 ^ 1'b0 ;
  assign n17983 = n8153 ^ n5775 ^ n5649 ;
  assign n17984 = ( ~n1318 & n17982 ) | ( ~n1318 & n17983 ) | ( n17982 & n17983 ) ;
  assign n17985 = ( x188 & n9295 ) | ( x188 & ~n17984 ) | ( n9295 & ~n17984 ) ;
  assign n17993 = n17992 ^ n17987 ^ n17985 ;
  assign n17994 = ( n3680 & n3972 ) | ( n3680 & ~n17289 ) | ( n3972 & ~n17289 ) ;
  assign n17995 = ( n4761 & ~n16995 ) | ( n4761 & n17994 ) | ( ~n16995 & n17994 ) ;
  assign n17999 = ( ~n1601 & n6573 ) | ( ~n1601 & n9847 ) | ( n6573 & n9847 ) ;
  assign n17996 = n12202 ^ n5072 ^ n1024 ;
  assign n17997 = ( ~n1387 & n5104 ) | ( ~n1387 & n17996 ) | ( n5104 & n17996 ) ;
  assign n17998 = n15678 | n17997 ;
  assign n18000 = n17999 ^ n17998 ^ n10169 ;
  assign n18001 = n8630 ^ n7302 ^ n1987 ;
  assign n18002 = ( n436 & ~n11050 ) | ( n436 & n18001 ) | ( ~n11050 & n18001 ) ;
  assign n18003 = n18002 ^ n9475 ^ n3073 ;
  assign n18004 = x132 & ~n18003 ;
  assign n18007 = n16289 ^ n8884 ^ n2474 ;
  assign n18006 = n2826 & n14074 ;
  assign n18008 = n18007 ^ n18006 ^ 1'b0 ;
  assign n18005 = n8744 ^ n7539 ^ n6591 ;
  assign n18009 = n18008 ^ n18005 ^ 1'b0 ;
  assign n18010 = ( n7869 & ~n10633 ) | ( n7869 & n18009 ) | ( ~n10633 & n18009 ) ;
  assign n18011 = ( n2450 & n3135 ) | ( n2450 & n12739 ) | ( n3135 & n12739 ) ;
  assign n18012 = n17767 ^ n9784 ^ n3631 ;
  assign n18013 = ( ~n2439 & n15737 ) | ( ~n2439 & n18012 ) | ( n15737 & n18012 ) ;
  assign n18014 = ( ~n3167 & n5545 ) | ( ~n3167 & n16693 ) | ( n5545 & n16693 ) ;
  assign n18015 = n7165 ^ n1672 ^ 1'b0 ;
  assign n18016 = ( ~n558 & n14161 ) | ( ~n558 & n18015 ) | ( n14161 & n18015 ) ;
  assign n18017 = n1831 | n18016 ;
  assign n18018 = n18017 ^ n7646 ^ 1'b0 ;
  assign n18019 = ( n615 & ~n11216 ) | ( n615 & n18018 ) | ( ~n11216 & n18018 ) ;
  assign n18020 = ( n8151 & n18014 ) | ( n8151 & ~n18019 ) | ( n18014 & ~n18019 ) ;
  assign n18022 = ( ~n5920 & n7786 ) | ( ~n5920 & n12097 ) | ( n7786 & n12097 ) ;
  assign n18023 = n1901 | n18022 ;
  assign n18021 = n1056 & ~n1186 ;
  assign n18024 = n18023 ^ n18021 ^ 1'b0 ;
  assign n18025 = n1062 | n3241 ;
  assign n18026 = n18025 ^ n15483 ^ n5776 ;
  assign n18027 = n18026 ^ n12285 ^ n1465 ;
  assign n18028 = ( ~n9299 & n14967 ) | ( ~n9299 & n15026 ) | ( n14967 & n15026 ) ;
  assign n18029 = ~n1647 & n4265 ;
  assign n18030 = n14741 ^ n6127 ^ 1'b0 ;
  assign n18031 = ~n13884 & n18030 ;
  assign n18032 = ( n10223 & n18029 ) | ( n10223 & ~n18031 ) | ( n18029 & ~n18031 ) ;
  assign n18033 = n9645 ^ n633 ^ n323 ;
  assign n18034 = ( n7175 & n10523 ) | ( n7175 & ~n13164 ) | ( n10523 & ~n13164 ) ;
  assign n18035 = ( n5044 & n18033 ) | ( n5044 & ~n18034 ) | ( n18033 & ~n18034 ) ;
  assign n18036 = n5540 ^ n4775 ^ n1971 ;
  assign n18037 = n14462 ^ n14003 ^ n4911 ;
  assign n18046 = n7565 ^ n6162 ^ n3958 ;
  assign n18038 = ( n3534 & n9959 ) | ( n3534 & n13943 ) | ( n9959 & n13943 ) ;
  assign n18039 = n7147 | n11089 ;
  assign n18040 = n18039 ^ n2317 ^ n2262 ;
  assign n18041 = ( x203 & ~n18038 ) | ( x203 & n18040 ) | ( ~n18038 & n18040 ) ;
  assign n18042 = ( n4103 & n9440 ) | ( n4103 & n9846 ) | ( n9440 & n9846 ) ;
  assign n18043 = ( ~n1530 & n18041 ) | ( ~n1530 & n18042 ) | ( n18041 & n18042 ) ;
  assign n18044 = ( ~n6892 & n11155 ) | ( ~n6892 & n18043 ) | ( n11155 & n18043 ) ;
  assign n18045 = n18044 ^ n16802 ^ n9677 ;
  assign n18047 = n18046 ^ n18045 ^ n1360 ;
  assign n18048 = n17373 ^ n7672 ^ n6308 ;
  assign n18049 = ( ~n2591 & n15903 ) | ( ~n2591 & n18048 ) | ( n15903 & n18048 ) ;
  assign n18050 = n7690 ^ n7451 ^ n2458 ;
  assign n18051 = n18050 ^ n17474 ^ n9918 ;
  assign n18052 = n18051 ^ n4811 ^ 1'b0 ;
  assign n18053 = n2827 & n3538 ;
  assign n18054 = ( n2829 & ~n11214 ) | ( n2829 & n18053 ) | ( ~n11214 & n18053 ) ;
  assign n18055 = n13368 & n18054 ;
  assign n18056 = ( n4472 & n18052 ) | ( n4472 & ~n18055 ) | ( n18052 & ~n18055 ) ;
  assign n18057 = ( n3316 & n4656 ) | ( n3316 & n4974 ) | ( n4656 & n4974 ) ;
  assign n18058 = n5990 ^ n1388 ^ 1'b0 ;
  assign n18059 = ( n6557 & n18057 ) | ( n6557 & n18058 ) | ( n18057 & n18058 ) ;
  assign n18060 = n18059 ^ n13883 ^ n4228 ;
  assign n18061 = n18060 ^ n916 ^ 1'b0 ;
  assign n18062 = n300 | n18061 ;
  assign n18065 = n16610 ^ n8006 ^ n4028 ;
  assign n18063 = n11510 ^ n9382 ^ n4083 ;
  assign n18064 = x157 | n18063 ;
  assign n18066 = n18065 ^ n18064 ^ n5892 ;
  assign n18067 = ( n1971 & ~n16888 ) | ( n1971 & n18066 ) | ( ~n16888 & n18066 ) ;
  assign n18068 = ( ~n551 & n9983 ) | ( ~n551 & n13434 ) | ( n9983 & n13434 ) ;
  assign n18069 = n18068 ^ n7613 ^ n1155 ;
  assign n18070 = n11252 & n18069 ;
  assign n18071 = n10803 ^ n5615 ^ n365 ;
  assign n18072 = n18071 ^ n9605 ^ n6482 ;
  assign n18073 = n12657 ^ n6005 ^ 1'b0 ;
  assign n18074 = n3006 & n18073 ;
  assign n18075 = n18074 ^ n5748 ^ 1'b0 ;
  assign n18076 = n6808 & n18075 ;
  assign n18084 = n6616 & n7325 ;
  assign n18085 = n18084 ^ n8733 ^ n752 ;
  assign n18086 = n18085 ^ n6709 ^ n2358 ;
  assign n18082 = n5774 & ~n10642 ;
  assign n18077 = n1191 ^ n1031 ^ 1'b0 ;
  assign n18078 = ( n2305 & n3173 ) | ( n2305 & n3204 ) | ( n3173 & n3204 ) ;
  assign n18079 = ( n2589 & n18077 ) | ( n2589 & ~n18078 ) | ( n18077 & ~n18078 ) ;
  assign n18080 = n18079 ^ n9597 ^ n5339 ;
  assign n18081 = n18080 ^ n17881 ^ n3505 ;
  assign n18083 = n18082 ^ n18081 ^ 1'b0 ;
  assign n18087 = n18086 ^ n18083 ^ n2910 ;
  assign n18093 = ( ~n3930 & n5481 ) | ( ~n3930 & n12536 ) | ( n5481 & n12536 ) ;
  assign n18094 = ( n2128 & n2861 ) | ( n2128 & ~n18093 ) | ( n2861 & ~n18093 ) ;
  assign n18090 = ~n5838 & n9412 ;
  assign n18091 = n6931 & n18090 ;
  assign n18088 = n11307 | n14180 ;
  assign n18089 = n10818 | n18088 ;
  assign n18092 = n18091 ^ n18089 ^ 1'b0 ;
  assign n18095 = n18094 ^ n18092 ^ n752 ;
  assign n18096 = n8829 ^ n8285 ^ n1156 ;
  assign n18097 = n3105 ^ n3091 ^ n1063 ;
  assign n18098 = n18096 & n18097 ;
  assign n18099 = ~n14941 & n18098 ;
  assign n18105 = ( n959 & n1022 ) | ( n959 & ~n1414 ) | ( n1022 & ~n1414 ) ;
  assign n18106 = n18105 ^ n7060 ^ n5957 ;
  assign n18107 = n18106 ^ n16003 ^ x213 ;
  assign n18100 = ( ~n3288 & n8788 ) | ( ~n3288 & n13223 ) | ( n8788 & n13223 ) ;
  assign n18101 = ( n6903 & ~n7154 ) | ( n6903 & n18100 ) | ( ~n7154 & n18100 ) ;
  assign n18102 = ( n3887 & n6106 ) | ( n3887 & n18101 ) | ( n6106 & n18101 ) ;
  assign n18103 = n18102 ^ n7472 ^ n319 ;
  assign n18104 = n18103 ^ n8708 ^ n5108 ;
  assign n18108 = n18107 ^ n18104 ^ n4267 ;
  assign n18109 = ( ~n4690 & n5934 ) | ( ~n4690 & n10028 ) | ( n5934 & n10028 ) ;
  assign n18110 = ( n9427 & n17474 ) | ( n9427 & ~n18109 ) | ( n17474 & ~n18109 ) ;
  assign n18117 = n5191 ^ n2878 ^ n625 ;
  assign n18111 = ( n1823 & ~n1877 ) | ( n1823 & n2438 ) | ( ~n1877 & n2438 ) ;
  assign n18112 = ( n1982 & n4316 ) | ( n1982 & n18111 ) | ( n4316 & n18111 ) ;
  assign n18113 = ( n1242 & n7618 ) | ( n1242 & ~n18112 ) | ( n7618 & ~n18112 ) ;
  assign n18114 = n7813 | n15976 ;
  assign n18115 = n6780 | n18114 ;
  assign n18116 = ( n15775 & n18113 ) | ( n15775 & n18115 ) | ( n18113 & n18115 ) ;
  assign n18118 = n18117 ^ n18116 ^ n1803 ;
  assign n18119 = ( n4733 & ~n11890 ) | ( n4733 & n18118 ) | ( ~n11890 & n18118 ) ;
  assign n18120 = ( n3298 & n18110 ) | ( n3298 & ~n18119 ) | ( n18110 & ~n18119 ) ;
  assign n18121 = n17515 ^ n10772 ^ n5435 ;
  assign n18122 = n18121 ^ n8364 ^ 1'b0 ;
  assign n18123 = ( n11521 & n13330 ) | ( n11521 & n16846 ) | ( n13330 & n16846 ) ;
  assign n18124 = ( n3710 & n7930 ) | ( n3710 & ~n18123 ) | ( n7930 & ~n18123 ) ;
  assign n18129 = n11029 ^ n6540 ^ n3732 ;
  assign n18125 = ( ~n1772 & n6544 ) | ( ~n1772 & n12881 ) | ( n6544 & n12881 ) ;
  assign n18126 = n18125 ^ n7962 ^ n7712 ;
  assign n18127 = n18126 ^ n3337 ^ n2523 ;
  assign n18128 = n15988 & ~n18127 ;
  assign n18130 = n18129 ^ n18128 ^ 1'b0 ;
  assign n18132 = n14758 ^ n6066 ^ 1'b0 ;
  assign n18131 = ( n580 & n1711 ) | ( n580 & ~n5799 ) | ( n1711 & ~n5799 ) ;
  assign n18133 = n18132 ^ n18131 ^ x156 ;
  assign n18134 = ( n7966 & n17633 ) | ( n7966 & ~n18133 ) | ( n17633 & ~n18133 ) ;
  assign n18135 = n2392 ^ n814 ^ x55 ;
  assign n18136 = n14937 ^ n1286 ^ 1'b0 ;
  assign n18137 = n813 & n8345 ;
  assign n18138 = n18137 ^ n3243 ^ 1'b0 ;
  assign n18139 = n9773 ^ n6641 ^ n3580 ;
  assign n18140 = n17996 ^ n17180 ^ n16025 ;
  assign n18141 = ( n13657 & n18139 ) | ( n13657 & n18140 ) | ( n18139 & n18140 ) ;
  assign n18142 = ( n5560 & n10277 ) | ( n5560 & n17687 ) | ( n10277 & n17687 ) ;
  assign n18143 = n18142 ^ n6614 ^ n6300 ;
  assign n18144 = ( n2217 & n11405 ) | ( n2217 & ~n14185 ) | ( n11405 & ~n14185 ) ;
  assign n18145 = n10505 & ~n11869 ;
  assign n18146 = ~n6843 & n18145 ;
  assign n18147 = ( n12497 & n18144 ) | ( n12497 & ~n18146 ) | ( n18144 & ~n18146 ) ;
  assign n18148 = ( ~n6679 & n8153 ) | ( ~n6679 & n18147 ) | ( n8153 & n18147 ) ;
  assign n18149 = ( ~n3620 & n3700 ) | ( ~n3620 & n5527 ) | ( n3700 & n5527 ) ;
  assign n18150 = n18149 ^ n10152 ^ n357 ;
  assign n18162 = n10713 ^ n6814 ^ 1'b0 ;
  assign n18158 = n14950 ^ n2750 ^ n2134 ;
  assign n18157 = ( n1985 & n3547 ) | ( n1985 & ~n9733 ) | ( n3547 & ~n9733 ) ;
  assign n18159 = n18158 ^ n18157 ^ n10706 ;
  assign n18160 = ( n11515 & n13957 ) | ( n11515 & n18159 ) | ( n13957 & n18159 ) ;
  assign n18151 = ( n1064 & n3513 ) | ( n1064 & ~n10143 ) | ( n3513 & ~n10143 ) ;
  assign n18152 = ( n2268 & ~n4260 ) | ( n2268 & n18151 ) | ( ~n4260 & n18151 ) ;
  assign n18153 = n18152 ^ n12822 ^ n11307 ;
  assign n18154 = n18153 ^ n16400 ^ n5369 ;
  assign n18155 = n18154 ^ n11800 ^ n6618 ;
  assign n18156 = n18155 ^ n8300 ^ n3878 ;
  assign n18161 = n18160 ^ n18156 ^ n13345 ;
  assign n18163 = n18162 ^ n18161 ^ n2985 ;
  assign n18164 = ( n12836 & n18150 ) | ( n12836 & ~n18163 ) | ( n18150 & ~n18163 ) ;
  assign n18165 = ( ~n2108 & n2238 ) | ( ~n2108 & n13595 ) | ( n2238 & n13595 ) ;
  assign n18166 = ( n923 & ~n1468 ) | ( n923 & n15937 ) | ( ~n1468 & n15937 ) ;
  assign n18167 = n17456 ^ n5795 ^ n5375 ;
  assign n18168 = ( n2567 & n17333 ) | ( n2567 & n18167 ) | ( n17333 & n18167 ) ;
  assign n18169 = ( n18165 & n18166 ) | ( n18165 & n18168 ) | ( n18166 & n18168 ) ;
  assign n18171 = ( n7857 & ~n7906 ) | ( n7857 & n14365 ) | ( ~n7906 & n14365 ) ;
  assign n18172 = ( n418 & ~n760 ) | ( n418 & n18171 ) | ( ~n760 & n18171 ) ;
  assign n18173 = n18172 ^ n11340 ^ n7603 ;
  assign n18170 = n278 & ~n11443 ;
  assign n18174 = n18173 ^ n18170 ^ n6893 ;
  assign n18175 = ( x206 & ~n677 ) | ( x206 & n8437 ) | ( ~n677 & n8437 ) ;
  assign n18176 = ( n4074 & n17048 ) | ( n4074 & ~n18175 ) | ( n17048 & ~n18175 ) ;
  assign n18177 = ( x43 & n11098 ) | ( x43 & ~n11794 ) | ( n11098 & ~n11794 ) ;
  assign n18178 = ( ~n6357 & n9610 ) | ( ~n6357 & n11589 ) | ( n9610 & n11589 ) ;
  assign n18179 = ( n4950 & n18177 ) | ( n4950 & ~n18178 ) | ( n18177 & ~n18178 ) ;
  assign n18180 = n16136 ^ n13178 ^ 1'b0 ;
  assign n18181 = n6835 ^ n4205 ^ n1265 ;
  assign n18182 = n13012 & ~n13898 ;
  assign n18183 = n18181 & n18182 ;
  assign n18184 = n580 | n18183 ;
  assign n18185 = n18184 ^ n6008 ^ n1113 ;
  assign n18186 = n13936 ^ n13291 ^ 1'b0 ;
  assign n18187 = n16814 & n18186 ;
  assign n18188 = n18187 ^ n10904 ^ n5229 ;
  assign n18189 = n18188 ^ n14169 ^ n3409 ;
  assign n18190 = ( ~n8292 & n8942 ) | ( ~n8292 & n15637 ) | ( n8942 & n15637 ) ;
  assign n18191 = n14683 ^ n457 ^ 1'b0 ;
  assign n18192 = n18191 ^ n11098 ^ n6818 ;
  assign n18193 = n9935 & n16654 ;
  assign n18194 = n8309 & ~n18193 ;
  assign n18195 = ( ~n2394 & n2867 ) | ( ~n2394 & n13030 ) | ( n2867 & n13030 ) ;
  assign n18197 = ( n7558 & n9754 ) | ( n7558 & n15529 ) | ( n9754 & n15529 ) ;
  assign n18198 = n18197 ^ n858 ^ 1'b0 ;
  assign n18199 = n959 & n18198 ;
  assign n18196 = ( n1500 & ~n6731 ) | ( n1500 & n11264 ) | ( ~n6731 & n11264 ) ;
  assign n18200 = n18199 ^ n18196 ^ n9948 ;
  assign n18201 = ( n9866 & n18195 ) | ( n9866 & n18200 ) | ( n18195 & n18200 ) ;
  assign n18203 = n16764 ^ n3879 ^ n716 ;
  assign n18202 = ( n2021 & n7729 ) | ( n2021 & ~n8822 ) | ( n7729 & ~n8822 ) ;
  assign n18204 = n18203 ^ n18202 ^ n16770 ;
  assign n18205 = n1688 ^ n395 ^ 1'b0 ;
  assign n18206 = ( n11906 & ~n14353 ) | ( n11906 & n15154 ) | ( ~n14353 & n15154 ) ;
  assign n18207 = ( n4454 & ~n18205 ) | ( n4454 & n18206 ) | ( ~n18205 & n18206 ) ;
  assign n18208 = ( n3514 & n4680 ) | ( n3514 & n5209 ) | ( n4680 & n5209 ) ;
  assign n18209 = n13059 ^ n3254 ^ 1'b0 ;
  assign n18210 = ~n3107 & n18209 ;
  assign n18211 = n18210 ^ n11390 ^ n2184 ;
  assign n18212 = ( ~n8732 & n12396 ) | ( ~n8732 & n18211 ) | ( n12396 & n18211 ) ;
  assign n18213 = n11272 ^ n7872 ^ n396 ;
  assign n18214 = n1340 & n1841 ;
  assign n18215 = n1584 ^ n805 ^ x159 ;
  assign n18216 = ( ~n9614 & n9870 ) | ( ~n9614 & n18215 ) | ( n9870 & n18215 ) ;
  assign n18217 = n18216 ^ n17303 ^ n10160 ;
  assign n18218 = ( n8629 & n11818 ) | ( n8629 & ~n18217 ) | ( n11818 & ~n18217 ) ;
  assign n18219 = n18218 ^ n13441 ^ n5862 ;
  assign n18220 = ( n18213 & n18214 ) | ( n18213 & ~n18219 ) | ( n18214 & ~n18219 ) ;
  assign n18225 = ~n8622 & n15969 ;
  assign n18226 = n8831 & n18225 ;
  assign n18221 = n3803 ^ n1821 ^ n459 ;
  assign n18222 = n18221 ^ n3158 ^ n814 ;
  assign n18223 = n8361 | n18222 ;
  assign n18224 = n18223 ^ n16197 ^ n6911 ;
  assign n18227 = n18226 ^ n18224 ^ n6450 ;
  assign n18229 = n12931 ^ n5348 ^ n772 ;
  assign n18228 = n7722 | n8725 ;
  assign n18230 = n18229 ^ n18228 ^ 1'b0 ;
  assign n18231 = n5321 & n15579 ;
  assign n18232 = n18230 & n18231 ;
  assign n18233 = n18232 ^ n10826 ^ n2736 ;
  assign n18234 = n767 & ~n9845 ;
  assign n18235 = ( n2346 & ~n7752 ) | ( n2346 & n17983 ) | ( ~n7752 & n17983 ) ;
  assign n18236 = ( ~n3451 & n18234 ) | ( ~n3451 & n18235 ) | ( n18234 & n18235 ) ;
  assign n18239 = n6704 ^ n4889 ^ n1965 ;
  assign n18240 = ( n4042 & ~n11035 ) | ( n4042 & n15155 ) | ( ~n11035 & n15155 ) ;
  assign n18241 = n18240 ^ n15293 ^ 1'b0 ;
  assign n18242 = n18239 & n18241 ;
  assign n18237 = n8221 ^ n1915 ^ n1471 ;
  assign n18238 = n18237 ^ n1612 ^ n1354 ;
  assign n18243 = n18242 ^ n18238 ^ n6022 ;
  assign n18244 = n12542 ^ n5754 ^ n1835 ;
  assign n18245 = ( n4510 & n5126 ) | ( n4510 & n18244 ) | ( n5126 & n18244 ) ;
  assign n18246 = n18245 ^ n8494 ^ 1'b0 ;
  assign n18247 = n1537 & n18246 ;
  assign n18248 = n1551 & n18247 ;
  assign n18249 = n5988 ^ n3975 ^ 1'b0 ;
  assign n18250 = n16197 & ~n18249 ;
  assign n18253 = ( n3487 & ~n9775 ) | ( n3487 & n13768 ) | ( ~n9775 & n13768 ) ;
  assign n18251 = ( n1009 & ~n4459 ) | ( n1009 & n8272 ) | ( ~n4459 & n8272 ) ;
  assign n18252 = n18251 ^ n9153 ^ n3466 ;
  assign n18254 = n18253 ^ n18252 ^ n3109 ;
  assign n18256 = n16504 ^ n5084 ^ 1'b0 ;
  assign n18257 = ~n2203 & n18256 ;
  assign n18255 = ( ~n3891 & n7753 ) | ( ~n3891 & n14824 ) | ( n7753 & n14824 ) ;
  assign n18258 = n18257 ^ n18255 ^ n9894 ;
  assign n18259 = ( n2411 & n6122 ) | ( n2411 & ~n12360 ) | ( n6122 & ~n12360 ) ;
  assign n18260 = n18259 ^ n5149 ^ n3610 ;
  assign n18261 = n6711 | n7264 ;
  assign n18262 = n2062 & ~n4181 ;
  assign n18263 = n8826 & n18262 ;
  assign n18264 = ( ~n18260 & n18261 ) | ( ~n18260 & n18263 ) | ( n18261 & n18263 ) ;
  assign n18265 = n13405 ^ n12384 ^ n4588 ;
  assign n18266 = n15921 ^ n2644 ^ 1'b0 ;
  assign n18267 = ( n8755 & n16869 ) | ( n8755 & n18266 ) | ( n16869 & n18266 ) ;
  assign n18268 = n18267 ^ n13513 ^ n1406 ;
  assign n18269 = n8573 | n11521 ;
  assign n18270 = n18269 ^ n660 ^ 1'b0 ;
  assign n18271 = n18270 ^ n16322 ^ n2386 ;
  assign n18275 = ( n752 & n12806 ) | ( n752 & ~n17037 ) | ( n12806 & ~n17037 ) ;
  assign n18274 = n6886 ^ n5268 ^ 1'b0 ;
  assign n18272 = n6690 ^ n3089 ^ n812 ;
  assign n18273 = n18272 ^ n6848 ^ n631 ;
  assign n18276 = n18275 ^ n18274 ^ n18273 ;
  assign n18277 = ( n10563 & n18271 ) | ( n10563 & ~n18276 ) | ( n18271 & ~n18276 ) ;
  assign n18278 = ( ~x106 & n13788 ) | ( ~x106 & n18277 ) | ( n13788 & n18277 ) ;
  assign n18279 = n16411 ^ n14732 ^ n9446 ;
  assign n18280 = n2201 | n18279 ;
  assign n18281 = ( n2949 & ~n3024 ) | ( n2949 & n16631 ) | ( ~n3024 & n16631 ) ;
  assign n18282 = ( ~x80 & n5922 ) | ( ~x80 & n18033 ) | ( n5922 & n18033 ) ;
  assign n18283 = ( n512 & ~n4416 ) | ( n512 & n7552 ) | ( ~n4416 & n7552 ) ;
  assign n18284 = ( n10218 & n18282 ) | ( n10218 & n18283 ) | ( n18282 & n18283 ) ;
  assign n18285 = ( n1289 & ~n18281 ) | ( n1289 & n18284 ) | ( ~n18281 & n18284 ) ;
  assign n18286 = ( ~n11264 & n18280 ) | ( ~n11264 & n18285 ) | ( n18280 & n18285 ) ;
  assign n18287 = ( n8783 & ~n8870 ) | ( n8783 & n18286 ) | ( ~n8870 & n18286 ) ;
  assign n18288 = n17501 ^ n9823 ^ n4517 ;
  assign n18289 = ( n10821 & n11386 ) | ( n10821 & ~n18288 ) | ( n11386 & ~n18288 ) ;
  assign n18290 = n12459 ^ n4692 ^ x52 ;
  assign n18291 = n18290 ^ n14741 ^ n8050 ;
  assign n18294 = n5495 ^ n4463 ^ n2033 ;
  assign n18295 = n18294 ^ n16003 ^ n2258 ;
  assign n18296 = ( n6537 & ~n16001 ) | ( n6537 & n18295 ) | ( ~n16001 & n18295 ) ;
  assign n18293 = ( ~n3404 & n9173 ) | ( ~n3404 & n17026 ) | ( n9173 & n17026 ) ;
  assign n18292 = n14571 ^ n7088 ^ n5303 ;
  assign n18297 = n18296 ^ n18293 ^ n18292 ;
  assign n18301 = n18259 ^ n4640 ^ n2869 ;
  assign n18298 = n7526 ^ n2078 ^ 1'b0 ;
  assign n18299 = n18298 ^ n8727 ^ n4278 ;
  assign n18300 = ( n8971 & ~n10726 ) | ( n8971 & n18299 ) | ( ~n10726 & n18299 ) ;
  assign n18302 = n18301 ^ n18300 ^ 1'b0 ;
  assign n18306 = n8557 ^ n4097 ^ n3664 ;
  assign n18307 = ( n3828 & ~n9692 ) | ( n3828 & n18306 ) | ( ~n9692 & n18306 ) ;
  assign n18304 = n14914 ^ n8081 ^ n3114 ;
  assign n18303 = ( n1994 & n8386 ) | ( n1994 & ~n14213 ) | ( n8386 & ~n14213 ) ;
  assign n18305 = n18304 ^ n18303 ^ n6828 ;
  assign n18308 = n18307 ^ n18305 ^ n10079 ;
  assign n18309 = n14787 ^ n10769 ^ n7768 ;
  assign n18310 = n14633 ^ n8216 ^ n1158 ;
  assign n18311 = ( ~n1802 & n5783 ) | ( ~n1802 & n14556 ) | ( n5783 & n14556 ) ;
  assign n18312 = ( n18309 & ~n18310 ) | ( n18309 & n18311 ) | ( ~n18310 & n18311 ) ;
  assign n18313 = ( n1115 & ~n7480 ) | ( n1115 & n7517 ) | ( ~n7480 & n7517 ) ;
  assign n18314 = n18313 ^ n17307 ^ 1'b0 ;
  assign n18315 = n6189 & n18314 ;
  assign n18316 = ( n2670 & ~n17403 ) | ( n2670 & n18315 ) | ( ~n17403 & n18315 ) ;
  assign n18317 = n15395 ^ n8808 ^ n2130 ;
  assign n18318 = ( n889 & n1816 ) | ( n889 & n18317 ) | ( n1816 & n18317 ) ;
  assign n18319 = ( n5278 & n16095 ) | ( n5278 & ~n18318 ) | ( n16095 & ~n18318 ) ;
  assign n18320 = ~n419 & n18144 ;
  assign n18321 = n14511 ^ n4429 ^ n1119 ;
  assign n18322 = n18321 ^ n16344 ^ 1'b0 ;
  assign n18323 = ( n4278 & n14422 ) | ( n4278 & ~n15647 ) | ( n14422 & ~n15647 ) ;
  assign n18328 = n13790 ^ n11506 ^ n7980 ;
  assign n18329 = n18328 ^ n10565 ^ n5527 ;
  assign n18324 = n6469 ^ n5961 ^ n3580 ;
  assign n18325 = n14320 ^ n13229 ^ n9358 ;
  assign n18326 = ( n10190 & n18324 ) | ( n10190 & n18325 ) | ( n18324 & n18325 ) ;
  assign n18327 = n9923 | n18326 ;
  assign n18330 = n18329 ^ n18327 ^ 1'b0 ;
  assign n18333 = n10605 ^ n2117 ^ n427 ;
  assign n18334 = n18333 ^ n8154 ^ n3628 ;
  assign n18331 = n1011 & n11577 ;
  assign n18332 = n2203 & n18331 ;
  assign n18335 = n18334 ^ n18332 ^ n15500 ;
  assign n18336 = n5686 ^ n5614 ^ x18 ;
  assign n18337 = ~n1257 & n18336 ;
  assign n18338 = n13276 ^ n8313 ^ n4427 ;
  assign n18339 = ( n4456 & n18337 ) | ( n4456 & ~n18338 ) | ( n18337 & ~n18338 ) ;
  assign n18340 = ( ~n3345 & n11210 ) | ( ~n3345 & n14140 ) | ( n11210 & n14140 ) ;
  assign n18342 = ( ~n862 & n14085 ) | ( ~n862 & n16335 ) | ( n14085 & n16335 ) ;
  assign n18341 = ( n1822 & ~n6819 ) | ( n1822 & n7747 ) | ( ~n6819 & n7747 ) ;
  assign n18343 = n18342 ^ n18341 ^ n4231 ;
  assign n18344 = n17138 ^ n15444 ^ n574 ;
  assign n18345 = n18344 ^ n11230 ^ n280 ;
  assign n18346 = ( n921 & n18343 ) | ( n921 & ~n18345 ) | ( n18343 & ~n18345 ) ;
  assign n18347 = n4609 ^ n2951 ^ 1'b0 ;
  assign n18348 = n18347 ^ n13970 ^ n4118 ;
  assign n18349 = n18348 ^ n4861 ^ n1955 ;
  assign n18350 = ( ~n4542 & n15134 ) | ( ~n4542 & n18349 ) | ( n15134 & n18349 ) ;
  assign n18351 = n10962 ^ n9894 ^ n9702 ;
  assign n18352 = ( x96 & n3566 ) | ( x96 & n9823 ) | ( n3566 & n9823 ) ;
  assign n18353 = ~n14602 & n18352 ;
  assign n18354 = n13743 & n18353 ;
  assign n18355 = n11496 & ~n17805 ;
  assign n18356 = n7784 ^ n3108 ^ n2776 ;
  assign n18357 = ( x35 & n11514 ) | ( x35 & n18356 ) | ( n11514 & n18356 ) ;
  assign n18364 = n12201 ^ n2318 ^ n1077 ;
  assign n18358 = ( n3159 & ~n8348 ) | ( n3159 & n9391 ) | ( ~n8348 & n9391 ) ;
  assign n18359 = ~n2751 & n4665 ;
  assign n18360 = ~n10020 & n18359 ;
  assign n18361 = n11347 ^ n3475 ^ n3127 ;
  assign n18362 = ( n14376 & ~n18360 ) | ( n14376 & n18361 ) | ( ~n18360 & n18361 ) ;
  assign n18363 = ( n5300 & n18358 ) | ( n5300 & ~n18362 ) | ( n18358 & ~n18362 ) ;
  assign n18365 = n18364 ^ n18363 ^ n17992 ;
  assign n18366 = n16192 ^ n3687 ^ n3067 ;
  assign n18367 = n6087 ^ n1284 ^ 1'b0 ;
  assign n18368 = n995 | n18367 ;
  assign n18369 = ~n8541 & n9602 ;
  assign n18370 = n18369 ^ n13319 ^ 1'b0 ;
  assign n18371 = n18370 ^ n14689 ^ n14207 ;
  assign n18372 = n7135 ^ n4987 ^ 1'b0 ;
  assign n18373 = ~n2011 & n18372 ;
  assign n18374 = ( n18368 & ~n18371 ) | ( n18368 & n18373 ) | ( ~n18371 & n18373 ) ;
  assign n18375 = x93 & n3357 ;
  assign n18376 = n18375 ^ n2895 ^ 1'b0 ;
  assign n18377 = n18376 ^ n1038 ^ 1'b0 ;
  assign n18378 = n2704 | n18377 ;
  assign n18379 = n18378 ^ n15541 ^ n7290 ;
  assign n18380 = ( ~n2035 & n7815 ) | ( ~n2035 & n11209 ) | ( n7815 & n11209 ) ;
  assign n18381 = ( n4009 & n14132 ) | ( n4009 & ~n18380 ) | ( n14132 & ~n18380 ) ;
  assign n18382 = ( n6440 & ~n17289 ) | ( n6440 & n18381 ) | ( ~n17289 & n18381 ) ;
  assign n18383 = n18382 ^ n16927 ^ n10985 ;
  assign n18384 = ( n1551 & n18260 ) | ( n1551 & ~n18383 ) | ( n18260 & ~n18383 ) ;
  assign n18386 = n11198 ^ n5515 ^ n3631 ;
  assign n18385 = n6575 & n12268 ;
  assign n18387 = n18386 ^ n18385 ^ 1'b0 ;
  assign n18388 = x186 & ~n2932 ;
  assign n18389 = n2291 & n18388 ;
  assign n18390 = n7400 ^ n6738 ^ n4685 ;
  assign n18391 = n2643 & n10752 ;
  assign n18392 = ~n18390 & n18391 ;
  assign n18393 = ( n10165 & ~n12978 ) | ( n10165 & n14861 ) | ( ~n12978 & n14861 ) ;
  assign n18394 = n10193 & n18393 ;
  assign n18395 = ( n18389 & ~n18392 ) | ( n18389 & n18394 ) | ( ~n18392 & n18394 ) ;
  assign n18396 = n1936 & n4312 ;
  assign n18397 = n18396 ^ n12863 ^ 1'b0 ;
  assign n18398 = ( ~n9507 & n14462 ) | ( ~n9507 & n18397 ) | ( n14462 & n18397 ) ;
  assign n18399 = ( ~n3964 & n14708 ) | ( ~n3964 & n17530 ) | ( n14708 & n17530 ) ;
  assign n18400 = ( n4567 & ~n6115 ) | ( n4567 & n16857 ) | ( ~n6115 & n16857 ) ;
  assign n18401 = n14955 ^ n3838 ^ n3446 ;
  assign n18405 = n4922 ^ n3879 ^ n2563 ;
  assign n18402 = ( n6071 & n13047 ) | ( n6071 & ~n17356 ) | ( n13047 & ~n17356 ) ;
  assign n18403 = n18402 ^ n1596 ^ 1'b0 ;
  assign n18404 = n4992 | n18403 ;
  assign n18406 = n18405 ^ n18404 ^ n12619 ;
  assign n18407 = ( n3966 & ~n4467 ) | ( n3966 & n18406 ) | ( ~n4467 & n18406 ) ;
  assign n18408 = n9816 ^ n4472 ^ n3720 ;
  assign n18409 = ( ~n5965 & n12108 ) | ( ~n5965 & n18408 ) | ( n12108 & n18408 ) ;
  assign n18410 = n11094 ^ n5096 ^ n3483 ;
  assign n18411 = ( n359 & n12767 ) | ( n359 & n18410 ) | ( n12767 & n18410 ) ;
  assign n18412 = ( ~n3461 & n3725 ) | ( ~n3461 & n4672 ) | ( n3725 & n4672 ) ;
  assign n18413 = ( ~n866 & n2739 ) | ( ~n866 & n18412 ) | ( n2739 & n18412 ) ;
  assign n18414 = ( n856 & n1558 ) | ( n856 & ~n18413 ) | ( n1558 & ~n18413 ) ;
  assign n18415 = ( ~n15952 & n18411 ) | ( ~n15952 & n18414 ) | ( n18411 & n18414 ) ;
  assign n18416 = n18415 ^ n3567 ^ 1'b0 ;
  assign n18417 = n18409 & n18416 ;
  assign n18418 = n13204 ^ n888 ^ x73 ;
  assign n18419 = n18418 ^ n1064 ^ 1'b0 ;
  assign n18420 = n6878 & ~n18419 ;
  assign n18421 = n18420 ^ n9607 ^ 1'b0 ;
  assign n18422 = n8353 ^ n7487 ^ n3924 ;
  assign n18423 = ( n13586 & n14233 ) | ( n13586 & n18422 ) | ( n14233 & n18422 ) ;
  assign n18424 = n15003 ^ n4564 ^ n273 ;
  assign n18425 = ~n4799 & n17802 ;
  assign n18426 = n18425 ^ n12427 ^ 1'b0 ;
  assign n18427 = n17135 ^ n4783 ^ 1'b0 ;
  assign n18428 = n18427 ^ n14401 ^ n5591 ;
  assign n18429 = n17821 ^ n11389 ^ n8238 ;
  assign n18430 = n18429 ^ n15307 ^ n3147 ;
  assign n18433 = ( ~x138 & n4504 ) | ( ~x138 & n15119 ) | ( n4504 & n15119 ) ;
  assign n18434 = n18433 ^ n7454 ^ n6574 ;
  assign n18431 = n8067 ^ n917 ^ 1'b0 ;
  assign n18432 = n2686 | n18431 ;
  assign n18435 = n18434 ^ n18432 ^ n4796 ;
  assign n18436 = n18435 ^ n5514 ^ 1'b0 ;
  assign n18437 = n18436 ^ n11370 ^ n9738 ;
  assign n18438 = n18437 ^ n6929 ^ n6621 ;
  assign n18439 = ~n18430 & n18438 ;
  assign n18440 = ( n1937 & ~n16529 ) | ( n1937 & n18439 ) | ( ~n16529 & n18439 ) ;
  assign n18441 = ( n1313 & n13175 ) | ( n1313 & ~n18181 ) | ( n13175 & ~n18181 ) ;
  assign n18444 = ( x120 & n6386 ) | ( x120 & n7499 ) | ( n6386 & n7499 ) ;
  assign n18442 = ( n5035 & ~n12898 ) | ( n5035 & n16141 ) | ( ~n12898 & n16141 ) ;
  assign n18443 = ~n17276 & n18442 ;
  assign n18445 = n18444 ^ n18443 ^ 1'b0 ;
  assign n18446 = ( ~n18229 & n18441 ) | ( ~n18229 & n18445 ) | ( n18441 & n18445 ) ;
  assign n18447 = n8976 & n13602 ;
  assign n18448 = ~n12984 & n18447 ;
  assign n18449 = n18448 ^ n17676 ^ n15830 ;
  assign n18450 = n4514 ^ n2870 ^ n453 ;
  assign n18451 = ( n2273 & n9550 ) | ( n2273 & n18450 ) | ( n9550 & n18450 ) ;
  assign n18452 = ( ~n600 & n1704 ) | ( ~n600 & n18451 ) | ( n1704 & n18451 ) ;
  assign n18453 = n1893 & n3006 ;
  assign n18454 = n11054 & n18453 ;
  assign n18455 = n6791 ^ n3217 ^ x101 ;
  assign n18456 = ( n5103 & ~n16468 ) | ( n5103 & n18455 ) | ( ~n16468 & n18455 ) ;
  assign n18457 = ( n6049 & ~n18454 ) | ( n6049 & n18456 ) | ( ~n18454 & n18456 ) ;
  assign n18458 = n18457 ^ n18127 ^ 1'b0 ;
  assign n18460 = n2251 ^ n1333 ^ n658 ;
  assign n18461 = ( n3734 & n8279 ) | ( n3734 & n18460 ) | ( n8279 & n18460 ) ;
  assign n18462 = ( n2938 & n4792 ) | ( n2938 & ~n10957 ) | ( n4792 & ~n10957 ) ;
  assign n18463 = ( n2678 & n18461 ) | ( n2678 & ~n18462 ) | ( n18461 & ~n18462 ) ;
  assign n18464 = n588 & n18463 ;
  assign n18459 = n5106 | n15980 ;
  assign n18465 = n18464 ^ n18459 ^ 1'b0 ;
  assign n18468 = ( n4265 & ~n11066 ) | ( n4265 & n15587 ) | ( ~n11066 & n15587 ) ;
  assign n18469 = n18468 ^ n10428 ^ n3594 ;
  assign n18466 = n13222 ^ n8435 ^ 1'b0 ;
  assign n18467 = n18466 ^ n1803 ^ n1410 ;
  assign n18470 = n18469 ^ n18467 ^ n4650 ;
  assign n18474 = n6461 ^ n1980 ^ n1565 ;
  assign n18471 = n10907 ^ n5277 ^ n1797 ;
  assign n18472 = ( n4036 & ~n9624 ) | ( n4036 & n18471 ) | ( ~n9624 & n18471 ) ;
  assign n18473 = n18472 ^ n14322 ^ n7997 ;
  assign n18475 = n18474 ^ n18473 ^ n3942 ;
  assign n18476 = ( n1673 & n2920 ) | ( n1673 & ~n18475 ) | ( n2920 & ~n18475 ) ;
  assign n18477 = n14202 | n16751 ;
  assign n18480 = n5180 | n12680 ;
  assign n18478 = n5565 ^ n5438 ^ 1'b0 ;
  assign n18479 = n10659 & n18478 ;
  assign n18481 = n18480 ^ n18479 ^ n9565 ;
  assign n18482 = n2724 & ~n6625 ;
  assign n18483 = ~x87 & n18482 ;
  assign n18484 = ( n14224 & n15346 ) | ( n14224 & ~n18483 ) | ( n15346 & ~n18483 ) ;
  assign n18487 = n13669 ^ n12632 ^ n6662 ;
  assign n18486 = n13388 ^ n8293 ^ 1'b0 ;
  assign n18485 = ( n334 & n11891 ) | ( n334 & n12122 ) | ( n11891 & n12122 ) ;
  assign n18488 = n18487 ^ n18486 ^ n18485 ;
  assign n18489 = ( n9048 & n13236 ) | ( n9048 & ~n18488 ) | ( n13236 & ~n18488 ) ;
  assign n18492 = ( n2256 & ~n8239 ) | ( n2256 & n12120 ) | ( ~n8239 & n12120 ) ;
  assign n18493 = n18492 ^ n18126 ^ n346 ;
  assign n18494 = ( n2390 & n7389 ) | ( n2390 & n18493 ) | ( n7389 & n18493 ) ;
  assign n18490 = n12403 ^ n10134 ^ n9615 ;
  assign n18491 = ( n5234 & n10790 ) | ( n5234 & ~n18490 ) | ( n10790 & ~n18490 ) ;
  assign n18495 = n18494 ^ n18491 ^ n5184 ;
  assign n18496 = n18489 & ~n18495 ;
  assign n18497 = ~n903 & n18496 ;
  assign n18498 = n13428 ^ n7018 ^ n418 ;
  assign n18499 = n18498 ^ n2252 ^ n1142 ;
  assign n18500 = ( n2679 & n10589 ) | ( n2679 & ~n18405 ) | ( n10589 & ~n18405 ) ;
  assign n18501 = ( n1165 & n15436 ) | ( n1165 & ~n17420 ) | ( n15436 & ~n17420 ) ;
  assign n18502 = n18501 ^ n2225 ^ n1774 ;
  assign n18503 = ( n633 & n18500 ) | ( n633 & ~n18502 ) | ( n18500 & ~n18502 ) ;
  assign n18504 = n2126 & ~n18088 ;
  assign n18505 = ( n1905 & ~n10688 ) | ( n1905 & n18504 ) | ( ~n10688 & n18504 ) ;
  assign n18506 = ( n1334 & ~n15649 ) | ( n1334 & n17837 ) | ( ~n15649 & n17837 ) ;
  assign n18507 = ( n5908 & n11125 ) | ( n5908 & ~n18506 ) | ( n11125 & ~n18506 ) ;
  assign n18508 = ( n18503 & n18505 ) | ( n18503 & n18507 ) | ( n18505 & n18507 ) ;
  assign n18512 = n14633 ^ n5134 ^ n2544 ;
  assign n18510 = ( ~n935 & n6383 ) | ( ~n935 & n11382 ) | ( n6383 & n11382 ) ;
  assign n18509 = n4784 | n7218 ;
  assign n18511 = n18510 ^ n18509 ^ n13302 ;
  assign n18513 = n18512 ^ n18511 ^ n11201 ;
  assign n18514 = n14316 ^ n7749 ^ n4312 ;
  assign n18515 = n18514 ^ n10971 ^ n3127 ;
  assign n18522 = n1862 | n2968 ;
  assign n18516 = ( n1175 & n3963 ) | ( n1175 & ~n7790 ) | ( n3963 & ~n7790 ) ;
  assign n18517 = n18516 ^ n8839 ^ n8672 ;
  assign n18519 = ( n8396 & n9083 ) | ( n8396 & ~n17090 ) | ( n9083 & ~n17090 ) ;
  assign n18518 = ( ~n9053 & n10596 ) | ( ~n9053 & n10738 ) | ( n10596 & n10738 ) ;
  assign n18520 = n18519 ^ n18518 ^ n4804 ;
  assign n18521 = ( n13373 & n18517 ) | ( n13373 & ~n18520 ) | ( n18517 & ~n18520 ) ;
  assign n18523 = n18522 ^ n18521 ^ 1'b0 ;
  assign n18524 = n1609 & ~n18523 ;
  assign n18525 = n14501 ^ n7680 ^ n7083 ;
  assign n18539 = ( n8755 & ~n12164 ) | ( n8755 & n15965 ) | ( ~n12164 & n15965 ) ;
  assign n18531 = ( n1326 & n2902 ) | ( n1326 & ~n3333 ) | ( n2902 & ~n3333 ) ;
  assign n18528 = n2012 | n7545 ;
  assign n18529 = n1380 | n18528 ;
  assign n18530 = ( n7264 & n12519 ) | ( n7264 & n18529 ) | ( n12519 & n18529 ) ;
  assign n18532 = n18531 ^ n18530 ^ n13422 ;
  assign n18526 = n1904 ^ n746 ^ n711 ;
  assign n18527 = ( n5085 & ~n11648 ) | ( n5085 & n18526 ) | ( ~n11648 & n18526 ) ;
  assign n18533 = n18532 ^ n18527 ^ n9800 ;
  assign n18534 = n17946 ^ n16341 ^ n9655 ;
  assign n18535 = ( n1208 & n17762 ) | ( n1208 & ~n18534 ) | ( n17762 & ~n18534 ) ;
  assign n18536 = n3453 ^ n2652 ^ 1'b0 ;
  assign n18537 = ( n9131 & n18535 ) | ( n9131 & ~n18536 ) | ( n18535 & ~n18536 ) ;
  assign n18538 = ( ~n8058 & n18533 ) | ( ~n8058 & n18537 ) | ( n18533 & n18537 ) ;
  assign n18540 = n18539 ^ n18538 ^ n9747 ;
  assign n18541 = ( n10407 & n18525 ) | ( n10407 & n18540 ) | ( n18525 & n18540 ) ;
  assign n18542 = n13505 ^ n10973 ^ n7253 ;
  assign n18543 = n18542 ^ n15846 ^ n2784 ;
  assign n18544 = ( ~n18524 & n18541 ) | ( ~n18524 & n18543 ) | ( n18541 & n18543 ) ;
  assign n18549 = ( ~n2544 & n5066 ) | ( ~n2544 & n13478 ) | ( n5066 & n13478 ) ;
  assign n18550 = n18549 ^ n2150 ^ n501 ;
  assign n18547 = n2864 ^ n1767 ^ n1305 ;
  assign n18545 = x201 & ~n3772 ;
  assign n18546 = n18545 ^ n1739 ^ 1'b0 ;
  assign n18548 = n18547 ^ n18546 ^ n6762 ;
  assign n18551 = n18550 ^ n18548 ^ n11948 ;
  assign n18552 = n7047 ^ n6356 ^ 1'b0 ;
  assign n18553 = n18179 & ~n18552 ;
  assign n18554 = ~n16190 & n18553 ;
  assign n18555 = n18203 ^ n18007 ^ n6567 ;
  assign n18556 = n15101 ^ n12473 ^ n10682 ;
  assign n18557 = n9892 ^ n2978 ^ 1'b0 ;
  assign n18558 = ( x133 & n272 ) | ( x133 & ~n7873 ) | ( n272 & ~n7873 ) ;
  assign n18559 = ( n17840 & n18557 ) | ( n17840 & n18558 ) | ( n18557 & n18558 ) ;
  assign n18560 = n15589 ^ n10119 ^ 1'b0 ;
  assign n18561 = ~n1323 & n18560 ;
  assign n18562 = ( n5188 & ~n16824 ) | ( n5188 & n18561 ) | ( ~n16824 & n18561 ) ;
  assign n18563 = n12429 ^ n5472 ^ n5263 ;
  assign n18564 = ( x170 & ~n829 ) | ( x170 & n17095 ) | ( ~n829 & n17095 ) ;
  assign n18565 = ( n2884 & ~n18563 ) | ( n2884 & n18564 ) | ( ~n18563 & n18564 ) ;
  assign n18566 = n18565 ^ n16105 ^ n13568 ;
  assign n18567 = ( n667 & n18562 ) | ( n667 & ~n18566 ) | ( n18562 & ~n18566 ) ;
  assign n18568 = x55 & n18197 ;
  assign n18572 = n14074 ^ n7221 ^ n2612 ;
  assign n18569 = n12079 ^ n10444 ^ n2865 ;
  assign n18570 = n18569 ^ n8307 ^ n4629 ;
  assign n18571 = n18570 ^ n15128 ^ n5523 ;
  assign n18573 = n18572 ^ n18571 ^ n2249 ;
  assign n18578 = n9449 ^ n7426 ^ n5064 ;
  assign n18574 = ( n2036 & n6808 ) | ( n2036 & n7060 ) | ( n6808 & n7060 ) ;
  assign n18575 = n16251 ^ n11303 ^ n2658 ;
  assign n18576 = n18575 ^ n17122 ^ n12199 ;
  assign n18577 = ( n14032 & n18574 ) | ( n14032 & ~n18576 ) | ( n18574 & ~n18576 ) ;
  assign n18579 = n18578 ^ n18577 ^ n9778 ;
  assign n18580 = n17887 ^ n11215 ^ n3356 ;
  assign n18585 = ( n2225 & ~n5660 ) | ( n2225 & n10964 ) | ( ~n5660 & n10964 ) ;
  assign n18583 = ( n6672 & n9131 ) | ( n6672 & ~n17501 ) | ( n9131 & ~n17501 ) ;
  assign n18581 = n11282 ^ x13 ^ 1'b0 ;
  assign n18582 = n18581 ^ n17524 ^ n8939 ;
  assign n18584 = n18583 ^ n18582 ^ n6702 ;
  assign n18586 = n18585 ^ n18584 ^ n3367 ;
  assign n18587 = n14584 ^ n8979 ^ n7383 ;
  assign n18591 = n15413 ^ n9776 ^ n3690 ;
  assign n18592 = ( x49 & ~x196 ) | ( x49 & n18591 ) | ( ~x196 & n18591 ) ;
  assign n18593 = ( n8966 & ~n13792 ) | ( n8966 & n18592 ) | ( ~n13792 & n18592 ) ;
  assign n18588 = n4549 & n15478 ;
  assign n18589 = ( n363 & n5867 ) | ( n363 & ~n9584 ) | ( n5867 & ~n9584 ) ;
  assign n18590 = ( n12682 & ~n18588 ) | ( n12682 & n18589 ) | ( ~n18588 & n18589 ) ;
  assign n18594 = n18593 ^ n18590 ^ x74 ;
  assign n18595 = ( ~n6080 & n18587 ) | ( ~n6080 & n18594 ) | ( n18587 & n18594 ) ;
  assign n18596 = ( ~n18580 & n18586 ) | ( ~n18580 & n18595 ) | ( n18586 & n18595 ) ;
  assign n18597 = ( ~n406 & n2239 ) | ( ~n406 & n14410 ) | ( n2239 & n14410 ) ;
  assign n18598 = ( n1991 & ~n6759 ) | ( n1991 & n18597 ) | ( ~n6759 & n18597 ) ;
  assign n18599 = n18598 ^ n7576 ^ 1'b0 ;
  assign n18600 = n15911 ^ n15659 ^ n6513 ;
  assign n18608 = ( n774 & n9805 ) | ( n774 & ~n12881 ) | ( n9805 & ~n12881 ) ;
  assign n18609 = ( ~x244 & n6819 ) | ( ~x244 & n18608 ) | ( n6819 & n18608 ) ;
  assign n18610 = n17602 & ~n18609 ;
  assign n18601 = n13987 ^ n7021 ^ n4095 ;
  assign n18602 = ( n10672 & n10979 ) | ( n10672 & ~n16565 ) | ( n10979 & ~n16565 ) ;
  assign n18603 = ( n2325 & n6454 ) | ( n2325 & n17818 ) | ( n6454 & n17818 ) ;
  assign n18604 = n18603 ^ n11663 ^ n5680 ;
  assign n18605 = ~n18602 & n18604 ;
  assign n18606 = n18605 ^ n8822 ^ 1'b0 ;
  assign n18607 = n18601 & n18606 ;
  assign n18611 = n18610 ^ n18607 ^ 1'b0 ;
  assign n18612 = ( n4886 & n12336 ) | ( n4886 & ~n16969 ) | ( n12336 & ~n16969 ) ;
  assign n18613 = ( ~n16255 & n16785 ) | ( ~n16255 & n18612 ) | ( n16785 & n18612 ) ;
  assign n18614 = n7694 ^ n7015 ^ n3995 ;
  assign n18615 = ( n3652 & n8618 ) | ( n3652 & n18614 ) | ( n8618 & n18614 ) ;
  assign n18616 = ( n4029 & ~n10599 ) | ( n4029 & n15269 ) | ( ~n10599 & n15269 ) ;
  assign n18617 = ( n13719 & n14467 ) | ( n13719 & n18616 ) | ( n14467 & n18616 ) ;
  assign n18621 = n16056 ^ n12849 ^ n6173 ;
  assign n18619 = n11497 ^ n4109 ^ n1606 ;
  assign n18618 = ~n875 & n2817 ;
  assign n18620 = n18619 ^ n18618 ^ n6264 ;
  assign n18622 = n18621 ^ n18620 ^ n3983 ;
  assign n18623 = n15494 ^ n13731 ^ n2485 ;
  assign n18624 = n11936 ^ n8434 ^ n979 ;
  assign n18625 = n16783 ^ n7102 ^ n451 ;
  assign n18626 = n18581 ^ n16842 ^ n16746 ;
  assign n18627 = n18626 ^ n11215 ^ 1'b0 ;
  assign n18628 = n18625 | n18627 ;
  assign n18629 = n14074 ^ n4586 ^ n3852 ;
  assign n18630 = ( ~n18624 & n18628 ) | ( ~n18624 & n18629 ) | ( n18628 & n18629 ) ;
  assign n18631 = n17837 ^ n8512 ^ n7094 ;
  assign n18637 = n13140 ^ n3948 ^ 1'b0 ;
  assign n18636 = n11395 ^ n7635 ^ n4019 ;
  assign n18634 = ~n4776 & n10774 ;
  assign n18632 = ( n3690 & n4214 ) | ( n3690 & n6481 ) | ( n4214 & n6481 ) ;
  assign n18633 = n13347 | n18632 ;
  assign n18635 = n18634 ^ n18633 ^ n12895 ;
  assign n18638 = n18637 ^ n18636 ^ n18635 ;
  assign n18639 = n11873 ^ n2536 ^ n641 ;
  assign n18643 = n16428 ^ n10667 ^ n2706 ;
  assign n18640 = ( x91 & ~n1534 ) | ( x91 & n3367 ) | ( ~n1534 & n3367 ) ;
  assign n18641 = n17947 ^ n3022 ^ 1'b0 ;
  assign n18642 = ( n13481 & n18640 ) | ( n13481 & ~n18641 ) | ( n18640 & ~n18641 ) ;
  assign n18644 = n18643 ^ n18642 ^ n11912 ;
  assign n18648 = n11924 ^ n5164 ^ n3576 ;
  assign n18645 = ( n599 & n1217 ) | ( n599 & ~n4096 ) | ( n1217 & ~n4096 ) ;
  assign n18646 = ( n10988 & ~n15884 ) | ( n10988 & n18645 ) | ( ~n15884 & n18645 ) ;
  assign n18647 = ( n5178 & n18516 ) | ( n5178 & n18646 ) | ( n18516 & n18646 ) ;
  assign n18649 = n18648 ^ n18647 ^ n8531 ;
  assign n18650 = n4284 & ~n4714 ;
  assign n18651 = n18650 ^ n14751 ^ 1'b0 ;
  assign n18652 = n18651 ^ n16797 ^ n10230 ;
  assign n18653 = ( n981 & n4501 ) | ( n981 & ~n5225 ) | ( n4501 & ~n5225 ) ;
  assign n18654 = ( n4036 & n8227 ) | ( n4036 & ~n18653 ) | ( n8227 & ~n18653 ) ;
  assign n18655 = n18654 ^ n6536 ^ 1'b0 ;
  assign n18656 = n3390 & n5766 ;
  assign n18657 = ( ~n15385 & n16876 ) | ( ~n15385 & n18656 ) | ( n16876 & n18656 ) ;
  assign n18658 = n12398 ^ n10857 ^ n3446 ;
  assign n18659 = n4309 | n5654 ;
  assign n18660 = n18659 ^ n3098 ^ 1'b0 ;
  assign n18661 = ( ~n11327 & n18658 ) | ( ~n11327 & n18660 ) | ( n18658 & n18660 ) ;
  assign n18662 = n1663 & ~n14600 ;
  assign n18663 = n18662 ^ n13974 ^ n4358 ;
  assign n18664 = n18663 ^ n10516 ^ n3829 ;
  assign n18665 = n2646 ^ n991 ^ n567 ;
  assign n18666 = n18665 ^ n6200 ^ 1'b0 ;
  assign n18667 = ~n10853 & n18666 ;
  assign n18668 = ~n1939 & n18667 ;
  assign n18669 = ~n13474 & n18668 ;
  assign n18671 = n2015 & n11826 ;
  assign n18670 = ( n4787 & ~n5648 ) | ( n4787 & n8700 ) | ( ~n5648 & n8700 ) ;
  assign n18672 = n18671 ^ n18670 ^ n8912 ;
  assign n18677 = ( n7202 & ~n12698 ) | ( n7202 & n13288 ) | ( ~n12698 & n13288 ) ;
  assign n18678 = x69 & ~n12323 ;
  assign n18679 = n18678 ^ n3105 ^ 1'b0 ;
  assign n18680 = n18679 ^ n17581 ^ n6365 ;
  assign n18681 = ( n4843 & n18677 ) | ( n4843 & n18680 ) | ( n18677 & n18680 ) ;
  assign n18673 = n14769 ^ n1695 ^ 1'b0 ;
  assign n18674 = n18673 ^ n13342 ^ n5007 ;
  assign n18675 = n18040 ^ n16142 ^ n7988 ;
  assign n18676 = ( n14967 & n18674 ) | ( n14967 & n18675 ) | ( n18674 & n18675 ) ;
  assign n18682 = n18681 ^ n18676 ^ n5988 ;
  assign n18683 = ( n2114 & n5453 ) | ( n2114 & ~n13085 ) | ( n5453 & ~n13085 ) ;
  assign n18684 = n18683 ^ n13292 ^ n6258 ;
  assign n18685 = ( n18672 & n18682 ) | ( n18672 & n18684 ) | ( n18682 & n18684 ) ;
  assign n18692 = ( n3494 & n3832 ) | ( n3494 & n7352 ) | ( n3832 & n7352 ) ;
  assign n18690 = n10396 ^ n4445 ^ n2565 ;
  assign n18689 = ( ~n3154 & n6081 ) | ( ~n3154 & n9900 ) | ( n6081 & n9900 ) ;
  assign n18687 = ( n4447 & n5556 ) | ( n4447 & ~n12170 ) | ( n5556 & ~n12170 ) ;
  assign n18688 = n18687 ^ n9022 ^ n8272 ;
  assign n18691 = n18690 ^ n18689 ^ n18688 ;
  assign n18693 = n18692 ^ n18691 ^ n3597 ;
  assign n18686 = ( n1200 & ~n4587 ) | ( n1200 & n17897 ) | ( ~n4587 & n17897 ) ;
  assign n18694 = n18693 ^ n18686 ^ n9797 ;
  assign n18695 = ( n6638 & n8072 ) | ( n6638 & ~n16504 ) | ( n8072 & ~n16504 ) ;
  assign n18696 = ( ~n1567 & n11613 ) | ( ~n1567 & n18695 ) | ( n11613 & n18695 ) ;
  assign n18697 = n18696 ^ n10819 ^ n5832 ;
  assign n18698 = ( n3781 & n8403 ) | ( n3781 & ~n9996 ) | ( n8403 & ~n9996 ) ;
  assign n18699 = ( n4782 & n6996 ) | ( n4782 & n18077 ) | ( n6996 & n18077 ) ;
  assign n18700 = ( n1586 & n3986 ) | ( n1586 & n9841 ) | ( n3986 & n9841 ) ;
  assign n18701 = n17108 ^ n16270 ^ n15630 ;
  assign n18702 = ( n12564 & n15894 ) | ( n12564 & ~n18701 ) | ( n15894 & ~n18701 ) ;
  assign n18703 = n18702 ^ n5894 ^ n5631 ;
  assign n18704 = ( n18102 & n18700 ) | ( n18102 & ~n18703 ) | ( n18700 & ~n18703 ) ;
  assign n18705 = ( n741 & n10744 ) | ( n741 & n16489 ) | ( n10744 & n16489 ) ;
  assign n18707 = ( ~n8383 & n10050 ) | ( ~n8383 & n17887 ) | ( n10050 & n17887 ) ;
  assign n18706 = ( ~n3118 & n7675 ) | ( ~n3118 & n17571 ) | ( n7675 & n17571 ) ;
  assign n18708 = n18707 ^ n18706 ^ n3871 ;
  assign n18709 = n16522 ^ n7613 ^ n4515 ;
  assign n18710 = n18709 ^ n3979 ^ 1'b0 ;
  assign n18711 = n8350 ^ n6543 ^ n5071 ;
  assign n18712 = n18711 ^ n6203 ^ 1'b0 ;
  assign n18715 = n10378 ^ n9891 ^ n4294 ;
  assign n18713 = ( n3908 & n7537 ) | ( n3908 & ~n18591 ) | ( n7537 & ~n18591 ) ;
  assign n18714 = ( n9860 & ~n13841 ) | ( n9860 & n18713 ) | ( ~n13841 & n18713 ) ;
  assign n18716 = n18715 ^ n18714 ^ n14891 ;
  assign n18730 = n10647 ^ n5900 ^ n291 ;
  assign n18726 = ( n606 & n3667 ) | ( n606 & ~n9483 ) | ( n3667 & ~n9483 ) ;
  assign n18727 = ( n8020 & ~n13511 ) | ( n8020 & n15444 ) | ( ~n13511 & n15444 ) ;
  assign n18728 = n13711 & ~n18727 ;
  assign n18729 = n18726 & n18728 ;
  assign n18717 = n9406 ^ n3890 ^ 1'b0 ;
  assign n18718 = n5714 & n9336 ;
  assign n18719 = n18718 ^ n11571 ^ 1'b0 ;
  assign n18720 = n18719 ^ n3508 ^ 1'b0 ;
  assign n18721 = n18717 | n18720 ;
  assign n18722 = ( n2849 & n2952 ) | ( n2849 & n18721 ) | ( n2952 & n18721 ) ;
  assign n18723 = ( n3378 & ~n3902 ) | ( n3378 & n18722 ) | ( ~n3902 & n18722 ) ;
  assign n18724 = n18723 ^ n14384 ^ n13568 ;
  assign n18725 = ( n4243 & n12595 ) | ( n4243 & ~n18724 ) | ( n12595 & ~n18724 ) ;
  assign n18731 = n18730 ^ n18729 ^ n18725 ;
  assign n18732 = n7655 ^ n5669 ^ 1'b0 ;
  assign n18733 = ( n384 & n5876 ) | ( n384 & ~n18732 ) | ( n5876 & ~n18732 ) ;
  assign n18734 = ( ~n1800 & n3517 ) | ( ~n1800 & n6451 ) | ( n3517 & n6451 ) ;
  assign n18735 = n18734 ^ n12896 ^ n11076 ;
  assign n18736 = ( n18005 & n18733 ) | ( n18005 & n18735 ) | ( n18733 & n18735 ) ;
  assign n18737 = n8115 & n8394 ;
  assign n18738 = n18737 ^ n4823 ^ 1'b0 ;
  assign n18739 = n15870 ^ n734 ^ n615 ;
  assign n18740 = ( n548 & n18738 ) | ( n548 & n18739 ) | ( n18738 & n18739 ) ;
  assign n18741 = n9953 ^ n6045 ^ 1'b0 ;
  assign n18742 = ( n4791 & ~n17053 ) | ( n4791 & n18714 ) | ( ~n17053 & n18714 ) ;
  assign n18743 = n16129 ^ n4896 ^ 1'b0 ;
  assign n18744 = n3454 | n18743 ;
  assign n18745 = n12473 ^ n10192 ^ n2019 ;
  assign n18746 = ( n9605 & n18744 ) | ( n9605 & ~n18745 ) | ( n18744 & ~n18745 ) ;
  assign n18747 = ( ~n16710 & n18742 ) | ( ~n16710 & n18746 ) | ( n18742 & n18746 ) ;
  assign n18748 = ( n18740 & n18741 ) | ( n18740 & ~n18747 ) | ( n18741 & ~n18747 ) ;
  assign n18751 = n2165 | n14787 ;
  assign n18752 = n8739 & ~n18751 ;
  assign n18753 = n18752 ^ n10667 ^ n6885 ;
  assign n18749 = n10708 ^ n5503 ^ n4215 ;
  assign n18750 = n18749 ^ n5608 ^ n866 ;
  assign n18754 = n18753 ^ n18750 ^ n14332 ;
  assign n18755 = ( ~n2122 & n6997 ) | ( ~n2122 & n7931 ) | ( n6997 & n7931 ) ;
  assign n18756 = n513 & ~n8239 ;
  assign n18757 = n18755 & n18756 ;
  assign n18758 = ( n4103 & n13340 ) | ( n4103 & ~n16320 ) | ( n13340 & ~n16320 ) ;
  assign n18759 = n18758 ^ n16894 ^ n4016 ;
  assign n18760 = n12518 ^ n3849 ^ 1'b0 ;
  assign n18761 = ( ~n5132 & n15769 ) | ( ~n5132 & n18760 ) | ( n15769 & n18760 ) ;
  assign n18762 = n17237 ^ n15603 ^ n1856 ;
  assign n18763 = n10922 ^ n6198 ^ 1'b0 ;
  assign n18764 = n17108 ^ n4640 ^ n1048 ;
  assign n18765 = x35 & ~n18764 ;
  assign n18768 = n4661 ^ n3939 ^ n433 ;
  assign n18769 = n18768 ^ n11337 ^ 1'b0 ;
  assign n18766 = ( x20 & ~n1114 ) | ( x20 & n3345 ) | ( ~n1114 & n3345 ) ;
  assign n18767 = ( ~n10248 & n18471 ) | ( ~n10248 & n18766 ) | ( n18471 & n18766 ) ;
  assign n18770 = n18769 ^ n18767 ^ n2898 ;
  assign n18771 = n7922 ^ n7233 ^ n483 ;
  assign n18772 = n18771 ^ n18766 ^ 1'b0 ;
  assign n18773 = n12525 & ~n18772 ;
  assign n18774 = ( n4564 & ~n6232 ) | ( n4564 & n18773 ) | ( ~n6232 & n18773 ) ;
  assign n18775 = n18774 ^ n3202 ^ n938 ;
  assign n18776 = ( ~n3443 & n4840 ) | ( ~n3443 & n18775 ) | ( n4840 & n18775 ) ;
  assign n18782 = ( n12791 & n13954 ) | ( n12791 & ~n14683 ) | ( n13954 & ~n14683 ) ;
  assign n18777 = n794 ^ x90 ^ 1'b0 ;
  assign n18778 = ~n4544 & n18038 ;
  assign n18779 = n18778 ^ n4883 ^ 1'b0 ;
  assign n18780 = n18779 ^ n14680 ^ n9267 ;
  assign n18781 = ( n17585 & n18777 ) | ( n17585 & ~n18780 ) | ( n18777 & ~n18780 ) ;
  assign n18783 = n18782 ^ n18781 ^ n16524 ;
  assign n18785 = n2915 | n8563 ;
  assign n18786 = ( ~n4147 & n16411 ) | ( ~n4147 & n18785 ) | ( n16411 & n18785 ) ;
  assign n18784 = n8243 ^ x191 ^ 1'b0 ;
  assign n18787 = n18786 ^ n18784 ^ n3488 ;
  assign n18788 = n1423 | n18787 ;
  assign n18789 = n488 | n18788 ;
  assign n18790 = n8919 | n15100 ;
  assign n18791 = ( n8037 & ~n8740 ) | ( n8037 & n12078 ) | ( ~n8740 & n12078 ) ;
  assign n18792 = n896 & n18791 ;
  assign n18793 = ~n18790 & n18792 ;
  assign n18794 = n8700 & ~n17949 ;
  assign n18795 = ( n4141 & ~n8819 ) | ( n4141 & n9347 ) | ( ~n8819 & n9347 ) ;
  assign n18796 = n18795 ^ n11195 ^ n4445 ;
  assign n18797 = ( n8738 & n9736 ) | ( n8738 & n18796 ) | ( n9736 & n18796 ) ;
  assign n18798 = ( n10908 & n18158 ) | ( n10908 & ~n18797 ) | ( n18158 & ~n18797 ) ;
  assign n18799 = ( n497 & ~n2367 ) | ( n497 & n3047 ) | ( ~n2367 & n3047 ) ;
  assign n18800 = n18799 ^ n487 ^ 1'b0 ;
  assign n18801 = ( n3464 & n17364 ) | ( n3464 & n18800 ) | ( n17364 & n18800 ) ;
  assign n18802 = ( n998 & n1598 ) | ( n998 & n1998 ) | ( n1598 & n1998 ) ;
  assign n18803 = n18802 ^ n10401 ^ n8701 ;
  assign n18804 = n18803 ^ n8458 ^ n4581 ;
  assign n18805 = ( n11659 & n13206 ) | ( n11659 & ~n18804 ) | ( n13206 & ~n18804 ) ;
  assign n18806 = n18805 ^ n16221 ^ n5503 ;
  assign n18807 = ( ~n16115 & n18801 ) | ( ~n16115 & n18806 ) | ( n18801 & n18806 ) ;
  assign n18808 = ( ~n389 & n5872 ) | ( ~n389 & n6799 ) | ( n5872 & n6799 ) ;
  assign n18809 = n18808 ^ n13916 ^ n5962 ;
  assign n18810 = ( n15085 & n16468 ) | ( n15085 & n18809 ) | ( n16468 & n18809 ) ;
  assign n18811 = ( x194 & ~n3383 ) | ( x194 & n18115 ) | ( ~n3383 & n18115 ) ;
  assign n18812 = n12333 ^ n11913 ^ n10411 ;
  assign n18813 = n18812 ^ n7087 ^ n6935 ;
  assign n18814 = n18813 ^ n8964 ^ n1804 ;
  assign n18815 = n5193 ^ n4492 ^ n3887 ;
  assign n18825 = ( ~n13574 & n14167 ) | ( ~n13574 & n17644 ) | ( n14167 & n17644 ) ;
  assign n18816 = n15064 ^ n3752 ^ n1025 ;
  assign n18817 = n1262 | n10762 ;
  assign n18818 = n18817 ^ n15460 ^ n8555 ;
  assign n18819 = ( n8045 & n18816 ) | ( n8045 & n18818 ) | ( n18816 & n18818 ) ;
  assign n18820 = ( ~n5544 & n7907 ) | ( ~n5544 & n16512 ) | ( n7907 & n16512 ) ;
  assign n18821 = n4651 ^ n2296 ^ n1661 ;
  assign n18822 = n18821 ^ n15712 ^ n7795 ;
  assign n18823 = n18820 & n18822 ;
  assign n18824 = ( n6581 & ~n18819 ) | ( n6581 & n18823 ) | ( ~n18819 & n18823 ) ;
  assign n18826 = n18825 ^ n18824 ^ n551 ;
  assign n18832 = n4142 & n10724 ;
  assign n18829 = n5833 ^ n2699 ^ n1258 ;
  assign n18830 = n18829 ^ n12443 ^ n9268 ;
  assign n18831 = ( n8151 & n14406 ) | ( n8151 & ~n18830 ) | ( n14406 & ~n18830 ) ;
  assign n18827 = n14869 ^ n13353 ^ 1'b0 ;
  assign n18828 = ( n3883 & n6491 ) | ( n3883 & ~n18827 ) | ( n6491 & ~n18827 ) ;
  assign n18833 = n18832 ^ n18831 ^ n18828 ;
  assign n18834 = n5994 ^ n1395 ^ n968 ;
  assign n18835 = n5864 | n11275 ;
  assign n18836 = n18835 ^ n3331 ^ 1'b0 ;
  assign n18837 = ( n2365 & n7205 ) | ( n2365 & n18836 ) | ( n7205 & n18836 ) ;
  assign n18838 = ~n11652 & n18837 ;
  assign n18839 = ~n18834 & n18838 ;
  assign n18840 = n18839 ^ n16059 ^ n2829 ;
  assign n18841 = ( n10770 & n12152 ) | ( n10770 & n12975 ) | ( n12152 & n12975 ) ;
  assign n18842 = ( ~n3327 & n5231 ) | ( ~n3327 & n6589 ) | ( n5231 & n6589 ) ;
  assign n18843 = n15861 ^ n15733 ^ 1'b0 ;
  assign n18844 = n18842 & n18843 ;
  assign n18845 = ( n334 & n897 ) | ( n334 & n5301 ) | ( n897 & n5301 ) ;
  assign n18846 = n9233 ^ n5468 ^ n3632 ;
  assign n18847 = ( n4478 & ~n11038 ) | ( n4478 & n18846 ) | ( ~n11038 & n18846 ) ;
  assign n18848 = ( n953 & ~n5943 ) | ( n953 & n12470 ) | ( ~n5943 & n12470 ) ;
  assign n18849 = n18848 ^ n5699 ^ n5120 ;
  assign n18850 = ~n6998 & n18849 ;
  assign n18851 = n18850 ^ n6086 ^ 1'b0 ;
  assign n18852 = ( n511 & ~n4067 ) | ( n511 & n18851 ) | ( ~n4067 & n18851 ) ;
  assign n18855 = ( ~n2461 & n2796 ) | ( ~n2461 & n11263 ) | ( n2796 & n11263 ) ;
  assign n18856 = ~n2559 & n18855 ;
  assign n18853 = n8640 ^ n2929 ^ 1'b0 ;
  assign n18854 = n17581 & n18853 ;
  assign n18857 = n18856 ^ n18854 ^ 1'b0 ;
  assign n18858 = ( ~n6098 & n16094 ) | ( ~n6098 & n18857 ) | ( n16094 & n18857 ) ;
  assign n18859 = ~n7159 & n7541 ;
  assign n18860 = n1334 & n18859 ;
  assign n18861 = n9262 | n18860 ;
  assign n18862 = n18861 ^ n3598 ^ 1'b0 ;
  assign n18863 = ~n14790 & n18862 ;
  assign n18864 = ( n7471 & n10542 ) | ( n7471 & ~n11891 ) | ( n10542 & ~n11891 ) ;
  assign n18865 = ( n4737 & n9383 ) | ( n4737 & ~n18864 ) | ( n9383 & ~n18864 ) ;
  assign n18866 = ( n5763 & n15855 ) | ( n5763 & n16483 ) | ( n15855 & n16483 ) ;
  assign n18867 = ( n1360 & ~n10089 ) | ( n1360 & n11923 ) | ( ~n10089 & n11923 ) ;
  assign n18868 = ( n1512 & n3488 ) | ( n1512 & n11115 ) | ( n3488 & n11115 ) ;
  assign n18869 = n18868 ^ n7876 ^ n4531 ;
  assign n18870 = ( n7816 & n7830 ) | ( n7816 & ~n8409 ) | ( n7830 & ~n8409 ) ;
  assign n18871 = n18870 ^ n6584 ^ n6062 ;
  assign n18872 = ( n3685 & ~n11587 ) | ( n3685 & n18871 ) | ( ~n11587 & n18871 ) ;
  assign n18873 = ( n16641 & n18869 ) | ( n16641 & ~n18872 ) | ( n18869 & ~n18872 ) ;
  assign n18874 = n12731 ^ n5527 ^ n1411 ;
  assign n18875 = ( n3188 & ~n10070 ) | ( n3188 & n10892 ) | ( ~n10070 & n10892 ) ;
  assign n18876 = n18875 ^ n8741 ^ n3472 ;
  assign n18877 = ( n7468 & n17728 ) | ( n7468 & n18876 ) | ( n17728 & n18876 ) ;
  assign n18878 = n6339 & ~n18877 ;
  assign n18879 = n18874 & n18878 ;
  assign n18880 = n8065 ^ n7897 ^ n7433 ;
  assign n18881 = n18880 ^ n14704 ^ n14306 ;
  assign n18882 = ~n1019 & n9680 ;
  assign n18883 = n18881 & n18882 ;
  assign n18884 = n16039 ^ n3087 ^ n2788 ;
  assign n18885 = n18884 ^ n6122 ^ n1005 ;
  assign n18886 = n13755 ^ n3964 ^ n374 ;
  assign n18887 = n3259 & ~n4788 ;
  assign n18888 = n409 & n18887 ;
  assign n18889 = ( ~n9713 & n11823 ) | ( ~n9713 & n18888 ) | ( n11823 & n18888 ) ;
  assign n18890 = ( n10929 & n18886 ) | ( n10929 & n18889 ) | ( n18886 & n18889 ) ;
  assign n18892 = n17132 ^ n9858 ^ n1841 ;
  assign n18891 = ( x178 & ~n7348 ) | ( x178 & n14364 ) | ( ~n7348 & n14364 ) ;
  assign n18893 = n18892 ^ n18891 ^ n16152 ;
  assign n18894 = n8341 ^ n5196 ^ n997 ;
  assign n18895 = ( n2029 & ~n6808 ) | ( n2029 & n10504 ) | ( ~n6808 & n10504 ) ;
  assign n18896 = n18894 & ~n18895 ;
  assign n18897 = n18893 & n18896 ;
  assign n18898 = n18897 ^ n13503 ^ n5688 ;
  assign n18899 = ( n6964 & ~n14294 ) | ( n6964 & n18898 ) | ( ~n14294 & n18898 ) ;
  assign n18900 = n4452 | n9466 ;
  assign n18901 = ( n8816 & ~n12109 ) | ( n8816 & n18900 ) | ( ~n12109 & n18900 ) ;
  assign n18902 = ~n17517 & n18901 ;
  assign n18903 = n18902 ^ n13982 ^ n9956 ;
  assign n18906 = n3663 | n10528 ;
  assign n18907 = ~n8816 & n18906 ;
  assign n18908 = n18907 ^ n1542 ^ 1'b0 ;
  assign n18904 = n7127 ^ n5465 ^ n467 ;
  assign n18905 = n283 & n18904 ;
  assign n18909 = n18908 ^ n18905 ^ 1'b0 ;
  assign n18910 = ( ~n3610 & n4720 ) | ( ~n3610 & n9848 ) | ( n4720 & n9848 ) ;
  assign n18911 = ( n6213 & n6399 ) | ( n6213 & n18910 ) | ( n6399 & n18910 ) ;
  assign n18912 = n5947 ^ n869 ^ n434 ;
  assign n18913 = n18912 ^ n7981 ^ n4723 ;
  assign n18914 = n18913 ^ n16190 ^ n6452 ;
  assign n18920 = n14623 ^ n1856 ^ n433 ;
  assign n18915 = n3101 | n5077 ;
  assign n18916 = n18915 ^ n11056 ^ n2013 ;
  assign n18917 = ( ~n8627 & n12760 ) | ( ~n8627 & n18916 ) | ( n12760 & n18916 ) ;
  assign n18918 = n15837 & n18917 ;
  assign n18919 = n18918 ^ n9322 ^ 1'b0 ;
  assign n18921 = n18920 ^ n18919 ^ n17580 ;
  assign n18922 = ( ~n6574 & n14004 ) | ( ~n6574 & n18921 ) | ( n14004 & n18921 ) ;
  assign n18934 = n17959 ^ n9898 ^ n7418 ;
  assign n18932 = n9459 ^ n4984 ^ n690 ;
  assign n18931 = n5630 & n13048 ;
  assign n18933 = n18932 ^ n18931 ^ n438 ;
  assign n18935 = n18934 ^ n18933 ^ n9702 ;
  assign n18923 = n15349 ^ n5332 ^ n3002 ;
  assign n18924 = n8238 & ~n11396 ;
  assign n18925 = n18924 ^ n304 ^ 1'b0 ;
  assign n18926 = ( n3409 & n5282 ) | ( n3409 & ~n18925 ) | ( n5282 & ~n18925 ) ;
  assign n18927 = n6166 & n9343 ;
  assign n18928 = n12066 & n18927 ;
  assign n18929 = ( x181 & n18926 ) | ( x181 & ~n18928 ) | ( n18926 & ~n18928 ) ;
  assign n18930 = ( n9613 & n18923 ) | ( n9613 & n18929 ) | ( n18923 & n18929 ) ;
  assign n18936 = n18935 ^ n18930 ^ n15729 ;
  assign n18953 = ( n10192 & n12049 ) | ( n10192 & ~n14039 ) | ( n12049 & ~n14039 ) ;
  assign n18937 = n6213 ^ n5683 ^ n4520 ;
  assign n18938 = n18937 ^ n15053 ^ n3571 ;
  assign n18940 = n3129 | n3184 ;
  assign n18941 = n9040 | n18940 ;
  assign n18939 = ( ~n3638 & n6307 ) | ( ~n3638 & n6325 ) | ( n6307 & n6325 ) ;
  assign n18942 = n18941 ^ n18939 ^ n8414 ;
  assign n18943 = ( ~n7587 & n18938 ) | ( ~n7587 & n18942 ) | ( n18938 & n18942 ) ;
  assign n18944 = n18943 ^ n13992 ^ n1830 ;
  assign n18949 = ( n10120 & ~n11869 ) | ( n10120 & n15673 ) | ( ~n11869 & n15673 ) ;
  assign n18946 = ( n2389 & ~n4661 ) | ( n2389 & n10866 ) | ( ~n4661 & n10866 ) ;
  assign n18947 = n18946 ^ n6465 ^ n5730 ;
  assign n18948 = n18947 ^ n7663 ^ 1'b0 ;
  assign n18945 = ( n3468 & n3537 ) | ( n3468 & n9121 ) | ( n3537 & n9121 ) ;
  assign n18950 = n18949 ^ n18948 ^ n18945 ;
  assign n18951 = ~n15577 & n18950 ;
  assign n18952 = ~n18944 & n18951 ;
  assign n18954 = n18953 ^ n18952 ^ n1072 ;
  assign n18955 = ( n15295 & n18936 ) | ( n15295 & n18954 ) | ( n18936 & n18954 ) ;
  assign n18956 = ( n562 & n2304 ) | ( n562 & n18829 ) | ( n2304 & n18829 ) ;
  assign n18957 = n18956 ^ n9912 ^ n4921 ;
  assign n18973 = n5017 ^ n2722 ^ 1'b0 ;
  assign n18974 = n18973 ^ n6264 ^ n3869 ;
  assign n18975 = ( n943 & n12182 ) | ( n943 & ~n18974 ) | ( n12182 & ~n18974 ) ;
  assign n18976 = n18975 ^ n18674 ^ n4300 ;
  assign n18971 = ( n579 & n1870 ) | ( n579 & n4275 ) | ( n1870 & n4275 ) ;
  assign n18965 = n10737 ^ n5709 ^ n3932 ;
  assign n18966 = n18965 ^ n12184 ^ n3054 ;
  assign n18967 = n18966 ^ n3309 ^ n1893 ;
  assign n18968 = n18341 | n18967 ;
  assign n18969 = n7515 & ~n18968 ;
  assign n18970 = n577 | n18969 ;
  assign n18972 = n18971 ^ n18970 ^ 1'b0 ;
  assign n18958 = ( n1548 & ~n5719 ) | ( n1548 & n10110 ) | ( ~n5719 & n10110 ) ;
  assign n18959 = ( ~n2025 & n7650 ) | ( ~n2025 & n18958 ) | ( n7650 & n18958 ) ;
  assign n18960 = ( n296 & n5972 ) | ( n296 & n6807 ) | ( n5972 & n6807 ) ;
  assign n18961 = n18960 ^ n14102 ^ n10445 ;
  assign n18962 = ( ~n3628 & n8040 ) | ( ~n3628 & n18658 ) | ( n8040 & n18658 ) ;
  assign n18963 = ( ~n17670 & n18961 ) | ( ~n17670 & n18962 ) | ( n18961 & n18962 ) ;
  assign n18964 = n18959 & n18963 ;
  assign n18977 = n18976 ^ n18972 ^ n18964 ;
  assign n18978 = n14942 ^ n14702 ^ n4042 ;
  assign n18979 = n17203 & n18978 ;
  assign n18980 = ~n17554 & n18979 ;
  assign n18984 = n10142 & ~n12705 ;
  assign n18983 = ( n7324 & n7484 ) | ( n7324 & ~n9267 ) | ( n7484 & ~n9267 ) ;
  assign n18981 = ( n1336 & n2102 ) | ( n1336 & n5633 ) | ( n2102 & n5633 ) ;
  assign n18982 = n18981 ^ n17346 ^ n3979 ;
  assign n18985 = n18984 ^ n18983 ^ n18982 ;
  assign n18986 = n15895 ^ n2174 ^ n1456 ;
  assign n18990 = n11485 & ~n11620 ;
  assign n18987 = ( n5271 & n10021 ) | ( n5271 & n15407 ) | ( n10021 & n15407 ) ;
  assign n18988 = ( n3648 & ~n5598 ) | ( n3648 & n18987 ) | ( ~n5598 & n18987 ) ;
  assign n18989 = n15317 & n18988 ;
  assign n18991 = n18990 ^ n18989 ^ 1'b0 ;
  assign n18992 = ~n13130 & n17155 ;
  assign n18993 = ( ~n1204 & n1586 ) | ( ~n1204 & n8336 ) | ( n1586 & n8336 ) ;
  assign n18994 = ( n1121 & n4382 ) | ( n1121 & n10741 ) | ( n4382 & n10741 ) ;
  assign n18995 = n18994 ^ n12399 ^ 1'b0 ;
  assign n18996 = ( ~n3263 & n11058 ) | ( ~n3263 & n18995 ) | ( n11058 & n18995 ) ;
  assign n18997 = ( n18944 & n18993 ) | ( n18944 & ~n18996 ) | ( n18993 & ~n18996 ) ;
  assign n18998 = n1991 ^ n352 ^ 1'b0 ;
  assign n18999 = n12065 ^ n10825 ^ n10036 ;
  assign n19000 = ( n4749 & n17665 ) | ( n4749 & n18999 ) | ( n17665 & n18999 ) ;
  assign n19001 = ~n18998 & n19000 ;
  assign n19002 = ~n7636 & n19001 ;
  assign n19003 = n12443 ^ n4829 ^ x21 ;
  assign n19004 = n19003 ^ n12150 ^ n10583 ;
  assign n19005 = ( n8325 & n15872 ) | ( n8325 & ~n19004 ) | ( n15872 & ~n19004 ) ;
  assign n19006 = ( ~n1446 & n5491 ) | ( ~n1446 & n19005 ) | ( n5491 & n19005 ) ;
  assign n19007 = n12590 ^ n3303 ^ n2930 ;
  assign n19008 = n19007 ^ n3881 ^ 1'b0 ;
  assign n19010 = ( n3106 & ~n5233 ) | ( n3106 & n5376 ) | ( ~n5233 & n5376 ) ;
  assign n19009 = n9230 ^ n9143 ^ n1729 ;
  assign n19011 = n19010 ^ n19009 ^ n16420 ;
  assign n19012 = n15678 ^ n12578 ^ n371 ;
  assign n19013 = n11289 ^ n4431 ^ n1605 ;
  assign n19014 = n15493 ^ n10178 ^ 1'b0 ;
  assign n19015 = n15388 & ~n19014 ;
  assign n19016 = ( x211 & n19013 ) | ( x211 & ~n19015 ) | ( n19013 & ~n19015 ) ;
  assign n19018 = ( n2454 & n11275 ) | ( n2454 & n15333 ) | ( n11275 & n15333 ) ;
  assign n19019 = ( n8026 & n8680 ) | ( n8026 & ~n19018 ) | ( n8680 & ~n19018 ) ;
  assign n19017 = ( n1961 & ~n4315 ) | ( n1961 & n4746 ) | ( ~n4315 & n4746 ) ;
  assign n19020 = n19019 ^ n19017 ^ n6173 ;
  assign n19021 = ( n1538 & n6787 ) | ( n1538 & ~n8646 ) | ( n6787 & ~n8646 ) ;
  assign n19022 = ( n2256 & n13005 ) | ( n2256 & n15188 ) | ( n13005 & n15188 ) ;
  assign n19023 = ( n3508 & n6150 ) | ( n3508 & n15350 ) | ( n6150 & n15350 ) ;
  assign n19024 = ( n19021 & n19022 ) | ( n19021 & n19023 ) | ( n19022 & n19023 ) ;
  assign n19027 = n2585 & ~n3779 ;
  assign n19025 = ( n6930 & n12493 ) | ( n6930 & ~n14853 ) | ( n12493 & ~n14853 ) ;
  assign n19026 = ( n1513 & n16685 ) | ( n1513 & n19025 ) | ( n16685 & n19025 ) ;
  assign n19028 = n19027 ^ n19026 ^ n5216 ;
  assign n19029 = n19028 ^ n6106 ^ n1223 ;
  assign n19030 = n11397 ^ n7178 ^ n5519 ;
  assign n19031 = n19030 ^ n6450 ^ n1089 ;
  assign n19032 = ( ~n16631 & n19029 ) | ( ~n16631 & n19031 ) | ( n19029 & n19031 ) ;
  assign n19033 = n13342 ^ n3042 ^ n2295 ;
  assign n19038 = ~n4836 & n7019 ;
  assign n19039 = ~n8152 & n19038 ;
  assign n19034 = n12482 ^ n791 ^ 1'b0 ;
  assign n19035 = n13893 & n19034 ;
  assign n19036 = ( ~n2220 & n2731 ) | ( ~n2220 & n4470 ) | ( n2731 & n4470 ) ;
  assign n19037 = ( n2600 & n19035 ) | ( n2600 & n19036 ) | ( n19035 & n19036 ) ;
  assign n19040 = n19039 ^ n19037 ^ n13086 ;
  assign n19041 = ( n7107 & n9893 ) | ( n7107 & ~n16919 ) | ( n9893 & ~n16919 ) ;
  assign n19042 = n19041 ^ n3592 ^ n571 ;
  assign n19043 = ( ~n6058 & n8121 ) | ( ~n6058 & n19042 ) | ( n8121 & n19042 ) ;
  assign n19044 = n3547 ^ x56 ^ 1'b0 ;
  assign n19045 = ~n19043 & n19044 ;
  assign n19046 = n3240 & ~n11245 ;
  assign n19047 = n2431 & n19046 ;
  assign n19048 = n19047 ^ n17484 ^ n2598 ;
  assign n19049 = ( n15301 & ~n17076 ) | ( n15301 & n19048 ) | ( ~n17076 & n19048 ) ;
  assign n19055 = ( n2495 & ~n5750 ) | ( n2495 & n10246 ) | ( ~n5750 & n10246 ) ;
  assign n19056 = n19055 ^ n17799 ^ n1539 ;
  assign n19054 = n18588 ^ n17707 ^ n7683 ;
  assign n19050 = n18048 ^ n13662 ^ n7010 ;
  assign n19051 = ~n9370 & n17470 ;
  assign n19052 = ~n621 & n19051 ;
  assign n19053 = ( n11425 & ~n19050 ) | ( n11425 & n19052 ) | ( ~n19050 & n19052 ) ;
  assign n19057 = n19056 ^ n19054 ^ n19053 ;
  assign n19058 = n19057 ^ n18317 ^ n2670 ;
  assign n19059 = ( n2028 & ~n10309 ) | ( n2028 & n15806 ) | ( ~n10309 & n15806 ) ;
  assign n19060 = ( n2483 & ~n7416 ) | ( n2483 & n8171 ) | ( ~n7416 & n8171 ) ;
  assign n19069 = ( x188 & n410 ) | ( x188 & ~n3939 ) | ( n410 & ~n3939 ) ;
  assign n19066 = n8646 ^ n5614 ^ n1000 ;
  assign n19065 = n5180 ^ n1609 ^ x157 ;
  assign n19067 = n19066 ^ n19065 ^ n10102 ;
  assign n19064 = n16976 ^ n12004 ^ n3404 ;
  assign n19068 = n19067 ^ n19064 ^ n2433 ;
  assign n19070 = n19069 ^ n19068 ^ n13663 ;
  assign n19061 = n4123 ^ n1579 ^ 1'b0 ;
  assign n19062 = n4308 & ~n19061 ;
  assign n19063 = n19062 ^ n14158 ^ n7333 ;
  assign n19071 = n19070 ^ n19063 ^ n15469 ;
  assign n19072 = ( n11928 & ~n19060 ) | ( n11928 & n19071 ) | ( ~n19060 & n19071 ) ;
  assign n19073 = ( n4016 & n5319 ) | ( n4016 & ~n8117 ) | ( n5319 & ~n8117 ) ;
  assign n19074 = ( n1246 & ~n5220 ) | ( n1246 & n19073 ) | ( ~n5220 & n19073 ) ;
  assign n19075 = ( ~n3805 & n17318 ) | ( ~n3805 & n19074 ) | ( n17318 & n19074 ) ;
  assign n19076 = n19075 ^ n2840 ^ 1'b0 ;
  assign n19077 = n8025 & ~n19076 ;
  assign n19078 = n19077 ^ n4263 ^ 1'b0 ;
  assign n19082 = n2097 & ~n9486 ;
  assign n19080 = ( ~n785 & n8380 ) | ( ~n785 & n18779 ) | ( n8380 & n18779 ) ;
  assign n19079 = n9608 ^ n7260 ^ n916 ;
  assign n19081 = n19080 ^ n19079 ^ n5848 ;
  assign n19083 = n19082 ^ n19081 ^ n16346 ;
  assign n19086 = n14136 ^ n11666 ^ n3152 ;
  assign n19084 = n13958 ^ n13804 ^ n1817 ;
  assign n19085 = ( n497 & n16757 ) | ( n497 & ~n19084 ) | ( n16757 & ~n19084 ) ;
  assign n19087 = n19086 ^ n19085 ^ n15047 ;
  assign n19106 = x146 & ~n16068 ;
  assign n19107 = n19106 ^ x19 ^ 1'b0 ;
  assign n19108 = ( ~n3130 & n10467 ) | ( ~n3130 & n19107 ) | ( n10467 & n19107 ) ;
  assign n19088 = n12466 ^ n11046 ^ n2106 ;
  assign n19089 = n5843 & ~n19088 ;
  assign n19090 = ( n7952 & n14285 ) | ( n7952 & n19089 ) | ( n14285 & n19089 ) ;
  assign n19091 = n15775 ^ n10690 ^ n5406 ;
  assign n19092 = ~n8739 & n19091 ;
  assign n19093 = n10932 ^ n10628 ^ n724 ;
  assign n19094 = ( n5164 & ~n10624 ) | ( n5164 & n19093 ) | ( ~n10624 & n19093 ) ;
  assign n19095 = ~n3915 & n19094 ;
  assign n19096 = n19095 ^ n456 ^ 1'b0 ;
  assign n19098 = n10899 ^ n3910 ^ n2624 ;
  assign n19099 = n3105 & n19098 ;
  assign n19100 = n3333 & n19099 ;
  assign n19097 = n11653 ^ n10173 ^ n5150 ;
  assign n19101 = n19100 ^ n19097 ^ n10650 ;
  assign n19102 = ( ~n12121 & n17788 ) | ( ~n12121 & n19101 ) | ( n17788 & n19101 ) ;
  assign n19103 = n19102 ^ n9227 ^ n4944 ;
  assign n19104 = ( ~n9485 & n19096 ) | ( ~n9485 & n19103 ) | ( n19096 & n19103 ) ;
  assign n19105 = ( n19090 & n19092 ) | ( n19090 & ~n19104 ) | ( n19092 & ~n19104 ) ;
  assign n19109 = n19108 ^ n19105 ^ n15247 ;
  assign n19110 = x32 & ~n4967 ;
  assign n19111 = n19110 ^ n18039 ^ n529 ;
  assign n19112 = n19111 ^ n17534 ^ n16452 ;
  assign n19113 = ( n7603 & ~n8199 ) | ( n7603 & n19112 ) | ( ~n8199 & n19112 ) ;
  assign n19114 = ( n2578 & ~n4300 ) | ( n2578 & n13468 ) | ( ~n4300 & n13468 ) ;
  assign n19115 = n12684 ^ n3243 ^ 1'b0 ;
  assign n19116 = n12251 & n19115 ;
  assign n19117 = n2738 & n19116 ;
  assign n19118 = ( ~n9142 & n12103 ) | ( ~n9142 & n19117 ) | ( n12103 & n19117 ) ;
  assign n19119 = n17065 ^ n5154 ^ 1'b0 ;
  assign n19120 = ( n2727 & n4474 ) | ( n2727 & ~n19119 ) | ( n4474 & ~n19119 ) ;
  assign n19121 = ( ~n5113 & n7072 ) | ( ~n5113 & n8903 ) | ( n7072 & n8903 ) ;
  assign n19122 = n9594 ^ n4159 ^ n3234 ;
  assign n19123 = n19122 ^ n15898 ^ n3723 ;
  assign n19124 = ( n7649 & n19121 ) | ( n7649 & ~n19123 ) | ( n19121 & ~n19123 ) ;
  assign n19125 = ( n11220 & ~n19120 ) | ( n11220 & n19124 ) | ( ~n19120 & n19124 ) ;
  assign n19126 = n8204 ^ n6684 ^ 1'b0 ;
  assign n19127 = n632 & ~n2489 ;
  assign n19128 = ( n10730 & n16894 ) | ( n10730 & ~n19127 ) | ( n16894 & ~n19127 ) ;
  assign n19129 = n12151 ^ n12044 ^ n2637 ;
  assign n19130 = ( n2775 & ~n9280 ) | ( n2775 & n19129 ) | ( ~n9280 & n19129 ) ;
  assign n19131 = ( n5885 & ~n6082 ) | ( n5885 & n7396 ) | ( ~n6082 & n7396 ) ;
  assign n19132 = n3960 & ~n6537 ;
  assign n19133 = n19132 ^ n10598 ^ 1'b0 ;
  assign n19134 = ( n4471 & ~n19131 ) | ( n4471 & n19133 ) | ( ~n19131 & n19133 ) ;
  assign n19135 = ( ~n4447 & n19130 ) | ( ~n4447 & n19134 ) | ( n19130 & n19134 ) ;
  assign n19136 = n15934 ^ n12454 ^ 1'b0 ;
  assign n19137 = n14069 | n19136 ;
  assign n19138 = ( n15047 & n19135 ) | ( n15047 & n19137 ) | ( n19135 & n19137 ) ;
  assign n19139 = ( x176 & n740 ) | ( x176 & n1094 ) | ( n740 & n1094 ) ;
  assign n19140 = ( x49 & ~x110 ) | ( x49 & n19139 ) | ( ~x110 & n19139 ) ;
  assign n19141 = n19140 ^ n5574 ^ n4889 ;
  assign n19142 = ( n2392 & n13124 ) | ( n2392 & ~n19141 ) | ( n13124 & ~n19141 ) ;
  assign n19143 = n19142 ^ n1838 ^ n881 ;
  assign n19153 = ( n3530 & n5706 ) | ( n3530 & ~n7095 ) | ( n5706 & ~n7095 ) ;
  assign n19144 = ( n762 & ~n5338 ) | ( n762 & n7289 ) | ( ~n5338 & n7289 ) ;
  assign n19145 = n14213 ^ n2377 ^ 1'b0 ;
  assign n19146 = n17503 & n19145 ;
  assign n19147 = ( n11686 & n19144 ) | ( n11686 & ~n19146 ) | ( n19144 & ~n19146 ) ;
  assign n19148 = n702 | n971 ;
  assign n19149 = n7234 | n19148 ;
  assign n19150 = n1228 & n19149 ;
  assign n19151 = n19150 ^ n16319 ^ 1'b0 ;
  assign n19152 = ( ~n14818 & n19147 ) | ( ~n14818 & n19151 ) | ( n19147 & n19151 ) ;
  assign n19154 = n19153 ^ n19152 ^ n378 ;
  assign n19155 = n11585 ^ n11311 ^ n2303 ;
  assign n19156 = n17937 ^ n3095 ^ n1131 ;
  assign n19157 = ( ~n2641 & n13067 ) | ( ~n2641 & n19156 ) | ( n13067 & n19156 ) ;
  assign n19163 = ( n7088 & n10719 ) | ( n7088 & n12520 ) | ( n10719 & n12520 ) ;
  assign n19158 = ( n987 & ~n8255 ) | ( n987 & n17026 ) | ( ~n8255 & n17026 ) ;
  assign n19159 = n6863 ^ x14 ^ 1'b0 ;
  assign n19160 = n19159 ^ n7352 ^ n4914 ;
  assign n19161 = ( ~n13894 & n19158 ) | ( ~n13894 & n19160 ) | ( n19158 & n19160 ) ;
  assign n19162 = ( n3461 & n3550 ) | ( n3461 & n19161 ) | ( n3550 & n19161 ) ;
  assign n19164 = n19163 ^ n19162 ^ n5095 ;
  assign n19165 = ( n1660 & n2694 ) | ( n1660 & n7407 ) | ( n2694 & n7407 ) ;
  assign n19166 = n8083 ^ n3278 ^ n2655 ;
  assign n19167 = ( n9256 & n10428 ) | ( n9256 & ~n19166 ) | ( n10428 & ~n19166 ) ;
  assign n19168 = n19167 ^ n18619 ^ 1'b0 ;
  assign n19169 = n6898 | n19168 ;
  assign n19170 = ( n19164 & ~n19165 ) | ( n19164 & n19169 ) | ( ~n19165 & n19169 ) ;
  assign n19171 = n10217 ^ n4992 ^ n1666 ;
  assign n19172 = n6762 ^ n2700 ^ 1'b0 ;
  assign n19173 = n2213 | n19172 ;
  assign n19174 = n19173 ^ n17162 ^ n14887 ;
  assign n19175 = ( n4648 & ~n4965 ) | ( n4648 & n9729 ) | ( ~n4965 & n9729 ) ;
  assign n19176 = n19175 ^ n5468 ^ n4877 ;
  assign n19177 = n13153 ^ n10314 ^ x217 ;
  assign n19178 = ( n4521 & ~n10341 ) | ( n4521 & n18480 ) | ( ~n10341 & n18480 ) ;
  assign n19181 = ( ~n3829 & n5876 ) | ( ~n3829 & n7361 ) | ( n5876 & n7361 ) ;
  assign n19182 = ( ~n2025 & n3500 ) | ( ~n2025 & n19181 ) | ( n3500 & n19181 ) ;
  assign n19183 = n19182 ^ n4153 ^ n2803 ;
  assign n19179 = ( n2100 & ~n10689 ) | ( n2100 & n11821 ) | ( ~n10689 & n11821 ) ;
  assign n19180 = n6706 & ~n19179 ;
  assign n19184 = n19183 ^ n19180 ^ n7599 ;
  assign n19185 = n19184 ^ x137 ^ x67 ;
  assign n19186 = ( n12640 & ~n19178 ) | ( n12640 & n19185 ) | ( ~n19178 & n19185 ) ;
  assign n19187 = n18522 ^ n12731 ^ 1'b0 ;
  assign n19188 = n12082 ^ n9576 ^ n2225 ;
  assign n19189 = ( n10072 & n13169 ) | ( n10072 & n19188 ) | ( n13169 & n19188 ) ;
  assign n19190 = n17953 ^ n7216 ^ n4102 ;
  assign n19191 = ( n8849 & n10637 ) | ( n8849 & n19190 ) | ( n10637 & n19190 ) ;
  assign n19192 = n9259 ^ n8937 ^ x131 ;
  assign n19193 = ( n8350 & ~n12564 ) | ( n8350 & n17084 ) | ( ~n12564 & n17084 ) ;
  assign n19194 = ( n5456 & n19192 ) | ( n5456 & n19193 ) | ( n19192 & n19193 ) ;
  assign n19195 = n19194 ^ n4042 ^ n2758 ;
  assign n19198 = ( n4579 & n9605 ) | ( n4579 & ~n18152 ) | ( n9605 & ~n18152 ) ;
  assign n19196 = ( n3206 & ~n3649 ) | ( n3206 & n10544 ) | ( ~n3649 & n10544 ) ;
  assign n19197 = n19196 ^ n17006 ^ n3244 ;
  assign n19199 = n19198 ^ n19197 ^ 1'b0 ;
  assign n19200 = n19199 ^ n5503 ^ n1283 ;
  assign n19201 = n5782 ^ n4967 ^ n4041 ;
  assign n19204 = ( n1744 & n6272 ) | ( n1744 & n9299 ) | ( n6272 & n9299 ) ;
  assign n19202 = n5584 & n11891 ;
  assign n19203 = n19202 ^ n11168 ^ 1'b0 ;
  assign n19205 = n19204 ^ n19203 ^ 1'b0 ;
  assign n19206 = n12783 & n19205 ;
  assign n19207 = ( ~n18223 & n19201 ) | ( ~n18223 & n19206 ) | ( n19201 & n19206 ) ;
  assign n19208 = n4322 ^ n1511 ^ n1500 ;
  assign n19209 = ( n479 & n6988 ) | ( n479 & n10300 ) | ( n6988 & n10300 ) ;
  assign n19210 = n19209 ^ n11962 ^ x186 ;
  assign n19211 = n19210 ^ n9275 ^ x173 ;
  assign n19212 = ( n5520 & ~n8321 ) | ( n5520 & n8472 ) | ( ~n8321 & n8472 ) ;
  assign n19213 = ~n1848 & n19212 ;
  assign n19214 = n19213 ^ n9365 ^ 1'b0 ;
  assign n19215 = ( n10046 & n19211 ) | ( n10046 & ~n19214 ) | ( n19211 & ~n19214 ) ;
  assign n19216 = ( ~n6894 & n13834 ) | ( ~n6894 & n18721 ) | ( n13834 & n18721 ) ;
  assign n19217 = ( ~n3522 & n14447 ) | ( ~n3522 & n17831 ) | ( n14447 & n17831 ) ;
  assign n19218 = n19217 ^ n13744 ^ n3677 ;
  assign n19219 = n10282 ^ n9560 ^ n6226 ;
  assign n19220 = n19219 ^ n13957 ^ n3801 ;
  assign n19221 = ( n498 & ~n2590 ) | ( n498 & n19220 ) | ( ~n2590 & n19220 ) ;
  assign n19222 = n9557 ^ n3601 ^ 1'b0 ;
  assign n19223 = ( ~n1971 & n8987 ) | ( ~n1971 & n9826 ) | ( n8987 & n9826 ) ;
  assign n19224 = n17647 ^ n14970 ^ n10721 ;
  assign n19225 = n18190 ^ n2586 ^ 1'b0 ;
  assign n19226 = n5566 | n19225 ;
  assign n19227 = ( n1167 & n9121 ) | ( n1167 & ~n12200 ) | ( n9121 & ~n12200 ) ;
  assign n19228 = n11959 ^ n6940 ^ x102 ;
  assign n19229 = ( ~n5653 & n11641 ) | ( ~n5653 & n19228 ) | ( n11641 & n19228 ) ;
  assign n19230 = n1015 & ~n14939 ;
  assign n19231 = ~n14026 & n19230 ;
  assign n19232 = n19231 ^ n16956 ^ n11154 ;
  assign n19233 = n19232 ^ n16790 ^ n11490 ;
  assign n19234 = ( n9434 & n19229 ) | ( n9434 & ~n19233 ) | ( n19229 & ~n19233 ) ;
  assign n19235 = ( n407 & ~n10862 ) | ( n407 & n14796 ) | ( ~n10862 & n14796 ) ;
  assign n19236 = ( n1653 & n6823 ) | ( n1653 & n19235 ) | ( n6823 & n19235 ) ;
  assign n19238 = n14997 ^ n12338 ^ n1299 ;
  assign n19239 = ( n1151 & ~n7524 ) | ( n1151 & n19238 ) | ( ~n7524 & n19238 ) ;
  assign n19237 = ~n688 & n4284 ;
  assign n19240 = n19239 ^ n19237 ^ 1'b0 ;
  assign n19241 = ( n1988 & ~n8951 ) | ( n1988 & n19240 ) | ( ~n8951 & n19240 ) ;
  assign n19242 = ( n524 & n12904 ) | ( n524 & n17604 ) | ( n12904 & n17604 ) ;
  assign n19243 = ( ~n13681 & n16969 ) | ( ~n13681 & n19242 ) | ( n16969 & n19242 ) ;
  assign n19244 = ( n6468 & n17408 ) | ( n6468 & n19243 ) | ( n17408 & n19243 ) ;
  assign n19245 = n19244 ^ n16468 ^ n11679 ;
  assign n19246 = ( ~n6828 & n7098 ) | ( ~n6828 & n8327 ) | ( n7098 & n8327 ) ;
  assign n19247 = ( ~n5194 & n18074 ) | ( ~n5194 & n19246 ) | ( n18074 & n19246 ) ;
  assign n19248 = ( n5628 & n19245 ) | ( n5628 & ~n19247 ) | ( n19245 & ~n19247 ) ;
  assign n19250 = n2362 & ~n6194 ;
  assign n19251 = n19250 ^ n13744 ^ n1795 ;
  assign n19252 = ( ~n328 & n17990 ) | ( ~n328 & n19251 ) | ( n17990 & n19251 ) ;
  assign n19253 = n19252 ^ n13436 ^ n384 ;
  assign n19249 = ( n7369 & n12481 ) | ( n7369 & ~n14725 ) | ( n12481 & ~n14725 ) ;
  assign n19254 = n19253 ^ n19249 ^ n710 ;
  assign n19255 = ( x50 & n5476 ) | ( x50 & n11845 ) | ( n5476 & n11845 ) ;
  assign n19256 = ( n11291 & ~n18974 ) | ( n11291 & n19255 ) | ( ~n18974 & n19255 ) ;
  assign n19257 = ( n4346 & n18257 ) | ( n4346 & n19256 ) | ( n18257 & n19256 ) ;
  assign n19258 = n17445 ^ n560 ^ 1'b0 ;
  assign n19259 = n19258 ^ n12916 ^ n3449 ;
  assign n19260 = n16824 ^ n11562 ^ n5863 ;
  assign n19261 = n9697 & n19260 ;
  assign n19265 = ( n4888 & ~n6172 ) | ( n4888 & n6659 ) | ( ~n6172 & n6659 ) ;
  assign n19266 = n19265 ^ n4020 ^ n896 ;
  assign n19264 = n5776 ^ n1420 ^ 1'b0 ;
  assign n19267 = n19266 ^ n19264 ^ n2169 ;
  assign n19262 = n12929 ^ n1397 ^ n936 ;
  assign n19263 = n19262 ^ n8891 ^ n8430 ;
  assign n19268 = n19267 ^ n19263 ^ 1'b0 ;
  assign n19269 = n16589 & n19268 ;
  assign n19270 = ( n3520 & ~n4637 ) | ( n3520 & n7113 ) | ( ~n4637 & n7113 ) ;
  assign n19271 = n9076 ^ n2683 ^ 1'b0 ;
  assign n19272 = n19270 & ~n19271 ;
  assign n19273 = n8994 & n19272 ;
  assign n19274 = ( x112 & n10390 ) | ( x112 & ~n19273 ) | ( n10390 & ~n19273 ) ;
  assign n19275 = n17562 ^ n6304 ^ n498 ;
  assign n19276 = n11913 & n19275 ;
  assign n19277 = ( ~n5821 & n19274 ) | ( ~n5821 & n19276 ) | ( n19274 & n19276 ) ;
  assign n19278 = n8308 & n14558 ;
  assign n19279 = n2291 & n19278 ;
  assign n19280 = ( n2662 & n5618 ) | ( n2662 & ~n15073 ) | ( n5618 & ~n15073 ) ;
  assign n19281 = n19280 ^ n11045 ^ n5182 ;
  assign n19282 = ( n1780 & n5045 ) | ( n1780 & n19281 ) | ( n5045 & n19281 ) ;
  assign n19283 = ( n11771 & n19279 ) | ( n11771 & n19282 ) | ( n19279 & n19282 ) ;
  assign n19293 = n5178 ^ n2532 ^ n830 ;
  assign n19294 = n19293 ^ n8257 ^ n6375 ;
  assign n19295 = n19294 ^ n7698 ^ n6116 ;
  assign n19284 = ( n2129 & n3109 ) | ( n2129 & n4408 ) | ( n3109 & n4408 ) ;
  assign n19285 = n7681 ^ n1663 ^ n1069 ;
  assign n19286 = ( n4341 & ~n19284 ) | ( n4341 & n19285 ) | ( ~n19284 & n19285 ) ;
  assign n19287 = ( n971 & ~n10200 ) | ( n971 & n19286 ) | ( ~n10200 & n19286 ) ;
  assign n19290 = ( n2459 & n3395 ) | ( n2459 & ~n12455 ) | ( n3395 & ~n12455 ) ;
  assign n19288 = ( n3577 & ~n5809 ) | ( n3577 & n10605 ) | ( ~n5809 & n10605 ) ;
  assign n19289 = ( n419 & ~n18205 ) | ( n419 & n19288 ) | ( ~n18205 & n19288 ) ;
  assign n19291 = n19290 ^ n19289 ^ n6416 ;
  assign n19292 = ( n17348 & ~n19287 ) | ( n17348 & n19291 ) | ( ~n19287 & n19291 ) ;
  assign n19296 = n19295 ^ n19292 ^ n3035 ;
  assign n19297 = n5207 & ~n12068 ;
  assign n19298 = ~n13344 & n19297 ;
  assign n19299 = n12765 ^ n7325 ^ 1'b0 ;
  assign n19300 = n5358 & n19299 ;
  assign n19301 = ( n2112 & n17841 ) | ( n2112 & ~n19300 ) | ( n17841 & ~n19300 ) ;
  assign n19302 = n15048 ^ n8453 ^ x151 ;
  assign n19303 = n19302 ^ n8144 ^ 1'b0 ;
  assign n19304 = n9629 | n19303 ;
  assign n19305 = n4862 ^ n3863 ^ n2890 ;
  assign n19306 = ( n3365 & ~n12120 ) | ( n3365 & n19305 ) | ( ~n12120 & n19305 ) ;
  assign n19307 = ( n9882 & ~n10938 ) | ( n9882 & n19306 ) | ( ~n10938 & n19306 ) ;
  assign n19308 = ( n2853 & n10110 ) | ( n2853 & ~n12260 ) | ( n10110 & ~n12260 ) ;
  assign n19309 = ( n4571 & n4653 ) | ( n4571 & ~n19308 ) | ( n4653 & ~n19308 ) ;
  assign n19310 = ( n12625 & n19307 ) | ( n12625 & n19309 ) | ( n19307 & n19309 ) ;
  assign n19311 = ( n4913 & ~n7059 ) | ( n4913 & n14235 ) | ( ~n7059 & n14235 ) ;
  assign n19312 = n15582 ^ n15156 ^ n4623 ;
  assign n19315 = ( ~x15 & n2341 ) | ( ~x15 & n7462 ) | ( n2341 & n7462 ) ;
  assign n19313 = n6931 ^ n5013 ^ n3059 ;
  assign n19314 = ( x88 & n4329 ) | ( x88 & n19313 ) | ( n4329 & n19313 ) ;
  assign n19316 = n19315 ^ n19314 ^ n8904 ;
  assign n19317 = n12138 & ~n19316 ;
  assign n19318 = ( n16523 & ~n19312 ) | ( n16523 & n19317 ) | ( ~n19312 & n19317 ) ;
  assign n19324 = n4949 ^ n3780 ^ n2618 ;
  assign n19325 = ( n9905 & n15030 ) | ( n9905 & n19324 ) | ( n15030 & n19324 ) ;
  assign n19326 = n19325 ^ n8141 ^ n2449 ;
  assign n19320 = n11388 ^ n2580 ^ 1'b0 ;
  assign n19321 = n19320 ^ n3587 ^ n3201 ;
  assign n19322 = n16650 | n19321 ;
  assign n19319 = n3460 | n9587 ;
  assign n19323 = n19322 ^ n19319 ^ n10686 ;
  assign n19327 = n19326 ^ n19323 ^ n7128 ;
  assign n19331 = n12079 ^ n7740 ^ n4609 ;
  assign n19332 = n19331 ^ n11232 ^ n10476 ;
  assign n19328 = n12295 ^ n6573 ^ n1595 ;
  assign n19329 = ( n2821 & n3197 ) | ( n2821 & ~n6738 ) | ( n3197 & ~n6738 ) ;
  assign n19330 = ( n18286 & ~n19328 ) | ( n18286 & n19329 ) | ( ~n19328 & n19329 ) ;
  assign n19333 = n19332 ^ n19330 ^ n9746 ;
  assign n19334 = n12109 ^ n7554 ^ n3142 ;
  assign n19335 = n12807 & n19334 ;
  assign n19336 = ~n7476 & n19335 ;
  assign n19337 = ~n9026 & n19336 ;
  assign n19338 = ( n8179 & n8608 ) | ( n8179 & n10650 ) | ( n8608 & n10650 ) ;
  assign n19342 = n9796 & ~n16730 ;
  assign n19343 = n19342 ^ n6875 ^ 1'b0 ;
  assign n19344 = ( n1303 & n9575 ) | ( n1303 & ~n19343 ) | ( n9575 & ~n19343 ) ;
  assign n19345 = n19344 ^ n5670 ^ 1'b0 ;
  assign n19346 = n3352 & ~n19345 ;
  assign n19347 = ( n4874 & ~n16280 ) | ( n4874 & n19346 ) | ( ~n16280 & n19346 ) ;
  assign n19339 = ( ~n6199 & n7691 ) | ( ~n6199 & n14244 ) | ( n7691 & n14244 ) ;
  assign n19340 = ( n10341 & ~n18959 ) | ( n10341 & n19339 ) | ( ~n18959 & n19339 ) ;
  assign n19341 = ( n13950 & n17573 ) | ( n13950 & n19340 ) | ( n17573 & n19340 ) ;
  assign n19348 = n19347 ^ n19341 ^ n942 ;
  assign n19356 = n11306 ^ n5581 ^ n1390 ;
  assign n19357 = n19356 ^ n10461 ^ n2497 ;
  assign n19352 = n537 & ~n4217 ;
  assign n19353 = n19352 ^ n1460 ^ 1'b0 ;
  assign n19354 = ( ~n2101 & n6827 ) | ( ~n2101 & n8286 ) | ( n6827 & n8286 ) ;
  assign n19355 = n19353 & ~n19354 ;
  assign n19358 = n19357 ^ n19355 ^ 1'b0 ;
  assign n19349 = n3833 | n6031 ;
  assign n19350 = n9337 ^ n5196 ^ n1726 ;
  assign n19351 = ( n9946 & ~n19349 ) | ( n9946 & n19350 ) | ( ~n19349 & n19350 ) ;
  assign n19359 = n19358 ^ n19351 ^ n15960 ;
  assign n19360 = ( n16243 & ~n17958 ) | ( n16243 & n19359 ) | ( ~n17958 & n19359 ) ;
  assign n19361 = ( n365 & n1684 ) | ( n365 & ~n7122 ) | ( n1684 & ~n7122 ) ;
  assign n19362 = ( n1112 & ~n1473 ) | ( n1112 & n19361 ) | ( ~n1473 & n19361 ) ;
  assign n19363 = n16138 ^ n11806 ^ n2953 ;
  assign n19364 = n16868 ^ n8347 ^ n4434 ;
  assign n19365 = n8579 & n19364 ;
  assign n19366 = ( n9443 & n19363 ) | ( n9443 & n19365 ) | ( n19363 & n19365 ) ;
  assign n19367 = n12892 ^ n1507 ^ n1058 ;
  assign n19368 = n19367 ^ n9449 ^ n5189 ;
  assign n19369 = ( n7678 & n9894 ) | ( n7678 & n13846 ) | ( n9894 & n13846 ) ;
  assign n19370 = ( ~x157 & n7914 ) | ( ~x157 & n19369 ) | ( n7914 & n19369 ) ;
  assign n19371 = n19370 ^ n10986 ^ n7222 ;
  assign n19372 = ( n10536 & n11503 ) | ( n10536 & n18475 ) | ( n11503 & n18475 ) ;
  assign n19373 = n14901 ^ n13155 ^ n5414 ;
  assign n19374 = ( x118 & n19372 ) | ( x118 & ~n19373 ) | ( n19372 & ~n19373 ) ;
  assign n19375 = n16068 ^ n15270 ^ n7227 ;
  assign n19376 = ( n8421 & ~n8660 ) | ( n8421 & n19375 ) | ( ~n8660 & n19375 ) ;
  assign n19377 = n19376 ^ n12677 ^ n2944 ;
  assign n19378 = n9395 | n13553 ;
  assign n19379 = n19377 | n19378 ;
  assign n19380 = n6197 ^ n5965 ^ n4558 ;
  assign n19381 = n19380 ^ n17322 ^ n10474 ;
  assign n19382 = ( n812 & n15614 ) | ( n812 & ~n19381 ) | ( n15614 & ~n19381 ) ;
  assign n19386 = n1966 & n7672 ;
  assign n19383 = n1850 ^ n1566 ^ n1300 ;
  assign n19384 = ~n5272 & n19383 ;
  assign n19385 = n19384 ^ n8378 ^ 1'b0 ;
  assign n19387 = n19386 ^ n19385 ^ n7184 ;
  assign n19388 = n13603 ^ x168 ^ x151 ;
  assign n19389 = ( n8448 & n16090 ) | ( n8448 & n18252 ) | ( n16090 & n18252 ) ;
  assign n19390 = n19389 ^ n3281 ^ 1'b0 ;
  assign n19391 = n19388 & ~n19390 ;
  assign n19392 = n8930 | n9062 ;
  assign n19393 = n19392 ^ n763 ^ 1'b0 ;
  assign n19394 = ( n7095 & ~n8882 ) | ( n7095 & n19393 ) | ( ~n8882 & n19393 ) ;
  assign n19395 = n19394 ^ n17860 ^ n8682 ;
  assign n19396 = ( n4067 & ~n6693 ) | ( n4067 & n11397 ) | ( ~n6693 & n11397 ) ;
  assign n19411 = ( n1621 & ~n5126 ) | ( n1621 & n12470 ) | ( ~n5126 & n12470 ) ;
  assign n19409 = n7764 ^ n4116 ^ n3656 ;
  assign n19410 = n19409 ^ n17185 ^ n15744 ;
  assign n19412 = n19411 ^ n19410 ^ n10875 ;
  assign n19397 = n2624 ^ n873 ^ n367 ;
  assign n19398 = ( ~n8622 & n16636 ) | ( ~n8622 & n19397 ) | ( n16636 & n19397 ) ;
  assign n19399 = ( n1800 & ~n3271 ) | ( n1800 & n19398 ) | ( ~n3271 & n19398 ) ;
  assign n19400 = n12698 ^ n10150 ^ n9591 ;
  assign n19401 = ( n6659 & n10377 ) | ( n6659 & n11820 ) | ( n10377 & n11820 ) ;
  assign n19402 = n16965 | n19401 ;
  assign n19403 = n19402 ^ x82 ^ 1'b0 ;
  assign n19404 = ( n464 & ~n19400 ) | ( n464 & n19403 ) | ( ~n19400 & n19403 ) ;
  assign n19405 = ( n5308 & n19399 ) | ( n5308 & n19404 ) | ( n19399 & n19404 ) ;
  assign n19406 = ( n293 & n2044 ) | ( n293 & ~n17524 ) | ( n2044 & ~n17524 ) ;
  assign n19407 = n19406 ^ n5475 ^ 1'b0 ;
  assign n19408 = n19405 | n19407 ;
  assign n19413 = n19412 ^ n19408 ^ n5891 ;
  assign n19414 = n2223 ^ x170 ^ 1'b0 ;
  assign n19415 = ( n8515 & n11144 ) | ( n8515 & ~n12386 ) | ( n11144 & ~n12386 ) ;
  assign n19416 = ( ~n19142 & n19414 ) | ( ~n19142 & n19415 ) | ( n19414 & n19415 ) ;
  assign n19417 = n19416 ^ n15923 ^ n9950 ;
  assign n19418 = ( n8553 & n11056 ) | ( n8553 & n13992 ) | ( n11056 & n13992 ) ;
  assign n19420 = n19389 ^ n16251 ^ n5590 ;
  assign n19419 = n9627 ^ n2712 ^ n1238 ;
  assign n19421 = n19420 ^ n19419 ^ n10677 ;
  assign n19422 = ( ~n5631 & n19418 ) | ( ~n5631 & n19421 ) | ( n19418 & n19421 ) ;
  assign n19423 = ( n3991 & n16970 ) | ( n3991 & ~n18688 ) | ( n16970 & ~n18688 ) ;
  assign n19425 = n379 & n9894 ;
  assign n19426 = ( n3262 & n3408 ) | ( n3262 & n10672 ) | ( n3408 & n10672 ) ;
  assign n19427 = ( n839 & n19425 ) | ( n839 & ~n19426 ) | ( n19425 & ~n19426 ) ;
  assign n19424 = ( n3937 & ~n11411 ) | ( n3937 & n16070 ) | ( ~n11411 & n16070 ) ;
  assign n19428 = n19427 ^ n19424 ^ n1307 ;
  assign n19429 = n6447 ^ n2513 ^ n1245 ;
  assign n19430 = ( n6079 & ~n7606 ) | ( n6079 & n14593 ) | ( ~n7606 & n14593 ) ;
  assign n19431 = ( n16043 & ~n19429 ) | ( n16043 & n19430 ) | ( ~n19429 & n19430 ) ;
  assign n19432 = n10454 ^ n10327 ^ n4502 ;
  assign n19433 = ( ~n11169 & n18310 ) | ( ~n11169 & n19432 ) | ( n18310 & n19432 ) ;
  assign n19437 = n7759 ^ n6982 ^ 1'b0 ;
  assign n19438 = n4404 & n19437 ;
  assign n19434 = ( n368 & ~n12747 ) | ( n368 & n19411 ) | ( ~n12747 & n19411 ) ;
  assign n19435 = ( n8338 & n17937 ) | ( n8338 & n19434 ) | ( n17937 & n19434 ) ;
  assign n19436 = ( ~n511 & n8939 ) | ( ~n511 & n19435 ) | ( n8939 & n19435 ) ;
  assign n19439 = n19438 ^ n19436 ^ n6175 ;
  assign n19441 = n589 | n3857 ;
  assign n19442 = n2195 & ~n19441 ;
  assign n19440 = ( n688 & n2228 ) | ( n688 & n16939 ) | ( n2228 & n16939 ) ;
  assign n19443 = n19442 ^ n19440 ^ x10 ;
  assign n19444 = ( n407 & ~n2635 ) | ( n407 & n19443 ) | ( ~n2635 & n19443 ) ;
  assign n19445 = n506 & ~n4802 ;
  assign n19446 = ( n7903 & n10180 ) | ( n7903 & n19445 ) | ( n10180 & n19445 ) ;
  assign n19455 = n5074 ^ n2742 ^ n1757 ;
  assign n19456 = n19455 ^ n4109 ^ 1'b0 ;
  assign n19457 = x236 & n19456 ;
  assign n19453 = ( n3622 & n6864 ) | ( n3622 & n15615 ) | ( n6864 & n15615 ) ;
  assign n19454 = n19453 ^ n1732 ^ n1389 ;
  assign n19447 = ( ~n2257 & n9624 ) | ( ~n2257 & n17954 ) | ( n9624 & n17954 ) ;
  assign n19448 = n19447 ^ n13085 ^ 1'b0 ;
  assign n19449 = n6768 | n15014 ;
  assign n19450 = ( ~n950 & n2064 ) | ( ~n950 & n18077 ) | ( n2064 & n18077 ) ;
  assign n19451 = n19449 & ~n19450 ;
  assign n19452 = ( ~n19228 & n19448 ) | ( ~n19228 & n19451 ) | ( n19448 & n19451 ) ;
  assign n19458 = n19457 ^ n19454 ^ n19452 ;
  assign n19459 = n7780 ^ n6847 ^ n3302 ;
  assign n19460 = n19459 ^ n7894 ^ x235 ;
  assign n19461 = n14998 & ~n19460 ;
  assign n19462 = n11716 ^ n7784 ^ n1226 ;
  assign n19463 = ~n6045 & n19462 ;
  assign n19464 = n2059 & n19463 ;
  assign n19465 = n16114 ^ n7290 ^ n6592 ;
  assign n19466 = n16567 ^ n4446 ^ n679 ;
  assign n19467 = n19466 ^ n16726 ^ n9578 ;
  assign n19468 = ( n4452 & n17265 ) | ( n4452 & ~n19467 ) | ( n17265 & ~n19467 ) ;
  assign n19469 = n3152 & ~n4693 ;
  assign n19470 = n19469 ^ n2680 ^ 1'b0 ;
  assign n19471 = ( ~n537 & n9747 ) | ( ~n537 & n19470 ) | ( n9747 & n19470 ) ;
  assign n19472 = n19471 ^ n10108 ^ 1'b0 ;
  assign n19473 = n11710 | n19472 ;
  assign n19474 = x105 & n8591 ;
  assign n19475 = ( n917 & ~n6169 ) | ( n917 & n16114 ) | ( ~n6169 & n16114 ) ;
  assign n19476 = n19475 ^ n15255 ^ n8271 ;
  assign n19477 = ( ~n6121 & n6195 ) | ( ~n6121 & n12357 ) | ( n6195 & n12357 ) ;
  assign n19478 = n7287 ^ n3186 ^ n1233 ;
  assign n19479 = n19478 ^ n4400 ^ n3156 ;
  assign n19480 = ( n9337 & n9856 ) | ( n9337 & n19479 ) | ( n9856 & n19479 ) ;
  assign n19483 = n9917 ^ n6786 ^ n6609 ;
  assign n19484 = n19483 ^ n4851 ^ 1'b0 ;
  assign n19485 = ( ~n1809 & n19158 ) | ( ~n1809 & n19484 ) | ( n19158 & n19484 ) ;
  assign n19481 = n10085 & n16591 ;
  assign n19482 = ~n16298 & n19481 ;
  assign n19486 = n19485 ^ n19482 ^ n1160 ;
  assign n19487 = ( n19477 & n19480 ) | ( n19477 & ~n19486 ) | ( n19480 & ~n19486 ) ;
  assign n19488 = n10494 ^ n8348 ^ n2059 ;
  assign n19489 = ( ~n12365 & n15038 ) | ( ~n12365 & n19488 ) | ( n15038 & n19488 ) ;
  assign n19490 = n19343 ^ n17871 ^ n2829 ;
  assign n19494 = ( n519 & n4238 ) | ( n519 & ~n14690 ) | ( n4238 & ~n14690 ) ;
  assign n19492 = ( n1160 & n7114 ) | ( n1160 & ~n14940 ) | ( n7114 & ~n14940 ) ;
  assign n19493 = ( x170 & ~n18376 ) | ( x170 & n19492 ) | ( ~n18376 & n19492 ) ;
  assign n19491 = ( n7381 & n10938 ) | ( n7381 & ~n12546 ) | ( n10938 & ~n12546 ) ;
  assign n19495 = n19494 ^ n19493 ^ n19491 ;
  assign n19496 = ( n2542 & n19490 ) | ( n2542 & n19495 ) | ( n19490 & n19495 ) ;
  assign n19500 = ( n4123 & n6066 ) | ( n4123 & ~n10105 ) | ( n6066 & ~n10105 ) ;
  assign n19501 = n19500 ^ n11346 ^ n1861 ;
  assign n19499 = n6599 ^ n2250 ^ 1'b0 ;
  assign n19502 = n19501 ^ n19499 ^ n1837 ;
  assign n19497 = n16997 ^ n14243 ^ n4054 ;
  assign n19498 = n19497 ^ n3131 ^ n872 ;
  assign n19503 = n19502 ^ n19498 ^ n548 ;
  assign n19504 = n10997 ^ n7685 ^ n6025 ;
  assign n19505 = ( n2179 & n3692 ) | ( n2179 & ~n5951 ) | ( n3692 & ~n5951 ) ;
  assign n19506 = n19505 ^ n4832 ^ n2376 ;
  assign n19507 = n19506 ^ n7921 ^ 1'b0 ;
  assign n19508 = n19504 & ~n19507 ;
  assign n19514 = n12757 ^ n5321 ^ n2920 ;
  assign n19510 = ( ~n856 & n9607 ) | ( ~n856 & n9843 ) | ( n9607 & n9843 ) ;
  assign n19509 = ( n320 & ~n12525 ) | ( n320 & n16172 ) | ( ~n12525 & n16172 ) ;
  assign n19511 = n19510 ^ n19509 ^ n11257 ;
  assign n19512 = n19019 ^ n5408 ^ 1'b0 ;
  assign n19513 = ( ~n297 & n19511 ) | ( ~n297 & n19512 ) | ( n19511 & n19512 ) ;
  assign n19515 = n19514 ^ n19513 ^ n15892 ;
  assign n19516 = ( n430 & n2316 ) | ( n430 & ~n3282 ) | ( n2316 & ~n3282 ) ;
  assign n19517 = n14350 ^ n12858 ^ n648 ;
  assign n19518 = ( n6462 & ~n19516 ) | ( n6462 & n19517 ) | ( ~n19516 & n19517 ) ;
  assign n19519 = n6093 & n8733 ;
  assign n19520 = n12962 ^ n8056 ^ 1'b0 ;
  assign n19521 = ( n1191 & n12552 ) | ( n1191 & ~n19520 ) | ( n12552 & ~n19520 ) ;
  assign n19522 = ( n6186 & n12912 ) | ( n6186 & ~n19521 ) | ( n12912 & ~n19521 ) ;
  assign n19523 = n19522 ^ n11383 ^ 1'b0 ;
  assign n19524 = n19519 | n19523 ;
  assign n19525 = n4187 ^ n3541 ^ n3527 ;
  assign n19526 = ( n8803 & n16733 ) | ( n8803 & n19525 ) | ( n16733 & n19525 ) ;
  assign n19527 = n5616 ^ n2277 ^ 1'b0 ;
  assign n19528 = n19527 ^ n9449 ^ n8699 ;
  assign n19529 = n4350 & n6150 ;
  assign n19530 = ~n19528 & n19529 ;
  assign n19531 = ( ~n8912 & n9084 ) | ( ~n8912 & n19530 ) | ( n9084 & n19530 ) ;
  assign n19532 = n1482 & n11998 ;
  assign n19533 = n19532 ^ n15737 ^ n14503 ;
  assign n19534 = ( n3332 & ~n9576 ) | ( n3332 & n13943 ) | ( ~n9576 & n13943 ) ;
  assign n19535 = n19534 ^ n11804 ^ n6203 ;
  assign n19536 = n19535 ^ n17996 ^ n16164 ;
  assign n19537 = ( n1427 & ~n9513 ) | ( n1427 & n14984 ) | ( ~n9513 & n14984 ) ;
  assign n19538 = n19537 ^ n18448 ^ n6330 ;
  assign n19539 = n19538 ^ n16474 ^ n6490 ;
  assign n19540 = ~n13795 & n13882 ;
  assign n19543 = n7354 ^ n5035 ^ 1'b0 ;
  assign n19544 = n1073 | n19543 ;
  assign n19545 = ( n10167 & ~n10181 ) | ( n10167 & n19544 ) | ( ~n10181 & n19544 ) ;
  assign n19541 = n6164 ^ n2908 ^ n389 ;
  assign n19542 = n19541 ^ n15624 ^ n15150 ;
  assign n19546 = n19545 ^ n19542 ^ n5470 ;
  assign n19547 = ( n2877 & ~n9611 ) | ( n2877 & n19546 ) | ( ~n9611 & n19546 ) ;
  assign n19548 = ( n1747 & n10036 ) | ( n1747 & n18871 ) | ( n10036 & n18871 ) ;
  assign n19549 = n19548 ^ n8406 ^ n1677 ;
  assign n19550 = ( n19540 & n19547 ) | ( n19540 & n19549 ) | ( n19547 & n19549 ) ;
  assign n19551 = n489 | n16451 ;
  assign n19552 = n19551 ^ n7367 ^ 1'b0 ;
  assign n19553 = n19552 ^ n6048 ^ n1841 ;
  assign n19554 = ( n14489 & ~n14509 ) | ( n14489 & n19553 ) | ( ~n14509 & n19553 ) ;
  assign n19555 = n11314 & ~n16039 ;
  assign n19556 = n1985 & n19555 ;
  assign n19557 = n7939 & ~n16322 ;
  assign n19558 = n19556 & n19557 ;
  assign n19559 = n19558 ^ n6710 ^ n4656 ;
  assign n19560 = n19559 ^ n12769 ^ n4261 ;
  assign n19561 = ( n5837 & n8877 ) | ( n5837 & ~n12489 ) | ( n8877 & ~n12489 ) ;
  assign n19562 = ( ~n756 & n4805 ) | ( ~n756 & n19561 ) | ( n4805 & n19561 ) ;
  assign n19563 = ( ~n15029 & n16741 ) | ( ~n15029 & n19562 ) | ( n16741 & n19562 ) ;
  assign n19564 = n8824 ^ n499 ^ 1'b0 ;
  assign n19565 = n7258 & ~n19564 ;
  assign n19566 = n19565 ^ n2082 ^ 1'b0 ;
  assign n19567 = n16522 & n19566 ;
  assign n19568 = n15991 | n19567 ;
  assign n19569 = n19568 ^ n19249 ^ 1'b0 ;
  assign n19570 = n14558 ^ n6171 ^ n4407 ;
  assign n19571 = n19570 ^ n18301 ^ n1670 ;
  assign n19572 = ( n11703 & ~n15286 ) | ( n11703 & n18773 ) | ( ~n15286 & n18773 ) ;
  assign n19573 = n16242 ^ n13909 ^ n4820 ;
  assign n19574 = ( n4021 & ~n19572 ) | ( n4021 & n19573 ) | ( ~n19572 & n19573 ) ;
  assign n19575 = n5782 | n14634 ;
  assign n19576 = n12951 | n19575 ;
  assign n19577 = ( n2147 & n8260 ) | ( n2147 & n9966 ) | ( n8260 & n9966 ) ;
  assign n19578 = ( ~n909 & n5920 ) | ( ~n909 & n11020 ) | ( n5920 & n11020 ) ;
  assign n19579 = ( n9918 & ~n15398 ) | ( n9918 & n19578 ) | ( ~n15398 & n19578 ) ;
  assign n19580 = ( n6567 & n19577 ) | ( n6567 & ~n19579 ) | ( n19577 & ~n19579 ) ;
  assign n19581 = n18619 ^ n9665 ^ n8140 ;
  assign n19582 = n11723 ^ n5646 ^ 1'b0 ;
  assign n19583 = n19582 ^ n11649 ^ n10179 ;
  assign n19584 = n280 & n19583 ;
  assign n19585 = ( n2338 & n2502 ) | ( n2338 & n6300 ) | ( n2502 & n6300 ) ;
  assign n19586 = n19585 ^ n13509 ^ n995 ;
  assign n19587 = n14423 & ~n19586 ;
  assign n19597 = n7863 ^ n7152 ^ 1'b0 ;
  assign n19598 = n1962 | n19597 ;
  assign n19588 = n10781 ^ n1778 ^ n1304 ;
  assign n19589 = n7325 & n19588 ;
  assign n19590 = n19589 ^ n11916 ^ 1'b0 ;
  assign n19591 = n19590 ^ n12182 ^ n7523 ;
  assign n19592 = n10482 ^ n2136 ^ 1'b0 ;
  assign n19593 = n4846 & n19592 ;
  assign n19594 = n19591 & n19593 ;
  assign n19595 = ~n15213 & n19594 ;
  assign n19596 = ( n7385 & n19485 ) | ( n7385 & n19595 ) | ( n19485 & n19595 ) ;
  assign n19599 = n19598 ^ n19596 ^ n18390 ;
  assign n19602 = ( n950 & n5106 ) | ( n950 & ~n5229 ) | ( n5106 & ~n5229 ) ;
  assign n19600 = n17407 ^ n3511 ^ 1'b0 ;
  assign n19601 = n6688 & n19600 ;
  assign n19603 = n19602 ^ n19601 ^ 1'b0 ;
  assign n19604 = n6160 & n13036 ;
  assign n19605 = ~n1775 & n19604 ;
  assign n19606 = ( n5422 & n7683 ) | ( n5422 & ~n18576 ) | ( n7683 & ~n18576 ) ;
  assign n19607 = n7262 & n7654 ;
  assign n19608 = ( n6392 & ~n7046 ) | ( n6392 & n19607 ) | ( ~n7046 & n19607 ) ;
  assign n19609 = n19606 & ~n19608 ;
  assign n19610 = n527 & n12674 ;
  assign n19611 = n19610 ^ n1047 ^ x251 ;
  assign n19612 = n13835 ^ n1911 ^ n1247 ;
  assign n19613 = n19612 ^ n5077 ^ 1'b0 ;
  assign n19614 = n3922 & n19613 ;
  assign n19615 = n13450 ^ n12463 ^ n8942 ;
  assign n19616 = ~n7913 & n19615 ;
  assign n19617 = ( ~n6901 & n19614 ) | ( ~n6901 & n19616 ) | ( n19614 & n19616 ) ;
  assign n19618 = n3822 ^ n3496 ^ n1184 ;
  assign n19619 = ( n1057 & n3897 ) | ( n1057 & n8537 ) | ( n3897 & n8537 ) ;
  assign n19620 = n19619 ^ n19219 ^ n4611 ;
  assign n19621 = ( n4505 & n12188 ) | ( n4505 & n19620 ) | ( n12188 & n19620 ) ;
  assign n19622 = ( n5288 & n19618 ) | ( n5288 & n19621 ) | ( n19618 & n19621 ) ;
  assign n19630 = ( n4744 & n5591 ) | ( n4744 & n6683 ) | ( n5591 & n6683 ) ;
  assign n19631 = n13212 & ~n19630 ;
  assign n19632 = ~n16207 & n19590 ;
  assign n19633 = n19632 ^ n11071 ^ 1'b0 ;
  assign n19634 = ( n12183 & ~n19631 ) | ( n12183 & n19633 ) | ( ~n19631 & n19633 ) ;
  assign n19629 = ( ~n4051 & n8125 ) | ( ~n4051 & n13037 ) | ( n8125 & n13037 ) ;
  assign n19635 = n19634 ^ n19629 ^ n2680 ;
  assign n19623 = n17005 ^ n8943 ^ 1'b0 ;
  assign n19624 = n1917 & ~n8220 ;
  assign n19625 = n19624 ^ n13896 ^ 1'b0 ;
  assign n19626 = n19625 ^ n8661 ^ n1425 ;
  assign n19627 = n19626 ^ n19425 ^ 1'b0 ;
  assign n19628 = ~n19623 & n19627 ;
  assign n19636 = n19635 ^ n19628 ^ 1'b0 ;
  assign n19637 = n5007 & ~n9418 ;
  assign n19638 = ~n7319 & n19637 ;
  assign n19639 = ( n1759 & n7176 ) | ( n1759 & ~n12310 ) | ( n7176 & ~n12310 ) ;
  assign n19640 = ( n4055 & n10156 ) | ( n4055 & n19639 ) | ( n10156 & n19639 ) ;
  assign n19641 = n11357 ^ n11000 ^ n7380 ;
  assign n19642 = ( n11705 & n19640 ) | ( n11705 & n19641 ) | ( n19640 & n19641 ) ;
  assign n19643 = ( n3548 & ~n4538 ) | ( n3548 & n16904 ) | ( ~n4538 & n16904 ) ;
  assign n19644 = ( n7834 & ~n17631 ) | ( n7834 & n19643 ) | ( ~n17631 & n19643 ) ;
  assign n19645 = ( ~n3898 & n12936 ) | ( ~n3898 & n14418 ) | ( n12936 & n14418 ) ;
  assign n19646 = n13140 ^ n5475 ^ n865 ;
  assign n19647 = n19646 ^ n10874 ^ n261 ;
  assign n19648 = n3653 | n11252 ;
  assign n19649 = ( n2114 & n2790 ) | ( n2114 & n10762 ) | ( n2790 & n10762 ) ;
  assign n19650 = n19649 ^ n1266 ^ 1'b0 ;
  assign n19651 = n19650 ^ n12979 ^ n9169 ;
  assign n19652 = ~n4917 & n12169 ;
  assign n19653 = ~n6411 & n19652 ;
  assign n19654 = ( ~n2260 & n5984 ) | ( ~n2260 & n19653 ) | ( n5984 & n19653 ) ;
  assign n19657 = n2851 & ~n8116 ;
  assign n19658 = n19657 ^ n13684 ^ 1'b0 ;
  assign n19659 = ( n1749 & ~n8291 ) | ( n1749 & n19658 ) | ( ~n8291 & n19658 ) ;
  assign n19655 = n7934 ^ n4974 ^ n1284 ;
  assign n19656 = ( n12714 & n17739 ) | ( n12714 & ~n19655 ) | ( n17739 & ~n19655 ) ;
  assign n19660 = n19659 ^ n19656 ^ n8939 ;
  assign n19664 = ( n2275 & n6884 ) | ( n2275 & ~n13670 ) | ( n6884 & ~n13670 ) ;
  assign n19665 = ( ~n7655 & n11084 ) | ( ~n7655 & n19664 ) | ( n11084 & n19664 ) ;
  assign n19666 = ~n13381 & n18454 ;
  assign n19667 = ( n2389 & n19665 ) | ( n2389 & ~n19666 ) | ( n19665 & ~n19666 ) ;
  assign n19661 = n13160 ^ n12262 ^ n5548 ;
  assign n19662 = n260 & n19661 ;
  assign n19663 = n19662 ^ n11928 ^ 1'b0 ;
  assign n19668 = n19667 ^ n19663 ^ 1'b0 ;
  assign n19669 = ( n19654 & ~n19660 ) | ( n19654 & n19668 ) | ( ~n19660 & n19668 ) ;
  assign n19670 = n9164 ^ n815 ^ 1'b0 ;
  assign n19671 = ( ~n478 & n9817 ) | ( ~n478 & n19670 ) | ( n9817 & n19670 ) ;
  assign n19672 = n7631 ^ n5896 ^ n718 ;
  assign n19677 = n9296 ^ n8341 ^ n4509 ;
  assign n19673 = n6183 ^ n1767 ^ n1243 ;
  assign n19674 = ~n19484 & n19673 ;
  assign n19675 = n19674 ^ n12975 ^ n3198 ;
  assign n19676 = ( n3791 & n10282 ) | ( n3791 & ~n19675 ) | ( n10282 & ~n19675 ) ;
  assign n19678 = n19677 ^ n19676 ^ 1'b0 ;
  assign n19679 = ~n19672 & n19678 ;
  assign n19683 = ( ~n1735 & n5083 ) | ( ~n1735 & n5624 ) | ( n5083 & n5624 ) ;
  assign n19684 = ( n9682 & n13780 ) | ( n9682 & ~n19683 ) | ( n13780 & ~n19683 ) ;
  assign n19685 = ( n8629 & n16105 ) | ( n8629 & ~n19684 ) | ( n16105 & ~n19684 ) ;
  assign n19686 = ( ~n7198 & n18645 ) | ( ~n7198 & n19685 ) | ( n18645 & n19685 ) ;
  assign n19681 = ( n2593 & n3595 ) | ( n2593 & n6471 ) | ( n3595 & n6471 ) ;
  assign n19680 = n15585 | n18058 ;
  assign n19682 = n19681 ^ n19680 ^ n7286 ;
  assign n19687 = n19686 ^ n19682 ^ n15398 ;
  assign n19691 = ( ~n334 & n3225 ) | ( ~n334 & n3244 ) | ( n3225 & n3244 ) ;
  assign n19692 = ( n2569 & ~n14012 ) | ( n2569 & n19691 ) | ( ~n14012 & n19691 ) ;
  assign n19688 = n365 & ~n1632 ;
  assign n19689 = n17942 & n19688 ;
  assign n19690 = n19689 ^ n11759 ^ n1437 ;
  assign n19693 = n19692 ^ n19690 ^ n4610 ;
  assign n19694 = ( n5809 & n6361 ) | ( n5809 & n19693 ) | ( n6361 & n19693 ) ;
  assign n19695 = ( ~n1648 & n8237 ) | ( ~n1648 & n11354 ) | ( n8237 & n11354 ) ;
  assign n19696 = ( n5462 & ~n14637 ) | ( n5462 & n19695 ) | ( ~n14637 & n19695 ) ;
  assign n19697 = ( ~n11114 & n19694 ) | ( ~n11114 & n19696 ) | ( n19694 & n19696 ) ;
  assign n19698 = n1571 & n2393 ;
  assign n19699 = ~n2101 & n19698 ;
  assign n19700 = n4647 ^ n3947 ^ n627 ;
  assign n19701 = n19700 ^ n14026 ^ n2377 ;
  assign n19703 = n17602 ^ n4436 ^ 1'b0 ;
  assign n19704 = ~n18270 & n19703 ;
  assign n19702 = ( n5834 & n7688 ) | ( n5834 & ~n17215 ) | ( n7688 & ~n17215 ) ;
  assign n19705 = n19704 ^ n19702 ^ n13764 ;
  assign n19706 = n7756 ^ n3484 ^ n787 ;
  assign n19707 = n16638 ^ n9783 ^ n5607 ;
  assign n19708 = ( n18549 & n19706 ) | ( n18549 & ~n19707 ) | ( n19706 & ~n19707 ) ;
  assign n19709 = ( n2717 & ~n8159 ) | ( n2717 & n18998 ) | ( ~n8159 & n18998 ) ;
  assign n19710 = n16415 ^ n8771 ^ 1'b0 ;
  assign n19711 = n16821 | n19710 ;
  assign n19712 = ( n19708 & n19709 ) | ( n19708 & n19711 ) | ( n19709 & n19711 ) ;
  assign n19713 = n19712 ^ n13770 ^ n5686 ;
  assign n19714 = ( n2332 & n4610 ) | ( n2332 & ~n7588 ) | ( n4610 & ~n7588 ) ;
  assign n19715 = n10980 & ~n19714 ;
  assign n19716 = ( ~n2766 & n2777 ) | ( ~n2766 & n16288 ) | ( n2777 & n16288 ) ;
  assign n19717 = ( n8842 & ~n16140 ) | ( n8842 & n19716 ) | ( ~n16140 & n19716 ) ;
  assign n19718 = n15262 ^ n9218 ^ n1952 ;
  assign n19719 = ( n12757 & n13705 ) | ( n12757 & n19718 ) | ( n13705 & n19718 ) ;
  assign n19720 = n2319 ^ n1835 ^ n858 ;
  assign n19721 = ~n4638 & n19720 ;
  assign n19722 = n19721 ^ n8134 ^ n5845 ;
  assign n19723 = ( n1776 & n19719 ) | ( n1776 & n19722 ) | ( n19719 & n19722 ) ;
  assign n19724 = ( n11693 & ~n19717 ) | ( n11693 & n19723 ) | ( ~n19717 & n19723 ) ;
  assign n19725 = n8565 ^ n537 ^ 1'b0 ;
  assign n19726 = ( n856 & n1243 ) | ( n856 & n3619 ) | ( n1243 & n3619 ) ;
  assign n19727 = n19726 ^ n13063 ^ n7031 ;
  assign n19728 = n10525 ^ n9740 ^ n4574 ;
  assign n19729 = n19728 ^ n19607 ^ n12260 ;
  assign n19730 = ( n8128 & ~n15737 ) | ( n8128 & n19729 ) | ( ~n15737 & n19729 ) ;
  assign n19731 = n11129 ^ n7136 ^ n6648 ;
  assign n19732 = ( n19727 & ~n19730 ) | ( n19727 & n19731 ) | ( ~n19730 & n19731 ) ;
  assign n19734 = n5647 | n6912 ;
  assign n19735 = n19734 ^ n3742 ^ 1'b0 ;
  assign n19733 = ( n290 & ~n2163 ) | ( n290 & n5060 ) | ( ~n2163 & n5060 ) ;
  assign n19736 = n19735 ^ n19733 ^ n9177 ;
  assign n19737 = n14154 ^ n12330 ^ n11807 ;
  assign n19738 = ( ~n6833 & n19736 ) | ( ~n6833 & n19737 ) | ( n19736 & n19737 ) ;
  assign n19742 = n1852 ^ n574 ^ 1'b0 ;
  assign n19740 = n9135 ^ n8959 ^ n6901 ;
  assign n19739 = ( n7501 & n9427 ) | ( n7501 & n17565 ) | ( n9427 & n17565 ) ;
  assign n19741 = n19740 ^ n19739 ^ n3610 ;
  assign n19743 = n19742 ^ n19741 ^ n4400 ;
  assign n19745 = n5793 ^ n1766 ^ 1'b0 ;
  assign n19746 = ~n15368 & n19745 ;
  assign n19747 = ( n9807 & n15422 ) | ( n9807 & n19746 ) | ( n15422 & n19746 ) ;
  assign n19748 = n10249 & ~n19747 ;
  assign n19749 = n19748 ^ n2145 ^ 1'b0 ;
  assign n19744 = n8555 & n17443 ;
  assign n19750 = n19749 ^ n19744 ^ 1'b0 ;
  assign n19751 = n561 | n15374 ;
  assign n19752 = n7926 ^ n7824 ^ n6455 ;
  assign n19753 = n19752 ^ n9633 ^ n4620 ;
  assign n19754 = n19753 ^ x199 ^ 1'b0 ;
  assign n19755 = ( n7357 & n7587 ) | ( n7357 & ~n19754 ) | ( n7587 & ~n19754 ) ;
  assign n19756 = ( n3343 & n8109 ) | ( n3343 & n13545 ) | ( n8109 & n13545 ) ;
  assign n19757 = ( ~n10474 & n12668 ) | ( ~n10474 & n15400 ) | ( n12668 & n15400 ) ;
  assign n19758 = ( n14227 & n19756 ) | ( n14227 & ~n19757 ) | ( n19756 & ~n19757 ) ;
  assign n19763 = n15664 ^ n13521 ^ 1'b0 ;
  assign n19762 = n7995 ^ n4240 ^ 1'b0 ;
  assign n19759 = n13265 ^ n9585 ^ n9352 ;
  assign n19760 = ~n18321 & n19759 ;
  assign n19761 = n5941 & n19760 ;
  assign n19764 = n19763 ^ n19762 ^ n19761 ;
  assign n19765 = ( n1350 & ~n6645 ) | ( n1350 & n12789 ) | ( ~n6645 & n12789 ) ;
  assign n19766 = n13420 | n18653 ;
  assign n19767 = ( x231 & ~n6873 ) | ( x231 & n19766 ) | ( ~n6873 & n19766 ) ;
  assign n19768 = ( n9677 & n18490 ) | ( n9677 & n19767 ) | ( n18490 & n19767 ) ;
  assign n19772 = ~n5623 & n6264 ;
  assign n19773 = n19772 ^ n9576 ^ 1'b0 ;
  assign n19774 = n14763 ^ n14485 ^ n8595 ;
  assign n19775 = n19774 ^ n4329 ^ 1'b0 ;
  assign n19776 = n19773 & n19775 ;
  assign n19769 = n11358 ^ n6934 ^ n4872 ;
  assign n19770 = n10377 ^ n5721 ^ n407 ;
  assign n19771 = ( ~n3354 & n19769 ) | ( ~n3354 & n19770 ) | ( n19769 & n19770 ) ;
  assign n19777 = n19776 ^ n19771 ^ n18181 ;
  assign n19778 = ( ~n3121 & n19768 ) | ( ~n3121 & n19777 ) | ( n19768 & n19777 ) ;
  assign n19779 = ~n18873 & n19778 ;
  assign n19780 = n19765 & n19779 ;
  assign n19781 = n4111 ^ n3819 ^ n1336 ;
  assign n19782 = ( n7857 & ~n15602 ) | ( n7857 & n19674 ) | ( ~n15602 & n19674 ) ;
  assign n19783 = ( n3969 & n19781 ) | ( n3969 & ~n19782 ) | ( n19781 & ~n19782 ) ;
  assign n19784 = ( n8607 & n16250 ) | ( n8607 & ~n19783 ) | ( n16250 & ~n19783 ) ;
  assign n19790 = n13213 ^ n1747 ^ n1724 ;
  assign n19791 = ( n5070 & n6521 ) | ( n5070 & n19790 ) | ( n6521 & n19790 ) ;
  assign n19785 = n14788 ^ n3759 ^ 1'b0 ;
  assign n19786 = ( n302 & n3062 ) | ( n302 & n19785 ) | ( n3062 & n19785 ) ;
  assign n19787 = ( n2033 & ~n5625 ) | ( n2033 & n19786 ) | ( ~n5625 & n19786 ) ;
  assign n19788 = n17240 & n19787 ;
  assign n19789 = ~n18370 & n19788 ;
  assign n19792 = n19791 ^ n19789 ^ n11162 ;
  assign n19793 = ( ~x243 & n9138 ) | ( ~x243 & n13271 ) | ( n9138 & n13271 ) ;
  assign n19794 = n19793 ^ n16511 ^ n6324 ;
  assign n19795 = ( n9773 & n18854 ) | ( n9773 & n19794 ) | ( n18854 & n19794 ) ;
  assign n19796 = n8523 ^ n4796 ^ 1'b0 ;
  assign n19797 = n19796 ^ n10883 ^ n9770 ;
  assign n19798 = ~n3260 & n19797 ;
  assign n19799 = ( n4206 & n17718 ) | ( n4206 & n19798 ) | ( n17718 & n19798 ) ;
  assign n19800 = ( n11101 & n12463 ) | ( n11101 & ~n19799 ) | ( n12463 & ~n19799 ) ;
  assign n19801 = n19800 ^ n17997 ^ n11088 ;
  assign n19802 = ( ~x154 & n1900 ) | ( ~x154 & n7227 ) | ( n1900 & n7227 ) ;
  assign n19803 = n9310 & ~n19802 ;
  assign n19804 = ( n6878 & n11535 ) | ( n6878 & ~n19803 ) | ( n11535 & ~n19803 ) ;
  assign n19805 = n3749 & n19091 ;
  assign n19806 = n19804 & n19805 ;
  assign n19807 = n19806 ^ n19105 ^ n18862 ;
  assign n19808 = ( n1954 & n10541 ) | ( n1954 & n11452 ) | ( n10541 & n11452 ) ;
  assign n19809 = ( ~n1286 & n4904 ) | ( ~n1286 & n13034 ) | ( n4904 & n13034 ) ;
  assign n19810 = n19809 ^ n16866 ^ 1'b0 ;
  assign n19811 = ~n4406 & n19810 ;
  assign n19812 = ( n4687 & ~n13999 ) | ( n4687 & n17452 ) | ( ~n13999 & n17452 ) ;
  assign n19813 = n19812 ^ n6934 ^ n2696 ;
  assign n19814 = ( ~n4876 & n9731 ) | ( ~n4876 & n19813 ) | ( n9731 & n19813 ) ;
  assign n19815 = ( n268 & ~n3730 ) | ( n268 & n10727 ) | ( ~n3730 & n10727 ) ;
  assign n19816 = n19815 ^ n17040 ^ n5433 ;
  assign n19817 = ( n5110 & n18079 ) | ( n5110 & n19816 ) | ( n18079 & n19816 ) ;
  assign n19818 = ( n3375 & ~n5546 ) | ( n3375 & n19817 ) | ( ~n5546 & n19817 ) ;
  assign n19819 = ( ~n19811 & n19814 ) | ( ~n19811 & n19818 ) | ( n19814 & n19818 ) ;
  assign n19820 = ( ~n4633 & n7064 ) | ( ~n4633 & n16029 ) | ( n7064 & n16029 ) ;
  assign n19821 = n19820 ^ n10180 ^ n1818 ;
  assign n19822 = ( n19808 & ~n19819 ) | ( n19808 & n19821 ) | ( ~n19819 & n19821 ) ;
  assign n19834 = n17710 ^ n3986 ^ n3588 ;
  assign n19829 = ( ~n7093 & n17252 ) | ( ~n7093 & n17866 ) | ( n17252 & n17866 ) ;
  assign n19830 = ( ~n2157 & n8629 ) | ( ~n2157 & n19829 ) | ( n8629 & n19829 ) ;
  assign n19831 = ( n2433 & n8128 ) | ( n2433 & ~n19830 ) | ( n8128 & ~n19830 ) ;
  assign n19832 = n6827 | n19831 ;
  assign n19833 = n19832 ^ n1644 ^ 1'b0 ;
  assign n19835 = n19834 ^ n19833 ^ n14280 ;
  assign n19825 = n12533 ^ n11095 ^ n4333 ;
  assign n19826 = x236 & ~n19825 ;
  assign n19827 = ~n7619 & n19826 ;
  assign n19823 = n1188 & ~n13633 ;
  assign n19824 = ( n2291 & ~n19482 ) | ( n2291 & n19823 ) | ( ~n19482 & n19823 ) ;
  assign n19828 = n19827 ^ n19824 ^ x122 ;
  assign n19836 = n19835 ^ n19828 ^ n12901 ;
  assign n19837 = n19836 ^ n6828 ^ n6025 ;
  assign n19838 = ~n9654 & n17515 ;
  assign n19839 = n669 ^ x230 ^ x19 ;
  assign n19840 = n6031 | n19839 ;
  assign n19841 = ( n15431 & ~n19838 ) | ( n15431 & n19840 ) | ( ~n19838 & n19840 ) ;
  assign n19842 = ~n6221 & n19841 ;
  assign n19843 = n7257 ^ n3925 ^ n889 ;
  assign n19844 = ( n5888 & n14132 ) | ( n5888 & n19843 ) | ( n14132 & n19843 ) ;
  assign n19845 = n17613 ^ n15468 ^ n1425 ;
  assign n19846 = n3857 ^ n1733 ^ n1596 ;
  assign n19847 = n16775 ^ n5863 ^ n4061 ;
  assign n19848 = n15586 ^ n10197 ^ n8044 ;
  assign n19849 = n8096 & ~n19848 ;
  assign n19850 = ( n19846 & n19847 ) | ( n19846 & n19849 ) | ( n19847 & n19849 ) ;
  assign n19851 = ( n12090 & n19845 ) | ( n12090 & ~n19850 ) | ( n19845 & ~n19850 ) ;
  assign n19852 = n19844 & n19851 ;
  assign n19853 = ( n2239 & n9140 ) | ( n2239 & n9198 ) | ( n9140 & n9198 ) ;
  assign n19854 = ( n6600 & n6689 ) | ( n6600 & n19853 ) | ( n6689 & n19853 ) ;
  assign n19855 = ( ~n5944 & n7191 ) | ( ~n5944 & n19854 ) | ( n7191 & n19854 ) ;
  assign n19856 = n8281 ^ n6132 ^ n1740 ;
  assign n19857 = ( n9588 & ~n11786 ) | ( n9588 & n19449 ) | ( ~n11786 & n19449 ) ;
  assign n19862 = n10523 ^ n5399 ^ 1'b0 ;
  assign n19863 = n14668 & n19862 ;
  assign n19860 = ( n317 & ~n3695 ) | ( n317 & n10650 ) | ( ~n3695 & n10650 ) ;
  assign n19861 = n19860 ^ n18500 ^ n3897 ;
  assign n19858 = ( n3067 & n4886 ) | ( n3067 & n6724 ) | ( n4886 & n6724 ) ;
  assign n19859 = ~n4692 & n19858 ;
  assign n19864 = n19863 ^ n19861 ^ n19859 ;
  assign n19865 = ( n8635 & n19857 ) | ( n8635 & ~n19864 ) | ( n19857 & ~n19864 ) ;
  assign n19869 = ~n1299 & n1584 ;
  assign n19867 = ( n6263 & n8973 ) | ( n6263 & n10675 ) | ( n8973 & n10675 ) ;
  assign n19868 = ( n15100 & n18547 ) | ( n15100 & n19867 ) | ( n18547 & n19867 ) ;
  assign n19870 = n19869 ^ n19868 ^ 1'b0 ;
  assign n19871 = n4918 & n19870 ;
  assign n19866 = n4209 & ~n15818 ;
  assign n19872 = n19871 ^ n19866 ^ 1'b0 ;
  assign n19873 = ( n15933 & n17184 ) | ( n15933 & n19872 ) | ( n17184 & n19872 ) ;
  assign n19875 = ( n2773 & n13566 ) | ( n2773 & n19073 ) | ( n13566 & n19073 ) ;
  assign n19874 = ( x167 & n2796 ) | ( x167 & ~n10843 ) | ( n2796 & ~n10843 ) ;
  assign n19876 = n19875 ^ n19874 ^ n14501 ;
  assign n19877 = n9173 & n10326 ;
  assign n19878 = ( n7568 & n19876 ) | ( n7568 & ~n19877 ) | ( n19876 & ~n19877 ) ;
  assign n19879 = n15134 ^ n14968 ^ n959 ;
  assign n19880 = n10402 ^ n9050 ^ n1512 ;
  assign n19881 = ( n1247 & ~n3126 ) | ( n1247 & n19880 ) | ( ~n3126 & n19880 ) ;
  assign n19882 = ( n1485 & n2725 ) | ( n1485 & n8885 ) | ( n2725 & n8885 ) ;
  assign n19883 = ~n1963 & n10374 ;
  assign n19884 = ( n3617 & n4621 ) | ( n3617 & ~n9860 ) | ( n4621 & ~n9860 ) ;
  assign n19885 = ( n3057 & ~n4128 ) | ( n3057 & n9524 ) | ( ~n4128 & n9524 ) ;
  assign n19886 = n18679 ^ n9349 ^ n1390 ;
  assign n19887 = ( n5317 & n5784 ) | ( n5317 & n19886 ) | ( n5784 & n19886 ) ;
  assign n19888 = ( n1889 & n19307 ) | ( n1889 & n19887 ) | ( n19307 & n19887 ) ;
  assign n19889 = ( ~n2796 & n17854 ) | ( ~n2796 & n19888 ) | ( n17854 & n19888 ) ;
  assign n19890 = ( n12415 & n18469 ) | ( n12415 & n19889 ) | ( n18469 & n19889 ) ;
  assign n19891 = ( n7666 & n8053 ) | ( n7666 & ~n12304 ) | ( n8053 & ~n12304 ) ;
  assign n19892 = n19891 ^ n14948 ^ n11022 ;
  assign n19893 = n5545 ^ n2782 ^ n704 ;
  assign n19894 = n19893 ^ n19818 ^ n11970 ;
  assign n19895 = ( n16668 & ~n19892 ) | ( n16668 & n19894 ) | ( ~n19892 & n19894 ) ;
  assign n19896 = n13657 ^ n7782 ^ n5192 ;
  assign n19897 = n11811 & n12523 ;
  assign n19898 = ( ~n944 & n11038 ) | ( ~n944 & n15011 ) | ( n11038 & n15011 ) ;
  assign n19899 = ( n3564 & n13633 ) | ( n3564 & n19898 ) | ( n13633 & n19898 ) ;
  assign n19900 = n13587 ^ n12832 ^ n5965 ;
  assign n19901 = n15190 ^ n12871 ^ n11821 ;
  assign n19902 = ( n7128 & ~n19252 ) | ( n7128 & n19901 ) | ( ~n19252 & n19901 ) ;
  assign n19903 = n6596 ^ n3154 ^ x193 ;
  assign n19904 = n19903 ^ n14067 ^ n4783 ;
  assign n19905 = ( n6226 & ~n6435 ) | ( n6226 & n19904 ) | ( ~n6435 & n19904 ) ;
  assign n19906 = n1268 | n16561 ;
  assign n19907 = n15422 & n19906 ;
  assign n19908 = ( n4726 & ~n12273 ) | ( n4726 & n19907 ) | ( ~n12273 & n19907 ) ;
  assign n19911 = ( n873 & ~n2703 ) | ( n873 & n17164 ) | ( ~n2703 & n17164 ) ;
  assign n19909 = n3808 & n9557 ;
  assign n19910 = n19909 ^ n19196 ^ 1'b0 ;
  assign n19912 = n19911 ^ n19910 ^ n2542 ;
  assign n19913 = n5795 ^ n5189 ^ n2493 ;
  assign n19914 = n19913 ^ n12166 ^ 1'b0 ;
  assign n19915 = n19914 ^ n18242 ^ n13647 ;
  assign n19926 = ( ~n473 & n1278 ) | ( ~n473 & n10618 ) | ( n1278 & n10618 ) ;
  assign n19921 = ( n1102 & n2497 ) | ( n1102 & n2793 ) | ( n2497 & n2793 ) ;
  assign n19922 = ( n8298 & n8396 ) | ( n8298 & n19921 ) | ( n8396 & n19921 ) ;
  assign n19920 = ~n2717 & n18371 ;
  assign n19923 = n19922 ^ n19920 ^ 1'b0 ;
  assign n19924 = n19923 ^ n10169 ^ n2163 ;
  assign n19917 = n16909 ^ n5464 ^ n794 ;
  assign n19916 = n13736 ^ n5728 ^ n2485 ;
  assign n19918 = n19917 ^ n19916 ^ n6554 ;
  assign n19919 = n19918 ^ n15048 ^ n10289 ;
  assign n19925 = n19924 ^ n19919 ^ n12130 ;
  assign n19927 = n19926 ^ n19925 ^ n2420 ;
  assign n19928 = n14732 ^ n13449 ^ n985 ;
  assign n19929 = ( ~n3711 & n3984 ) | ( ~n3711 & n12929 ) | ( n3984 & n12929 ) ;
  assign n19930 = ( ~n14774 & n17019 ) | ( ~n14774 & n19929 ) | ( n17019 & n19929 ) ;
  assign n19931 = n19930 ^ n19898 ^ n1595 ;
  assign n19932 = n6588 ^ n828 ^ 1'b0 ;
  assign n19933 = n14672 & ~n19932 ;
  assign n19936 = n8474 | n9789 ;
  assign n19937 = n4842 | n19936 ;
  assign n19934 = ~n13644 & n16091 ;
  assign n19935 = n19934 ^ n5047 ^ 1'b0 ;
  assign n19938 = n19937 ^ n19935 ^ n6830 ;
  assign n19939 = n19938 ^ n8334 ^ n5826 ;
  assign n19940 = ( ~n2765 & n3069 ) | ( ~n2765 & n19939 ) | ( n3069 & n19939 ) ;
  assign n19942 = n16248 ^ n1111 ^ 1'b0 ;
  assign n19941 = ( ~n3175 & n17123 ) | ( ~n3175 & n17593 ) | ( n17123 & n17593 ) ;
  assign n19943 = n19942 ^ n19941 ^ n569 ;
  assign n19945 = n4678 ^ n3772 ^ n1579 ;
  assign n19946 = n12744 ^ n6264 ^ x196 ;
  assign n19947 = n19946 ^ n5798 ^ 1'b0 ;
  assign n19948 = ~n19945 & n19947 ;
  assign n19944 = ( n4426 & n5064 ) | ( n4426 & n8498 ) | ( n5064 & n8498 ) ;
  assign n19949 = n19948 ^ n19944 ^ n2402 ;
  assign n19956 = n8415 & ~n14063 ;
  assign n19950 = ( n6925 & n12644 ) | ( n6925 & n17153 ) | ( n12644 & n17153 ) ;
  assign n19951 = ( n5921 & n10740 ) | ( n5921 & ~n11388 ) | ( n10740 & ~n11388 ) ;
  assign n19952 = n3159 ^ n2430 ^ x12 ;
  assign n19953 = n7812 & ~n19952 ;
  assign n19954 = ( ~n14902 & n19951 ) | ( ~n14902 & n19953 ) | ( n19951 & n19953 ) ;
  assign n19955 = ( ~n6464 & n19950 ) | ( ~n6464 & n19954 ) | ( n19950 & n19954 ) ;
  assign n19957 = n19956 ^ n19955 ^ 1'b0 ;
  assign n19958 = ~n8707 & n19957 ;
  assign n19959 = ~n5651 & n8564 ;
  assign n19960 = n19959 ^ n15871 ^ 1'b0 ;
  assign n19961 = n12874 ^ n9294 ^ n3467 ;
  assign n19965 = ( n3382 & ~n11907 ) | ( n3382 & n17286 ) | ( ~n11907 & n17286 ) ;
  assign n19962 = ~x230 & n400 ;
  assign n19963 = n1585 | n19962 ;
  assign n19964 = n19963 ^ n5842 ^ 1'b0 ;
  assign n19966 = n19965 ^ n19964 ^ n1783 ;
  assign n19967 = ( n19960 & ~n19961 ) | ( n19960 & n19966 ) | ( ~n19961 & n19966 ) ;
  assign n19968 = n6479 ^ n2838 ^ n1267 ;
  assign n19969 = n1318 | n2925 ;
  assign n19970 = n19968 | n19969 ;
  assign n19971 = n19970 ^ n7786 ^ n3594 ;
  assign n19972 = n19971 ^ n14880 ^ 1'b0 ;
  assign n19973 = ( ~n4464 & n14682 ) | ( ~n4464 & n19972 ) | ( n14682 & n19972 ) ;
  assign n19974 = n13445 ^ x173 ^ 1'b0 ;
  assign n19975 = n12445 ^ n10116 ^ n3934 ;
  assign n19976 = n19975 ^ n17280 ^ n13710 ;
  assign n19978 = n6452 ^ n1114 ^ 1'b0 ;
  assign n19977 = n6160 | n11270 ;
  assign n19979 = n19978 ^ n19977 ^ n6198 ;
  assign n19980 = ( ~n19974 & n19976 ) | ( ~n19974 & n19979 ) | ( n19976 & n19979 ) ;
  assign n19991 = ( ~x66 & n6593 ) | ( ~x66 & n16244 ) | ( n6593 & n16244 ) ;
  assign n19989 = n8857 ^ n5893 ^ n280 ;
  assign n19987 = ( n4413 & n7886 ) | ( n4413 & ~n9483 ) | ( n7886 & ~n9483 ) ;
  assign n19988 = ( n1744 & n8566 ) | ( n1744 & ~n19987 ) | ( n8566 & ~n19987 ) ;
  assign n19986 = n16543 ^ n15306 ^ n8499 ;
  assign n19990 = n19989 ^ n19988 ^ n19986 ;
  assign n19981 = n15154 ^ n9592 ^ n2039 ;
  assign n19982 = ( ~n6382 & n10808 ) | ( ~n6382 & n19981 ) | ( n10808 & n19981 ) ;
  assign n19983 = n19982 ^ n3991 ^ n1218 ;
  assign n19984 = n19983 ^ n7404 ^ n5284 ;
  assign n19985 = n19984 ^ n12001 ^ n604 ;
  assign n19992 = n19991 ^ n19990 ^ n19985 ;
  assign n19993 = ( ~n6112 & n6643 ) | ( ~n6112 & n9926 ) | ( n6643 & n9926 ) ;
  assign n19994 = ( n904 & ~n13049 ) | ( n904 & n19993 ) | ( ~n13049 & n19993 ) ;
  assign n19995 = ( n1479 & n6485 ) | ( n1479 & n7999 ) | ( n6485 & n7999 ) ;
  assign n19996 = n19995 ^ n2420 ^ n1874 ;
  assign n19997 = ( n1950 & n4565 ) | ( n1950 & n19996 ) | ( n4565 & n19996 ) ;
  assign n19998 = n19997 ^ n10049 ^ n7593 ;
  assign n19999 = ( n897 & ~n6576 ) | ( n897 & n14927 ) | ( ~n6576 & n14927 ) ;
  assign n20001 = ( ~n1572 & n3177 ) | ( ~n1572 & n3601 ) | ( n3177 & n3601 ) ;
  assign n20002 = n12797 ^ n11006 ^ n2181 ;
  assign n20003 = n2200 & ~n2675 ;
  assign n20004 = n20003 ^ n10862 ^ n3339 ;
  assign n20005 = n20004 ^ n10322 ^ 1'b0 ;
  assign n20006 = n17530 | n20005 ;
  assign n20007 = ( n8577 & ~n15911 ) | ( n8577 & n20006 ) | ( ~n15911 & n20006 ) ;
  assign n20008 = ( n8500 & n19649 ) | ( n8500 & n20007 ) | ( n19649 & n20007 ) ;
  assign n20009 = ( n14616 & n20002 ) | ( n14616 & ~n20008 ) | ( n20002 & ~n20008 ) ;
  assign n20010 = n14949 | n20009 ;
  assign n20011 = n20001 | n20010 ;
  assign n20000 = n12103 ^ n1229 ^ n744 ;
  assign n20012 = n20011 ^ n20000 ^ n16082 ;
  assign n20015 = n10158 ^ n4481 ^ 1'b0 ;
  assign n20014 = n12222 ^ n11032 ^ n9850 ;
  assign n20013 = n9041 | n15790 ;
  assign n20016 = n20015 ^ n20014 ^ n20013 ;
  assign n20017 = ( n4611 & ~n19522 ) | ( n4611 & n20016 ) | ( ~n19522 & n20016 ) ;
  assign n20018 = n11965 ^ n3273 ^ 1'b0 ;
  assign n20020 = ( ~n3879 & n6011 ) | ( ~n3879 & n10461 ) | ( n6011 & n10461 ) ;
  assign n20021 = n20020 ^ n7344 ^ n2854 ;
  assign n20019 = n4232 | n8072 ;
  assign n20022 = n20021 ^ n20019 ^ 1'b0 ;
  assign n20023 = ( n3816 & n20018 ) | ( n3816 & ~n20022 ) | ( n20018 & ~n20022 ) ;
  assign n20024 = n7115 & n8286 ;
  assign n20025 = ( n9759 & n14937 ) | ( n9759 & ~n20024 ) | ( n14937 & ~n20024 ) ;
  assign n20035 = ( ~x172 & n4226 ) | ( ~x172 & n5555 ) | ( n4226 & n5555 ) ;
  assign n20031 = ( n394 & ~n4295 ) | ( n394 & n6488 ) | ( ~n4295 & n6488 ) ;
  assign n20032 = n9365 & n20031 ;
  assign n20033 = n9485 & n20032 ;
  assign n20026 = ( n483 & n804 ) | ( n483 & n846 ) | ( n804 & n846 ) ;
  assign n20027 = n20026 ^ n7609 ^ n3401 ;
  assign n20028 = ( n2915 & n4585 ) | ( n2915 & ~n5494 ) | ( n4585 & ~n5494 ) ;
  assign n20029 = ( n1443 & n14553 ) | ( n1443 & n20028 ) | ( n14553 & n20028 ) ;
  assign n20030 = ( n3798 & ~n20027 ) | ( n3798 & n20029 ) | ( ~n20027 & n20029 ) ;
  assign n20034 = n20033 ^ n20030 ^ n17545 ;
  assign n20036 = n20035 ^ n20034 ^ n3106 ;
  assign n20037 = n18237 ^ n12884 ^ n3531 ;
  assign n20038 = ( n578 & n7114 ) | ( n578 & ~n20037 ) | ( n7114 & ~n20037 ) ;
  assign n20039 = n20038 ^ n2086 ^ 1'b0 ;
  assign n20040 = n7857 ^ n1509 ^ n278 ;
  assign n20041 = ( ~n11167 & n20039 ) | ( ~n11167 & n20040 ) | ( n20039 & n20040 ) ;
  assign n20042 = n7740 & ~n20041 ;
  assign n20043 = n20042 ^ n2408 ^ 1'b0 ;
  assign n20044 = ( n552 & n3849 ) | ( n552 & ~n6234 ) | ( n3849 & ~n6234 ) ;
  assign n20045 = n20044 ^ n8115 ^ n617 ;
  assign n20046 = n17122 ^ n15302 ^ n1052 ;
  assign n20047 = ( n19454 & n20045 ) | ( n19454 & n20046 ) | ( n20045 & n20046 ) ;
  assign n20048 = n20043 & ~n20047 ;
  assign n20049 = ~n18837 & n20048 ;
  assign n20054 = ( n497 & ~n3504 ) | ( n497 & n16963 ) | ( ~n3504 & n16963 ) ;
  assign n20055 = n20054 ^ n15552 ^ n1235 ;
  assign n20052 = n14803 ^ n13181 ^ n504 ;
  assign n20051 = ~n5067 & n17048 ;
  assign n20053 = n20052 ^ n20051 ^ 1'b0 ;
  assign n20050 = n18486 ^ n13575 ^ n13215 ;
  assign n20056 = n20055 ^ n20053 ^ n20050 ;
  assign n20057 = ( ~n1277 & n8547 ) | ( ~n1277 & n9129 ) | ( n8547 & n9129 ) ;
  assign n20058 = ( n6218 & n6516 ) | ( n6218 & ~n20057 ) | ( n6516 & ~n20057 ) ;
  assign n20059 = n15064 ^ n13943 ^ n4085 ;
  assign n20060 = n20059 ^ n15373 ^ n2019 ;
  assign n20061 = ( n400 & n16332 ) | ( n400 & n20060 ) | ( n16332 & n20060 ) ;
  assign n20062 = ~n1504 & n11244 ;
  assign n20063 = ( ~n7981 & n14387 ) | ( ~n7981 & n20062 ) | ( n14387 & n20062 ) ;
  assign n20064 = ( n262 & ~n20061 ) | ( n262 & n20063 ) | ( ~n20061 & n20063 ) ;
  assign n20065 = n16115 ^ n5977 ^ n5719 ;
  assign n20066 = n19735 ^ n17322 ^ 1'b0 ;
  assign n20067 = n18235 & n20066 ;
  assign n20068 = n3964 | n6999 ;
  assign n20069 = n20068 ^ n4585 ^ 1'b0 ;
  assign n20070 = n12385 ^ n11897 ^ n1167 ;
  assign n20071 = n548 | n20070 ;
  assign n20072 = n20071 ^ n8968 ^ n4935 ;
  assign n20073 = ( n1806 & ~n20069 ) | ( n1806 & n20072 ) | ( ~n20069 & n20072 ) ;
  assign n20074 = n20073 ^ n11820 ^ n9653 ;
  assign n20076 = ( ~n9701 & n13292 ) | ( ~n9701 & n19075 ) | ( n13292 & n19075 ) ;
  assign n20075 = n13665 ^ n11281 ^ n7164 ;
  assign n20077 = n20076 ^ n20075 ^ n5833 ;
  assign n20078 = ( ~n938 & n8913 ) | ( ~n938 & n16369 ) | ( n8913 & n16369 ) ;
  assign n20079 = n16971 ^ n9169 ^ n7077 ;
  assign n20080 = ( n1956 & n6910 ) | ( n1956 & n20079 ) | ( n6910 & n20079 ) ;
  assign n20081 = n3654 & n5297 ;
  assign n20082 = n20081 ^ n7837 ^ 1'b0 ;
  assign n20083 = n6369 ^ n6052 ^ 1'b0 ;
  assign n20084 = ~n7381 & n20083 ;
  assign n20085 = n20084 ^ n11345 ^ 1'b0 ;
  assign n20086 = x171 & n20085 ;
  assign n20087 = n13067 ^ n9567 ^ 1'b0 ;
  assign n20088 = n20086 & n20087 ;
  assign n20089 = ( n809 & n20082 ) | ( n809 & ~n20088 ) | ( n20082 & ~n20088 ) ;
  assign n20091 = ( n9409 & n16423 ) | ( n9409 & ~n18454 ) | ( n16423 & ~n18454 ) ;
  assign n20090 = n19880 ^ n2065 ^ n742 ;
  assign n20092 = n20091 ^ n20090 ^ n12862 ;
  assign n20093 = n20092 ^ n9156 ^ n3337 ;
  assign n20106 = n14014 ^ n11291 ^ n998 ;
  assign n20107 = n1290 | n4667 ;
  assign n20108 = n20107 ^ n18040 ^ 1'b0 ;
  assign n20109 = ( n10330 & n20106 ) | ( n10330 & n20108 ) | ( n20106 & n20108 ) ;
  assign n20103 = n7897 ^ n2066 ^ x217 ;
  assign n20102 = n14376 ^ n5037 ^ 1'b0 ;
  assign n20099 = ( n506 & n11785 ) | ( n506 & n13742 ) | ( n11785 & n13742 ) ;
  assign n20100 = n16335 & ~n20099 ;
  assign n20101 = ~n9350 & n20100 ;
  assign n20104 = n20103 ^ n20102 ^ n20101 ;
  assign n20094 = n3592 ^ n2358 ^ n1396 ;
  assign n20095 = ( ~n1193 & n5427 ) | ( ~n1193 & n14262 ) | ( n5427 & n14262 ) ;
  assign n20096 = n20094 & ~n20095 ;
  assign n20097 = n20096 ^ n14310 ^ 1'b0 ;
  assign n20098 = ( n13298 & n16917 ) | ( n13298 & n20097 ) | ( n16917 & n20097 ) ;
  assign n20105 = n20104 ^ n20098 ^ n7483 ;
  assign n20110 = n20109 ^ n20105 ^ n13649 ;
  assign n20111 = ( n1006 & n9560 ) | ( n1006 & ~n18973 ) | ( n9560 & ~n18973 ) ;
  assign n20112 = n19483 ^ n13345 ^ n11013 ;
  assign n20113 = ( n5429 & ~n18829 ) | ( n5429 & n19545 ) | ( ~n18829 & n19545 ) ;
  assign n20114 = ( n6982 & n20112 ) | ( n6982 & ~n20113 ) | ( n20112 & ~n20113 ) ;
  assign n20115 = ( ~n6414 & n20111 ) | ( ~n6414 & n20114 ) | ( n20111 & n20114 ) ;
  assign n20116 = ~n2770 & n5036 ;
  assign n20117 = n20116 ^ n2930 ^ 1'b0 ;
  assign n20118 = ( n12120 & ~n15275 ) | ( n12120 & n20117 ) | ( ~n15275 & n20117 ) ;
  assign n20119 = ~n4610 & n15127 ;
  assign n20120 = ~n9539 & n20119 ;
  assign n20121 = n18131 & ~n20120 ;
  assign n20122 = ~n20118 & n20121 ;
  assign n20123 = n4538 & ~n20122 ;
  assign n20124 = n20123 ^ n17874 ^ 1'b0 ;
  assign n20125 = n16249 ^ n12783 ^ n5814 ;
  assign n20126 = n20125 ^ n15965 ^ n11794 ;
  assign n20127 = ( n8347 & ~n20124 ) | ( n8347 & n20126 ) | ( ~n20124 & n20126 ) ;
  assign n20128 = ( n6128 & ~n6768 ) | ( n6128 & n17707 ) | ( ~n6768 & n17707 ) ;
  assign n20129 = n20128 ^ n16295 ^ n2122 ;
  assign n20130 = ( n1123 & n2890 ) | ( n1123 & ~n13848 ) | ( n2890 & ~n13848 ) ;
  assign n20131 = n8276 & ~n20130 ;
  assign n20132 = n20131 ^ n16102 ^ 1'b0 ;
  assign n20133 = ( n925 & n3331 ) | ( n925 & ~n4645 ) | ( n3331 & ~n4645 ) ;
  assign n20134 = n20133 ^ n15196 ^ n6102 ;
  assign n20137 = n5764 & n9473 ;
  assign n20138 = n20137 ^ n4430 ^ 1'b0 ;
  assign n20135 = n12642 & ~n18612 ;
  assign n20136 = n20135 ^ n2881 ^ 1'b0 ;
  assign n20139 = n20138 ^ n20136 ^ n15779 ;
  assign n20140 = ( n1647 & ~n7848 ) | ( n1647 & n9961 ) | ( ~n7848 & n9961 ) ;
  assign n20141 = n6808 ^ n6039 ^ x147 ;
  assign n20142 = ( n12375 & n20140 ) | ( n12375 & ~n20141 ) | ( n20140 & ~n20141 ) ;
  assign n20143 = n5340 ^ n3654 ^ n1267 ;
  assign n20144 = n20143 ^ n1793 ^ 1'b0 ;
  assign n20145 = n20144 ^ n6131 ^ 1'b0 ;
  assign n20146 = ( n2159 & n10976 ) | ( n2159 & n20145 ) | ( n10976 & n20145 ) ;
  assign n20147 = n3376 & ~n4922 ;
  assign n20149 = n873 | n1218 ;
  assign n20150 = n9362 | n20149 ;
  assign n20151 = ( n4224 & n7933 ) | ( n4224 & ~n20150 ) | ( n7933 & ~n20150 ) ;
  assign n20152 = n13447 & ~n20151 ;
  assign n20148 = n18235 ^ n11163 ^ n8749 ;
  assign n20153 = n20152 ^ n20148 ^ n9950 ;
  assign n20154 = n6922 ^ n961 ^ x252 ;
  assign n20155 = ( n7466 & n14984 ) | ( n7466 & n20154 ) | ( n14984 & n20154 ) ;
  assign n20157 = ( n6313 & n7585 ) | ( n6313 & n7997 ) | ( n7585 & n7997 ) ;
  assign n20156 = ( n885 & n7205 ) | ( n885 & ~n9155 ) | ( n7205 & ~n9155 ) ;
  assign n20158 = n20157 ^ n20156 ^ 1'b0 ;
  assign n20159 = n6104 & n20158 ;
  assign n20160 = n13775 ^ n6096 ^ n2505 ;
  assign n20161 = n20160 ^ n2064 ^ 1'b0 ;
  assign n20162 = ( ~n5392 & n8279 ) | ( ~n5392 & n11981 ) | ( n8279 & n11981 ) ;
  assign n20166 = ( n1089 & n2585 ) | ( n1089 & n5184 ) | ( n2585 & n5184 ) ;
  assign n20167 = ( n1766 & ~n3448 ) | ( n1766 & n20166 ) | ( ~n3448 & n20166 ) ;
  assign n20163 = n13973 ^ n5073 ^ n1033 ;
  assign n20164 = n464 & n20163 ;
  assign n20165 = n20164 ^ n14611 ^ 1'b0 ;
  assign n20168 = n20167 ^ n20165 ^ n13714 ;
  assign n20169 = ( n4746 & ~n20162 ) | ( n4746 & n20168 ) | ( ~n20162 & n20168 ) ;
  assign n20170 = n1571 & ~n6793 ;
  assign n20171 = ~n4127 & n20170 ;
  assign n20172 = n10915 & ~n20171 ;
  assign n20173 = ( n583 & n1494 ) | ( n583 & n20172 ) | ( n1494 & n20172 ) ;
  assign n20174 = ( n2600 & n3522 ) | ( n2600 & ~n12036 ) | ( n3522 & ~n12036 ) ;
  assign n20176 = ( n14769 & n16950 ) | ( n14769 & n19971 ) | ( n16950 & n19971 ) ;
  assign n20175 = n4391 & ~n12281 ;
  assign n20177 = n20176 ^ n20175 ^ 1'b0 ;
  assign n20178 = n20177 ^ n3570 ^ 1'b0 ;
  assign n20179 = n13792 ^ n12832 ^ 1'b0 ;
  assign n20183 = ( n1085 & n7540 ) | ( n1085 & n11802 ) | ( n7540 & n11802 ) ;
  assign n20180 = n9537 & n17900 ;
  assign n20181 = n5237 ^ n5225 ^ n463 ;
  assign n20182 = ( ~n9028 & n20180 ) | ( ~n9028 & n20181 ) | ( n20180 & n20181 ) ;
  assign n20184 = n20183 ^ n20182 ^ n9351 ;
  assign n20185 = n20184 ^ n1842 ^ n413 ;
  assign n20186 = n6311 | n9447 ;
  assign n20187 = n20186 ^ n8337 ^ 1'b0 ;
  assign n20188 = n1787 & ~n20187 ;
  assign n20189 = n13086 ^ n3035 ^ n2549 ;
  assign n20190 = n20188 & n20189 ;
  assign n20191 = n6914 & n20190 ;
  assign n20193 = n10063 | n12483 ;
  assign n20194 = n20193 ^ n7808 ^ 1'b0 ;
  assign n20195 = ~n7006 & n20194 ;
  assign n20196 = n20195 ^ n758 ^ 1'b0 ;
  assign n20192 = ( n1676 & n7882 ) | ( n1676 & n13207 ) | ( n7882 & n13207 ) ;
  assign n20197 = n20196 ^ n20192 ^ n14764 ;
  assign n20198 = ( n3639 & ~n10350 ) | ( n3639 & n16451 ) | ( ~n10350 & n16451 ) ;
  assign n20199 = n20198 ^ n12890 ^ 1'b0 ;
  assign n20203 = n7486 ^ n4503 ^ 1'b0 ;
  assign n20204 = ~n14731 & n20203 ;
  assign n20200 = ( n2742 & ~n2884 ) | ( n2742 & n5330 ) | ( ~n2884 & n5330 ) ;
  assign n20201 = n3186 ^ n3148 ^ n473 ;
  assign n20202 = ( n10195 & n20200 ) | ( n10195 & ~n20201 ) | ( n20200 & ~n20201 ) ;
  assign n20205 = n20204 ^ n20202 ^ n6879 ;
  assign n20206 = n11653 ^ n6545 ^ n2183 ;
  assign n20207 = n11725 ^ n3274 ^ n3157 ;
  assign n20208 = n8516 ^ n6800 ^ 1'b0 ;
  assign n20209 = n20207 | n20208 ;
  assign n20210 = n20209 ^ n12283 ^ 1'b0 ;
  assign n20211 = ( ~n9399 & n20206 ) | ( ~n9399 & n20210 ) | ( n20206 & n20210 ) ;
  assign n20213 = n903 | n1443 ;
  assign n20214 = n20213 ^ n5670 ^ 1'b0 ;
  assign n20212 = n20027 ^ n3405 ^ x13 ;
  assign n20215 = n20214 ^ n20212 ^ 1'b0 ;
  assign n20217 = ( n2774 & n4082 ) | ( n2774 & n7584 ) | ( n4082 & n7584 ) ;
  assign n20216 = n14510 ^ n5927 ^ 1'b0 ;
  assign n20218 = n20217 ^ n20216 ^ n2934 ;
  assign n20219 = ~n755 & n5545 ;
  assign n20220 = n20219 ^ n4578 ^ 1'b0 ;
  assign n20221 = ( ~n8369 & n17639 ) | ( ~n8369 & n20220 ) | ( n17639 & n20220 ) ;
  assign n20223 = n11614 ^ n6081 ^ n4985 ;
  assign n20222 = n9963 ^ n8951 ^ n4673 ;
  assign n20224 = n20223 ^ n20222 ^ n8976 ;
  assign n20226 = n4677 ^ n1394 ^ 1'b0 ;
  assign n20227 = n969 & ~n20226 ;
  assign n20228 = n20227 ^ n465 ^ 1'b0 ;
  assign n20225 = n4363 & n20091 ;
  assign n20229 = n20228 ^ n20225 ^ 1'b0 ;
  assign n20230 = n20229 ^ n5472 ^ n4685 ;
  assign n20231 = ( n2218 & ~n7698 ) | ( n2218 & n8300 ) | ( ~n7698 & n8300 ) ;
  assign n20234 = n10770 ^ n9263 ^ n2029 ;
  assign n20235 = ( n10294 & n15877 ) | ( n10294 & ~n20234 ) | ( n15877 & ~n20234 ) ;
  assign n20236 = n20235 ^ n8199 ^ n6301 ;
  assign n20232 = n8725 & n9289 ;
  assign n20233 = n20232 ^ n13639 ^ n1902 ;
  assign n20237 = n20236 ^ n20233 ^ n11462 ;
  assign n20238 = ( ~n645 & n11263 ) | ( ~n645 & n14026 ) | ( n11263 & n14026 ) ;
  assign n20239 = ( n9017 & n18656 ) | ( n9017 & ~n20238 ) | ( n18656 & ~n20238 ) ;
  assign n20240 = ( n2788 & ~n3815 ) | ( n2788 & n8404 ) | ( ~n3815 & n8404 ) ;
  assign n20241 = ( n6580 & n16284 ) | ( n6580 & ~n20240 ) | ( n16284 & ~n20240 ) ;
  assign n20242 = n18115 ^ n3268 ^ 1'b0 ;
  assign n20243 = n20241 & n20242 ;
  assign n20244 = n20243 ^ n14436 ^ 1'b0 ;
  assign n20245 = n16268 & ~n20244 ;
  assign n20246 = ( n7723 & n13082 ) | ( n7723 & n19791 ) | ( n13082 & n19791 ) ;
  assign n20247 = ( n855 & n3203 ) | ( n855 & ~n3230 ) | ( n3203 & ~n3230 ) ;
  assign n20248 = ( n10791 & n13157 ) | ( n10791 & ~n20247 ) | ( n13157 & ~n20247 ) ;
  assign n20249 = n20248 ^ n13393 ^ n9845 ;
  assign n20250 = n6142 & n20249 ;
  assign n20251 = n15028 ^ n3034 ^ n2091 ;
  assign n20252 = n14558 ^ n8689 ^ n863 ;
  assign n20253 = ( n15135 & n18390 ) | ( n15135 & n20252 ) | ( n18390 & n20252 ) ;
  assign n20254 = n20253 ^ n304 ^ x39 ;
  assign n20255 = ( ~n10203 & n20251 ) | ( ~n10203 & n20254 ) | ( n20251 & n20254 ) ;
  assign n20256 = ~n2280 & n5807 ;
  assign n20257 = n20256 ^ n6124 ^ 1'b0 ;
  assign n20258 = ~n3500 & n11187 ;
  assign n20259 = n14339 & n20258 ;
  assign n20260 = ( n557 & n20257 ) | ( n557 & ~n20259 ) | ( n20257 & ~n20259 ) ;
  assign n20261 = n3686 & n3783 ;
  assign n20262 = n8320 & ~n20261 ;
  assign n20263 = ( n4218 & ~n10719 ) | ( n4218 & n12268 ) | ( ~n10719 & n12268 ) ;
  assign n20264 = ( n2760 & ~n5098 ) | ( n2760 & n20263 ) | ( ~n5098 & n20263 ) ;
  assign n20265 = n1947 & ~n20264 ;
  assign n20266 = n3022 | n4424 ;
  assign n20267 = n20266 ^ n12517 ^ n9325 ;
  assign n20268 = n2380 ^ n1766 ^ n855 ;
  assign n20269 = ( ~n1668 & n4373 ) | ( ~n1668 & n20268 ) | ( n4373 & n20268 ) ;
  assign n20270 = ( n7780 & n9898 ) | ( n7780 & ~n20269 ) | ( n9898 & ~n20269 ) ;
  assign n20271 = n20270 ^ n2994 ^ 1'b0 ;
  assign n20272 = n10363 ^ n6484 ^ n996 ;
  assign n20273 = n20272 ^ n7657 ^ n1613 ;
  assign n20274 = n20273 ^ n12743 ^ n4683 ;
  assign n20275 = ( n8104 & n17574 ) | ( n8104 & n20274 ) | ( n17574 & n20274 ) ;
  assign n20276 = ( n3214 & n20271 ) | ( n3214 & n20275 ) | ( n20271 & n20275 ) ;
  assign n20277 = ( ~n11559 & n20267 ) | ( ~n11559 & n20276 ) | ( n20267 & n20276 ) ;
  assign n20278 = ( n1256 & n5703 ) | ( n1256 & ~n10304 ) | ( n5703 & ~n10304 ) ;
  assign n20279 = n20278 ^ n12980 ^ 1'b0 ;
  assign n20280 = ( x67 & n5183 ) | ( x67 & n9703 ) | ( n5183 & n9703 ) ;
  assign n20281 = n9204 ^ n5794 ^ n4149 ;
  assign n20282 = n20281 ^ n14321 ^ x94 ;
  assign n20283 = ( n4839 & n20280 ) | ( n4839 & ~n20282 ) | ( n20280 & ~n20282 ) ;
  assign n20284 = n1719 | n6807 ;
  assign n20285 = n1941 | n20284 ;
  assign n20286 = n11144 ^ n11068 ^ n4493 ;
  assign n20287 = n19991 & ~n20286 ;
  assign n20288 = ( x105 & n4610 ) | ( x105 & ~n13507 ) | ( n4610 & ~n13507 ) ;
  assign n20289 = ( n2623 & n15221 ) | ( n2623 & ~n20288 ) | ( n15221 & ~n20288 ) ;
  assign n20290 = n2043 & n20289 ;
  assign n20291 = ( ~n10406 & n11912 ) | ( ~n10406 & n14335 ) | ( n11912 & n14335 ) ;
  assign n20292 = n15380 ^ n7602 ^ 1'b0 ;
  assign n20298 = n17060 ^ n13636 ^ n9720 ;
  assign n20296 = n8356 & n14259 ;
  assign n20297 = n20296 ^ n805 ^ 1'b0 ;
  assign n20293 = n7499 ^ n3053 ^ n569 ;
  assign n20294 = n7316 | n12833 ;
  assign n20295 = n20293 | n20294 ;
  assign n20299 = n20298 ^ n20297 ^ n20295 ;
  assign n20300 = ( n20291 & n20292 ) | ( n20291 & n20299 ) | ( n20292 & n20299 ) ;
  assign n20301 = ( n13519 & n20290 ) | ( n13519 & ~n20300 ) | ( n20290 & ~n20300 ) ;
  assign n20302 = n18149 ^ n13816 ^ n12767 ;
  assign n20303 = ( n1482 & n7832 ) | ( n1482 & ~n20302 ) | ( n7832 & ~n20302 ) ;
  assign n20304 = n17407 ^ n13159 ^ 1'b0 ;
  assign n20305 = x186 & n20304 ;
  assign n20306 = n20305 ^ n11832 ^ n9641 ;
  assign n20310 = ( n2375 & n12116 ) | ( n2375 & ~n17026 ) | ( n12116 & ~n17026 ) ;
  assign n20311 = n20310 ^ n6223 ^ 1'b0 ;
  assign n20312 = n4529 | n20311 ;
  assign n20308 = ( n4234 & n4286 ) | ( n4234 & ~n5595 ) | ( n4286 & ~n5595 ) ;
  assign n20307 = n8676 ^ n6613 ^ n4949 ;
  assign n20309 = n20308 ^ n20307 ^ n15119 ;
  assign n20313 = n20312 ^ n20309 ^ n13926 ;
  assign n20314 = ( ~n3262 & n16022 ) | ( ~n3262 & n19398 ) | ( n16022 & n19398 ) ;
  assign n20315 = n18829 ^ n2543 ^ n1623 ;
  assign n20316 = n20315 ^ n8914 ^ n2760 ;
  assign n20317 = ( ~n9361 & n20314 ) | ( ~n9361 & n20316 ) | ( n20314 & n20316 ) ;
  assign n20318 = ( ~n653 & n5310 ) | ( ~n653 & n14599 ) | ( n5310 & n14599 ) ;
  assign n20319 = n19846 ^ n17723 ^ n1235 ;
  assign n20320 = ~n13853 & n20319 ;
  assign n20321 = n20320 ^ n7460 ^ 1'b0 ;
  assign n20322 = n6700 ^ n3631 ^ 1'b0 ;
  assign n20323 = ~n6091 & n20322 ;
  assign n20324 = n20323 ^ n7991 ^ n2752 ;
  assign n20325 = n20324 ^ n14933 ^ n1689 ;
  assign n20326 = ( n3186 & n7489 ) | ( n3186 & n13351 ) | ( n7489 & n13351 ) ;
  assign n20327 = ( n15435 & n20325 ) | ( n15435 & n20326 ) | ( n20325 & n20326 ) ;
  assign n20328 = ( ~n9646 & n17390 ) | ( ~n9646 & n20327 ) | ( n17390 & n20327 ) ;
  assign n20329 = ( ~n524 & n6665 ) | ( ~n524 & n6938 ) | ( n6665 & n6938 ) ;
  assign n20330 = ( n11144 & n14022 ) | ( n11144 & ~n20329 ) | ( n14022 & ~n20329 ) ;
  assign n20331 = n20330 ^ n12782 ^ n5303 ;
  assign n20332 = ( ~n2752 & n5496 ) | ( ~n2752 & n5618 ) | ( n5496 & n5618 ) ;
  assign n20333 = n8444 ^ n3586 ^ 1'b0 ;
  assign n20334 = n14113 & ~n20333 ;
  assign n20335 = ( n3018 & n20332 ) | ( n3018 & n20334 ) | ( n20332 & n20334 ) ;
  assign n20336 = n16235 ^ n7578 ^ n4988 ;
  assign n20337 = n8204 ^ n3484 ^ n2454 ;
  assign n20338 = ( n6594 & n9279 ) | ( n6594 & n16770 ) | ( n9279 & n16770 ) ;
  assign n20345 = n14739 ^ n2039 ^ n606 ;
  assign n20346 = ( n8500 & n9428 ) | ( n8500 & ~n10162 ) | ( n9428 & ~n10162 ) ;
  assign n20347 = ( n18642 & n20345 ) | ( n18642 & n20346 ) | ( n20345 & n20346 ) ;
  assign n20343 = n19179 ^ n504 ^ 1'b0 ;
  assign n20341 = ( n2305 & n6142 ) | ( n2305 & ~n8951 ) | ( n6142 & ~n8951 ) ;
  assign n20339 = n15674 ^ n5710 ^ n3170 ;
  assign n20340 = ( ~n7884 & n10882 ) | ( ~n7884 & n20339 ) | ( n10882 & n20339 ) ;
  assign n20342 = n20341 ^ n20340 ^ 1'b0 ;
  assign n20344 = n20343 ^ n20342 ^ n19906 ;
  assign n20348 = n20347 ^ n20344 ^ n7469 ;
  assign n20353 = ( ~n4576 & n13851 ) | ( ~n4576 & n20165 ) | ( n13851 & n20165 ) ;
  assign n20352 = n15900 ^ n11015 ^ n5913 ;
  assign n20354 = n20353 ^ n20352 ^ n12697 ;
  assign n20349 = ( ~n5896 & n7067 ) | ( ~n5896 & n10744 ) | ( n7067 & n10744 ) ;
  assign n20350 = ( n8109 & n12657 ) | ( n8109 & ~n20349 ) | ( n12657 & ~n20349 ) ;
  assign n20351 = ( n9183 & n14293 ) | ( n9183 & n20350 ) | ( n14293 & n20350 ) ;
  assign n20355 = n20354 ^ n20351 ^ n1423 ;
  assign n20356 = n15180 ^ n6176 ^ n1240 ;
  assign n20357 = n8471 & ~n13439 ;
  assign n20358 = n20357 ^ n9014 ^ 1'b0 ;
  assign n20359 = n16644 ^ n291 ^ 1'b0 ;
  assign n20360 = n16895 ^ n9227 ^ n8102 ;
  assign n20361 = n20360 ^ n12862 ^ n7685 ;
  assign n20362 = n20361 ^ n5892 ^ n4989 ;
  assign n20365 = ( ~n7626 & n12717 ) | ( ~n7626 & n15506 ) | ( n12717 & n15506 ) ;
  assign n20363 = ( n3103 & n7007 ) | ( n3103 & ~n11300 ) | ( n7007 & ~n11300 ) ;
  assign n20364 = n20363 ^ n17356 ^ n1377 ;
  assign n20366 = n20365 ^ n20364 ^ n15600 ;
  assign n20367 = ( n419 & n2064 ) | ( n419 & n9829 ) | ( n2064 & n9829 ) ;
  assign n20368 = ~n7974 & n20367 ;
  assign n20369 = n13427 & n20368 ;
  assign n20370 = ( ~n644 & n3712 ) | ( ~n644 & n20369 ) | ( n3712 & n20369 ) ;
  assign n20371 = n20370 ^ n15284 ^ n7308 ;
  assign n20372 = n17369 ^ n8861 ^ n5536 ;
  assign n20381 = n3386 ^ n818 ^ n411 ;
  assign n20377 = ( ~n853 & n4198 ) | ( ~n853 & n11198 ) | ( n4198 & n11198 ) ;
  assign n20378 = n14859 ^ n8622 ^ n2523 ;
  assign n20379 = ( n4299 & n20377 ) | ( n4299 & ~n20378 ) | ( n20377 & ~n20378 ) ;
  assign n20373 = n19329 ^ n4811 ^ 1'b0 ;
  assign n20374 = ( n1167 & n14044 ) | ( n1167 & ~n20373 ) | ( n14044 & ~n20373 ) ;
  assign n20375 = ( ~n13409 & n19769 ) | ( ~n13409 & n20374 ) | ( n19769 & n20374 ) ;
  assign n20376 = n20375 ^ n15366 ^ 1'b0 ;
  assign n20380 = n20379 ^ n20376 ^ n17530 ;
  assign n20382 = n20381 ^ n20380 ^ n10774 ;
  assign n20383 = n17497 ^ n13394 ^ n8777 ;
  assign n20384 = n13768 ^ n9318 ^ n2029 ;
  assign n20385 = n20384 ^ n15597 ^ n1207 ;
  assign n20386 = ( ~n1387 & n8309 ) | ( ~n1387 & n14229 ) | ( n8309 & n14229 ) ;
  assign n20387 = n3169 ^ n2817 ^ 1'b0 ;
  assign n20388 = n15219 & ~n20387 ;
  assign n20389 = n20388 ^ n12530 ^ 1'b0 ;
  assign n20390 = n7862 & n11063 ;
  assign n20391 = n15929 ^ n4831 ^ 1'b0 ;
  assign n20392 = ( n10953 & n12896 ) | ( n10953 & ~n20391 ) | ( n12896 & ~n20391 ) ;
  assign n20393 = n17877 ^ n11871 ^ n11646 ;
  assign n20394 = n17651 ^ n6661 ^ 1'b0 ;
  assign n20395 = n15903 | n20394 ;
  assign n20396 = n20395 ^ n19408 ^ 1'b0 ;
  assign n20397 = n16845 ^ n11563 ^ 1'b0 ;
  assign n20398 = ( n555 & n9983 ) | ( n555 & n20397 ) | ( n9983 & n20397 ) ;
  assign n20399 = n3076 | n20398 ;
  assign n20402 = n312 & n362 ;
  assign n20403 = n20402 ^ n3787 ^ n1526 ;
  assign n20400 = ( n2389 & ~n4593 ) | ( n2389 & n10345 ) | ( ~n4593 & n10345 ) ;
  assign n20401 = n20400 ^ n5794 ^ n2493 ;
  assign n20404 = n20403 ^ n20401 ^ n5376 ;
  assign n20405 = n14516 ^ n5510 ^ n5259 ;
  assign n20406 = n20405 ^ n11845 ^ n9343 ;
  assign n20407 = ( n4775 & n12403 ) | ( n4775 & n13020 ) | ( n12403 & n13020 ) ;
  assign n20408 = n20407 ^ n16142 ^ n10646 ;
  assign n20409 = ( ~n2620 & n5088 ) | ( ~n2620 & n5863 ) | ( n5088 & n5863 ) ;
  assign n20410 = n20409 ^ n17678 ^ n4002 ;
  assign n20411 = n20410 ^ n18085 ^ n12973 ;
  assign n20412 = n4291 ^ n4258 ^ n2262 ;
  assign n20413 = ( n2420 & n11839 ) | ( n2420 & ~n20412 ) | ( n11839 & ~n20412 ) ;
  assign n20414 = n16427 ^ n13600 ^ n10391 ;
  assign n20419 = n7357 ^ n3560 ^ n1083 ;
  assign n20417 = n10702 ^ n3657 ^ n2521 ;
  assign n20418 = n20417 ^ n2408 ^ n2156 ;
  assign n20420 = n20419 ^ n20418 ^ n18504 ;
  assign n20415 = n13058 ^ n4045 ^ 1'b0 ;
  assign n20416 = n20415 ^ n4918 ^ 1'b0 ;
  assign n20421 = n20420 ^ n20416 ^ n10502 ;
  assign n20422 = ( n1049 & ~n20414 ) | ( n1049 & n20421 ) | ( ~n20414 & n20421 ) ;
  assign n20427 = n5847 ^ n3034 ^ x30 ;
  assign n20426 = ( n1777 & n18257 ) | ( n1777 & ~n19874 ) | ( n18257 & ~n19874 ) ;
  assign n20423 = n1397 | n3703 ;
  assign n20424 = n16336 & ~n20423 ;
  assign n20425 = ( n7129 & n10724 ) | ( n7129 & n20424 ) | ( n10724 & n20424 ) ;
  assign n20428 = n20427 ^ n20426 ^ n20425 ;
  assign n20429 = ( ~n5958 & n8372 ) | ( ~n5958 & n14945 ) | ( n8372 & n14945 ) ;
  assign n20430 = n20429 ^ n19386 ^ 1'b0 ;
  assign n20434 = n15177 ^ n7111 ^ n699 ;
  assign n20431 = n13507 ^ n5307 ^ n628 ;
  assign n20432 = ( n11517 & ~n13361 ) | ( n11517 & n20431 ) | ( ~n13361 & n20431 ) ;
  assign n20433 = ( ~n632 & n8172 ) | ( ~n632 & n20432 ) | ( n8172 & n20432 ) ;
  assign n20435 = n20434 ^ n20433 ^ n14244 ;
  assign n20436 = n17922 ^ n2086 ^ 1'b0 ;
  assign n20437 = n9064 & n20436 ;
  assign n20438 = ( n13905 & ~n16252 ) | ( n13905 & n20437 ) | ( ~n16252 & n20437 ) ;
  assign n20439 = n12097 ^ n3019 ^ 1'b0 ;
  assign n20440 = ( n1845 & ~n14625 ) | ( n1845 & n20439 ) | ( ~n14625 & n20439 ) ;
  assign n20441 = n8896 | n11765 ;
  assign n20442 = n20440 & ~n20441 ;
  assign n20443 = ( ~n9960 & n16124 ) | ( ~n9960 & n20442 ) | ( n16124 & n20442 ) ;
  assign n20444 = n1651 & ~n3460 ;
  assign n20445 = n3763 & n20444 ;
  assign n20446 = n16698 ^ n11196 ^ n7612 ;
  assign n20447 = ( n1454 & n14347 ) | ( n1454 & n20446 ) | ( n14347 & n20446 ) ;
  assign n20448 = ( n18702 & n20445 ) | ( n18702 & n20447 ) | ( n20445 & n20447 ) ;
  assign n20449 = n20448 ^ n4173 ^ n4011 ;
  assign n20450 = n11436 ^ n8945 ^ n1318 ;
  assign n20451 = ( n940 & ~n4687 ) | ( n940 & n20450 ) | ( ~n4687 & n20450 ) ;
  assign n20452 = n18740 & n20451 ;
  assign n20453 = ( n7434 & n8873 ) | ( n7434 & ~n11752 ) | ( n8873 & ~n11752 ) ;
  assign n20454 = ~n13570 & n20453 ;
  assign n20455 = n20454 ^ n10848 ^ 1'b0 ;
  assign n20456 = n6457 ^ n1456 ^ 1'b0 ;
  assign n20457 = ~n20455 & n20456 ;
  assign n20460 = n10130 ^ n1249 ^ n1119 ;
  assign n20458 = ( x6 & n3255 ) | ( x6 & ~n5074 ) | ( n3255 & ~n5074 ) ;
  assign n20459 = n13244 | n20458 ;
  assign n20461 = n20460 ^ n20459 ^ n14653 ;
  assign n20462 = n20461 ^ n19162 ^ n1818 ;
  assign n20463 = n20280 ^ n10088 ^ n379 ;
  assign n20464 = ( n1303 & n1989 ) | ( n1303 & ~n20463 ) | ( n1989 & ~n20463 ) ;
  assign n20465 = n20464 ^ n6889 ^ n376 ;
  assign n20470 = n13976 ^ n6339 ^ n3442 ;
  assign n20466 = n6975 ^ n6838 ^ n4991 ;
  assign n20467 = n20466 ^ n9425 ^ n8185 ;
  assign n20468 = ( n293 & n6911 ) | ( n293 & ~n20467 ) | ( n6911 & ~n20467 ) ;
  assign n20469 = n13797 & ~n20468 ;
  assign n20471 = n20470 ^ n20469 ^ 1'b0 ;
  assign n20472 = ( ~n10144 & n11694 ) | ( ~n10144 & n13509 ) | ( n11694 & n13509 ) ;
  assign n20473 = ( n5586 & ~n15468 ) | ( n5586 & n20472 ) | ( ~n15468 & n20472 ) ;
  assign n20474 = n20473 ^ n9649 ^ n5393 ;
  assign n20475 = n20474 ^ n11081 ^ n2085 ;
  assign n20476 = n13016 ^ n12673 ^ n12407 ;
  assign n20477 = n20476 ^ n7253 ^ n4443 ;
  assign n20479 = n1647 ^ n1173 ^ 1'b0 ;
  assign n20480 = n5038 & ~n20479 ;
  assign n20478 = ( n6788 & n8127 ) | ( n6788 & ~n18434 ) | ( n8127 & ~n18434 ) ;
  assign n20481 = n20480 ^ n20478 ^ 1'b0 ;
  assign n20482 = ( n9742 & n17308 ) | ( n9742 & n20481 ) | ( n17308 & n20481 ) ;
  assign n20483 = n16376 ^ n7283 ^ 1'b0 ;
  assign n20484 = ( n3392 & ~n16471 ) | ( n3392 & n20483 ) | ( ~n16471 & n20483 ) ;
  assign n20485 = n11981 ^ n11924 ^ n2637 ;
  assign n20486 = n17180 ^ n12089 ^ n8307 ;
  assign n20487 = n20485 & ~n20486 ;
  assign n20488 = n20487 ^ n12513 ^ 1'b0 ;
  assign n20489 = ( n4812 & ~n20484 ) | ( n4812 & n20488 ) | ( ~n20484 & n20488 ) ;
  assign n20495 = n7719 ^ n2709 ^ n2317 ;
  assign n20490 = ( n2941 & ~n9560 ) | ( n2941 & n15065 ) | ( ~n9560 & n15065 ) ;
  assign n20491 = ( n8034 & n18916 ) | ( n8034 & ~n20490 ) | ( n18916 & ~n20490 ) ;
  assign n20492 = n20491 ^ n7522 ^ n7457 ;
  assign n20493 = n20492 ^ n17237 ^ n9076 ;
  assign n20494 = ( ~n3809 & n11415 ) | ( ~n3809 & n20493 ) | ( n11415 & n20493 ) ;
  assign n20496 = n20495 ^ n20494 ^ n17986 ;
  assign n20497 = n7251 ^ n3571 ^ n1235 ;
  assign n20498 = ( ~n14966 & n18512 ) | ( ~n14966 & n20497 ) | ( n18512 & n20497 ) ;
  assign n20499 = ( n7354 & n10285 ) | ( n7354 & n20498 ) | ( n10285 & n20498 ) ;
  assign n20500 = n1217 & n13933 ;
  assign n20501 = n13458 ^ n6109 ^ n3053 ;
  assign n20502 = n20501 ^ n8980 ^ n8396 ;
  assign n20503 = n12029 ^ n4585 ^ x182 ;
  assign n20504 = ( n16786 & n19812 ) | ( n16786 & ~n20503 ) | ( n19812 & ~n20503 ) ;
  assign n20505 = n8016 ^ n2687 ^ n2544 ;
  assign n20506 = ( n807 & n10105 ) | ( n807 & ~n20505 ) | ( n10105 & ~n20505 ) ;
  assign n20507 = n11955 ^ n3120 ^ n933 ;
  assign n20508 = n7044 ^ n2951 ^ n1838 ;
  assign n20509 = ( ~n5008 & n12733 ) | ( ~n5008 & n20508 ) | ( n12733 & n20508 ) ;
  assign n20510 = n20509 ^ n13684 ^ n3051 ;
  assign n20511 = ( n17157 & ~n20507 ) | ( n17157 & n20510 ) | ( ~n20507 & n20510 ) ;
  assign n20512 = ( n2713 & n11352 ) | ( n2713 & ~n12311 ) | ( n11352 & ~n12311 ) ;
  assign n20513 = n20511 & n20512 ;
  assign n20514 = ~n15179 & n20513 ;
  assign n20515 = n4638 | n20514 ;
  assign n20516 = n20506 & ~n20515 ;
  assign n20517 = n15373 ^ n4155 ^ n2289 ;
  assign n20518 = n1845 & n8133 ;
  assign n20519 = ( n3464 & ~n20517 ) | ( n3464 & n20518 ) | ( ~n20517 & n20518 ) ;
  assign n20520 = n14647 ^ n6775 ^ n6037 ;
  assign n20521 = n8369 ^ n6836 ^ n6071 ;
  assign n20522 = n20521 ^ n5867 ^ n4080 ;
  assign n20523 = n14690 | n20522 ;
  assign n20524 = n20523 ^ n4887 ^ 1'b0 ;
  assign n20525 = n20524 ^ n6129 ^ 1'b0 ;
  assign n20526 = ~n19424 & n20525 ;
  assign n20527 = ( x67 & n3466 ) | ( x67 & n11552 ) | ( n3466 & n11552 ) ;
  assign n20529 = n7509 & ~n8944 ;
  assign n20530 = n20529 ^ n10031 ^ 1'b0 ;
  assign n20531 = n11471 & ~n20530 ;
  assign n20532 = n8611 & n20531 ;
  assign n20528 = n17683 ^ n9783 ^ n6774 ;
  assign n20533 = n20532 ^ n20528 ^ n5429 ;
  assign n20534 = n20533 ^ n16599 ^ n11381 ;
  assign n20539 = n10642 | n11574 ;
  assign n20540 = n6255 & ~n20539 ;
  assign n20538 = ( n1461 & n6513 ) | ( n1461 & n7934 ) | ( n6513 & n7934 ) ;
  assign n20541 = n20540 ^ n20538 ^ 1'b0 ;
  assign n20535 = n12926 ^ n9862 ^ n1764 ;
  assign n20536 = n20535 ^ n5901 ^ 1'b0 ;
  assign n20537 = n20536 ^ n6009 ^ n1662 ;
  assign n20542 = n20541 ^ n20537 ^ n18051 ;
  assign n20543 = ( n13043 & ~n20534 ) | ( n13043 & n20542 ) | ( ~n20534 & n20542 ) ;
  assign n20550 = ( x94 & n462 ) | ( x94 & n11007 ) | ( n462 & n11007 ) ;
  assign n20551 = ( ~n4052 & n9542 ) | ( ~n4052 & n20550 ) | ( n9542 & n20550 ) ;
  assign n20548 = n15064 ^ n8007 ^ n1101 ;
  assign n20544 = n880 & ~n10999 ;
  assign n20545 = n20544 ^ n5910 ^ 1'b0 ;
  assign n20546 = ( ~n8359 & n9252 ) | ( ~n8359 & n20545 ) | ( n9252 & n20545 ) ;
  assign n20547 = n20546 ^ n13030 ^ n1250 ;
  assign n20549 = n20548 ^ n20547 ^ n18591 ;
  assign n20552 = n20551 ^ n20549 ^ n13704 ;
  assign n20558 = n1747 & ~n7244 ;
  assign n20559 = ~n6618 & n20558 ;
  assign n20555 = ~n4267 & n17501 ;
  assign n20556 = n15059 ^ n15002 ^ n1182 ;
  assign n20557 = ( n978 & n20555 ) | ( n978 & n20556 ) | ( n20555 & n20556 ) ;
  assign n20553 = n18900 ^ n962 ^ 1'b0 ;
  assign n20554 = n10487 & n20553 ;
  assign n20560 = n20559 ^ n20557 ^ n20554 ;
  assign n20561 = n16723 ^ n15574 ^ n8629 ;
  assign n20562 = n20561 ^ n16140 ^ n2062 ;
  assign n20563 = ( ~n8929 & n10809 ) | ( ~n8929 & n20562 ) | ( n10809 & n20562 ) ;
  assign n20564 = ~n7099 & n20563 ;
  assign n20565 = n20560 & n20564 ;
  assign n20566 = n11237 ^ n8390 ^ n6996 ;
  assign n20567 = ( n519 & n4653 ) | ( n519 & ~n5719 ) | ( n4653 & ~n5719 ) ;
  assign n20568 = ( n13311 & ~n13441 ) | ( n13311 & n20567 ) | ( ~n13441 & n20567 ) ;
  assign n20569 = ( n1988 & n3794 ) | ( n1988 & n15132 ) | ( n3794 & n15132 ) ;
  assign n20570 = n4880 | n12866 ;
  assign n20571 = ( n2835 & n20451 ) | ( n2835 & n20570 ) | ( n20451 & n20570 ) ;
  assign n20575 = n8008 ^ n5968 ^ n5932 ;
  assign n20576 = n20575 ^ n2945 ^ n946 ;
  assign n20577 = n6649 ^ n3162 ^ n2100 ;
  assign n20578 = ( n11756 & ~n20576 ) | ( n11756 & n20577 ) | ( ~n20576 & n20577 ) ;
  assign n20572 = ( n983 & n4914 ) | ( n983 & ~n20108 ) | ( n4914 & ~n20108 ) ;
  assign n20573 = n17398 ^ n16031 ^ n8305 ;
  assign n20574 = ( n16975 & n20572 ) | ( n16975 & n20573 ) | ( n20572 & n20573 ) ;
  assign n20579 = n20578 ^ n20574 ^ n16829 ;
  assign n20580 = n7430 ^ n3622 ^ n791 ;
  assign n20581 = n11714 ^ n9701 ^ n6679 ;
  assign n20582 = ( n7963 & ~n13051 ) | ( n7963 & n19203 ) | ( ~n13051 & n19203 ) ;
  assign n20583 = n20582 ^ n19350 ^ n4181 ;
  assign n20592 = ( n379 & n3137 ) | ( n379 & ~n11318 ) | ( n3137 & ~n11318 ) ;
  assign n20593 = n12806 ^ n10734 ^ n5057 ;
  assign n20594 = ( n16491 & n20592 ) | ( n16491 & ~n20593 ) | ( n20592 & ~n20593 ) ;
  assign n20589 = n12150 ^ n5066 ^ n3160 ;
  assign n20588 = ( n3127 & ~n3995 ) | ( n3127 & n5954 ) | ( ~n3995 & n5954 ) ;
  assign n20590 = n20589 ^ n20588 ^ n7933 ;
  assign n20586 = n11839 | n18732 ;
  assign n20584 = ( n2702 & ~n3791 ) | ( n2702 & n12323 ) | ( ~n3791 & n12323 ) ;
  assign n20585 = ( n1887 & n9869 ) | ( n1887 & n20584 ) | ( n9869 & n20584 ) ;
  assign n20587 = n20586 ^ n20585 ^ n2287 ;
  assign n20591 = n20590 ^ n20587 ^ n9354 ;
  assign n20595 = n20594 ^ n20591 ^ n8870 ;
  assign n20596 = n13541 ^ n10150 ^ n783 ;
  assign n20597 = ( ~n1623 & n6780 ) | ( ~n1623 & n14455 ) | ( n6780 & n14455 ) ;
  assign n20598 = n13357 ^ n9035 ^ n4418 ;
  assign n20599 = n20598 ^ n12153 ^ n10426 ;
  assign n20601 = ( ~n2300 & n7432 ) | ( ~n2300 & n15437 ) | ( n7432 & n15437 ) ;
  assign n20600 = ( n2312 & ~n4557 ) | ( n2312 & n6321 ) | ( ~n4557 & n6321 ) ;
  assign n20602 = n20601 ^ n20600 ^ n4799 ;
  assign n20603 = ( n20597 & ~n20599 ) | ( n20597 & n20602 ) | ( ~n20599 & n20602 ) ;
  assign n20605 = n6952 ^ n4080 ^ n3987 ;
  assign n20604 = n6892 & n19639 ;
  assign n20606 = n20605 ^ n20604 ^ 1'b0 ;
  assign n20607 = ( n433 & n14979 ) | ( n433 & n20606 ) | ( n14979 & n20606 ) ;
  assign n20608 = ( n641 & n5322 ) | ( n641 & n9587 ) | ( n5322 & n9587 ) ;
  assign n20609 = ( n6120 & ~n11615 ) | ( n6120 & n20608 ) | ( ~n11615 & n20608 ) ;
  assign n20610 = n20609 ^ n18002 ^ n6132 ;
  assign n20611 = n6095 & n20610 ;
  assign n20612 = ~n6144 & n20611 ;
  assign n20613 = n19446 ^ n18546 ^ n3039 ;
  assign n20614 = ( n10298 & n12775 ) | ( n10298 & ~n18454 ) | ( n12775 & ~n18454 ) ;
  assign n20615 = n20614 ^ n18974 ^ n8843 ;
  assign n20616 = ( n13939 & n15702 ) | ( n13939 & n20615 ) | ( n15702 & n20615 ) ;
  assign n20617 = n19797 ^ n11798 ^ n3318 ;
  assign n20625 = ( ~n659 & n733 ) | ( ~n659 & n11863 ) | ( n733 & n11863 ) ;
  assign n20626 = n18162 ^ n15608 ^ n9793 ;
  assign n20627 = n20626 ^ n14262 ^ n4463 ;
  assign n20628 = ( n8531 & n20625 ) | ( n8531 & ~n20627 ) | ( n20625 & ~n20627 ) ;
  assign n20618 = n15544 ^ n9481 ^ n2115 ;
  assign n20619 = ( n886 & n6711 ) | ( n886 & n20618 ) | ( n6711 & n20618 ) ;
  assign n20620 = n13906 ^ n12122 ^ n4488 ;
  assign n20621 = n4707 & ~n15505 ;
  assign n20622 = n20621 ^ n13625 ^ 1'b0 ;
  assign n20623 = ( n19848 & n20620 ) | ( n19848 & ~n20622 ) | ( n20620 & ~n20622 ) ;
  assign n20624 = ( n867 & ~n20619 ) | ( n867 & n20623 ) | ( ~n20619 & n20623 ) ;
  assign n20629 = n20628 ^ n20624 ^ n15447 ;
  assign n20630 = x163 & n20629 ;
  assign n20631 = ~n20617 & n20630 ;
  assign n20636 = n20584 ^ n14069 ^ n4580 ;
  assign n20632 = ( n2154 & n2621 ) | ( n2154 & n8327 ) | ( n2621 & n8327 ) ;
  assign n20633 = n10811 ^ n9140 ^ n8336 ;
  assign n20634 = n20633 ^ n10838 ^ n7075 ;
  assign n20635 = ( ~n3160 & n20632 ) | ( ~n3160 & n20634 ) | ( n20632 & n20634 ) ;
  assign n20637 = n20636 ^ n20635 ^ n11853 ;
  assign n20638 = n15626 ^ n6845 ^ 1'b0 ;
  assign n20639 = n2506 ^ n1751 ^ n765 ;
  assign n20640 = n20639 ^ n4329 ^ n1484 ;
  assign n20641 = n20640 ^ n20534 ^ n14629 ;
  assign n20642 = ( n5079 & n18386 ) | ( n5079 & n20641 ) | ( n18386 & n20641 ) ;
  assign n20643 = n11346 & ~n13130 ;
  assign n20644 = ~n5631 & n20643 ;
  assign n20645 = ( ~n3428 & n17777 ) | ( ~n3428 & n20644 ) | ( n17777 & n20644 ) ;
  assign n20646 = ( n1553 & ~n12516 ) | ( n1553 & n20645 ) | ( ~n12516 & n20645 ) ;
  assign n20647 = ( ~n1927 & n4056 ) | ( ~n1927 & n20646 ) | ( n4056 & n20646 ) ;
  assign n20648 = ( n2316 & n6528 ) | ( n2316 & ~n20647 ) | ( n6528 & ~n20647 ) ;
  assign n20649 = ~n10121 & n10217 ;
  assign n20650 = ~n5428 & n20649 ;
  assign n20651 = ( n1891 & n6631 ) | ( n1891 & ~n20650 ) | ( n6631 & ~n20650 ) ;
  assign n20653 = ( ~n536 & n10515 ) | ( ~n536 & n13112 ) | ( n10515 & n13112 ) ;
  assign n20652 = n11968 | n13358 ;
  assign n20654 = n20653 ^ n20652 ^ n10087 ;
  assign n20655 = ( n5798 & n20651 ) | ( n5798 & ~n20654 ) | ( n20651 & ~n20654 ) ;
  assign n20656 = ( n3361 & n3895 ) | ( n3361 & n7746 ) | ( n3895 & n7746 ) ;
  assign n20657 = n20656 ^ n9986 ^ 1'b0 ;
  assign n20658 = ( n555 & n961 ) | ( n555 & n20657 ) | ( n961 & n20657 ) ;
  assign n20659 = ~n2088 & n3154 ;
  assign n20660 = n20659 ^ n13779 ^ 1'b0 ;
  assign n20661 = ( n1446 & n4927 ) | ( n1446 & n19815 ) | ( n4927 & n19815 ) ;
  assign n20662 = ( n1785 & n3615 ) | ( n1785 & ~n3856 ) | ( n3615 & ~n3856 ) ;
  assign n20663 = n20662 ^ n13596 ^ n6373 ;
  assign n20664 = ( n20660 & n20661 ) | ( n20660 & n20663 ) | ( n20661 & n20663 ) ;
  assign n20665 = ( n4215 & n4968 ) | ( n4215 & n6150 ) | ( n4968 & n6150 ) ;
  assign n20666 = ( ~n3739 & n4460 ) | ( ~n3739 & n4732 ) | ( n4460 & n4732 ) ;
  assign n20667 = n20665 | n20666 ;
  assign n20668 = n12121 ^ n8603 ^ n5731 ;
  assign n20669 = ( n15048 & ~n19737 ) | ( n15048 & n20668 ) | ( ~n19737 & n20668 ) ;
  assign n20670 = ( n1402 & ~n2481 ) | ( n1402 & n3486 ) | ( ~n2481 & n3486 ) ;
  assign n20671 = n20670 ^ n10198 ^ n3933 ;
  assign n20672 = ( ~n5817 & n14825 ) | ( ~n5817 & n20671 ) | ( n14825 & n20671 ) ;
  assign n20673 = n20672 ^ n8267 ^ 1'b0 ;
  assign n20674 = n20673 ^ n13923 ^ n13261 ;
  assign n20675 = n20674 ^ n5495 ^ n2054 ;
  assign n20676 = ( n4031 & n5330 ) | ( n4031 & n7139 ) | ( n5330 & n7139 ) ;
  assign n20677 = n20676 ^ n18944 ^ n3768 ;
  assign n20678 = n5815 & ~n6787 ;
  assign n20679 = n5240 & n20678 ;
  assign n20680 = n12180 ^ n9320 ^ n5847 ;
  assign n20681 = n20680 ^ n20007 ^ n15734 ;
  assign n20682 = ( ~n18471 & n20679 ) | ( ~n18471 & n20681 ) | ( n20679 & n20681 ) ;
  assign n20683 = ( n11719 & ~n12682 ) | ( n11719 & n17623 ) | ( ~n12682 & n17623 ) ;
  assign n20684 = ( n12326 & n20682 ) | ( n12326 & ~n20683 ) | ( n20682 & ~n20683 ) ;
  assign n20685 = n20684 ^ n15557 ^ n8101 ;
  assign n20686 = n12557 ^ n1636 ^ 1'b0 ;
  assign n20687 = n15868 & ~n20686 ;
  assign n20688 = ( ~n5171 & n5809 ) | ( ~n5171 & n16338 ) | ( n5809 & n16338 ) ;
  assign n20689 = ( n2379 & ~n10642 ) | ( n2379 & n20688 ) | ( ~n10642 & n20688 ) ;
  assign n20690 = n6227 ^ n2556 ^ n2458 ;
  assign n20691 = n20690 ^ n6079 ^ 1'b0 ;
  assign n20692 = n3475 & ~n20691 ;
  assign n20693 = ( ~n2139 & n8601 ) | ( ~n2139 & n20692 ) | ( n8601 & n20692 ) ;
  assign n20694 = n19525 ^ n14025 ^ n1954 ;
  assign n20695 = n20694 ^ n17996 ^ n7125 ;
  assign n20696 = ( x45 & ~n13035 ) | ( x45 & n14106 ) | ( ~n13035 & n14106 ) ;
  assign n20697 = n15234 ^ n8349 ^ 1'b0 ;
  assign n20698 = n20697 ^ n12160 ^ n5128 ;
  assign n20699 = ( n5727 & n9357 ) | ( n5727 & n10725 ) | ( n9357 & n10725 ) ;
  assign n20700 = ( ~n740 & n4673 ) | ( ~n740 & n20699 ) | ( n4673 & n20699 ) ;
  assign n20701 = n20700 ^ n14274 ^ n5322 ;
  assign n20702 = n2664 | n16939 ;
  assign n20703 = n20702 ^ n4863 ^ 1'b0 ;
  assign n20704 = n4322 | n20703 ;
  assign n20705 = n15676 ^ n9003 ^ n8525 ;
  assign n20706 = ( n5470 & n14645 ) | ( n5470 & n15806 ) | ( n14645 & n15806 ) ;
  assign n20707 = n16985 ^ n10049 ^ 1'b0 ;
  assign n20708 = ( n5053 & n11113 ) | ( n5053 & ~n15041 ) | ( n11113 & ~n15041 ) ;
  assign n20709 = n20707 | n20708 ;
  assign n20710 = ( n2267 & n3329 ) | ( n2267 & n3667 ) | ( n3329 & n3667 ) ;
  assign n20711 = n14371 | n20710 ;
  assign n20712 = ( n4394 & n10570 ) | ( n4394 & n10636 ) | ( n10570 & n10636 ) ;
  assign n20713 = ( n10097 & ~n13749 ) | ( n10097 & n16091 ) | ( ~n13749 & n16091 ) ;
  assign n20719 = ( x41 & n1335 ) | ( x41 & ~n3273 ) | ( n1335 & ~n3273 ) ;
  assign n20714 = n11393 ^ n8844 ^ n1551 ;
  assign n20715 = ( n1636 & n2122 ) | ( n1636 & ~n20714 ) | ( n2122 & ~n20714 ) ;
  assign n20716 = ( n1132 & n10504 ) | ( n1132 & ~n19749 ) | ( n10504 & ~n19749 ) ;
  assign n20717 = ~n14127 & n20716 ;
  assign n20718 = n20715 & n20717 ;
  assign n20720 = n20719 ^ n20718 ^ 1'b0 ;
  assign n20721 = n5751 ^ n884 ^ x94 ;
  assign n20722 = n10396 ^ n3471 ^ n978 ;
  assign n20723 = ( n3569 & n8260 ) | ( n3569 & n19317 ) | ( n8260 & n19317 ) ;
  assign n20724 = ( n2728 & n20722 ) | ( n2728 & ~n20723 ) | ( n20722 & ~n20723 ) ;
  assign n20725 = ( n736 & n20721 ) | ( n736 & n20724 ) | ( n20721 & n20724 ) ;
  assign n20726 = n20725 ^ n5335 ^ n2703 ;
  assign n20727 = n20726 ^ n8342 ^ n1638 ;
  assign n20730 = ( ~n325 & n1224 ) | ( ~n325 & n1254 ) | ( n1224 & n1254 ) ;
  assign n20731 = ( n1987 & n11390 ) | ( n1987 & n20644 ) | ( n11390 & n20644 ) ;
  assign n20732 = n7640 & n20731 ;
  assign n20733 = ( ~n3065 & n20730 ) | ( ~n3065 & n20732 ) | ( n20730 & n20732 ) ;
  assign n20728 = ( n4460 & ~n10401 ) | ( n4460 & n19074 ) | ( ~n10401 & n19074 ) ;
  assign n20729 = n20728 ^ n11220 ^ n7690 ;
  assign n20734 = n20733 ^ n20729 ^ n13342 ;
  assign n20735 = ( n4232 & n8745 ) | ( n4232 & ~n16554 ) | ( n8745 & ~n16554 ) ;
  assign n20737 = ( n1012 & n3481 ) | ( n1012 & n4768 ) | ( n3481 & n4768 ) ;
  assign n20736 = n6639 ^ n5024 ^ 1'b0 ;
  assign n20738 = n20737 ^ n20736 ^ n18471 ;
  assign n20739 = ( n11464 & n20735 ) | ( n11464 & n20738 ) | ( n20735 & n20738 ) ;
  assign n20740 = ( n3028 & ~n5490 ) | ( n3028 & n19093 ) | ( ~n5490 & n19093 ) ;
  assign n20741 = n20740 ^ n10255 ^ n3859 ;
  assign n20742 = n8980 ^ n3822 ^ n2705 ;
  assign n20745 = n3725 & n11153 ;
  assign n20743 = n9232 ^ n1812 ^ n462 ;
  assign n20744 = n20743 ^ n5897 ^ n3921 ;
  assign n20746 = n20745 ^ n20744 ^ n7999 ;
  assign n20747 = n20746 ^ n8450 ^ n5081 ;
  assign n20753 = ( n1127 & n4040 ) | ( n1127 & ~n13509 ) | ( n4040 & ~n13509 ) ;
  assign n20754 = n20753 ^ n1473 ^ 1'b0 ;
  assign n20748 = n4781 ^ n3659 ^ 1'b0 ;
  assign n20749 = n8136 ^ n2251 ^ 1'b0 ;
  assign n20750 = n2513 | n20749 ;
  assign n20751 = ( n2074 & ~n20748 ) | ( n2074 & n20750 ) | ( ~n20748 & n20750 ) ;
  assign n20752 = n20751 ^ n19120 ^ n3759 ;
  assign n20755 = n20754 ^ n20752 ^ n1639 ;
  assign n20756 = n9966 ^ n5920 ^ n4553 ;
  assign n20757 = ( n8150 & n13521 ) | ( n8150 & ~n20756 ) | ( n13521 & ~n20756 ) ;
  assign n20758 = n15713 ^ n5491 ^ n5472 ;
  assign n20759 = ( n1670 & ~n13321 ) | ( n1670 & n14072 ) | ( ~n13321 & n14072 ) ;
  assign n20760 = ( n7187 & n15326 ) | ( n7187 & n20759 ) | ( n15326 & n20759 ) ;
  assign n20766 = n10906 ^ n10783 ^ n1837 ;
  assign n20761 = ( n456 & ~n8023 ) | ( n456 & n18510 ) | ( ~n8023 & n18510 ) ;
  assign n20762 = n11558 ^ x134 ^ 1'b0 ;
  assign n20763 = ( ~n3387 & n20761 ) | ( ~n3387 & n20762 ) | ( n20761 & n20762 ) ;
  assign n20764 = ( ~n6411 & n19438 ) | ( ~n6411 & n20763 ) | ( n19438 & n20763 ) ;
  assign n20765 = ( n8647 & n19736 ) | ( n8647 & ~n20764 ) | ( n19736 & ~n20764 ) ;
  assign n20767 = n20766 ^ n20765 ^ 1'b0 ;
  assign n20768 = ( ~n8557 & n9866 ) | ( ~n8557 & n10777 ) | ( n9866 & n10777 ) ;
  assign n20769 = n20768 ^ n14524 ^ n11027 ;
  assign n20770 = n13625 ^ n9399 ^ n8615 ;
  assign n20771 = ( n4310 & n4445 ) | ( n4310 & ~n20770 ) | ( n4445 & ~n20770 ) ;
  assign n20772 = n20771 ^ n18509 ^ n3600 ;
  assign n20773 = n20772 ^ n12647 ^ n6385 ;
  assign n20774 = n1808 | n7752 ;
  assign n20775 = n4678 | n20774 ;
  assign n20776 = ( ~n284 & n11503 ) | ( ~n284 & n12249 ) | ( n11503 & n12249 ) ;
  assign n20777 = ( ~n984 & n2687 ) | ( ~n984 & n20776 ) | ( n2687 & n20776 ) ;
  assign n20778 = n20777 ^ n19084 ^ n11529 ;
  assign n20779 = ( ~n20773 & n20775 ) | ( ~n20773 & n20778 ) | ( n20775 & n20778 ) ;
  assign n20780 = ( ~n1236 & n4952 ) | ( ~n1236 & n5748 ) | ( n4952 & n5748 ) ;
  assign n20781 = ( n3766 & n12754 ) | ( n3766 & ~n20780 ) | ( n12754 & ~n20780 ) ;
  assign n20782 = ( ~n3807 & n20033 ) | ( ~n3807 & n20781 ) | ( n20033 & n20781 ) ;
  assign n20783 = n9409 ^ n3639 ^ n663 ;
  assign n20784 = ( n14525 & ~n18050 ) | ( n14525 & n20783 ) | ( ~n18050 & n20783 ) ;
  assign n20785 = n2829 ^ n382 ^ 1'b0 ;
  assign n20786 = ( ~x192 & n2201 ) | ( ~x192 & n20785 ) | ( n2201 & n20785 ) ;
  assign n20787 = ( ~n20782 & n20784 ) | ( ~n20782 & n20786 ) | ( n20784 & n20786 ) ;
  assign n20788 = n20787 ^ n19682 ^ n16027 ;
  assign n20789 = n20551 ^ n11720 ^ n2183 ;
  assign n20790 = ( n19192 & n20788 ) | ( n19192 & ~n20789 ) | ( n20788 & ~n20789 ) ;
  assign n20791 = ( n5515 & n11574 ) | ( n5515 & n19401 ) | ( n11574 & n19401 ) ;
  assign n20792 = ( ~n4164 & n13447 ) | ( ~n4164 & n20791 ) | ( n13447 & n20791 ) ;
  assign n20793 = ( n5138 & n7542 ) | ( n5138 & n20792 ) | ( n7542 & n20792 ) ;
  assign n20797 = ( n5892 & n7768 ) | ( n5892 & n11854 ) | ( n7768 & n11854 ) ;
  assign n20794 = ( n2154 & n9464 ) | ( n2154 & ~n11207 ) | ( n9464 & ~n11207 ) ;
  assign n20795 = n20794 ^ n3332 ^ x65 ;
  assign n20796 = n20795 ^ n17797 ^ n7888 ;
  assign n20798 = n20797 ^ n20796 ^ n5765 ;
  assign n20799 = ( n3348 & n3558 ) | ( n3348 & n20798 ) | ( n3558 & n20798 ) ;
  assign n20800 = n17784 ^ n11259 ^ n6674 ;
  assign n20801 = n13664 & ~n20800 ;
  assign n20802 = ~n13460 & n20801 ;
  assign n20803 = ( n16640 & ~n18824 ) | ( n16640 & n20802 ) | ( ~n18824 & n20802 ) ;
  assign n20804 = n8839 & ~n11528 ;
  assign n20805 = n20803 & n20804 ;
  assign n20806 = ~n11752 & n19923 ;
  assign n20807 = n20806 ^ n1711 ^ 1'b0 ;
  assign n20808 = n1658 & n12473 ;
  assign n20810 = ( x126 & n2505 ) | ( x126 & ~n6679 ) | ( n2505 & ~n6679 ) ;
  assign n20811 = n20810 ^ n433 ^ x224 ;
  assign n20809 = n18846 ^ n18090 ^ n4482 ;
  assign n20812 = n20811 ^ n20809 ^ n15765 ;
  assign n20813 = n18973 ^ n10772 ^ n5704 ;
  assign n20814 = n20813 ^ n3585 ^ n593 ;
  assign n20815 = n20814 ^ n11822 ^ n9351 ;
  assign n20816 = n7044 ^ x208 ^ 1'b0 ;
  assign n20817 = n17623 ^ n13079 ^ n11689 ;
  assign n20818 = ( ~n19290 & n20816 ) | ( ~n19290 & n20817 ) | ( n20816 & n20817 ) ;
  assign n20819 = ( n1459 & n20815 ) | ( n1459 & ~n20818 ) | ( n20815 & ~n20818 ) ;
  assign n20820 = ( n20808 & n20812 ) | ( n20808 & ~n20819 ) | ( n20812 & ~n20819 ) ;
  assign n20821 = ( n711 & n7494 ) | ( n711 & ~n16071 ) | ( n7494 & ~n16071 ) ;
  assign n20822 = n20821 ^ n18605 ^ 1'b0 ;
  assign n20823 = n12521 ^ n7906 ^ n6122 ;
  assign n20824 = n20823 ^ n15546 ^ n11210 ;
  assign n20825 = ( n6052 & ~n6248 ) | ( n6052 & n20824 ) | ( ~n6248 & n20824 ) ;
  assign n20826 = n16832 ^ n10327 ^ n9165 ;
  assign n20827 = n20826 ^ n14090 ^ n289 ;
  assign n20828 = n5709 ^ n5493 ^ n4807 ;
  assign n20829 = n20828 ^ n16221 ^ n10515 ;
  assign n20830 = ~n6830 & n20829 ;
  assign n20831 = ( n20825 & n20827 ) | ( n20825 & ~n20830 ) | ( n20827 & ~n20830 ) ;
  assign n20832 = n20633 ^ n17939 ^ n7746 ;
  assign n20846 = n8364 & n17858 ;
  assign n20847 = n20846 ^ n9355 ^ 1'b0 ;
  assign n20848 = ( n6177 & n18211 ) | ( n6177 & ~n20847 ) | ( n18211 & ~n20847 ) ;
  assign n20840 = ~n1742 & n4725 ;
  assign n20841 = ~x189 & n20840 ;
  assign n20842 = ( n3422 & ~n16106 ) | ( n3422 & n20841 ) | ( ~n16106 & n20841 ) ;
  assign n20843 = ( ~n3910 & n5379 ) | ( ~n3910 & n10973 ) | ( n5379 & n10973 ) ;
  assign n20844 = n20843 ^ n18213 ^ n16095 ;
  assign n20845 = ( ~n15034 & n20842 ) | ( ~n15034 & n20844 ) | ( n20842 & n20844 ) ;
  assign n20833 = ( ~n1709 & n3420 ) | ( ~n1709 & n13114 ) | ( n3420 & n13114 ) ;
  assign n20834 = n3487 ^ n2254 ^ x234 ;
  assign n20835 = ( n6313 & n20833 ) | ( n6313 & n20834 ) | ( n20833 & n20834 ) ;
  assign n20836 = ( n4045 & ~n17242 ) | ( n4045 & n20835 ) | ( ~n17242 & n20835 ) ;
  assign n20837 = ~n11698 & n20836 ;
  assign n20838 = ( n14704 & n20508 ) | ( n14704 & ~n20837 ) | ( n20508 & ~n20837 ) ;
  assign n20839 = n20838 ^ n14134 ^ n1843 ;
  assign n20849 = n20848 ^ n20845 ^ n20839 ;
  assign n20850 = ( n8388 & n13300 ) | ( n8388 & ~n13910 ) | ( n13300 & ~n13910 ) ;
  assign n20851 = n8884 ^ n3279 ^ n2247 ;
  assign n20852 = ( n891 & ~n16082 ) | ( n891 & n20851 ) | ( ~n16082 & n20851 ) ;
  assign n20853 = ( n5107 & n9863 ) | ( n5107 & n14172 ) | ( n9863 & n14172 ) ;
  assign n20854 = ( ~n6167 & n11329 ) | ( ~n6167 & n20853 ) | ( n11329 & n20853 ) ;
  assign n20855 = ( n1288 & n12003 ) | ( n1288 & n17075 ) | ( n12003 & n17075 ) ;
  assign n20856 = n14150 ^ n12776 ^ n3370 ;
  assign n20857 = n14129 ^ n4413 ^ 1'b0 ;
  assign n20858 = n4292 ^ n1979 ^ 1'b0 ;
  assign n20859 = n20858 ^ n15369 ^ n8807 ;
  assign n20860 = n20859 ^ n16573 ^ 1'b0 ;
  assign n20861 = ( n3735 & ~n20857 ) | ( n3735 & n20860 ) | ( ~n20857 & n20860 ) ;
  assign n20864 = x32 & n20104 ;
  assign n20865 = n6251 & n20864 ;
  assign n20862 = n11102 ^ n9355 ^ n8293 ;
  assign n20863 = ( n393 & n13714 ) | ( n393 & ~n20862 ) | ( n13714 & ~n20862 ) ;
  assign n20866 = n20865 ^ n20863 ^ n10429 ;
  assign n20869 = n10544 ^ n9855 ^ n1598 ;
  assign n20870 = n20869 ^ n13916 ^ 1'b0 ;
  assign n20867 = n14246 | n14437 ;
  assign n20868 = n20867 ^ n14955 ^ 1'b0 ;
  assign n20871 = n20870 ^ n20868 ^ n6075 ;
  assign n20872 = n1988 ^ x230 ^ 1'b0 ;
  assign n20873 = n13806 ^ n12735 ^ n2909 ;
  assign n20874 = n17932 | n19664 ;
  assign n20875 = n18042 | n20874 ;
  assign n20876 = n8609 ^ n828 ^ n802 ;
  assign n20877 = ( n2197 & ~n20875 ) | ( n2197 & n20876 ) | ( ~n20875 & n20876 ) ;
  assign n20878 = n17942 ^ n11392 ^ n4474 ;
  assign n20879 = n4058 & n9846 ;
  assign n20880 = n19989 & n20879 ;
  assign n20881 = n20880 ^ n17580 ^ n6336 ;
  assign n20882 = n20881 ^ n16990 ^ n3734 ;
  assign n20883 = n10212 ^ n8155 ^ n6516 ;
  assign n20885 = ( ~n8908 & n9995 ) | ( ~n8908 & n18029 ) | ( n9995 & n18029 ) ;
  assign n20884 = n12739 ^ n6110 ^ 1'b0 ;
  assign n20886 = n20885 ^ n20884 ^ n3643 ;
  assign n20887 = ( n3685 & n12386 ) | ( n3685 & n20886 ) | ( n12386 & n20886 ) ;
  assign n20888 = ( n4271 & n15401 ) | ( n4271 & n20887 ) | ( n15401 & n20887 ) ;
  assign n20889 = ( ~n4213 & n20883 ) | ( ~n4213 & n20888 ) | ( n20883 & n20888 ) ;
  assign n20890 = n1298 & n11736 ;
  assign n20891 = n20890 ^ n8734 ^ 1'b0 ;
  assign n20895 = n2475 & ~n5275 ;
  assign n20896 = n6300 & n20895 ;
  assign n20897 = n20896 ^ n3582 ^ 1'b0 ;
  assign n20898 = n20897 ^ n11389 ^ n2374 ;
  assign n20894 = ( n5253 & n11863 ) | ( n5253 & n17603 ) | ( n11863 & n17603 ) ;
  assign n20892 = n5491 ^ n4840 ^ n2447 ;
  assign n20893 = ( n1022 & ~n12861 ) | ( n1022 & n20892 ) | ( ~n12861 & n20892 ) ;
  assign n20899 = n20898 ^ n20894 ^ n20893 ;
  assign n20900 = n12594 ^ n10578 ^ 1'b0 ;
  assign n20901 = n16636 ^ n11751 ^ n647 ;
  assign n20902 = n6028 ^ n4749 ^ 1'b0 ;
  assign n20903 = n20901 & n20902 ;
  assign n20904 = ( n14604 & n20900 ) | ( n14604 & n20903 ) | ( n20900 & n20903 ) ;
  assign n20905 = n20904 ^ n19482 ^ n16338 ;
  assign n20906 = n10811 ^ n394 ^ 1'b0 ;
  assign n20907 = n9855 & n20906 ;
  assign n20908 = ( n328 & n1605 ) | ( n328 & n9282 ) | ( n1605 & n9282 ) ;
  assign n20909 = ( ~n8152 & n20907 ) | ( ~n8152 & n20908 ) | ( n20907 & n20908 ) ;
  assign n20910 = n9136 ^ n3244 ^ n483 ;
  assign n20911 = n13724 ^ n6330 ^ n6088 ;
  assign n20912 = ( n20117 & n20910 ) | ( n20117 & ~n20911 ) | ( n20910 & ~n20911 ) ;
  assign n20913 = n5824 ^ n648 ^ n426 ;
  assign n20916 = n17871 ^ n3527 ^ 1'b0 ;
  assign n20915 = ( n4595 & ~n4606 ) | ( n4595 & n10777 ) | ( ~n4606 & n10777 ) ;
  assign n20917 = n20916 ^ n20915 ^ n11876 ;
  assign n20914 = ( n326 & n9806 ) | ( n326 & ~n11015 ) | ( n9806 & ~n11015 ) ;
  assign n20918 = n20917 ^ n20914 ^ 1'b0 ;
  assign n20919 = n20913 & n20918 ;
  assign n20920 = n10555 ^ n7314 ^ n2543 ;
  assign n20921 = ( n7598 & ~n12310 ) | ( n7598 & n20920 ) | ( ~n12310 & n20920 ) ;
  assign n20924 = n3135 ^ n1148 ^ n1078 ;
  assign n20922 = ( n6138 & ~n6377 ) | ( n6138 & n7756 ) | ( ~n6377 & n7756 ) ;
  assign n20923 = ( n2811 & n11566 ) | ( n2811 & n20922 ) | ( n11566 & n20922 ) ;
  assign n20925 = n20924 ^ n20923 ^ n12329 ;
  assign n20926 = n20925 ^ n17006 ^ n5546 ;
  assign n20927 = n4057 ^ n2587 ^ n2424 ;
  assign n20928 = n20927 ^ n3154 ^ n2272 ;
  assign n20929 = ~n2026 & n2348 ;
  assign n20930 = n9059 ^ n1997 ^ n1710 ;
  assign n20931 = ( ~n284 & n20929 ) | ( ~n284 & n20930 ) | ( n20929 & n20930 ) ;
  assign n20932 = ( n3952 & ~n20928 ) | ( n3952 & n20931 ) | ( ~n20928 & n20931 ) ;
  assign n20933 = n14204 ^ n12643 ^ n6509 ;
  assign n20934 = n3402 | n20933 ;
  assign n20935 = n6339 | n20934 ;
  assign n20936 = ( n8815 & n17877 ) | ( n8815 & n20935 ) | ( n17877 & n20935 ) ;
  assign n20943 = ( n7529 & n8296 ) | ( n7529 & n10466 ) | ( n8296 & n10466 ) ;
  assign n20939 = n9159 ^ n5286 ^ n1326 ;
  assign n20940 = n20939 ^ n8489 ^ n1351 ;
  assign n20941 = ( n3789 & n11786 ) | ( n3789 & n20940 ) | ( n11786 & n20940 ) ;
  assign n20942 = ~n11404 & n20941 ;
  assign n20937 = n13395 ^ n3197 ^ 1'b0 ;
  assign n20938 = n20937 ^ n19322 ^ n11281 ;
  assign n20944 = n20943 ^ n20942 ^ n20938 ;
  assign n20945 = ( n2139 & n5196 ) | ( n2139 & n16301 ) | ( n5196 & n16301 ) ;
  assign n20946 = ( n20936 & n20944 ) | ( n20936 & ~n20945 ) | ( n20944 & ~n20945 ) ;
  assign n20947 = ( n4828 & n11212 ) | ( n4828 & n20946 ) | ( n11212 & n20946 ) ;
  assign n20948 = n20947 ^ n18818 ^ n2572 ;
  assign n20949 = n14869 ^ n3681 ^ 1'b0 ;
  assign n20950 = n15310 & ~n20949 ;
  assign n20951 = ~n3182 & n3911 ;
  assign n20952 = n20951 ^ n1406 ^ 1'b0 ;
  assign n20953 = n20952 ^ n17309 ^ n14539 ;
  assign n20954 = ( n588 & ~n7075 ) | ( n588 & n20953 ) | ( ~n7075 & n20953 ) ;
  assign n20955 = ( x94 & n1026 ) | ( x94 & ~n20954 ) | ( n1026 & ~n20954 ) ;
  assign n20956 = ( n8535 & n20950 ) | ( n8535 & ~n20955 ) | ( n20950 & ~n20955 ) ;
  assign n20957 = ( ~n1922 & n8578 ) | ( ~n1922 & n9303 ) | ( n8578 & n9303 ) ;
  assign n20958 = ( n3763 & ~n19641 ) | ( n3763 & n20957 ) | ( ~n19641 & n20957 ) ;
  assign n20959 = n20299 ^ n11396 ^ n1183 ;
  assign n20963 = n1651 & n1935 ;
  assign n20964 = n2566 & n20963 ;
  assign n20965 = n20964 ^ n13065 ^ n10501 ;
  assign n20961 = ( n340 & ~n6498 ) | ( n340 & n8653 ) | ( ~n6498 & n8653 ) ;
  assign n20960 = ( ~n886 & n4782 ) | ( ~n886 & n13775 ) | ( n4782 & n13775 ) ;
  assign n20962 = n20961 ^ n20960 ^ n7627 ;
  assign n20966 = n20965 ^ n20962 ^ n11660 ;
  assign n20971 = n10444 ^ n9530 ^ n3453 ;
  assign n20972 = n13256 & n16569 ;
  assign n20973 = ~n9622 & n20972 ;
  assign n20974 = n20973 ^ n14135 ^ 1'b0 ;
  assign n20975 = n20971 & n20974 ;
  assign n20967 = n11095 ^ n2603 ^ 1'b0 ;
  assign n20968 = n18050 & n20967 ;
  assign n20969 = ~n8099 & n20968 ;
  assign n20970 = ~n2243 & n20969 ;
  assign n20976 = n20975 ^ n20970 ^ 1'b0 ;
  assign n20977 = ( x62 & n9466 ) | ( x62 & ~n16571 ) | ( n9466 & ~n16571 ) ;
  assign n20978 = ( n8292 & n10484 ) | ( n8292 & n16845 ) | ( n10484 & n16845 ) ;
  assign n20979 = n20977 & n20978 ;
  assign n20980 = ( n4018 & n5651 ) | ( n4018 & n8408 ) | ( n5651 & n8408 ) ;
  assign n20981 = ( ~n13023 & n15149 ) | ( ~n13023 & n20980 ) | ( n15149 & n20980 ) ;
  assign n20982 = n1601 & n9592 ;
  assign n20983 = n20982 ^ n19364 ^ n2727 ;
  assign n20984 = n6173 ^ n814 ^ 1'b0 ;
  assign n20985 = n17199 ^ n12694 ^ n4930 ;
  assign n20986 = n16242 ^ n5405 ^ x189 ;
  assign n20987 = n20986 ^ n4981 ^ n1169 ;
  assign n20988 = n20987 ^ n5871 ^ n2455 ;
  assign n20990 = ( n5309 & ~n6707 ) | ( n5309 & n14159 ) | ( ~n6707 & n14159 ) ;
  assign n20989 = ( n7179 & ~n15913 ) | ( n7179 & n16803 ) | ( ~n15913 & n16803 ) ;
  assign n20991 = n20990 ^ n20989 ^ n7515 ;
  assign n20992 = ( n1338 & ~n20988 ) | ( n1338 & n20991 ) | ( ~n20988 & n20991 ) ;
  assign n20993 = ( ~n18996 & n20985 ) | ( ~n18996 & n20992 ) | ( n20985 & n20992 ) ;
  assign n20999 = ( n7659 & ~n12366 ) | ( n7659 & n15247 ) | ( ~n12366 & n15247 ) ;
  assign n20996 = n10533 ^ n6617 ^ n3002 ;
  assign n20997 = n20996 ^ n10805 ^ n1621 ;
  assign n20994 = n11767 ^ n3062 ^ 1'b0 ;
  assign n20995 = n7873 & ~n20994 ;
  assign n20998 = n20997 ^ n20995 ^ n5565 ;
  assign n21000 = n20999 ^ n20998 ^ n17533 ;
  assign n21001 = ( n7003 & n7651 ) | ( n7003 & n14694 ) | ( n7651 & n14694 ) ;
  assign n21002 = ( n8265 & n18530 ) | ( n8265 & ~n18726 ) | ( n18530 & ~n18726 ) ;
  assign n21003 = ( n4611 & n16374 ) | ( n4611 & ~n21002 ) | ( n16374 & ~n21002 ) ;
  assign n21013 = n4191 ^ n3731 ^ n3203 ;
  assign n21011 = ( n8356 & n19505 ) | ( n8356 & ~n20234 ) | ( n19505 & ~n20234 ) ;
  assign n21010 = ( x78 & n10553 ) | ( x78 & n18474 ) | ( n10553 & n18474 ) ;
  assign n21004 = n11528 ^ n8978 ^ n2854 ;
  assign n21005 = ( n3688 & n8415 ) | ( n3688 & n17585 ) | ( n8415 & n17585 ) ;
  assign n21006 = ~n12451 & n21005 ;
  assign n21007 = n21006 ^ n17253 ^ n8885 ;
  assign n21008 = ( n2391 & n8425 ) | ( n2391 & ~n21007 ) | ( n8425 & ~n21007 ) ;
  assign n21009 = ( ~n3764 & n21004 ) | ( ~n3764 & n21008 ) | ( n21004 & n21008 ) ;
  assign n21012 = n21011 ^ n21010 ^ n21009 ;
  assign n21014 = n21013 ^ n21012 ^ n9643 ;
  assign n21015 = n15977 ^ n11084 ^ n4807 ;
  assign n21029 = ( ~n5970 & n6349 ) | ( ~n5970 & n14244 ) | ( n6349 & n14244 ) ;
  assign n21030 = n8318 & ~n21029 ;
  assign n21024 = n11083 ^ n9925 ^ n3980 ;
  assign n21025 = n21024 ^ n10973 ^ n972 ;
  assign n21026 = ( n484 & n1303 ) | ( n484 & n21025 ) | ( n1303 & n21025 ) ;
  assign n21022 = ( n2756 & ~n4229 ) | ( n2756 & n7521 ) | ( ~n4229 & n7521 ) ;
  assign n21021 = n8561 & n9455 ;
  assign n21023 = n21022 ^ n21021 ^ 1'b0 ;
  assign n21027 = n21026 ^ n21023 ^ n6886 ;
  assign n21028 = ( n7462 & ~n9537 ) | ( n7462 & n21027 ) | ( ~n9537 & n21027 ) ;
  assign n21016 = ( n716 & ~n725 ) | ( n716 & n3637 ) | ( ~n725 & n3637 ) ;
  assign n21017 = n21016 ^ n20811 ^ n1184 ;
  assign n21018 = n20071 & n21017 ;
  assign n21019 = n21018 ^ n11129 ^ n7711 ;
  assign n21020 = ( x3 & n5106 ) | ( x3 & n21019 ) | ( n5106 & n21019 ) ;
  assign n21031 = n21030 ^ n21028 ^ n21020 ;
  assign n21032 = ( n15691 & n18935 ) | ( n15691 & ~n21031 ) | ( n18935 & ~n21031 ) ;
  assign n21033 = n21032 ^ n19781 ^ x11 ;
  assign n21035 = n4917 ^ n3024 ^ n523 ;
  assign n21034 = n17215 ^ n5334 ^ n2349 ;
  assign n21036 = n21035 ^ n21034 ^ n18701 ;
  assign n21037 = n15674 & n21036 ;
  assign n21038 = n21037 ^ n1467 ^ 1'b0 ;
  assign n21039 = ( n1989 & n2978 ) | ( n1989 & ~n4005 ) | ( n2978 & ~n4005 ) ;
  assign n21040 = n21039 ^ n6714 ^ n2900 ;
  assign n21041 = ( ~n16125 & n16853 ) | ( ~n16125 & n21040 ) | ( n16853 & n21040 ) ;
  assign n21042 = ( n1598 & ~n5234 ) | ( n1598 & n11211 ) | ( ~n5234 & n11211 ) ;
  assign n21043 = ( n5361 & n9510 ) | ( n5361 & n21042 ) | ( n9510 & n21042 ) ;
  assign n21045 = n16438 ^ n7003 ^ n4236 ;
  assign n21044 = n10072 ^ n8374 ^ n6231 ;
  assign n21046 = n21045 ^ n21044 ^ n16129 ;
  assign n21050 = n8538 ^ n6427 ^ 1'b0 ;
  assign n21047 = ( n1549 & ~n1770 ) | ( n1549 & n5223 ) | ( ~n1770 & n5223 ) ;
  assign n21048 = n18532 ^ n7189 ^ n3680 ;
  assign n21049 = n21047 & n21048 ;
  assign n21051 = n21050 ^ n21049 ^ 1'b0 ;
  assign n21052 = n2385 & n11471 ;
  assign n21053 = n416 & n21052 ;
  assign n21054 = n21053 ^ n6747 ^ n3442 ;
  assign n21055 = n10535 | n11231 ;
  assign n21056 = n21055 ^ n13121 ^ n9750 ;
  assign n21057 = n21056 ^ n20717 ^ n16259 ;
  assign n21058 = ( n3379 & ~n9991 ) | ( n3379 & n11968 ) | ( ~n9991 & n11968 ) ;
  assign n21059 = ( n4663 & ~n4670 ) | ( n4663 & n9907 ) | ( ~n4670 & n9907 ) ;
  assign n21060 = n21059 ^ n11688 ^ 1'b0 ;
  assign n21063 = n8833 ^ n8761 ^ n3885 ;
  assign n21061 = ( n1204 & n4168 ) | ( n1204 & ~n7972 ) | ( n4168 & ~n7972 ) ;
  assign n21062 = n21061 ^ n18462 ^ n5809 ;
  assign n21064 = n21063 ^ n21062 ^ n4203 ;
  assign n21066 = ( ~n7793 & n11398 ) | ( ~n7793 & n17992 ) | ( n11398 & n17992 ) ;
  assign n21067 = ( n14238 & n16979 ) | ( n14238 & n21066 ) | ( n16979 & n21066 ) ;
  assign n21065 = n20597 ^ n17069 ^ n9854 ;
  assign n21068 = n21067 ^ n21065 ^ n16009 ;
  assign n21074 = n5025 | n5298 ;
  assign n21069 = ( ~n3367 & n4649 ) | ( ~n3367 & n17379 ) | ( n4649 & n17379 ) ;
  assign n21070 = ( n4769 & n12484 ) | ( n4769 & n21069 ) | ( n12484 & n21069 ) ;
  assign n21071 = ( ~n5766 & n19840 ) | ( ~n5766 & n21070 ) | ( n19840 & n21070 ) ;
  assign n21072 = ( n10316 & n17454 ) | ( n10316 & n21071 ) | ( n17454 & n21071 ) ;
  assign n21073 = ( n1837 & n19462 ) | ( n1837 & ~n21072 ) | ( n19462 & ~n21072 ) ;
  assign n21075 = n21074 ^ n21073 ^ n2217 ;
  assign n21076 = ( ~n2977 & n6275 ) | ( ~n2977 & n15059 ) | ( n6275 & n15059 ) ;
  assign n21077 = ( n7009 & n11673 ) | ( n7009 & n21076 ) | ( n11673 & n21076 ) ;
  assign n21078 = n3405 & ~n4925 ;
  assign n21079 = n21077 & n21078 ;
  assign n21080 = ( n16771 & n18660 ) | ( n16771 & n20825 ) | ( n18660 & n20825 ) ;
  assign n21081 = ( n3194 & ~n21079 ) | ( n3194 & n21080 ) | ( ~n21079 & n21080 ) ;
  assign n21082 = n15811 ^ n1355 ^ n538 ;
  assign n21083 = n21082 ^ n6039 ^ n5668 ;
  assign n21084 = ( n11991 & n12343 ) | ( n11991 & ~n21083 ) | ( n12343 & ~n21083 ) ;
  assign n21085 = n20606 ^ n14571 ^ 1'b0 ;
  assign n21086 = ~n18063 & n21085 ;
  assign n21087 = ( n950 & ~n10402 ) | ( n950 & n13242 ) | ( ~n10402 & n13242 ) ;
  assign n21088 = n21087 ^ n4243 ^ 1'b0 ;
  assign n21089 = n21088 ^ n13219 ^ n4989 ;
  assign n21090 = n21089 ^ n20289 ^ n19319 ;
  assign n21093 = ( n1620 & n3018 ) | ( n1620 & ~n6932 ) | ( n3018 & ~n6932 ) ;
  assign n21091 = n6637 ^ n3602 ^ n2595 ;
  assign n21092 = n10724 & n21091 ;
  assign n21094 = n21093 ^ n21092 ^ 1'b0 ;
  assign n21096 = ( n3457 & n7281 ) | ( n3457 & n16481 ) | ( n7281 & n16481 ) ;
  assign n21097 = ( ~n9494 & n17680 ) | ( ~n9494 & n21096 ) | ( n17680 & n21096 ) ;
  assign n21098 = ( n2728 & n3383 ) | ( n2728 & ~n8660 ) | ( n3383 & ~n8660 ) ;
  assign n21099 = ~n17284 & n21098 ;
  assign n21100 = ~n21097 & n21099 ;
  assign n21095 = n12669 ^ n12254 ^ n2954 ;
  assign n21101 = n21100 ^ n21095 ^ n4656 ;
  assign n21102 = n21101 ^ n13916 ^ n12512 ;
  assign n21103 = n2541 & n3828 ;
  assign n21104 = n13004 & n21103 ;
  assign n21105 = n1263 & n12190 ;
  assign n21106 = ( n6847 & n21104 ) | ( n6847 & ~n21105 ) | ( n21104 & ~n21105 ) ;
  assign n21107 = n21106 ^ n20810 ^ 1'b0 ;
  assign n21108 = n9543 | n21107 ;
  assign n21109 = ( n6801 & n19069 ) | ( n6801 & ~n21108 ) | ( n19069 & ~n21108 ) ;
  assign n21110 = ( n1408 & n4110 ) | ( n1408 & n6837 ) | ( n4110 & n6837 ) ;
  assign n21119 = ( x29 & n5083 ) | ( x29 & ~n5194 ) | ( n5083 & ~n5194 ) ;
  assign n21117 = ( n433 & n3106 ) | ( n433 & ~n5419 ) | ( n3106 & ~n5419 ) ;
  assign n21115 = n9472 ^ n5107 ^ n2945 ;
  assign n21111 = ( ~x28 & n2441 ) | ( ~x28 & n20589 ) | ( n2441 & n20589 ) ;
  assign n21112 = n21111 ^ n5624 ^ n2138 ;
  assign n21113 = n14769 | n21112 ;
  assign n21114 = n21113 ^ n3316 ^ 1'b0 ;
  assign n21116 = n21115 ^ n21114 ^ n1170 ;
  assign n21118 = n21117 ^ n21116 ^ n3689 ;
  assign n21120 = n21119 ^ n21118 ^ n18520 ;
  assign n21121 = ( n19501 & n21110 ) | ( n19501 & ~n21120 ) | ( n21110 & ~n21120 ) ;
  assign n21122 = n19537 ^ n12824 ^ 1'b0 ;
  assign n21123 = ~n10169 & n21122 ;
  assign n21124 = ~n7610 & n21123 ;
  assign n21125 = ( ~n985 & n5606 ) | ( ~n985 & n11513 ) | ( n5606 & n11513 ) ;
  assign n21126 = n4937 | n10379 ;
  assign n21127 = n21126 ^ n8231 ^ 1'b0 ;
  assign n21128 = ~n16660 & n20545 ;
  assign n21129 = n7554 & n21128 ;
  assign n21130 = ( n11420 & n21127 ) | ( n11420 & ~n21129 ) | ( n21127 & ~n21129 ) ;
  assign n21131 = n5878 ^ n1572 ^ x63 ;
  assign n21132 = ( n6297 & n7510 ) | ( n6297 & ~n21131 ) | ( n7510 & ~n21131 ) ;
  assign n21133 = n13898 ^ n6579 ^ n1537 ;
  assign n21134 = ( n6105 & ~n13987 ) | ( n6105 & n16243 ) | ( ~n13987 & n16243 ) ;
  assign n21135 = ( ~n21132 & n21133 ) | ( ~n21132 & n21134 ) | ( n21133 & n21134 ) ;
  assign n21136 = ( ~n21125 & n21130 ) | ( ~n21125 & n21135 ) | ( n21130 & n21135 ) ;
  assign n21137 = ( ~n7769 & n8387 ) | ( ~n7769 & n21136 ) | ( n8387 & n21136 ) ;
  assign n21139 = n7526 & ~n15087 ;
  assign n21140 = n21139 ^ n7607 ^ 1'b0 ;
  assign n21138 = n18753 ^ n11945 ^ n2609 ;
  assign n21141 = n21140 ^ n21138 ^ n20893 ;
  assign n21142 = ( n1805 & n2712 ) | ( n1805 & ~n5235 ) | ( n2712 & ~n5235 ) ;
  assign n21143 = ( n3469 & n9283 ) | ( n3469 & n21142 ) | ( n9283 & n21142 ) ;
  assign n21144 = n5575 & ~n6513 ;
  assign n21145 = ( n1448 & n5408 ) | ( n1448 & n21144 ) | ( n5408 & n21144 ) ;
  assign n21146 = ~n6722 & n21145 ;
  assign n21147 = ( ~n20862 & n21143 ) | ( ~n20862 & n21146 ) | ( n21143 & n21146 ) ;
  assign n21154 = n11490 ^ n1957 ^ 1'b0 ;
  assign n21148 = n3365 ^ n1831 ^ 1'b0 ;
  assign n21149 = n624 & n21148 ;
  assign n21150 = n5564 ^ n3811 ^ n2572 ;
  assign n21151 = ( n1060 & ~n9821 ) | ( n1060 & n21150 ) | ( ~n9821 & n21150 ) ;
  assign n21152 = n21151 ^ n13438 ^ 1'b0 ;
  assign n21153 = n21149 & ~n21152 ;
  assign n21155 = n21154 ^ n21153 ^ n19351 ;
  assign n21156 = n1210 ^ n1160 ^ n871 ;
  assign n21157 = n21156 ^ n21028 ^ n18378 ;
  assign n21160 = n13097 ^ n10814 ^ n5515 ;
  assign n21158 = ( n8935 & ~n14190 ) | ( n8935 & n15059 ) | ( ~n14190 & n15059 ) ;
  assign n21159 = ( x101 & ~n20702 ) | ( x101 & n21158 ) | ( ~n20702 & n21158 ) ;
  assign n21161 = n21160 ^ n21159 ^ n5940 ;
  assign n21163 = n8929 | n19893 ;
  assign n21164 = n6254 & ~n21163 ;
  assign n21162 = n17505 ^ n10478 ^ n2305 ;
  assign n21165 = n21164 ^ n21162 ^ n15993 ;
  assign n21170 = n4379 ^ n729 ^ 1'b0 ;
  assign n21171 = ~n3731 & n21170 ;
  assign n21172 = ( n9040 & n15852 ) | ( n9040 & ~n21171 ) | ( n15852 & ~n21171 ) ;
  assign n21168 = ( ~n2001 & n2543 ) | ( ~n2001 & n8561 ) | ( n2543 & n8561 ) ;
  assign n21166 = ( n7828 & ~n9668 ) | ( n7828 & n17276 ) | ( ~n9668 & n17276 ) ;
  assign n21167 = n21166 ^ n2106 ^ n590 ;
  assign n21169 = n21168 ^ n21167 ^ n6593 ;
  assign n21173 = n21172 ^ n21169 ^ n20584 ;
  assign n21174 = n13076 ^ n12207 ^ n2675 ;
  assign n21183 = n20968 ^ n2245 ^ n1267 ;
  assign n21184 = n21183 ^ n5195 ^ n1465 ;
  assign n21180 = n2342 ^ n1577 ^ n981 ;
  assign n21181 = n9384 ^ n5240 ^ n3112 ;
  assign n21182 = ( n12896 & n21180 ) | ( n12896 & n21181 ) | ( n21180 & n21181 ) ;
  assign n21185 = n21184 ^ n21182 ^ n17571 ;
  assign n21178 = ( n10292 & n12801 ) | ( n10292 & ~n18818 ) | ( n12801 & ~n18818 ) ;
  assign n21175 = n8603 ^ n3217 ^ n2943 ;
  assign n21176 = ( n513 & n868 ) | ( n513 & n14708 ) | ( n868 & n14708 ) ;
  assign n21177 = n21175 & n21176 ;
  assign n21179 = n21178 ^ n21177 ^ 1'b0 ;
  assign n21186 = n21185 ^ n21179 ^ n4309 ;
  assign n21187 = ( ~n989 & n8585 ) | ( ~n989 & n16524 ) | ( n8585 & n16524 ) ;
  assign n21188 = n21187 ^ n17312 ^ n6467 ;
  assign n21189 = n6733 ^ n6288 ^ n1298 ;
  assign n21190 = n12162 ^ n6508 ^ n473 ;
  assign n21191 = n15437 ^ x230 ^ 1'b0 ;
  assign n21192 = n7502 | n21191 ;
  assign n21193 = ( ~n1050 & n12013 ) | ( ~n1050 & n21192 ) | ( n12013 & n21192 ) ;
  assign n21194 = n21193 ^ n14748 ^ 1'b0 ;
  assign n21195 = n21190 | n21194 ;
  assign n21196 = n18288 ^ n5289 ^ n1881 ;
  assign n21197 = ( ~n2014 & n21195 ) | ( ~n2014 & n21196 ) | ( n21195 & n21196 ) ;
  assign n21199 = n21047 ^ n11814 ^ n9496 ;
  assign n21198 = n14363 ^ n6149 ^ x80 ;
  assign n21200 = n21199 ^ n21198 ^ n6040 ;
  assign n21201 = n21200 ^ n11430 ^ n10205 ;
  assign n21202 = n10466 ^ n7243 ^ n4989 ;
  assign n21203 = ( n4174 & n20931 ) | ( n4174 & n21202 ) | ( n20931 & n21202 ) ;
  assign n21204 = n16228 ^ n9574 ^ 1'b0 ;
  assign n21205 = ( n1755 & ~n6033 ) | ( n1755 & n11318 ) | ( ~n6033 & n11318 ) ;
  assign n21206 = n11205 ^ n6161 ^ n3801 ;
  assign n21207 = n15144 ^ n15034 ^ n9918 ;
  assign n21208 = n21207 ^ n10938 ^ n968 ;
  assign n21209 = ( n3616 & n4618 ) | ( n3616 & ~n21208 ) | ( n4618 & ~n21208 ) ;
  assign n21210 = n21209 ^ n15135 ^ n3326 ;
  assign n21211 = ( n4923 & n21206 ) | ( n4923 & ~n21210 ) | ( n21206 & ~n21210 ) ;
  assign n21212 = n9028 ^ n1896 ^ x116 ;
  assign n21213 = n21212 ^ n13391 ^ n2875 ;
  assign n21214 = ( x76 & n1484 ) | ( x76 & ~n21213 ) | ( n1484 & ~n21213 ) ;
  assign n21215 = ( n8272 & n12903 ) | ( n8272 & n21214 ) | ( n12903 & n21214 ) ;
  assign n21216 = n21215 ^ n17946 ^ n11508 ;
  assign n21217 = n8592 ^ n7930 ^ 1'b0 ;
  assign n21218 = ( n2035 & n8384 ) | ( n2035 & n10752 ) | ( n8384 & n10752 ) ;
  assign n21219 = n9757 ^ n4667 ^ n1188 ;
  assign n21220 = n7750 ^ n3477 ^ 1'b0 ;
  assign n21221 = n11614 ^ n3266 ^ x13 ;
  assign n21222 = n4895 & n14766 ;
  assign n21224 = n4921 | n12822 ;
  assign n21223 = n8772 ^ n3977 ^ n2190 ;
  assign n21225 = n21224 ^ n21223 ^ 1'b0 ;
  assign n21226 = n21222 | n21225 ;
  assign n21227 = ( ~n4686 & n21221 ) | ( ~n4686 & n21226 ) | ( n21221 & n21226 ) ;
  assign n21228 = ( n21219 & ~n21220 ) | ( n21219 & n21227 ) | ( ~n21220 & n21227 ) ;
  assign n21229 = ( n4621 & n21218 ) | ( n4621 & ~n21228 ) | ( n21218 & ~n21228 ) ;
  assign n21231 = ( ~n4635 & n4994 ) | ( ~n4635 & n6680 ) | ( n4994 & n6680 ) ;
  assign n21232 = ( ~n2859 & n13087 ) | ( ~n2859 & n21231 ) | ( n13087 & n21231 ) ;
  assign n21230 = n5040 | n7242 ;
  assign n21233 = n21232 ^ n21230 ^ 1'b0 ;
  assign n21234 = ( n835 & n12720 ) | ( n835 & n18430 ) | ( n12720 & n18430 ) ;
  assign n21235 = n21234 ^ n10625 ^ n7912 ;
  assign n21236 = n18239 ^ n4697 ^ 1'b0 ;
  assign n21237 = n6824 | n21236 ;
  assign n21238 = ( n1681 & n14292 ) | ( n1681 & ~n18713 ) | ( n14292 & ~n18713 ) ;
  assign n21239 = n8679 & n19500 ;
  assign n21240 = n12891 ^ n5909 ^ n2380 ;
  assign n21241 = n21239 | n21240 ;
  assign n21242 = n21241 ^ n20041 ^ n9096 ;
  assign n21243 = ( x191 & n2932 ) | ( x191 & ~n6550 ) | ( n2932 & ~n6550 ) ;
  assign n21244 = n2456 & n21243 ;
  assign n21245 = ~n11657 & n21244 ;
  assign n21246 = n21245 ^ n5489 ^ n1859 ;
  assign n21250 = n16337 ^ n9342 ^ n5722 ;
  assign n21252 = ( n567 & n2778 ) | ( n567 & n9780 ) | ( n2778 & n9780 ) ;
  assign n21253 = ( n1368 & n8388 ) | ( n1368 & ~n21252 ) | ( n8388 & ~n21252 ) ;
  assign n21251 = ( n546 & n10882 ) | ( n546 & ~n14539 ) | ( n10882 & ~n14539 ) ;
  assign n21254 = n21253 ^ n21251 ^ n3904 ;
  assign n21255 = ( n20536 & n21250 ) | ( n20536 & n21254 ) | ( n21250 & n21254 ) ;
  assign n21247 = n2586 ^ x194 ^ 1'b0 ;
  assign n21248 = n21210 & n21247 ;
  assign n21249 = ( n662 & ~n16576 ) | ( n662 & n21248 ) | ( ~n16576 & n21248 ) ;
  assign n21256 = n21255 ^ n21249 ^ n11663 ;
  assign n21257 = ( ~n12178 & n21246 ) | ( ~n12178 & n21256 ) | ( n21246 & n21256 ) ;
  assign n21258 = ( n21190 & n21242 ) | ( n21190 & n21257 ) | ( n21242 & n21257 ) ;
  assign n21259 = ( n9489 & ~n21238 ) | ( n9489 & n21258 ) | ( ~n21238 & n21258 ) ;
  assign n21260 = n14029 ^ n5943 ^ n343 ;
  assign n21261 = n21260 ^ n17079 ^ n5779 ;
  assign n21262 = n7658 ^ n6022 ^ n5279 ;
  assign n21263 = ( n644 & n8159 ) | ( n644 & n21262 ) | ( n8159 & n21262 ) ;
  assign n21264 = n19844 ^ n13714 ^ n2084 ;
  assign n21266 = n4123 ^ n1295 ^ n766 ;
  assign n21265 = ( ~x161 & n7223 ) | ( ~x161 & n18734 ) | ( n7223 & n18734 ) ;
  assign n21267 = n21266 ^ n21265 ^ n8335 ;
  assign n21268 = ( ~n13178 & n21264 ) | ( ~n13178 & n21267 ) | ( n21264 & n21267 ) ;
  assign n21289 = ( ~n2219 & n2705 ) | ( ~n2219 & n5587 ) | ( n2705 & n5587 ) ;
  assign n21287 = n15189 ^ n10065 ^ n580 ;
  assign n21282 = ( ~x226 & n2844 ) | ( ~x226 & n19706 ) | ( n2844 & n19706 ) ;
  assign n21283 = n16802 ^ n10495 ^ n3417 ;
  assign n21284 = ( n16332 & n21282 ) | ( n16332 & n21283 ) | ( n21282 & n21283 ) ;
  assign n21285 = n21284 ^ n16312 ^ 1'b0 ;
  assign n21286 = n13226 & ~n21285 ;
  assign n21288 = n21287 ^ n21286 ^ n4100 ;
  assign n21279 = n569 | n11095 ;
  assign n21280 = ( n12108 & ~n13443 ) | ( n12108 & n21279 ) | ( ~n13443 & n21279 ) ;
  assign n21274 = n6348 ^ n5056 ^ n308 ;
  assign n21275 = ~n17436 & n21274 ;
  assign n21276 = n21275 ^ n8725 ^ n3502 ;
  assign n21277 = n10234 & ~n21276 ;
  assign n21278 = n21277 ^ n7247 ^ 1'b0 ;
  assign n21269 = n3925 & n6191 ;
  assign n21270 = ~n4792 & n21269 ;
  assign n21271 = ( n6007 & n8000 ) | ( n6007 & n21270 ) | ( n8000 & n21270 ) ;
  assign n21272 = n21271 ^ n6193 ^ 1'b0 ;
  assign n21273 = n3461 & ~n21272 ;
  assign n21281 = n21280 ^ n21278 ^ n21273 ;
  assign n21290 = n21289 ^ n21288 ^ n21281 ;
  assign n21291 = ( ~n1348 & n12571 ) | ( ~n1348 & n14238 ) | ( n12571 & n14238 ) ;
  assign n21292 = n21291 ^ n12690 ^ n3471 ;
  assign n21293 = n21292 ^ n18535 ^ n10910 ;
  assign n21294 = n4331 | n21293 ;
  assign n21295 = n5073 ^ n3008 ^ 1'b0 ;
  assign n21296 = ~n5940 & n8412 ;
  assign n21297 = n21296 ^ n18237 ^ 1'b0 ;
  assign n21298 = ( ~n2214 & n16326 ) | ( ~n2214 & n21297 ) | ( n16326 & n21297 ) ;
  assign n21299 = ( n4358 & n4703 ) | ( n4358 & n8289 ) | ( n4703 & n8289 ) ;
  assign n21300 = ( n5077 & n10394 ) | ( n5077 & n19989 ) | ( n10394 & n19989 ) ;
  assign n21301 = ( n16109 & n21299 ) | ( n16109 & n21300 ) | ( n21299 & n21300 ) ;
  assign n21302 = ( ~n17343 & n21298 ) | ( ~n17343 & n21301 ) | ( n21298 & n21301 ) ;
  assign n21303 = n17816 ^ n12664 ^ n3828 ;
  assign n21304 = ( n8403 & n17659 ) | ( n8403 & ~n21303 ) | ( n17659 & ~n21303 ) ;
  assign n21305 = ( ~n3358 & n11672 ) | ( ~n3358 & n12093 ) | ( n11672 & n12093 ) ;
  assign n21306 = n8707 & n19306 ;
  assign n21307 = n21287 ^ n15438 ^ 1'b0 ;
  assign n21308 = n10244 ^ n5988 ^ 1'b0 ;
  assign n21309 = n21307 | n21308 ;
  assign n21310 = n19525 & ~n21309 ;
  assign n21311 = n21310 ^ n12519 ^ n4021 ;
  assign n21313 = ( n5662 & ~n6324 ) | ( n5662 & n11406 ) | ( ~n6324 & n11406 ) ;
  assign n21314 = n5141 ^ n4564 ^ n1927 ;
  assign n21315 = n21314 ^ n20020 ^ n6524 ;
  assign n21316 = n21315 ^ n13885 ^ n6983 ;
  assign n21317 = ( n20503 & n21313 ) | ( n20503 & n21316 ) | ( n21313 & n21316 ) ;
  assign n21312 = n11524 ^ n3339 ^ 1'b0 ;
  assign n21318 = n21317 ^ n21312 ^ n16915 ;
  assign n21319 = n3691 & n3809 ;
  assign n21320 = ~n3471 & n21319 ;
  assign n21321 = n16610 ^ n11575 ^ n6952 ;
  assign n21322 = ( n19272 & n21320 ) | ( n19272 & n21321 ) | ( n21320 & n21321 ) ;
  assign n21323 = n21322 ^ n3799 ^ n2407 ;
  assign n21324 = ( n8752 & n8811 ) | ( n8752 & n11398 ) | ( n8811 & n11398 ) ;
  assign n21325 = n18876 ^ n18448 ^ n9298 ;
  assign n21326 = ( n745 & ~n888 ) | ( n745 & n4846 ) | ( ~n888 & n4846 ) ;
  assign n21327 = n21326 ^ n10524 ^ n1225 ;
  assign n21328 = n10884 | n21327 ;
  assign n21329 = n21325 & ~n21328 ;
  assign n21330 = n21329 ^ n17221 ^ n6984 ;
  assign n21331 = ( n15937 & ~n21324 ) | ( n15937 & n21330 ) | ( ~n21324 & n21330 ) ;
  assign n21335 = n18344 ^ n16505 ^ n2668 ;
  assign n21336 = ( n2275 & ~n9530 ) | ( n2275 & n21335 ) | ( ~n9530 & n21335 ) ;
  assign n21337 = n8628 ^ n2526 ^ x146 ;
  assign n21338 = ( n17044 & n20104 ) | ( n17044 & ~n21337 ) | ( n20104 & ~n21337 ) ;
  assign n21339 = n21338 ^ n20144 ^ n8618 ;
  assign n21340 = n21339 ^ n9220 ^ 1'b0 ;
  assign n21341 = ( n16397 & ~n21336 ) | ( n16397 & n21340 ) | ( ~n21336 & n21340 ) ;
  assign n21332 = x51 & ~n4652 ;
  assign n21333 = n21332 ^ n17458 ^ 1'b0 ;
  assign n21334 = ( n2000 & n17413 ) | ( n2000 & ~n21333 ) | ( n17413 & ~n21333 ) ;
  assign n21342 = n21341 ^ n21334 ^ 1'b0 ;
  assign n21343 = n3522 ^ n1448 ^ n1148 ;
  assign n21344 = ( n6812 & ~n13120 ) | ( n6812 & n21343 ) | ( ~n13120 & n21343 ) ;
  assign n21345 = n4259 ^ n3263 ^ n3016 ;
  assign n21346 = n4842 & n8288 ;
  assign n21347 = ( n18612 & ~n21345 ) | ( n18612 & n21346 ) | ( ~n21345 & n21346 ) ;
  assign n21348 = n2856 ^ n2379 ^ n294 ;
  assign n21349 = n21348 ^ n2399 ^ 1'b0 ;
  assign n21350 = ~n14109 & n21349 ;
  assign n21351 = ( x238 & n7527 ) | ( x238 & ~n11424 ) | ( n7527 & ~n11424 ) ;
  assign n21352 = n21351 ^ n18492 ^ n2333 ;
  assign n21353 = ( n1874 & n2305 ) | ( n1874 & ~n12453 ) | ( n2305 & ~n12453 ) ;
  assign n21354 = ~n3022 & n12901 ;
  assign n21355 = n18474 & n21354 ;
  assign n21356 = ( n10849 & n21353 ) | ( n10849 & n21355 ) | ( n21353 & n21355 ) ;
  assign n21357 = n21356 ^ n8500 ^ n7549 ;
  assign n21358 = n21357 ^ n19650 ^ n16985 ;
  assign n21365 = ( n475 & n1329 ) | ( n475 & n11199 ) | ( n1329 & n11199 ) ;
  assign n21366 = n21365 ^ n11662 ^ 1'b0 ;
  assign n21367 = n7992 & ~n21366 ;
  assign n21368 = n21367 ^ n7233 ^ n2805 ;
  assign n21362 = n13209 & n17364 ;
  assign n21363 = n2104 & n21362 ;
  assign n21364 = ( n4588 & n11919 ) | ( n4588 & n21363 ) | ( n11919 & n21363 ) ;
  assign n21360 = ( n10267 & ~n18500 ) | ( n10267 & n19110 ) | ( ~n18500 & n19110 ) ;
  assign n21359 = ( n3962 & n5951 ) | ( n3962 & ~n9355 ) | ( n5951 & ~n9355 ) ;
  assign n21361 = n21360 ^ n21359 ^ n17913 ;
  assign n21369 = n21368 ^ n21364 ^ n21361 ;
  assign n21370 = n13612 ^ n5633 ^ n5609 ;
  assign n21371 = n21370 ^ n11357 ^ n4677 ;
  assign n21372 = n8984 & ~n21371 ;
  assign n21373 = n5667 ^ n3886 ^ n1519 ;
  assign n21374 = ( n2234 & n3213 ) | ( n2234 & ~n8269 ) | ( n3213 & ~n8269 ) ;
  assign n21375 = ( n9781 & n21373 ) | ( n9781 & n21374 ) | ( n21373 & n21374 ) ;
  assign n21376 = ( n4122 & n13270 ) | ( n4122 & n21375 ) | ( n13270 & n21375 ) ;
  assign n21377 = ( n4220 & ~n5347 ) | ( n4220 & n9886 ) | ( ~n5347 & n9886 ) ;
  assign n21378 = n21377 ^ n4549 ^ n4289 ;
  assign n21381 = n828 & ~n12035 ;
  assign n21382 = n21381 ^ n5489 ^ 1'b0 ;
  assign n21379 = n21142 ^ n9375 ^ n3541 ;
  assign n21380 = n1818 | n21379 ;
  assign n21383 = n21382 ^ n21380 ^ 1'b0 ;
  assign n21384 = n9958 & n21383 ;
  assign n21385 = n15821 & n21384 ;
  assign n21386 = ( n1182 & n7627 ) | ( n1182 & n13132 ) | ( n7627 & n13132 ) ;
  assign n21387 = ( n5705 & n11810 ) | ( n5705 & n21386 ) | ( n11810 & n21386 ) ;
  assign n21393 = ~n1098 & n3524 ;
  assign n21394 = ( n1033 & n1170 ) | ( n1033 & ~n16320 ) | ( n1170 & ~n16320 ) ;
  assign n21395 = ( n1864 & ~n21393 ) | ( n1864 & n21394 ) | ( ~n21393 & n21394 ) ;
  assign n21388 = n16038 ^ n9382 ^ n5885 ;
  assign n21390 = n12505 ^ n2852 ^ n2373 ;
  assign n21389 = n9274 & ~n19820 ;
  assign n21391 = n21390 ^ n21389 ^ 1'b0 ;
  assign n21392 = ( n741 & n21388 ) | ( n741 & n21391 ) | ( n21388 & n21391 ) ;
  assign n21396 = n21395 ^ n21392 ^ n7100 ;
  assign n21397 = ( n9685 & ~n14384 ) | ( n9685 & n21396 ) | ( ~n14384 & n21396 ) ;
  assign n21398 = n16250 ^ n2865 ^ 1'b0 ;
  assign n21399 = n5185 | n21398 ;
  assign n21400 = n21399 ^ n16825 ^ n4643 ;
  assign n21401 = n17631 ^ n12074 ^ n3332 ;
  assign n21402 = ~n5680 & n12324 ;
  assign n21403 = n19343 ^ n9251 ^ n773 ;
  assign n21404 = ( n9174 & n15022 ) | ( n9174 & n21403 ) | ( n15022 & n21403 ) ;
  assign n21405 = ( n3309 & ~n6951 ) | ( n3309 & n14876 ) | ( ~n6951 & n14876 ) ;
  assign n21406 = ( n21402 & n21404 ) | ( n21402 & ~n21405 ) | ( n21404 & ~n21405 ) ;
  assign n21409 = n18461 ^ n4161 ^ n740 ;
  assign n21410 = n18832 ^ n8029 ^ 1'b0 ;
  assign n21411 = ~n699 & n21410 ;
  assign n21412 = ( ~n4055 & n12818 ) | ( ~n4055 & n21411 ) | ( n12818 & n21411 ) ;
  assign n21413 = ~n21409 & n21412 ;
  assign n21407 = ( n5151 & ~n5670 ) | ( n5151 & n6621 ) | ( ~n5670 & n6621 ) ;
  assign n21408 = n21407 ^ n10195 ^ n3073 ;
  assign n21414 = n21413 ^ n21408 ^ 1'b0 ;
  assign n21415 = ( n1246 & n14867 ) | ( n1246 & ~n16288 ) | ( n14867 & ~n16288 ) ;
  assign n21416 = ( n11007 & n12655 ) | ( n11007 & n21415 ) | ( n12655 & n21415 ) ;
  assign n21417 = n21416 ^ n18281 ^ n3097 ;
  assign n21418 = n8109 & ~n15447 ;
  assign n21419 = ( n4592 & n12395 ) | ( n4592 & n14726 ) | ( n12395 & n14726 ) ;
  assign n21420 = ( n2336 & n18296 ) | ( n2336 & ~n21419 ) | ( n18296 & ~n21419 ) ;
  assign n21422 = n13012 ^ n9025 ^ n4665 ;
  assign n21423 = n6767 ^ n1213 ^ 1'b0 ;
  assign n21424 = n21422 & ~n21423 ;
  assign n21421 = ( n4115 & n4622 ) | ( n4115 & n9206 ) | ( n4622 & n9206 ) ;
  assign n21425 = n21424 ^ n21421 ^ 1'b0 ;
  assign n21426 = ( n7296 & n16192 ) | ( n7296 & ~n18557 ) | ( n16192 & ~n18557 ) ;
  assign n21427 = n5971 & n18433 ;
  assign n21428 = ( ~n1937 & n16289 ) | ( ~n1937 & n21427 ) | ( n16289 & n21427 ) ;
  assign n21429 = n21428 ^ n3781 ^ n2700 ;
  assign n21430 = n11596 ^ n6665 ^ n4562 ;
  assign n21431 = ( n14041 & n16764 ) | ( n14041 & ~n21430 ) | ( n16764 & ~n21430 ) ;
  assign n21432 = ( n8699 & n19313 ) | ( n8699 & ~n21431 ) | ( n19313 & ~n21431 ) ;
  assign n21433 = ( n2391 & ~n3140 ) | ( n2391 & n10305 ) | ( ~n3140 & n10305 ) ;
  assign n21434 = ~n21432 & n21433 ;
  assign n21435 = x19 & n21434 ;
  assign n21436 = n14287 ^ n2051 ^ n687 ;
  assign n21437 = n18956 ^ n18764 ^ n2822 ;
  assign n21438 = n19404 ^ n6766 ^ 1'b0 ;
  assign n21439 = ( n21436 & ~n21437 ) | ( n21436 & n21438 ) | ( ~n21437 & n21438 ) ;
  assign n21440 = n9155 ^ n2140 ^ 1'b0 ;
  assign n21441 = n15847 & ~n21440 ;
  assign n21442 = n20818 ^ n15313 ^ 1'b0 ;
  assign n21443 = ( ~n9423 & n21441 ) | ( ~n9423 & n21442 ) | ( n21441 & n21442 ) ;
  assign n21449 = n4965 ^ n4371 ^ n810 ;
  assign n21445 = ( n4091 & ~n4373 ) | ( n4091 & n14365 ) | ( ~n4373 & n14365 ) ;
  assign n21446 = n13484 ^ n2408 ^ 1'b0 ;
  assign n21447 = ( n4892 & n21445 ) | ( n4892 & ~n21446 ) | ( n21445 & ~n21446 ) ;
  assign n21448 = n21447 ^ n20369 ^ n16805 ;
  assign n21450 = n21449 ^ n21448 ^ n6367 ;
  assign n21444 = n2899 & n20835 ;
  assign n21451 = n21450 ^ n21444 ^ 1'b0 ;
  assign n21452 = n7270 & n9149 ;
  assign n21453 = ~n21451 & n21452 ;
  assign n21454 = n9611 & ~n10904 ;
  assign n21455 = n21454 ^ n12575 ^ n8353 ;
  assign n21458 = n19270 ^ n4720 ^ n3962 ;
  assign n21456 = n6809 ^ n669 ^ 1'b0 ;
  assign n21457 = n11290 & ~n21456 ;
  assign n21459 = n21458 ^ n21457 ^ n20708 ;
  assign n21460 = n1263 & n3392 ;
  assign n21461 = n21460 ^ n14533 ^ 1'b0 ;
  assign n21462 = n13786 & n16189 ;
  assign n21463 = ( n690 & n3564 ) | ( n690 & n8056 ) | ( n3564 & n8056 ) ;
  assign n21464 = n21463 ^ n17051 ^ n9141 ;
  assign n21465 = n5592 ^ n4615 ^ n3868 ;
  assign n21466 = ( n6973 & n12003 ) | ( n6973 & ~n15101 ) | ( n12003 & ~n15101 ) ;
  assign n21467 = n21466 ^ n12685 ^ 1'b0 ;
  assign n21468 = n21465 | n21467 ;
  assign n21469 = n21468 ^ n18700 ^ n11007 ;
  assign n21470 = n16002 ^ n4810 ^ n3705 ;
  assign n21471 = n21470 ^ n8257 ^ n5221 ;
  assign n21472 = ( n720 & ~n1122 ) | ( n720 & n9541 ) | ( ~n1122 & n9541 ) ;
  assign n21473 = ( ~n13719 & n21471 ) | ( ~n13719 & n21472 ) | ( n21471 & n21472 ) ;
  assign n21474 = ( ~n3954 & n4300 ) | ( ~n3954 & n7511 ) | ( n4300 & n7511 ) ;
  assign n21475 = ( n1822 & ~n3054 ) | ( n1822 & n21474 ) | ( ~n3054 & n21474 ) ;
  assign n21476 = ( ~n14710 & n15093 ) | ( ~n14710 & n20572 ) | ( n15093 & n20572 ) ;
  assign n21477 = ( ~n261 & n5862 ) | ( ~n261 & n15711 ) | ( n5862 & n15711 ) ;
  assign n21478 = n6891 & ~n19312 ;
  assign n21479 = n19961 ^ n14654 ^ x35 ;
  assign n21480 = ( n21477 & n21478 ) | ( n21477 & ~n21479 ) | ( n21478 & ~n21479 ) ;
  assign n21481 = ( ~n3768 & n4934 ) | ( ~n3768 & n9213 ) | ( n4934 & n9213 ) ;
  assign n21482 = ( n4983 & n6639 ) | ( n4983 & n10228 ) | ( n6639 & n10228 ) ;
  assign n21483 = n21482 ^ n13729 ^ n1016 ;
  assign n21485 = ( n4127 & n5903 ) | ( n4127 & n10482 ) | ( n5903 & n10482 ) ;
  assign n21484 = n3762 | n11740 ;
  assign n21486 = n21485 ^ n21484 ^ 1'b0 ;
  assign n21487 = n7846 & n10705 ;
  assign n21488 = n21487 ^ n18125 ^ 1'b0 ;
  assign n21489 = n21488 ^ n15223 ^ 1'b0 ;
  assign n21490 = ( n2157 & n6259 ) | ( n2157 & ~n21489 ) | ( n6259 & ~n21489 ) ;
  assign n21491 = ( n21483 & n21486 ) | ( n21483 & n21490 ) | ( n21486 & n21490 ) ;
  assign n21492 = ( n2976 & n9572 ) | ( n2976 & ~n10809 ) | ( n9572 & ~n10809 ) ;
  assign n21500 = n18263 ^ n9905 ^ 1'b0 ;
  assign n21501 = n5525 & ~n21500 ;
  assign n21502 = ( ~n12470 & n17893 ) | ( ~n12470 & n21501 ) | ( n17893 & n21501 ) ;
  assign n21503 = n8182 ^ n5203 ^ n758 ;
  assign n21504 = ~n12973 & n21503 ;
  assign n21505 = ~n21502 & n21504 ;
  assign n21493 = ( n10355 & n18892 ) | ( n10355 & n19026 ) | ( n18892 & n19026 ) ;
  assign n21494 = n21493 ^ n7459 ^ n3641 ;
  assign n21495 = n13175 | n21494 ;
  assign n21496 = n1794 & ~n21495 ;
  assign n21497 = ( n4586 & ~n6076 ) | ( n4586 & n14405 ) | ( ~n6076 & n14405 ) ;
  assign n21498 = n21497 ^ n20101 ^ n2585 ;
  assign n21499 = ~n21496 & n21498 ;
  assign n21506 = n21505 ^ n21499 ^ 1'b0 ;
  assign n21507 = n20829 ^ n10147 ^ n10130 ;
  assign n21508 = n21507 ^ n10115 ^ n9911 ;
  assign n21509 = ( n4275 & ~n5458 ) | ( n4275 & n21508 ) | ( ~n5458 & n21508 ) ;
  assign n21510 = n16411 ^ n13843 ^ n2731 ;
  assign n21511 = ( n7573 & n13962 ) | ( n7573 & ~n19825 ) | ( n13962 & ~n19825 ) ;
  assign n21512 = ( n16002 & ~n21326 ) | ( n16002 & n21511 ) | ( ~n21326 & n21511 ) ;
  assign n21513 = n922 | n6347 ;
  assign n21514 = n21513 ^ n14274 ^ n4070 ;
  assign n21515 = ( n266 & ~n13612 ) | ( n266 & n13984 ) | ( ~n13612 & n13984 ) ;
  assign n21516 = n21515 ^ n12474 ^ n12205 ;
  assign n21517 = n2222 & n21516 ;
  assign n21518 = ~n21514 & n21517 ;
  assign n21519 = ( n1464 & n2871 ) | ( n1464 & ~n21518 ) | ( n2871 & ~n21518 ) ;
  assign n21520 = n20052 ^ n19112 ^ n13340 ;
  assign n21521 = ( n2331 & ~n9625 ) | ( n2331 & n10134 ) | ( ~n9625 & n10134 ) ;
  assign n21523 = n3596 ^ n3210 ^ n3164 ;
  assign n21524 = ( n16595 & n20676 ) | ( n16595 & ~n21523 ) | ( n20676 & ~n21523 ) ;
  assign n21522 = n2992 | n7124 ;
  assign n21525 = n21524 ^ n21522 ^ n12789 ;
  assign n21526 = n21525 ^ n18937 ^ n10079 ;
  assign n21527 = ( n6519 & n21521 ) | ( n6519 & n21526 ) | ( n21521 & n21526 ) ;
  assign n21528 = ( n2125 & n17658 ) | ( n2125 & ~n20521 ) | ( n17658 & ~n20521 ) ;
  assign n21529 = n19320 ^ n5329 ^ 1'b0 ;
  assign n21530 = ( n4674 & n6579 ) | ( n4674 & n21529 ) | ( n6579 & n21529 ) ;
  assign n21531 = ( n2258 & n8104 ) | ( n2258 & n13566 ) | ( n8104 & n13566 ) ;
  assign n21532 = ( n15001 & ~n20780 ) | ( n15001 & n21531 ) | ( ~n20780 & n21531 ) ;
  assign n21533 = ( n2000 & ~n7596 ) | ( n2000 & n16048 ) | ( ~n7596 & n16048 ) ;
  assign n21534 = n8313 ^ n3685 ^ 1'b0 ;
  assign n21535 = n7979 & ~n21534 ;
  assign n21536 = ( ~n4979 & n13491 ) | ( ~n4979 & n21535 ) | ( n13491 & n21535 ) ;
  assign n21537 = n21536 ^ n9079 ^ n3829 ;
  assign n21538 = n21537 ^ n1984 ^ 1'b0 ;
  assign n21539 = ~n21533 & n21538 ;
  assign n21540 = ( n2031 & ~n2667 ) | ( n2031 & n15648 ) | ( ~n2667 & n15648 ) ;
  assign n21541 = ~n6363 & n21540 ;
  assign n21542 = ( n10885 & n19816 ) | ( n10885 & ~n21541 ) | ( n19816 & ~n21541 ) ;
  assign n21543 = n14399 & ~n21542 ;
  assign n21544 = n21543 ^ n6885 ^ 1'b0 ;
  assign n21545 = ( n355 & n9565 ) | ( n355 & ~n21409 ) | ( n9565 & ~n21409 ) ;
  assign n21546 = ( n10392 & ~n13536 ) | ( n10392 & n21545 ) | ( ~n13536 & n21545 ) ;
  assign n21547 = ( ~n5682 & n6170 ) | ( ~n5682 & n16890 ) | ( n6170 & n16890 ) ;
  assign n21548 = ( n4528 & n16369 ) | ( n4528 & n21547 ) | ( n16369 & n21547 ) ;
  assign n21549 = n21548 ^ n3591 ^ n2923 ;
  assign n21550 = ( n2948 & n6029 ) | ( n2948 & ~n7806 ) | ( n6029 & ~n7806 ) ;
  assign n21551 = n10785 ^ n3306 ^ n397 ;
  assign n21552 = n21550 | n21551 ;
  assign n21553 = n7770 & ~n21552 ;
  assign n21554 = n21553 ^ n15842 ^ n9353 ;
  assign n21555 = n6792 & n12466 ;
  assign n21556 = n21554 & n21555 ;
  assign n21557 = n11343 ^ n5471 ^ n4074 ;
  assign n21558 = n21557 ^ n3610 ^ 1'b0 ;
  assign n21559 = n2314 & n21558 ;
  assign n21560 = ( n660 & n11416 ) | ( n660 & n21559 ) | ( n11416 & n21559 ) ;
  assign n21561 = ( n7444 & n9770 ) | ( n7444 & ~n21560 ) | ( n9770 & ~n21560 ) ;
  assign n21562 = ( n3432 & ~n12510 ) | ( n3432 & n17989 ) | ( ~n12510 & n17989 ) ;
  assign n21563 = n21562 ^ n13141 ^ n6895 ;
  assign n21564 = n21563 ^ n10396 ^ 1'b0 ;
  assign n21566 = n2438 | n6835 ;
  assign n21567 = n2344 | n21566 ;
  assign n21568 = n21567 ^ n8908 ^ n7646 ;
  assign n21565 = n515 | n6859 ;
  assign n21569 = n21568 ^ n21565 ^ 1'b0 ;
  assign n21570 = n20875 ^ n12336 ^ n1383 ;
  assign n21578 = ~n5941 & n11994 ;
  assign n21579 = n21578 ^ n13777 ^ 1'b0 ;
  assign n21580 = ( n2089 & n8766 ) | ( n2089 & ~n21579 ) | ( n8766 & ~n21579 ) ;
  assign n21573 = n7621 & ~n9301 ;
  assign n21574 = ~n19718 & n21573 ;
  assign n21571 = n8869 ^ n4917 ^ n332 ;
  assign n21572 = ( n4738 & n14098 ) | ( n4738 & n21571 ) | ( n14098 & n21571 ) ;
  assign n21575 = n21574 ^ n21572 ^ n8283 ;
  assign n21576 = ( n4257 & n19250 ) | ( n4257 & ~n21575 ) | ( n19250 & ~n21575 ) ;
  assign n21577 = ~n4143 & n21576 ;
  assign n21581 = n21580 ^ n21577 ^ 1'b0 ;
  assign n21582 = n12002 & n20907 ;
  assign n21583 = n21582 ^ n12706 ^ 1'b0 ;
  assign n21584 = n10564 & n21583 ;
  assign n21585 = n21584 ^ n15561 ^ 1'b0 ;
  assign n21586 = x0 & ~n21585 ;
  assign n21587 = ~n4233 & n21586 ;
  assign n21595 = ( n4794 & n7533 ) | ( n4794 & ~n8401 ) | ( n7533 & ~n8401 ) ;
  assign n21592 = n15855 ^ n6822 ^ n3925 ;
  assign n21588 = n6843 & n11075 ;
  assign n21589 = ( n416 & n3498 ) | ( n416 & n9901 ) | ( n3498 & n9901 ) ;
  assign n21590 = n3825 & n4384 ;
  assign n21591 = ( n21588 & ~n21589 ) | ( n21588 & n21590 ) | ( ~n21589 & n21590 ) ;
  assign n21593 = n21592 ^ n21591 ^ 1'b0 ;
  assign n21594 = n6481 | n21593 ;
  assign n21596 = n21595 ^ n21594 ^ n15430 ;
  assign n21597 = ( n2374 & n8408 ) | ( n2374 & n14920 ) | ( n8408 & n14920 ) ;
  assign n21598 = n16004 ^ n6795 ^ n5428 ;
  assign n21599 = n21598 ^ n14868 ^ n2429 ;
  assign n21600 = n21599 ^ n13764 ^ n9965 ;
  assign n21601 = n21600 ^ n5093 ^ n2136 ;
  assign n21602 = n13632 ^ n10583 ^ x131 ;
  assign n21603 = ( n12996 & n16835 ) | ( n12996 & ~n21602 ) | ( n16835 & ~n21602 ) ;
  assign n21604 = n21603 ^ n14998 ^ 1'b0 ;
  assign n21605 = n3284 | n21604 ;
  assign n21606 = ( n6579 & n10540 ) | ( n6579 & ~n16535 ) | ( n10540 & ~n16535 ) ;
  assign n21607 = ~n15952 & n21606 ;
  assign n21608 = n21607 ^ n21465 ^ n15269 ;
  assign n21609 = ( n8608 & n12029 ) | ( n8608 & n21608 ) | ( n12029 & n21608 ) ;
  assign n21610 = n7051 & ~n8593 ;
  assign n21611 = ( n482 & ~n15596 ) | ( n482 & n21610 ) | ( ~n15596 & n21610 ) ;
  assign n21612 = ( ~n16140 & n17388 ) | ( ~n16140 & n21611 ) | ( n17388 & n21611 ) ;
  assign n21613 = n8474 ^ n2389 ^ n436 ;
  assign n21614 = ( n15965 & ~n18604 ) | ( n15965 & n21613 ) | ( ~n18604 & n21613 ) ;
  assign n21615 = n21614 ^ n15189 ^ n8727 ;
  assign n21616 = ( n1491 & n7262 ) | ( n1491 & ~n8531 ) | ( n7262 & ~n8531 ) ;
  assign n21617 = ( n904 & n3896 ) | ( n904 & n15057 ) | ( n3896 & n15057 ) ;
  assign n21618 = n16466 ^ n12091 ^ n7090 ;
  assign n21619 = n21618 ^ n20429 ^ n460 ;
  assign n21621 = n9091 ^ n8434 ^ 1'b0 ;
  assign n21622 = ~n13244 & n21621 ;
  assign n21620 = n5125 & ~n10836 ;
  assign n21623 = n21622 ^ n21620 ^ 1'b0 ;
  assign n21624 = n21623 ^ n13649 ^ n430 ;
  assign n21625 = ( n2755 & n21619 ) | ( n2755 & ~n21624 ) | ( n21619 & ~n21624 ) ;
  assign n21626 = n16027 ^ n11497 ^ n7739 ;
  assign n21627 = ( n21617 & n21625 ) | ( n21617 & n21626 ) | ( n21625 & n21626 ) ;
  assign n21628 = n6805 ^ n3393 ^ n907 ;
  assign n21629 = ( n429 & n7176 ) | ( n429 & ~n21628 ) | ( n7176 & ~n21628 ) ;
  assign n21640 = n9606 ^ n9171 ^ n7838 ;
  assign n21641 = n21640 ^ n8641 ^ 1'b0 ;
  assign n21639 = n2323 & n20980 ;
  assign n21642 = n21641 ^ n21639 ^ 1'b0 ;
  assign n21643 = ( n7239 & ~n9459 ) | ( n7239 & n21642 ) | ( ~n9459 & n21642 ) ;
  assign n21630 = n2762 ^ n1971 ^ 1'b0 ;
  assign n21631 = ( n1415 & ~n7345 ) | ( n1415 & n21630 ) | ( ~n7345 & n21630 ) ;
  assign n21634 = n8210 ^ n3627 ^ 1'b0 ;
  assign n21635 = n17818 & n21634 ;
  assign n21636 = n21635 ^ n393 ^ 1'b0 ;
  assign n21632 = ( n559 & ~n10190 ) | ( n559 & n12585 ) | ( ~n10190 & n12585 ) ;
  assign n21633 = n21632 ^ n13386 ^ n3080 ;
  assign n21637 = n21636 ^ n21633 ^ n1665 ;
  assign n21638 = n21631 | n21637 ;
  assign n21644 = n21643 ^ n21638 ^ 1'b0 ;
  assign n21647 = ( ~n419 & n13636 ) | ( ~n419 & n17158 ) | ( n13636 & n17158 ) ;
  assign n21648 = n21647 ^ n1904 ^ n1372 ;
  assign n21645 = n21130 ^ n12659 ^ n3711 ;
  assign n21646 = n21645 ^ n19798 ^ n10256 ;
  assign n21649 = n21648 ^ n21646 ^ n15464 ;
  assign n21650 = ( ~n4086 & n8548 ) | ( ~n4086 & n17135 ) | ( n8548 & n17135 ) ;
  assign n21651 = n2027 & n16208 ;
  assign n21652 = n21651 ^ n14948 ^ n14407 ;
  assign n21653 = n21652 ^ n9763 ^ n4670 ;
  assign n21654 = ( n5178 & ~n21650 ) | ( n5178 & n21653 ) | ( ~n21650 & n21653 ) ;
  assign n21655 = n12152 ^ n7588 ^ n5919 ;
  assign n21656 = n21655 ^ n15329 ^ n7719 ;
  assign n21657 = n2649 ^ n888 ^ 1'b0 ;
  assign n21658 = ~n21656 & n21657 ;
  assign n21669 = n21061 ^ n18257 ^ n7775 ;
  assign n21668 = ( n4520 & ~n17165 ) | ( n4520 & n20589 ) | ( ~n17165 & n20589 ) ;
  assign n21670 = n21669 ^ n21668 ^ 1'b0 ;
  assign n21659 = n6418 ^ n4545 ^ n2169 ;
  assign n21664 = n11094 & ~n14043 ;
  assign n21665 = ~n14512 & n21664 ;
  assign n21662 = n20969 ^ n9249 ^ n4396 ;
  assign n21660 = n6410 & n7789 ;
  assign n21661 = ( n6843 & n13177 ) | ( n6843 & ~n21660 ) | ( n13177 & ~n21660 ) ;
  assign n21663 = n21662 ^ n21661 ^ n19806 ;
  assign n21666 = n21665 ^ n21663 ^ n959 ;
  assign n21667 = n21659 | n21666 ;
  assign n21671 = n21670 ^ n21667 ^ 1'b0 ;
  assign n21672 = ( n298 & n9659 ) | ( n298 & ~n12578 ) | ( n9659 & ~n12578 ) ;
  assign n21673 = n21672 ^ n18432 ^ n16771 ;
  assign n21674 = n11078 ^ n10493 ^ 1'b0 ;
  assign n21675 = n21674 ^ n6859 ^ x35 ;
  assign n21676 = n21675 ^ x55 ^ 1'b0 ;
  assign n21677 = ( n15315 & n21673 ) | ( n15315 & n21676 ) | ( n21673 & n21676 ) ;
  assign n21682 = n21265 ^ n11269 ^ n5300 ;
  assign n21678 = n18949 ^ n10232 ^ 1'b0 ;
  assign n21679 = n13961 & ~n21678 ;
  assign n21680 = ( n1833 & n14320 ) | ( n1833 & ~n21679 ) | ( n14320 & ~n21679 ) ;
  assign n21681 = ( n15429 & ~n16640 ) | ( n15429 & n21680 ) | ( ~n16640 & n21680 ) ;
  assign n21683 = n21682 ^ n21681 ^ n20669 ;
  assign n21686 = n1376 & n5511 ;
  assign n21687 = n21686 ^ n624 ^ 1'b0 ;
  assign n21688 = n21687 ^ n2059 ^ n1507 ;
  assign n21689 = ( n3350 & n21535 ) | ( n3350 & n21688 ) | ( n21535 & n21688 ) ;
  assign n21690 = n21689 ^ n13578 ^ n7472 ;
  assign n21691 = ( ~n574 & n12680 ) | ( ~n574 & n21690 ) | ( n12680 & n21690 ) ;
  assign n21685 = ( ~n985 & n11182 ) | ( ~n985 & n12244 ) | ( n11182 & n12244 ) ;
  assign n21684 = n17237 ^ n8698 ^ n7673 ;
  assign n21692 = n21691 ^ n21685 ^ n21684 ;
  assign n21693 = n21692 ^ n13982 ^ n5445 ;
  assign n21694 = n19621 ^ n8351 ^ n4913 ;
  assign n21706 = n3504 ^ n315 ^ 1'b0 ;
  assign n21707 = n10993 & ~n21706 ;
  assign n21695 = ( ~n2174 & n6896 ) | ( ~n2174 & n16895 ) | ( n6896 & n16895 ) ;
  assign n21698 = n7283 ^ n2275 ^ n1683 ;
  assign n21697 = n7100 ^ n5101 ^ n4218 ;
  assign n21696 = ( n1176 & ~n4755 ) | ( n1176 & n8294 ) | ( ~n4755 & n8294 ) ;
  assign n21699 = n21698 ^ n21697 ^ n21696 ;
  assign n21702 = n10118 ^ n7164 ^ 1'b0 ;
  assign n21700 = ( n10256 & n14486 ) | ( n10256 & ~n14997 ) | ( n14486 & ~n14997 ) ;
  assign n21701 = n5556 & ~n21700 ;
  assign n21703 = n21702 ^ n21701 ^ 1'b0 ;
  assign n21704 = ~n21699 & n21703 ;
  assign n21705 = ~n21695 & n21704 ;
  assign n21708 = n21707 ^ n21705 ^ n7155 ;
  assign n21712 = x105 & n2766 ;
  assign n21709 = n15879 ^ n11701 ^ n1211 ;
  assign n21710 = n21709 ^ n17418 ^ 1'b0 ;
  assign n21711 = n7658 & ~n21710 ;
  assign n21713 = n21712 ^ n21711 ^ n13162 ;
  assign n21714 = n16562 ^ n16167 ^ 1'b0 ;
  assign n21715 = n21714 ^ n8890 ^ n967 ;
  assign n21716 = n21715 ^ n12848 ^ n1895 ;
  assign n21717 = ( n8143 & n8787 ) | ( n8143 & ~n18414 ) | ( n8787 & ~n18414 ) ;
  assign n21718 = n19664 ^ n8393 ^ n6931 ;
  assign n21719 = ( n11200 & n21717 ) | ( n11200 & ~n21718 ) | ( n21717 & ~n21718 ) ;
  assign n21721 = n4322 ^ n4185 ^ 1'b0 ;
  assign n21722 = n3453 & n21721 ;
  assign n21720 = n5512 ^ n4835 ^ n2310 ;
  assign n21723 = n21722 ^ n21720 ^ n9106 ;
  assign n21724 = ( n5851 & ~n8686 ) | ( n5851 & n14602 ) | ( ~n8686 & n14602 ) ;
  assign n21725 = ( n8561 & n9671 ) | ( n8561 & n21724 ) | ( n9671 & n21724 ) ;
  assign n21726 = n8405 & n21725 ;
  assign n21727 = ~n14609 & n21726 ;
  assign n21735 = n10354 ^ x166 ^ 1'b0 ;
  assign n21736 = ( n604 & n10467 ) | ( n604 & ~n21735 ) | ( n10467 & ~n21735 ) ;
  assign n21728 = ( ~n1030 & n4195 ) | ( ~n1030 & n14191 ) | ( n4195 & n14191 ) ;
  assign n21729 = ~n8033 & n21728 ;
  assign n21730 = n21729 ^ n10788 ^ 1'b0 ;
  assign n21731 = n5672 ^ n4395 ^ n2664 ;
  assign n21732 = ( n3971 & ~n7641 ) | ( n3971 & n14401 ) | ( ~n7641 & n14401 ) ;
  assign n21733 = ( n3019 & n21731 ) | ( n3019 & n21732 ) | ( n21731 & n21732 ) ;
  assign n21734 = ( n18363 & n21730 ) | ( n18363 & ~n21733 ) | ( n21730 & ~n21733 ) ;
  assign n21737 = n21736 ^ n21734 ^ 1'b0 ;
  assign n21738 = n21488 ^ n16372 ^ n6546 ;
  assign n21739 = ( n5082 & ~n5247 ) | ( n5082 & n16152 ) | ( ~n5247 & n16152 ) ;
  assign n21740 = ( n4362 & n4407 ) | ( n4362 & n9315 ) | ( n4407 & n9315 ) ;
  assign n21741 = n21740 ^ n12178 ^ 1'b0 ;
  assign n21742 = n21379 | n21741 ;
  assign n21744 = ~n339 & n16863 ;
  assign n21743 = ( n4581 & n12837 ) | ( n4581 & n18589 ) | ( n12837 & n18589 ) ;
  assign n21745 = n21744 ^ n21743 ^ n1405 ;
  assign n21748 = n7653 ^ n5106 ^ n1677 ;
  assign n21749 = n14106 ^ n6243 ^ n325 ;
  assign n21750 = ( n18900 & n21748 ) | ( n18900 & ~n21749 ) | ( n21748 & ~n21749 ) ;
  assign n21746 = n8446 ^ n4653 ^ n3272 ;
  assign n21747 = n21746 ^ n14365 ^ n1674 ;
  assign n21751 = n21750 ^ n21747 ^ n10103 ;
  assign n21754 = n2515 | n5490 ;
  assign n21752 = n10403 ^ n10127 ^ 1'b0 ;
  assign n21753 = ( n10462 & n14440 ) | ( n10462 & n21752 ) | ( n14440 & n21752 ) ;
  assign n21755 = n21754 ^ n21753 ^ n15818 ;
  assign n21756 = ( ~n5725 & n9596 ) | ( ~n5725 & n21755 ) | ( n9596 & n21755 ) ;
  assign n21757 = n1652 & n2190 ;
  assign n21758 = n21757 ^ n1881 ^ 1'b0 ;
  assign n21759 = n21758 ^ n3270 ^ n1488 ;
  assign n21760 = n14032 ^ n7044 ^ n1297 ;
  assign n21761 = ( n11689 & n21759 ) | ( n11689 & ~n21760 ) | ( n21759 & ~n21760 ) ;
  assign n21762 = n4481 & ~n11332 ;
  assign n21763 = n21762 ^ n8935 ^ n5017 ;
  assign n21765 = ( n2153 & ~n13509 ) | ( n2153 & n15811 ) | ( ~n13509 & n15811 ) ;
  assign n21764 = n16007 ^ n3886 ^ 1'b0 ;
  assign n21766 = n21765 ^ n21764 ^ n19572 ;
  assign n21767 = ~n13117 & n19929 ;
  assign n21768 = n2289 ^ n2167 ^ 1'b0 ;
  assign n21769 = ~n783 & n21768 ;
  assign n21770 = n14437 ^ n13418 ^ n6473 ;
  assign n21771 = n5498 & ~n17107 ;
  assign n21772 = ( n21769 & n21770 ) | ( n21769 & ~n21771 ) | ( n21770 & ~n21771 ) ;
  assign n21773 = n15735 | n21772 ;
  assign n21776 = n599 & ~n1956 ;
  assign n21777 = n10652 & n21776 ;
  assign n21778 = n8082 & ~n21777 ;
  assign n21774 = n12220 ^ n8539 ^ 1'b0 ;
  assign n21775 = ~n12841 & n21774 ;
  assign n21779 = n21778 ^ n21775 ^ n1795 ;
  assign n21780 = ( n611 & n5303 ) | ( n611 & ~n12491 ) | ( n5303 & ~n12491 ) ;
  assign n21781 = n4724 ^ n3399 ^ 1'b0 ;
  assign n21782 = n21780 & n21781 ;
  assign n21783 = n21782 ^ n17952 ^ n5731 ;
  assign n21784 = ( ~n780 & n7506 ) | ( ~n780 & n12849 ) | ( n7506 & n12849 ) ;
  assign n21785 = n21784 ^ n12399 ^ n6971 ;
  assign n21786 = n21785 ^ n20961 ^ n9414 ;
  assign n21787 = ( n6010 & ~n21783 ) | ( n6010 & n21786 ) | ( ~n21783 & n21786 ) ;
  assign n21788 = n3813 & n9375 ;
  assign n21789 = ~n8040 & n21788 ;
  assign n21793 = n16659 ^ n14229 ^ n7071 ;
  assign n21794 = n21793 ^ n12342 ^ n8621 ;
  assign n21795 = n16954 ^ n5564 ^ n3022 ;
  assign n21796 = ( n16709 & n21794 ) | ( n16709 & ~n21795 ) | ( n21794 & ~n21795 ) ;
  assign n21790 = n6158 ^ n5414 ^ x1 ;
  assign n21791 = n21790 ^ n6680 ^ n3497 ;
  assign n21792 = n21791 ^ n13890 ^ n11878 ;
  assign n21797 = n21796 ^ n21792 ^ n5348 ;
  assign n21798 = n21789 | n21797 ;
  assign n21799 = n3347 & ~n4625 ;
  assign n21800 = n21799 ^ n3761 ^ 1'b0 ;
  assign n21801 = n11262 ^ n2609 ^ x41 ;
  assign n21802 = n21801 ^ n3484 ^ n409 ;
  assign n21803 = n10659 & ~n21802 ;
  assign n21804 = n21803 ^ n21327 ^ 1'b0 ;
  assign n21805 = ( n8874 & ~n10076 ) | ( n8874 & n21454 ) | ( ~n10076 & n21454 ) ;
  assign n21806 = n21805 ^ n11770 ^ n2234 ;
  assign n21807 = ( ~n6471 & n21804 ) | ( ~n6471 & n21806 ) | ( n21804 & n21806 ) ;
  assign n21808 = ( n2517 & n3247 ) | ( n2517 & n4180 ) | ( n3247 & n4180 ) ;
  assign n21809 = ( ~n1944 & n7073 ) | ( ~n1944 & n9311 ) | ( n7073 & n9311 ) ;
  assign n21810 = ( n18983 & n21808 ) | ( n18983 & n21809 ) | ( n21808 & n21809 ) ;
  assign n21811 = n8185 ^ n5006 ^ n2643 ;
  assign n21812 = n10988 ^ n8015 ^ 1'b0 ;
  assign n21813 = ~n21811 & n21812 ;
  assign n21817 = ( n2602 & n5984 ) | ( n2602 & n6740 ) | ( n5984 & n6740 ) ;
  assign n21815 = ( n5878 & ~n6353 ) | ( n5878 & n15387 ) | ( ~n6353 & n15387 ) ;
  assign n21816 = n21815 ^ n13335 ^ n7714 ;
  assign n21818 = n21817 ^ n21816 ^ n18915 ;
  assign n21814 = ( n2004 & n3191 ) | ( n2004 & ~n12857 ) | ( n3191 & ~n12857 ) ;
  assign n21819 = n21818 ^ n21814 ^ n12247 ;
  assign n21824 = n11413 ^ n8090 ^ n6014 ;
  assign n21823 = n16909 ^ n10495 ^ n3188 ;
  assign n21820 = ( n522 & n7501 ) | ( n522 & n16091 ) | ( n7501 & n16091 ) ;
  assign n21821 = n4933 | n21820 ;
  assign n21822 = ( ~n10650 & n17998 ) | ( ~n10650 & n21821 ) | ( n17998 & n21821 ) ;
  assign n21825 = n21824 ^ n21823 ^ n21822 ;
  assign n21826 = n8167 & ~n16626 ;
  assign n21827 = n21826 ^ n12091 ^ x197 ;
  assign n21828 = n21827 ^ n19572 ^ 1'b0 ;
  assign n21829 = n7524 ^ n5148 ^ 1'b0 ;
  assign n21830 = n21829 ^ n19905 ^ n16626 ;
  assign n21831 = ( n819 & ~n6985 ) | ( n819 & n13743 ) | ( ~n6985 & n13743 ) ;
  assign n21832 = n19874 ^ n5298 ^ n2333 ;
  assign n21834 = ( n1861 & ~n2968 ) | ( n1861 & n7396 ) | ( ~n2968 & n7396 ) ;
  assign n21833 = ( ~n1761 & n4231 ) | ( ~n1761 & n8106 ) | ( n4231 & n8106 ) ;
  assign n21835 = n21834 ^ n21833 ^ n16907 ;
  assign n21836 = ( n1250 & ~n6339 ) | ( n1250 & n17713 ) | ( ~n6339 & n17713 ) ;
  assign n21837 = n9877 ^ n3963 ^ n888 ;
  assign n21838 = ( n7312 & n17188 ) | ( n7312 & n21837 ) | ( n17188 & n21837 ) ;
  assign n21839 = n8331 ^ n3790 ^ n1374 ;
  assign n21840 = n21839 ^ n13308 ^ n5819 ;
  assign n21841 = ( n4150 & ~n8387 ) | ( n4150 & n18919 ) | ( ~n8387 & n18919 ) ;
  assign n21842 = ( n10290 & n11358 ) | ( n10290 & n11987 ) | ( n11358 & n11987 ) ;
  assign n21843 = ( n1123 & ~n9673 ) | ( n1123 & n21842 ) | ( ~n9673 & n21842 ) ;
  assign n21845 = ( ~n10734 & n11736 ) | ( ~n10734 & n12889 ) | ( n11736 & n12889 ) ;
  assign n21844 = n6101 ^ n2932 ^ n1518 ;
  assign n21846 = n21845 ^ n21844 ^ n3927 ;
  assign n21847 = n11331 & n21846 ;
  assign n21848 = ~n8637 & n21847 ;
  assign n21849 = n13684 ^ n8854 ^ n5235 ;
  assign n21850 = n16140 ^ n9083 ^ n4674 ;
  assign n21852 = n9600 ^ n6081 ^ n2923 ;
  assign n21851 = n5369 | n6281 ;
  assign n21853 = n21852 ^ n21851 ^ 1'b0 ;
  assign n21854 = ( n18702 & n19179 ) | ( n18702 & ~n21853 ) | ( n19179 & ~n21853 ) ;
  assign n21855 = ( n11511 & n21850 ) | ( n11511 & n21854 ) | ( n21850 & n21854 ) ;
  assign n21856 = ( n359 & n5174 ) | ( n359 & n6042 ) | ( n5174 & n6042 ) ;
  assign n21857 = n21856 ^ n11202 ^ n8827 ;
  assign n21858 = n21857 ^ n16617 ^ n2822 ;
  assign n21860 = ( ~n3534 & n4776 ) | ( ~n3534 & n9895 ) | ( n4776 & n9895 ) ;
  assign n21861 = n9508 | n21860 ;
  assign n21862 = n3248 | n21861 ;
  assign n21863 = n21862 ^ n6875 ^ n5751 ;
  assign n21864 = ( n9917 & ~n15045 ) | ( n9917 & n21863 ) | ( ~n15045 & n21863 ) ;
  assign n21859 = ( ~n5884 & n15669 ) | ( ~n5884 & n18953 ) | ( n15669 & n18953 ) ;
  assign n21865 = n21864 ^ n21859 ^ n13998 ;
  assign n21866 = ( n4244 & n9251 ) | ( n4244 & n14974 ) | ( n9251 & n14974 ) ;
  assign n21867 = x65 & ~n4723 ;
  assign n21868 = ~n14064 & n21867 ;
  assign n21869 = n18527 ^ n11951 ^ 1'b0 ;
  assign n21874 = ~n6981 & n10267 ;
  assign n21875 = n21874 ^ n20737 ^ 1'b0 ;
  assign n21871 = n9856 ^ n7673 ^ n5277 ;
  assign n21870 = n10493 ^ n7619 ^ n5468 ;
  assign n21872 = n21871 ^ n21870 ^ n1528 ;
  assign n21873 = n11792 & ~n21872 ;
  assign n21876 = n21875 ^ n21873 ^ n19649 ;
  assign n21878 = ( n2250 & ~n3576 ) | ( n2250 & n11470 ) | ( ~n3576 & n11470 ) ;
  assign n21877 = n6720 & n11596 ;
  assign n21879 = n21878 ^ n21877 ^ 1'b0 ;
  assign n21880 = ( n1129 & ~n10420 ) | ( n1129 & n16643 ) | ( ~n10420 & n16643 ) ;
  assign n21881 = n15800 ^ n6799 ^ n4304 ;
  assign n21882 = ( n6926 & ~n21880 ) | ( n6926 & n21881 ) | ( ~n21880 & n21881 ) ;
  assign n21883 = n8312 ^ n5628 ^ 1'b0 ;
  assign n21884 = n20069 & n21883 ;
  assign n21885 = n12082 | n15326 ;
  assign n21886 = n2397 | n21885 ;
  assign n21887 = ~n3247 & n14100 ;
  assign n21888 = ( n1621 & ~n2922 ) | ( n1621 & n8618 ) | ( ~n2922 & n8618 ) ;
  assign n21889 = ( ~n21886 & n21887 ) | ( ~n21886 & n21888 ) | ( n21887 & n21888 ) ;
  assign n21890 = n21245 ^ n7080 ^ 1'b0 ;
  assign n21891 = n21890 ^ n15674 ^ 1'b0 ;
  assign n21893 = n11617 ^ n1084 ^ 1'b0 ;
  assign n21894 = ( ~x244 & n9200 ) | ( ~x244 & n21893 ) | ( n9200 & n21893 ) ;
  assign n21892 = n17986 ^ n10783 ^ n7904 ;
  assign n21895 = n21894 ^ n21892 ^ n2003 ;
  assign n21896 = ~n671 & n1822 ;
  assign n21897 = n16846 ^ n9650 ^ n4443 ;
  assign n21898 = ~n969 & n17565 ;
  assign n21899 = n21897 | n21898 ;
  assign n21900 = ( n7802 & n21896 ) | ( n7802 & n21899 ) | ( n21896 & n21899 ) ;
  assign n21901 = ( n4685 & n7509 ) | ( n4685 & n18983 ) | ( n7509 & n18983 ) ;
  assign n21902 = ( n10159 & ~n19722 ) | ( n10159 & n21901 ) | ( ~n19722 & n21901 ) ;
  assign n21903 = n21902 ^ n9690 ^ n3079 ;
  assign n21904 = ( x130 & n4140 ) | ( x130 & n12880 ) | ( n4140 & n12880 ) ;
  assign n21905 = n2591 | n2907 ;
  assign n21906 = n21905 ^ n454 ^ 1'b0 ;
  assign n21907 = n3210 ^ n2424 ^ 1'b0 ;
  assign n21908 = n2775 & n21907 ;
  assign n21909 = ~n12818 & n21908 ;
  assign n21910 = n14167 & n21909 ;
  assign n21911 = ( n20070 & n21906 ) | ( n20070 & ~n21910 ) | ( n21906 & ~n21910 ) ;
  assign n21912 = ( ~n669 & n6308 ) | ( ~n669 & n20582 ) | ( n6308 & n20582 ) ;
  assign n21913 = n10494 ^ n4216 ^ 1'b0 ;
  assign n21914 = ( ~n2571 & n21912 ) | ( ~n2571 & n21913 ) | ( n21912 & n21913 ) ;
  assign n21915 = ( n11454 & n18255 ) | ( n11454 & n20013 ) | ( n18255 & n20013 ) ;
  assign n21923 = n1496 & n3461 ;
  assign n21921 = n5470 ^ x216 ^ x107 ;
  assign n21922 = n21921 ^ n2348 ^ n1784 ;
  assign n21916 = n6669 ^ n1855 ^ 1'b0 ;
  assign n21917 = n21916 ^ n8138 ^ n5330 ;
  assign n21918 = n12832 | n15539 ;
  assign n21919 = n21917 | n21918 ;
  assign n21920 = ( n14927 & n20893 ) | ( n14927 & ~n21919 ) | ( n20893 & ~n21919 ) ;
  assign n21924 = n21923 ^ n21922 ^ n21920 ;
  assign n21925 = ( ~n418 & n13371 ) | ( ~n418 & n17833 ) | ( n13371 & n17833 ) ;
  assign n21926 = n21925 ^ n19820 ^ n16448 ;
  assign n21927 = ( ~n4095 & n5693 ) | ( ~n4095 & n18530 ) | ( n5693 & n18530 ) ;
  assign n21928 = n8396 & ~n21927 ;
  assign n21929 = ~n17288 & n21928 ;
  assign n21930 = n21929 ^ n20247 ^ n15840 ;
  assign n21931 = n777 | n9756 ;
  assign n21932 = n11491 & ~n21931 ;
  assign n21933 = n9234 ^ n8783 ^ n782 ;
  assign n21934 = n21933 ^ n11704 ^ n3272 ;
  assign n21935 = ( n2780 & n21932 ) | ( n2780 & n21934 ) | ( n21932 & n21934 ) ;
  assign n21936 = n2780 & ~n4551 ;
  assign n21937 = n21936 ^ n14084 ^ n4583 ;
  assign n21938 = n6039 & ~n7202 ;
  assign n21939 = n8398 | n21938 ;
  assign n21940 = ( ~n3869 & n21937 ) | ( ~n3869 & n21939 ) | ( n21937 & n21939 ) ;
  assign n21941 = n701 | n16090 ;
  assign n21942 = n21941 ^ n3403 ^ 1'b0 ;
  assign n21943 = n21942 ^ n17821 ^ n9854 ;
  assign n21944 = n20526 & n21943 ;
  assign n21945 = n21944 ^ n17959 ^ 1'b0 ;
  assign n21946 = n6211 ^ n4308 ^ 1'b0 ;
  assign n21947 = ( n4787 & n13267 ) | ( n4787 & n21946 ) | ( n13267 & n21946 ) ;
  assign n21948 = n12136 ^ n11694 ^ n6147 ;
  assign n21953 = n15705 ^ n7071 ^ x112 ;
  assign n21952 = n5148 ^ n2041 ^ x232 ;
  assign n21954 = n21953 ^ n21952 ^ n19708 ;
  assign n21949 = n9784 ^ n1955 ^ n779 ;
  assign n21950 = n21949 ^ x54 ^ 1'b0 ;
  assign n21951 = ( ~n2611 & n2813 ) | ( ~n2611 & n21950 ) | ( n2813 & n21950 ) ;
  assign n21955 = n21954 ^ n21951 ^ n8041 ;
  assign n21956 = n14430 ^ n10304 ^ n5459 ;
  assign n21957 = ( n739 & n4500 ) | ( n739 & n12288 ) | ( n4500 & n12288 ) ;
  assign n21958 = ( n4181 & n8035 ) | ( n4181 & n10025 ) | ( n8035 & n10025 ) ;
  assign n21959 = n5573 ^ n1812 ^ n281 ;
  assign n21960 = n21959 ^ n19062 ^ 1'b0 ;
  assign n21961 = n3800 & n21960 ;
  assign n21962 = ( n21957 & n21958 ) | ( n21957 & ~n21961 ) | ( n21958 & ~n21961 ) ;
  assign n21963 = n2076 & ~n3042 ;
  assign n21964 = ~n2341 & n16018 ;
  assign n21965 = ( n10331 & n21963 ) | ( n10331 & ~n21964 ) | ( n21963 & ~n21964 ) ;
  assign n21966 = n3764 ^ n3415 ^ 1'b0 ;
  assign n21967 = n10820 ^ n9755 ^ 1'b0 ;
  assign n21968 = n21966 | n21967 ;
  assign n21969 = ~n21965 & n21968 ;
  assign n21970 = n11091 ^ n10110 ^ n7933 ;
  assign n21971 = n21970 ^ n5934 ^ 1'b0 ;
  assign n21972 = n14933 ^ n7592 ^ n4476 ;
  assign n21973 = ( n3240 & n11029 ) | ( n3240 & n21972 ) | ( n11029 & n21972 ) ;
  assign n21974 = ( x81 & n967 ) | ( x81 & ~n6062 ) | ( n967 & ~n6062 ) ;
  assign n21975 = ( ~n14898 & n21973 ) | ( ~n14898 & n21974 ) | ( n21973 & n21974 ) ;
  assign n21976 = n18537 ^ n14195 ^ n2585 ;
  assign n21977 = ( n4604 & ~n9003 ) | ( n4604 & n10506 ) | ( ~n9003 & n10506 ) ;
  assign n21978 = n13240 ^ n8761 ^ n5439 ;
  assign n21979 = n16133 ^ n8208 ^ n5609 ;
  assign n21980 = n9970 & ~n21979 ;
  assign n21981 = n21980 ^ n7146 ^ 1'b0 ;
  assign n21982 = ( n13294 & n21978 ) | ( n13294 & ~n21981 ) | ( n21978 & ~n21981 ) ;
  assign n21986 = ( ~n4824 & n5334 ) | ( ~n4824 & n12295 ) | ( n5334 & n12295 ) ;
  assign n21983 = ~n12201 & n12551 ;
  assign n21984 = ( n13402 & ~n19538 ) | ( n13402 & n21983 ) | ( ~n19538 & n21983 ) ;
  assign n21985 = n21984 ^ n17634 ^ 1'b0 ;
  assign n21987 = n21986 ^ n21985 ^ n14006 ;
  assign n21988 = n5502 ^ n3628 ^ n3376 ;
  assign n21989 = ~n12963 & n20375 ;
  assign n21990 = n9545 ^ n1949 ^ 1'b0 ;
  assign n21991 = n3058 | n21990 ;
  assign n21993 = ( ~n4655 & n9475 ) | ( ~n4655 & n13354 ) | ( n9475 & n13354 ) ;
  assign n21994 = ( n9222 & n10492 ) | ( n9222 & ~n21993 ) | ( n10492 & ~n21993 ) ;
  assign n21992 = n7731 & n8712 ;
  assign n21995 = n21994 ^ n21992 ^ n14658 ;
  assign n21996 = n10620 ^ n9487 ^ n8618 ;
  assign n21997 = n2125 ^ n1549 ^ n511 ;
  assign n21998 = ( ~n9599 & n21996 ) | ( ~n9599 & n21997 ) | ( n21996 & n21997 ) ;
  assign n21999 = ( n6608 & ~n8903 ) | ( n6608 & n16053 ) | ( ~n8903 & n16053 ) ;
  assign n22002 = n12330 ^ n7722 ^ n7714 ;
  assign n22000 = n15615 ^ n10361 ^ x247 ;
  assign n22001 = ( n9902 & n14556 ) | ( n9902 & ~n22000 ) | ( n14556 & ~n22000 ) ;
  assign n22003 = n22002 ^ n22001 ^ n7238 ;
  assign n22004 = ( n2078 & n13112 ) | ( n2078 & n17271 ) | ( n13112 & n17271 ) ;
  assign n22011 = n21953 ^ n19159 ^ n3242 ;
  assign n22012 = n14420 ^ n8052 ^ n3422 ;
  assign n22013 = n16455 ^ n6724 ^ n2021 ;
  assign n22014 = ( ~n22011 & n22012 ) | ( ~n22011 & n22013 ) | ( n22012 & n22013 ) ;
  assign n22005 = n5718 ^ n2781 ^ n2249 ;
  assign n22006 = n9328 & ~n22005 ;
  assign n22007 = ~n11090 & n22006 ;
  assign n22008 = n22007 ^ n16827 ^ n1151 ;
  assign n22009 = n16164 | n22008 ;
  assign n22010 = n22009 ^ n9166 ^ 1'b0 ;
  assign n22015 = n22014 ^ n22010 ^ 1'b0 ;
  assign n22016 = n22004 & n22015 ;
  assign n22017 = n13219 ^ n9198 ^ 1'b0 ;
  assign n22019 = ( n854 & ~n6648 ) | ( n854 & n13141 ) | ( ~n6648 & n13141 ) ;
  assign n22018 = ( n3830 & n5924 ) | ( n3830 & n9677 ) | ( n5924 & n9677 ) ;
  assign n22020 = n22019 ^ n22018 ^ n14069 ;
  assign n22021 = ( n15682 & n22017 ) | ( n15682 & n22020 ) | ( n22017 & n22020 ) ;
  assign n22023 = n8233 ^ n953 ^ 1'b0 ;
  assign n22024 = n836 & ~n22023 ;
  assign n22022 = n14183 ^ n5421 ^ 1'b0 ;
  assign n22025 = n22024 ^ n22022 ^ n4282 ;
  assign n22028 = ( n1291 & ~n1556 ) | ( n1291 & n1665 ) | ( ~n1556 & n1665 ) ;
  assign n22026 = x249 & ~n4009 ;
  assign n22027 = n14602 & n22026 ;
  assign n22029 = n22028 ^ n22027 ^ n2471 ;
  assign n22030 = n8439 & n18301 ;
  assign n22031 = n22029 & n22030 ;
  assign n22032 = n22031 ^ n18978 ^ 1'b0 ;
  assign n22033 = n1309 ^ x56 ^ 1'b0 ;
  assign n22034 = n4948 & ~n8370 ;
  assign n22035 = n16763 & n22034 ;
  assign n22036 = ( n20117 & ~n22033 ) | ( n20117 & n22035 ) | ( ~n22033 & n22035 ) ;
  assign n22037 = n22036 ^ n21394 ^ n12623 ;
  assign n22038 = n22037 ^ n21168 ^ n13411 ;
  assign n22039 = n17331 ^ n15557 ^ n11056 ;
  assign n22040 = ( n3298 & ~n10498 ) | ( n3298 & n22039 ) | ( ~n10498 & n22039 ) ;
  assign n22041 = ( n20117 & ~n22038 ) | ( n20117 & n22040 ) | ( ~n22038 & n22040 ) ;
  assign n22042 = n7214 ^ n4207 ^ 1'b0 ;
  assign n22043 = ( n1145 & n7067 ) | ( n1145 & ~n8044 ) | ( n7067 & ~n8044 ) ;
  assign n22044 = ( ~n7054 & n22042 ) | ( ~n7054 & n22043 ) | ( n22042 & n22043 ) ;
  assign n22048 = ( ~n1571 & n12578 ) | ( ~n1571 & n15420 ) | ( n12578 & n15420 ) ;
  assign n22045 = n14410 ^ n13768 ^ n10123 ;
  assign n22046 = ( n1142 & n2056 ) | ( n1142 & ~n22045 ) | ( n2056 & ~n22045 ) ;
  assign n22047 = n22046 ^ n5277 ^ n4065 ;
  assign n22049 = n22048 ^ n22047 ^ n16534 ;
  assign n22050 = ( n632 & n11926 ) | ( n632 & n13613 ) | ( n11926 & n13613 ) ;
  assign n22051 = ( ~n7164 & n18290 ) | ( ~n7164 & n21446 ) | ( n18290 & n21446 ) ;
  assign n22052 = ( ~n1402 & n6156 ) | ( ~n1402 & n22051 ) | ( n6156 & n22051 ) ;
  assign n22053 = n22052 ^ n9421 ^ 1'b0 ;
  assign n22054 = n3856 & ~n22053 ;
  assign n22055 = ~n5152 & n8485 ;
  assign n22056 = n22055 ^ n3310 ^ 1'b0 ;
  assign n22057 = ( n16538 & n16988 ) | ( n16538 & ~n22056 ) | ( n16988 & ~n22056 ) ;
  assign n22058 = ( n371 & n12784 ) | ( n371 & n22057 ) | ( n12784 & n22057 ) ;
  assign n22059 = ( n13717 & n14288 ) | ( n13717 & n17277 ) | ( n14288 & n17277 ) ;
  assign n22060 = n12288 & ~n22059 ;
  assign n22061 = n12595 ^ n11265 ^ n1670 ;
  assign n22062 = ( n8518 & n17166 ) | ( n8518 & n22061 ) | ( n17166 & n22061 ) ;
  assign n22066 = ( n9441 & n10207 ) | ( n9441 & n17155 ) | ( n10207 & n17155 ) ;
  assign n22063 = ~n7024 & n14174 ;
  assign n22064 = n4141 & ~n9488 ;
  assign n22065 = ~n22063 & n22064 ;
  assign n22067 = n22066 ^ n22065 ^ n17331 ;
  assign n22077 = n16466 ^ n13312 ^ n10779 ;
  assign n22071 = n1285 | n6736 ;
  assign n22072 = n4650 & ~n22071 ;
  assign n22073 = ( n3074 & n6848 ) | ( n3074 & n22072 ) | ( n6848 & n22072 ) ;
  assign n22069 = n11817 ^ n4783 ^ 1'b0 ;
  assign n22070 = ~n2103 & n22069 ;
  assign n22074 = n22073 ^ n22070 ^ n5914 ;
  assign n22068 = n3725 & n10170 ;
  assign n22075 = n22074 ^ n22068 ^ 1'b0 ;
  assign n22076 = n22075 ^ n18721 ^ n3552 ;
  assign n22078 = n22077 ^ n22076 ^ n16158 ;
  assign n22079 = ( ~n2356 & n10777 ) | ( ~n2356 & n22078 ) | ( n10777 & n22078 ) ;
  assign n22080 = ( n667 & n14293 ) | ( n667 & n17499 ) | ( n14293 & n17499 ) ;
  assign n22081 = ( ~n3036 & n10180 ) | ( ~n3036 & n22080 ) | ( n10180 & n22080 ) ;
  assign n22082 = n13700 ^ n7855 ^ n910 ;
  assign n22083 = n2006 & n22082 ;
  assign n22084 = ~n22081 & n22083 ;
  assign n22085 = n11863 ^ n794 ^ x65 ;
  assign n22086 = n2576 | n22085 ;
  assign n22087 = n12492 & ~n22086 ;
  assign n22088 = ( n16742 & n16987 ) | ( n16742 & ~n22087 ) | ( n16987 & ~n22087 ) ;
  assign n22089 = ( n614 & n22084 ) | ( n614 & ~n22088 ) | ( n22084 & ~n22088 ) ;
  assign n22091 = n10194 ^ n7898 ^ 1'b0 ;
  assign n22090 = ( n1565 & ~n1747 ) | ( n1565 & n3159 ) | ( ~n1747 & n3159 ) ;
  assign n22092 = n22091 ^ n22090 ^ n15048 ;
  assign n22093 = n22092 ^ n18882 ^ n13160 ;
  assign n22094 = ( n2374 & n9318 ) | ( n2374 & n17978 ) | ( n9318 & n17978 ) ;
  assign n22095 = n17989 ^ n1228 ^ 1'b0 ;
  assign n22096 = ( n3344 & ~n6007 ) | ( n3344 & n9370 ) | ( ~n6007 & n9370 ) ;
  assign n22097 = ( ~n4865 & n22095 ) | ( ~n4865 & n22096 ) | ( n22095 & n22096 ) ;
  assign n22098 = n22097 ^ n14887 ^ n7896 ;
  assign n22099 = n3423 & ~n22098 ;
  assign n22100 = n20133 ^ n13637 ^ n13302 ;
  assign n22101 = n9066 ^ n7488 ^ n2450 ;
  assign n22102 = n22101 ^ n20106 ^ n15870 ;
  assign n22103 = n1330 | n12996 ;
  assign n22104 = n22102 | n22103 ;
  assign n22105 = n22104 ^ n17214 ^ n9489 ;
  assign n22106 = n13123 ^ n8232 ^ n3592 ;
  assign n22107 = ~n8221 & n15168 ;
  assign n22108 = ( ~n18082 & n22106 ) | ( ~n18082 & n22107 ) | ( n22106 & n22107 ) ;
  assign n22109 = n2645 ^ n2290 ^ n1603 ;
  assign n22110 = n5365 & n22109 ;
  assign n22111 = ~n17602 & n22110 ;
  assign n22112 = n15655 ^ n8236 ^ n6139 ;
  assign n22113 = n22112 ^ n14808 ^ n933 ;
  assign n22114 = ( n10466 & ~n12492 ) | ( n10466 & n12739 ) | ( ~n12492 & n12739 ) ;
  assign n22115 = ( ~n747 & n12474 ) | ( ~n747 & n22114 ) | ( n12474 & n22114 ) ;
  assign n22116 = n6637 ^ n2012 ^ 1'b0 ;
  assign n22117 = ~n1197 & n22116 ;
  assign n22118 = n12110 ^ n2377 ^ n1084 ;
  assign n22119 = n22118 ^ n11995 ^ 1'b0 ;
  assign n22120 = n821 & ~n22119 ;
  assign n22121 = ( n4876 & n13164 ) | ( n4876 & ~n22120 ) | ( n13164 & ~n22120 ) ;
  assign n22122 = ( n1412 & n19993 ) | ( n1412 & n22121 ) | ( n19993 & n22121 ) ;
  assign n22123 = ( ~n3567 & n22117 ) | ( ~n3567 & n22122 ) | ( n22117 & n22122 ) ;
  assign n22124 = n2534 ^ n1267 ^ 1'b0 ;
  assign n22125 = n10354 ^ x25 ^ 1'b0 ;
  assign n22126 = ( n13967 & n22124 ) | ( n13967 & ~n22125 ) | ( n22124 & ~n22125 ) ;
  assign n22133 = n8912 ^ n2742 ^ x156 ;
  assign n22127 = n10902 | n13110 ;
  assign n22128 = n2335 & ~n22127 ;
  assign n22129 = n6663 ^ n678 ^ 1'b0 ;
  assign n22130 = n14144 ^ n5514 ^ 1'b0 ;
  assign n22131 = ( n22128 & n22129 ) | ( n22128 & n22130 ) | ( n22129 & n22130 ) ;
  assign n22132 = ( n2471 & n3681 ) | ( n2471 & ~n22131 ) | ( n3681 & ~n22131 ) ;
  assign n22134 = n22133 ^ n22132 ^ n17058 ;
  assign n22138 = ( n2364 & n15974 ) | ( n2364 & ~n16344 ) | ( n15974 & ~n16344 ) ;
  assign n22135 = n9377 ^ n1067 ^ n779 ;
  assign n22136 = ( n3514 & n6718 ) | ( n3514 & n22135 ) | ( n6718 & n22135 ) ;
  assign n22137 = ( n1827 & n4907 ) | ( n1827 & ~n22136 ) | ( n4907 & ~n22136 ) ;
  assign n22139 = n22138 ^ n22137 ^ 1'b0 ;
  assign n22140 = n5208 ^ n4706 ^ n507 ;
  assign n22141 = ( x40 & n22139 ) | ( x40 & ~n22140 ) | ( n22139 & ~n22140 ) ;
  assign n22142 = n14008 ^ n6279 ^ x250 ;
  assign n22143 = n22142 ^ n18588 ^ 1'b0 ;
  assign n22144 = ( n9632 & ~n16355 ) | ( n9632 & n22143 ) | ( ~n16355 & n22143 ) ;
  assign n22145 = ( n3436 & n9097 ) | ( n3436 & ~n17509 ) | ( n9097 & ~n17509 ) ;
  assign n22146 = ( n1747 & n13773 ) | ( n1747 & n22145 ) | ( n13773 & n22145 ) ;
  assign n22147 = n22146 ^ n18746 ^ n6838 ;
  assign n22148 = ( n14213 & n17418 ) | ( n14213 & ~n22147 ) | ( n17418 & ~n22147 ) ;
  assign n22149 = n22148 ^ n20494 ^ n14867 ;
  assign n22150 = n19721 | n22149 ;
  assign n22151 = ( ~n3051 & n3992 ) | ( ~n3051 & n18251 ) | ( n3992 & n18251 ) ;
  assign n22152 = n20910 ^ n19190 ^ 1'b0 ;
  assign n22153 = n4693 | n22152 ;
  assign n22155 = ( n512 & n4020 ) | ( n512 & n8268 ) | ( n4020 & n8268 ) ;
  assign n22154 = n4638 | n11632 ;
  assign n22156 = n22155 ^ n22154 ^ 1'b0 ;
  assign n22157 = n22156 ^ n8414 ^ 1'b0 ;
  assign n22158 = n22157 ^ n11131 ^ n6593 ;
  assign n22159 = ( ~n22151 & n22153 ) | ( ~n22151 & n22158 ) | ( n22153 & n22158 ) ;
  assign n22160 = ( n1281 & ~n10902 ) | ( n1281 & n16730 ) | ( ~n10902 & n16730 ) ;
  assign n22161 = ( ~n6431 & n16607 ) | ( ~n6431 & n22160 ) | ( n16607 & n22160 ) ;
  assign n22162 = n10116 ^ n9898 ^ n3690 ;
  assign n22163 = ~n10583 & n22162 ;
  assign n22164 = ( n2379 & ~n9882 ) | ( n2379 & n22163 ) | ( ~n9882 & n22163 ) ;
  assign n22165 = n22164 ^ n1781 ^ x58 ;
  assign n22166 = ( n1582 & n15988 ) | ( n1582 & n22165 ) | ( n15988 & n22165 ) ;
  assign n22167 = n22161 | n22166 ;
  assign n22168 = n22167 ^ n8433 ^ 1'b0 ;
  assign n22169 = n19181 | n22168 ;
  assign n22170 = n20737 ^ n13539 ^ n4458 ;
  assign n22171 = ~n7377 & n18641 ;
  assign n22172 = ( n6905 & n22170 ) | ( n6905 & ~n22171 ) | ( n22170 & ~n22171 ) ;
  assign n22173 = n19267 ^ n2277 ^ n435 ;
  assign n22174 = ( ~n14936 & n16855 ) | ( ~n14936 & n22173 ) | ( n16855 & n22173 ) ;
  assign n22175 = ( n1136 & n16481 ) | ( n1136 & n22174 ) | ( n16481 & n22174 ) ;
  assign n22176 = ( ~n666 & n13296 ) | ( ~n666 & n22175 ) | ( n13296 & n22175 ) ;
  assign n22177 = ( n10884 & ~n22172 ) | ( n10884 & n22176 ) | ( ~n22172 & n22176 ) ;
  assign n22180 = ~n7886 & n12298 ;
  assign n22181 = n916 & n22180 ;
  assign n22179 = ( n6960 & ~n11268 ) | ( n6960 & n13549 ) | ( ~n11268 & n13549 ) ;
  assign n22178 = n18288 ^ n17987 ^ n16166 ;
  assign n22182 = n22181 ^ n22179 ^ n22178 ;
  assign n22183 = ( n4771 & ~n13957 ) | ( n4771 & n16179 ) | ( ~n13957 & n16179 ) ;
  assign n22184 = n20650 ^ n12453 ^ n10786 ;
  assign n22185 = n22184 ^ n12420 ^ n8309 ;
  assign n22186 = ( n11209 & n18157 ) | ( n11209 & n22185 ) | ( n18157 & n22185 ) ;
  assign n22187 = ( x160 & n22183 ) | ( x160 & ~n22186 ) | ( n22183 & ~n22186 ) ;
  assign n22188 = ( n4147 & ~n10743 ) | ( n4147 & n21824 ) | ( ~n10743 & n21824 ) ;
  assign n22189 = n18821 ^ n18609 ^ 1'b0 ;
  assign n22190 = ( n7936 & n15872 ) | ( n7936 & ~n22189 ) | ( n15872 & ~n22189 ) ;
  assign n22191 = ( n3701 & ~n22188 ) | ( n3701 & n22190 ) | ( ~n22188 & n22190 ) ;
  assign n22192 = n22191 ^ n14589 ^ 1'b0 ;
  assign n22193 = n19641 | n22192 ;
  assign n22194 = n21222 ^ n9931 ^ n6180 ;
  assign n22195 = n10286 ^ n4973 ^ 1'b0 ;
  assign n22196 = n5792 & n22195 ;
  assign n22197 = n22196 ^ n10055 ^ n7375 ;
  assign n22198 = ( n3546 & n8920 ) | ( n3546 & n22197 ) | ( n8920 & n22197 ) ;
  assign n22199 = ( n4946 & n22194 ) | ( n4946 & ~n22198 ) | ( n22194 & ~n22198 ) ;
  assign n22200 = ~n1381 & n19250 ;
  assign n22201 = n18591 & n22200 ;
  assign n22202 = n22117 ^ n21749 ^ n10667 ;
  assign n22203 = ( n2384 & n22201 ) | ( n2384 & n22202 ) | ( n22201 & n22202 ) ;
  assign n22204 = n6055 ^ n4745 ^ n4132 ;
  assign n22205 = n4219 ^ n4207 ^ 1'b0 ;
  assign n22206 = ( x199 & ~n22204 ) | ( x199 & n22205 ) | ( ~n22204 & n22205 ) ;
  assign n22211 = n13707 ^ n10410 ^ n8011 ;
  assign n22207 = n10778 ^ n10504 ^ 1'b0 ;
  assign n22208 = n16628 ^ n5578 ^ n2388 ;
  assign n22209 = x132 & n22208 ;
  assign n22210 = n22207 & n22209 ;
  assign n22212 = n22211 ^ n22210 ^ n11120 ;
  assign n22213 = n22039 ^ n21689 ^ n14987 ;
  assign n22214 = n14246 ^ n3663 ^ 1'b0 ;
  assign n22215 = ( n7293 & n7529 ) | ( n7293 & n22214 ) | ( n7529 & n22214 ) ;
  assign n22216 = ( n11068 & n12588 ) | ( n11068 & ~n22215 ) | ( n12588 & ~n22215 ) ;
  assign n22217 = ~n1967 & n1997 ;
  assign n22218 = ~n2388 & n22217 ;
  assign n22219 = ( n1901 & n2310 ) | ( n1901 & n5300 ) | ( n2310 & n5300 ) ;
  assign n22220 = ( n13943 & n21343 ) | ( n13943 & ~n22219 ) | ( n21343 & ~n22219 ) ;
  assign n22221 = n22220 ^ n3058 ^ 1'b0 ;
  assign n22222 = n22221 ^ n13549 ^ n1442 ;
  assign n22223 = ( n15508 & ~n22218 ) | ( n15508 & n22222 ) | ( ~n22218 & n22222 ) ;
  assign n22224 = ~n19217 & n20530 ;
  assign n22225 = n13003 ^ n5063 ^ 1'b0 ;
  assign n22226 = n9922 | n22225 ;
  assign n22227 = n22224 & ~n22226 ;
  assign n22228 = n9567 ^ n1591 ^ 1'b0 ;
  assign n22229 = n372 | n22228 ;
  assign n22230 = n19938 ^ n3188 ^ n883 ;
  assign n22231 = ( ~n768 & n13577 ) | ( ~n768 & n22230 ) | ( n13577 & n22230 ) ;
  assign n22240 = n4789 ^ n3298 ^ 1'b0 ;
  assign n22232 = n11617 ^ n1471 ^ 1'b0 ;
  assign n22233 = n7277 & ~n22232 ;
  assign n22234 = ( n5504 & n11263 ) | ( n5504 & ~n22233 ) | ( n11263 & ~n22233 ) ;
  assign n22235 = n7324 ^ n7172 ^ n1733 ;
  assign n22236 = ( ~n10010 & n21579 ) | ( ~n10010 & n22235 ) | ( n21579 & n22235 ) ;
  assign n22237 = n22234 & ~n22236 ;
  assign n22238 = ~n11347 & n22237 ;
  assign n22239 = ( n18973 & n19573 ) | ( n18973 & n22238 ) | ( n19573 & n22238 ) ;
  assign n22241 = n22240 ^ n22239 ^ n16410 ;
  assign n22254 = n11821 ^ n7459 ^ n1057 ;
  assign n22255 = ( n1346 & n14854 ) | ( n1346 & n22254 ) | ( n14854 & n22254 ) ;
  assign n22256 = n22255 ^ n14357 ^ n2162 ;
  assign n22257 = ( n6233 & ~n19520 ) | ( n6233 & n22256 ) | ( ~n19520 & n22256 ) ;
  assign n22242 = n1935 & n19314 ;
  assign n22250 = ~n1000 & n3075 ;
  assign n22251 = n22250 ^ n1527 ^ 1'b0 ;
  assign n22244 = ( n3749 & n5028 ) | ( n3749 & n10110 ) | ( n5028 & n10110 ) ;
  assign n22245 = n22244 ^ n657 ^ 1'b0 ;
  assign n22246 = n7040 & n22245 ;
  assign n22243 = n3425 | n8872 ;
  assign n22247 = n22246 ^ n22243 ^ 1'b0 ;
  assign n22248 = n22247 ^ n19787 ^ n540 ;
  assign n22249 = n8171 & n22248 ;
  assign n22252 = n22251 ^ n22249 ^ 1'b0 ;
  assign n22253 = ~n22242 & n22252 ;
  assign n22258 = n22257 ^ n22253 ^ 1'b0 ;
  assign n22259 = ( x0 & n3309 ) | ( x0 & ~n11464 ) | ( n3309 & ~n11464 ) ;
  assign n22264 = n2778 & ~n2840 ;
  assign n22265 = n1865 & n22264 ;
  assign n22262 = n4824 | n17771 ;
  assign n22260 = x17 & n8302 ;
  assign n22261 = n12733 & n22260 ;
  assign n22263 = n22262 ^ n22261 ^ 1'b0 ;
  assign n22266 = n22265 ^ n22263 ^ n12760 ;
  assign n22268 = n21313 ^ n17568 ^ n7455 ;
  assign n22269 = n22268 ^ n13057 ^ n6286 ;
  assign n22267 = n10947 & n17749 ;
  assign n22270 = n22269 ^ n22267 ^ 1'b0 ;
  assign n22271 = ( ~n2021 & n4194 ) | ( ~n2021 & n11576 ) | ( n4194 & n11576 ) ;
  assign n22272 = n22271 ^ n18798 ^ n18016 ;
  assign n22275 = n13081 ^ n11718 ^ n2851 ;
  assign n22273 = n18912 ^ n7287 ^ n3736 ;
  assign n22274 = ~n2505 & n22273 ;
  assign n22276 = n22275 ^ n22274 ^ 1'b0 ;
  assign n22277 = n22276 ^ n18034 ^ n16034 ;
  assign n22278 = n7842 ^ n3991 ^ n2322 ;
  assign n22279 = ( n1289 & ~n21802 ) | ( n1289 & n22278 ) | ( ~n21802 & n22278 ) ;
  assign n22280 = ( n3030 & ~n15002 ) | ( n3030 & n22279 ) | ( ~n15002 & n22279 ) ;
  assign n22281 = ( n3666 & n5829 ) | ( n3666 & n16861 ) | ( n5829 & n16861 ) ;
  assign n22282 = n10152 & ~n22281 ;
  assign n22283 = n22282 ^ n19243 ^ 1'b0 ;
  assign n22284 = n1053 & ~n22283 ;
  assign n22285 = ( n5253 & n6149 ) | ( n5253 & ~n20794 ) | ( n6149 & ~n20794 ) ;
  assign n22286 = n11260 & ~n22285 ;
  assign n22287 = n7685 & n22286 ;
  assign n22288 = ( n6973 & n9444 ) | ( n6973 & n13715 ) | ( n9444 & n13715 ) ;
  assign n22289 = n22288 ^ n22136 ^ n12337 ;
  assign n22290 = n16446 ^ n2444 ^ x224 ;
  assign n22291 = ( n9177 & n21032 ) | ( n9177 & ~n22290 ) | ( n21032 & ~n22290 ) ;
  assign n22293 = n11529 ^ n8441 ^ n3436 ;
  assign n22292 = n8891 ^ n6410 ^ 1'b0 ;
  assign n22294 = n22293 ^ n22292 ^ n13915 ;
  assign n22295 = ( n6923 & n10979 ) | ( n6923 & ~n22294 ) | ( n10979 & ~n22294 ) ;
  assign n22296 = n20898 ^ n14976 ^ n544 ;
  assign n22297 = n19839 & ~n22296 ;
  assign n22298 = n22297 ^ n17254 ^ n11579 ;
  assign n22303 = n21997 ^ n16693 ^ n10087 ;
  assign n22299 = ( ~n959 & n5874 ) | ( ~n959 & n6207 ) | ( n5874 & n6207 ) ;
  assign n22300 = n22299 ^ n19839 ^ n15867 ;
  assign n22301 = n6795 ^ n546 ^ 1'b0 ;
  assign n22302 = n22300 & n22301 ;
  assign n22304 = n22303 ^ n22302 ^ n11332 ;
  assign n22307 = n18723 ^ n11015 ^ n1274 ;
  assign n22308 = ( ~n12893 & n14742 ) | ( ~n12893 & n22307 ) | ( n14742 & n22307 ) ;
  assign n22305 = n5125 ^ n5101 ^ 1'b0 ;
  assign n22306 = n16135 & ~n22305 ;
  assign n22309 = n22308 ^ n22306 ^ n9940 ;
  assign n22310 = n5890 ^ n4316 ^ n1412 ;
  assign n22311 = ( n3748 & ~n5252 ) | ( n3748 & n22310 ) | ( ~n5252 & n22310 ) ;
  assign n22312 = ( ~n2178 & n4310 ) | ( ~n2178 & n22311 ) | ( n4310 & n22311 ) ;
  assign n22313 = n11674 | n22312 ;
  assign n22314 = n22313 ^ n3347 ^ n1311 ;
  assign n22315 = ( n1197 & n9461 ) | ( n1197 & ~n18976 ) | ( n9461 & ~n18976 ) ;
  assign n22319 = n9689 & ~n11396 ;
  assign n22320 = n22319 ^ n21059 ^ n4921 ;
  assign n22316 = ( n4300 & ~n5312 ) | ( n4300 & n6424 ) | ( ~n5312 & n6424 ) ;
  assign n22317 = n22316 ^ n17732 ^ 1'b0 ;
  assign n22318 = ( n11711 & ~n12065 ) | ( n11711 & n22317 ) | ( ~n12065 & n22317 ) ;
  assign n22321 = n22320 ^ n22318 ^ n10843 ;
  assign n22322 = n2099 & n11048 ;
  assign n22323 = n22322 ^ n4998 ^ 1'b0 ;
  assign n22324 = n22323 ^ n11433 ^ n6600 ;
  assign n22325 = n22324 ^ n7903 ^ n5421 ;
  assign n22326 = n10927 ^ n4401 ^ 1'b0 ;
  assign n22327 = n7918 & n11284 ;
  assign n22328 = n12494 ^ n7064 ^ n6609 ;
  assign n22329 = ( x156 & ~n2629 ) | ( x156 & n22328 ) | ( ~n2629 & n22328 ) ;
  assign n22330 = n22329 ^ n10950 ^ n4745 ;
  assign n22331 = n22330 ^ n7808 ^ n855 ;
  assign n22332 = ~n8674 & n16219 ;
  assign n22333 = ( n9094 & n21647 ) | ( n9094 & ~n22332 ) | ( n21647 & ~n22332 ) ;
  assign n22334 = n11270 ^ n2027 ^ 1'b0 ;
  assign n22335 = ( n17794 & n19193 ) | ( n17794 & ~n22334 ) | ( n19193 & ~n22334 ) ;
  assign n22336 = n3075 & n5352 ;
  assign n22337 = n22336 ^ n9366 ^ 1'b0 ;
  assign n22338 = ( n6041 & ~n21860 ) | ( n6041 & n22337 ) | ( ~n21860 & n22337 ) ;
  assign n22339 = ( n1510 & n2051 ) | ( n1510 & ~n22027 ) | ( n2051 & ~n22027 ) ;
  assign n22340 = ( n8215 & ~n22338 ) | ( n8215 & n22339 ) | ( ~n22338 & n22339 ) ;
  assign n22341 = n22340 ^ n4307 ^ n2144 ;
  assign n22342 = ( x236 & ~n3685 ) | ( x236 & n11645 ) | ( ~n3685 & n11645 ) ;
  assign n22343 = n2133 & ~n15098 ;
  assign n22344 = n22342 & n22343 ;
  assign n22345 = ( n820 & n1183 ) | ( n820 & n7578 ) | ( n1183 & n7578 ) ;
  assign n22346 = ( n5115 & ~n6523 ) | ( n5115 & n9689 ) | ( ~n6523 & n9689 ) ;
  assign n22349 = n3711 | n20833 ;
  assign n22347 = n15990 ^ n11771 ^ n6648 ;
  assign n22348 = ( n6200 & n10429 ) | ( n6200 & ~n22347 ) | ( n10429 & ~n22347 ) ;
  assign n22350 = n22349 ^ n22348 ^ x244 ;
  assign n22351 = ( n22345 & n22346 ) | ( n22345 & ~n22350 ) | ( n22346 & ~n22350 ) ;
  assign n22352 = n20582 ^ n15615 ^ n6341 ;
  assign n22353 = ~n14861 & n22352 ;
  assign n22354 = n11754 ^ n9445 ^ n825 ;
  assign n22355 = n10947 ^ n483 ^ 1'b0 ;
  assign n22356 = n22355 ^ n16371 ^ 1'b0 ;
  assign n22363 = ( n665 & ~n8916 ) | ( n665 & n12743 ) | ( ~n8916 & n12743 ) ;
  assign n22359 = n9591 & n20310 ;
  assign n22360 = n22359 ^ n21529 ^ 1'b0 ;
  assign n22357 = n1839 | n12084 ;
  assign n22358 = n22357 ^ n4395 ^ 1'b0 ;
  assign n22361 = n22360 ^ n22358 ^ n4968 ;
  assign n22362 = ( n4490 & n15102 ) | ( n4490 & n22361 ) | ( n15102 & n22361 ) ;
  assign n22364 = n22363 ^ n22362 ^ n2836 ;
  assign n22365 = ( n11760 & n12425 ) | ( n11760 & ~n12874 ) | ( n12425 & ~n12874 ) ;
  assign n22366 = n22365 ^ n9342 ^ 1'b0 ;
  assign n22367 = ~n7987 & n22366 ;
  assign n22368 = n12803 ^ n11444 ^ n2557 ;
  assign n22369 = n15072 ^ n6088 ^ n2785 ;
  assign n22370 = ( n3627 & n22368 ) | ( n3627 & ~n22369 ) | ( n22368 & ~n22369 ) ;
  assign n22371 = ( ~n20259 & n20941 ) | ( ~n20259 & n21180 ) | ( n20941 & n21180 ) ;
  assign n22372 = ( n5594 & ~n6875 ) | ( n5594 & n9728 ) | ( ~n6875 & n9728 ) ;
  assign n22373 = n17362 ^ n8978 ^ n7611 ;
  assign n22374 = n22373 ^ n4772 ^ n2938 ;
  assign n22375 = n22374 ^ n13058 ^ 1'b0 ;
  assign n22376 = n22372 | n22375 ;
  assign n22377 = ( n5418 & n14711 ) | ( n5418 & ~n14889 ) | ( n14711 & ~n14889 ) ;
  assign n22378 = n6028 & ~n22377 ;
  assign n22379 = n22378 ^ n4513 ^ 1'b0 ;
  assign n22380 = n16336 ^ n3277 ^ 1'b0 ;
  assign n22381 = n22380 ^ n17594 ^ n3911 ;
  assign n22382 = ( n2256 & ~n5622 ) | ( n2256 & n20001 ) | ( ~n5622 & n20001 ) ;
  assign n22383 = ( ~n3448 & n4091 ) | ( ~n3448 & n7810 ) | ( n4091 & n7810 ) ;
  assign n22384 = x175 & n2901 ;
  assign n22385 = n22383 & n22384 ;
  assign n22386 = n1057 & n3643 ;
  assign n22387 = n22386 ^ n8533 ^ 1'b0 ;
  assign n22388 = ( ~n2813 & n5618 ) | ( ~n2813 & n15562 ) | ( n5618 & n15562 ) ;
  assign n22389 = ( n16916 & n19253 ) | ( n16916 & n22388 ) | ( n19253 & n22388 ) ;
  assign n22390 = n22389 ^ n13804 ^ 1'b0 ;
  assign n22391 = n6703 & ~n22390 ;
  assign n22392 = n22391 ^ n21047 ^ n17467 ;
  assign n22393 = ( ~n3862 & n22387 ) | ( ~n3862 & n22392 ) | ( n22387 & n22392 ) ;
  assign n22394 = n4145 ^ n2224 ^ 1'b0 ;
  assign n22395 = ( ~n2521 & n13040 ) | ( ~n2521 & n22394 ) | ( n13040 & n22394 ) ;
  assign n22396 = ( ~n12294 & n22393 ) | ( ~n12294 & n22395 ) | ( n22393 & n22395 ) ;
  assign n22397 = n12961 ^ n5837 ^ n3255 ;
  assign n22398 = n19991 & ~n22397 ;
  assign n22399 = n12248 & n22398 ;
  assign n22400 = n16028 ^ n6699 ^ n312 ;
  assign n22401 = n22400 ^ n18450 ^ n3850 ;
  assign n22402 = n22401 ^ n5977 ^ 1'b0 ;
  assign n22403 = ( n19525 & n22399 ) | ( n19525 & ~n22402 ) | ( n22399 & ~n22402 ) ;
  assign n22404 = n3199 & n11405 ;
  assign n22405 = n22404 ^ n21270 ^ 1'b0 ;
  assign n22406 = n4341 & n7866 ;
  assign n22407 = n19197 ^ n6254 ^ n1656 ;
  assign n22408 = n22407 ^ n19577 ^ n1266 ;
  assign n22409 = ( ~n22405 & n22406 ) | ( ~n22405 & n22408 ) | ( n22406 & n22408 ) ;
  assign n22410 = n8928 ^ n3879 ^ n2382 ;
  assign n22411 = n22410 ^ n11526 ^ n1469 ;
  assign n22412 = n22411 ^ n9026 ^ n2322 ;
  assign n22413 = ( n3117 & n12564 ) | ( n3117 & n22412 ) | ( n12564 & n22412 ) ;
  assign n22415 = n2736 & ~n21483 ;
  assign n22414 = n18342 ^ n10594 ^ n9351 ;
  assign n22416 = n22415 ^ n22414 ^ n3636 ;
  assign n22417 = n10071 ^ n6887 ^ n6433 ;
  assign n22418 = ( n4760 & ~n6913 ) | ( n4760 & n22417 ) | ( ~n6913 & n22417 ) ;
  assign n22419 = ~n22416 & n22418 ;
  assign n22420 = n22413 & n22419 ;
  assign n22421 = n16652 ^ n11202 ^ n3567 ;
  assign n22426 = n21320 ^ n1219 ^ 1'b0 ;
  assign n22423 = n5742 & n16819 ;
  assign n22424 = n22423 ^ n6342 ^ 1'b0 ;
  assign n22425 = ( n9502 & n14339 ) | ( n9502 & ~n22424 ) | ( n14339 & ~n22424 ) ;
  assign n22422 = n11605 ^ n8452 ^ n7886 ;
  assign n22427 = n22426 ^ n22425 ^ n22422 ;
  assign n22428 = n22427 ^ n17832 ^ n7650 ;
  assign n22429 = n11057 ^ n5464 ^ n5297 ;
  assign n22430 = ( n6158 & ~n14094 ) | ( n6158 & n22429 ) | ( ~n14094 & n22429 ) ;
  assign n22431 = ( n281 & n9060 ) | ( n281 & ~n10189 ) | ( n9060 & ~n10189 ) ;
  assign n22432 = n269 | n20290 ;
  assign n22433 = n22431 & ~n22432 ;
  assign n22434 = n22430 | n22433 ;
  assign n22435 = n22434 ^ n3975 ^ 1'b0 ;
  assign n22436 = n5019 ^ n2355 ^ 1'b0 ;
  assign n22437 = n22435 & n22436 ;
  assign n22438 = n18296 ^ n9737 ^ n8624 ;
  assign n22439 = n12931 & n17758 ;
  assign n22440 = n22439 ^ n8690 ^ 1'b0 ;
  assign n22441 = n9279 ^ n547 ^ 1'b0 ;
  assign n22442 = n17177 ^ n12097 ^ n2486 ;
  assign n22443 = ( ~n3109 & n8111 ) | ( ~n3109 & n8555 ) | ( n8111 & n8555 ) ;
  assign n22444 = ( n8706 & n9688 ) | ( n8706 & n22443 ) | ( n9688 & n22443 ) ;
  assign n22447 = n19097 ^ n14982 ^ n6554 ;
  assign n22445 = n20839 ^ n12323 ^ n3923 ;
  assign n22446 = n22445 ^ n15960 ^ n15613 ;
  assign n22448 = n22447 ^ n22446 ^ n734 ;
  assign n22449 = n12731 ^ n1774 ^ n1180 ;
  assign n22450 = ( n3148 & n10241 ) | ( n3148 & n22449 ) | ( n10241 & n22449 ) ;
  assign n22454 = n9020 ^ n6458 ^ n4126 ;
  assign n22452 = ( n321 & n369 ) | ( n321 & n15313 ) | ( n369 & n15313 ) ;
  assign n22451 = n9453 ^ n5172 ^ n4643 ;
  assign n22453 = n22452 ^ n22451 ^ n21025 ;
  assign n22455 = n22454 ^ n22453 ^ n12477 ;
  assign n22468 = n16058 ^ n10906 ^ n5629 ;
  assign n22469 = n3920 & ~n22468 ;
  assign n22464 = n13418 ^ n7384 ^ n2101 ;
  assign n22465 = n22464 ^ n4291 ^ 1'b0 ;
  assign n22466 = n7748 & n22465 ;
  assign n22461 = ( n1352 & ~n17110 ) | ( n1352 & n17710 ) | ( ~n17110 & n17710 ) ;
  assign n22462 = n2956 & n8045 ;
  assign n22463 = ~n22461 & n22462 ;
  assign n22460 = n14008 ^ n8945 ^ n1974 ;
  assign n22467 = n22466 ^ n22463 ^ n22460 ;
  assign n22456 = n2905 & ~n10130 ;
  assign n22457 = ~n6878 & n22456 ;
  assign n22458 = ( n9333 & ~n9823 ) | ( n9333 & n22457 ) | ( ~n9823 & n22457 ) ;
  assign n22459 = n22458 ^ n5675 ^ n1698 ;
  assign n22470 = n22469 ^ n22467 ^ n22459 ;
  assign n22471 = n7227 | n8924 ;
  assign n22472 = n22471 ^ n17565 ^ n4465 ;
  assign n22473 = ( n1443 & n16917 ) | ( n1443 & n22472 ) | ( n16917 & n22472 ) ;
  assign n22474 = ( n11323 & ~n20041 ) | ( n11323 & n22473 ) | ( ~n20041 & n22473 ) ;
  assign n22475 = ( n7958 & n20904 ) | ( n7958 & ~n22474 ) | ( n20904 & ~n22474 ) ;
  assign n22476 = ( n13868 & n16423 ) | ( n13868 & n17261 ) | ( n16423 & n17261 ) ;
  assign n22477 = n20458 ^ n8335 ^ 1'b0 ;
  assign n22478 = ~n22476 & n22477 ;
  assign n22482 = ( ~n7940 & n9730 ) | ( ~n7940 & n15648 ) | ( n9730 & n15648 ) ;
  assign n22479 = n8841 ^ n6491 ^ 1'b0 ;
  assign n22480 = n2458 & n22479 ;
  assign n22481 = n22480 ^ n12902 ^ n5782 ;
  assign n22483 = n22482 ^ n22481 ^ n3723 ;
  assign n22484 = n19625 ^ n14174 ^ n7788 ;
  assign n22485 = n3057 ^ n1849 ^ 1'b0 ;
  assign n22486 = n22485 ^ n7789 ^ n5498 ;
  assign n22487 = ( x77 & n22484 ) | ( x77 & ~n22486 ) | ( n22484 & ~n22486 ) ;
  assign n22488 = ( n12992 & n19232 ) | ( n12992 & n20152 ) | ( n19232 & n20152 ) ;
  assign n22489 = n22488 ^ n7789 ^ n7559 ;
  assign n22490 = n7107 & n15758 ;
  assign n22491 = ( ~n8989 & n13812 ) | ( ~n8989 & n22490 ) | ( n13812 & n22490 ) ;
  assign n22492 = n17781 & ~n22491 ;
  assign n22493 = n12006 & n22492 ;
  assign n22494 = n7650 ^ n3724 ^ n3070 ;
  assign n22495 = n20584 ^ n17327 ^ n2972 ;
  assign n22496 = ( n8777 & ~n22494 ) | ( n8777 & n22495 ) | ( ~n22494 & n22495 ) ;
  assign n22497 = n22496 ^ n2568 ^ 1'b0 ;
  assign n22498 = ~n4164 & n22497 ;
  assign n22499 = ( ~n7066 & n22493 ) | ( ~n7066 & n22498 ) | ( n22493 & n22498 ) ;
  assign n22500 = n4920 ^ n1131 ^ x134 ;
  assign n22501 = ( n12946 & n13356 ) | ( n12946 & n22500 ) | ( n13356 & n22500 ) ;
  assign n22503 = ( n1008 & ~n6615 ) | ( n1008 & n8525 ) | ( ~n6615 & n8525 ) ;
  assign n22504 = n14132 ^ n5261 ^ 1'b0 ;
  assign n22505 = n22504 ^ n12623 ^ n2405 ;
  assign n22506 = ( ~n7254 & n22503 ) | ( ~n7254 & n22505 ) | ( n22503 & n22505 ) ;
  assign n22502 = n21844 ^ n5295 ^ n3622 ;
  assign n22507 = n22506 ^ n22502 ^ n1028 ;
  assign n22508 = n10358 | n21628 ;
  assign n22511 = ( n4031 & n4263 ) | ( n4031 & n7492 ) | ( n4263 & n7492 ) ;
  assign n22510 = n17815 ^ n15438 ^ n7002 ;
  assign n22512 = n22511 ^ n22510 ^ n10392 ;
  assign n22509 = n4098 ^ x29 ^ 1'b0 ;
  assign n22513 = n22512 ^ n22509 ^ n15647 ;
  assign n22517 = ( n4371 & n6019 ) | ( n4371 & ~n15505 ) | ( n6019 & ~n15505 ) ;
  assign n22514 = ( n6477 & n6574 ) | ( n6477 & n10738 ) | ( n6574 & n10738 ) ;
  assign n22515 = ( n5820 & n9050 ) | ( n5820 & n12502 ) | ( n9050 & n12502 ) ;
  assign n22516 = ( n1262 & ~n22514 ) | ( n1262 & n22515 ) | ( ~n22514 & n22515 ) ;
  assign n22518 = n22517 ^ n22516 ^ n5852 ;
  assign n22519 = n16828 ^ n8500 ^ n5736 ;
  assign n22520 = n22519 ^ n16037 ^ n1085 ;
  assign n22521 = n18823 ^ n15393 ^ n3720 ;
  assign n22522 = ~n17482 & n22521 ;
  assign n22523 = n22522 ^ n1783 ^ 1'b0 ;
  assign n22524 = n6999 ^ n5401 ^ n3329 ;
  assign n22525 = n7612 | n7877 ;
  assign n22526 = ( n5618 & ~n22524 ) | ( n5618 & n22525 ) | ( ~n22524 & n22525 ) ;
  assign n22527 = n14356 ^ n5546 ^ n752 ;
  assign n22528 = ~n12042 & n18025 ;
  assign n22529 = ~n1407 & n8718 ;
  assign n22537 = ( n1499 & n4740 ) | ( n1499 & ~n13258 ) | ( n4740 & ~n13258 ) ;
  assign n22535 = n18744 ^ n2767 ^ 1'b0 ;
  assign n22534 = ~n8613 & n11987 ;
  assign n22536 = n22535 ^ n22534 ^ n15860 ;
  assign n22538 = n22537 ^ n22536 ^ n14352 ;
  assign n22530 = n20409 ^ n9318 ^ n2602 ;
  assign n22531 = n22530 ^ n11307 ^ n609 ;
  assign n22532 = n3579 & ~n7368 ;
  assign n22533 = n22531 & n22532 ;
  assign n22539 = n22538 ^ n22533 ^ n20363 ;
  assign n22540 = ( n22528 & ~n22529 ) | ( n22528 & n22539 ) | ( ~n22529 & n22539 ) ;
  assign n22541 = ( n1822 & n7046 ) | ( n1822 & ~n16098 ) | ( n7046 & ~n16098 ) ;
  assign n22542 = n13219 & ~n18358 ;
  assign n22543 = n22541 | n22542 ;
  assign n22544 = ( n6502 & ~n8166 ) | ( n6502 & n9386 ) | ( ~n8166 & n9386 ) ;
  assign n22545 = n22544 ^ n21626 ^ n7581 ;
  assign n22551 = n2444 ^ n1034 ^ x37 ;
  assign n22548 = n8853 ^ n3718 ^ x21 ;
  assign n22546 = n4593 | n14974 ;
  assign n22547 = n22546 ^ n5312 ^ 1'b0 ;
  assign n22549 = n22548 ^ n22547 ^ n4533 ;
  assign n22550 = n22549 ^ n13329 ^ n814 ;
  assign n22552 = n22551 ^ n22550 ^ n17713 ;
  assign n22553 = ( n4254 & n9181 ) | ( n4254 & ~n13460 ) | ( n9181 & ~n13460 ) ;
  assign n22554 = n12286 ^ n11306 ^ n8330 ;
  assign n22555 = ( n2478 & n3947 ) | ( n2478 & n6293 ) | ( n3947 & n6293 ) ;
  assign n22556 = ( n1361 & n22554 ) | ( n1361 & ~n22555 ) | ( n22554 & ~n22555 ) ;
  assign n22557 = n22556 ^ n850 ^ 1'b0 ;
  assign n22558 = ~n1495 & n22557 ;
  assign n22567 = ( x105 & n1262 ) | ( x105 & ~n1289 ) | ( n1262 & ~n1289 ) ;
  assign n22568 = ( ~n836 & n10565 ) | ( ~n836 & n22567 ) | ( n10565 & n22567 ) ;
  assign n22569 = ( n8291 & n10883 ) | ( n8291 & n22568 ) | ( n10883 & n22568 ) ;
  assign n22563 = n2051 ^ n584 ^ 1'b0 ;
  assign n22564 = ~n6772 & n22563 ;
  assign n22565 = n11633 | n22564 ;
  assign n22559 = n11017 ^ n8470 ^ x74 ;
  assign n22560 = n20217 ^ n16810 ^ x103 ;
  assign n22561 = ( n2477 & ~n16802 ) | ( n2477 & n22560 ) | ( ~n16802 & n22560 ) ;
  assign n22562 = ( ~n16842 & n22559 ) | ( ~n16842 & n22561 ) | ( n22559 & n22561 ) ;
  assign n22566 = n22565 ^ n22562 ^ n6337 ;
  assign n22570 = n22569 ^ n22566 ^ n15947 ;
  assign n22572 = ( ~n4798 & n6042 ) | ( ~n4798 & n8312 ) | ( n6042 & n8312 ) ;
  assign n22573 = ( ~n6317 & n6997 ) | ( ~n6317 & n17180 ) | ( n6997 & n17180 ) ;
  assign n22574 = ( n4699 & n22073 ) | ( n4699 & n22573 ) | ( n22073 & n22573 ) ;
  assign n22575 = ( ~n4523 & n12211 ) | ( ~n4523 & n22574 ) | ( n12211 & n22574 ) ;
  assign n22576 = n18334 | n22575 ;
  assign n22577 = n22572 | n22576 ;
  assign n22578 = ( n693 & n7270 ) | ( n693 & ~n22577 ) | ( n7270 & ~n22577 ) ;
  assign n22571 = ( ~n4961 & n5140 ) | ( ~n4961 & n6237 ) | ( n5140 & n6237 ) ;
  assign n22579 = n22578 ^ n22571 ^ n4277 ;
  assign n22588 = ( n1892 & n3091 ) | ( n1892 & ~n19117 ) | ( n3091 & ~n19117 ) ;
  assign n22583 = n8205 & n13479 ;
  assign n22581 = n3015 ^ n281 ^ 1'b0 ;
  assign n22580 = n15778 ^ n11591 ^ 1'b0 ;
  assign n22582 = n22581 ^ n22580 ^ n20540 ;
  assign n22584 = n22583 ^ n22582 ^ n15063 ;
  assign n22585 = ( n7196 & n12857 ) | ( n7196 & ~n22484 ) | ( n12857 & ~n22484 ) ;
  assign n22586 = n22585 ^ n17037 ^ n15029 ;
  assign n22587 = ( n21357 & ~n22584 ) | ( n21357 & n22586 ) | ( ~n22584 & n22586 ) ;
  assign n22589 = n22588 ^ n22587 ^ n1660 ;
  assign n22591 = ( n3452 & ~n5858 ) | ( n3452 & n11341 ) | ( ~n5858 & n11341 ) ;
  assign n22590 = n19295 ^ n18422 ^ 1'b0 ;
  assign n22592 = n22591 ^ n22590 ^ n4091 ;
  assign n22593 = n11267 ^ n3737 ^ n2668 ;
  assign n22594 = n22593 ^ n10314 ^ 1'b0 ;
  assign n22595 = n3175 & ~n11485 ;
  assign n22596 = n8600 & n10671 ;
  assign n22597 = n22510 ^ n21234 ^ n11946 ;
  assign n22598 = ( n1303 & ~n3439 ) | ( n1303 & n21390 ) | ( ~n3439 & n21390 ) ;
  assign n22599 = ( n2437 & n7316 ) | ( n2437 & n22598 ) | ( n7316 & n22598 ) ;
  assign n22600 = n5681 | n21802 ;
  assign n22601 = n1416 ^ n685 ^ n345 ;
  assign n22602 = ( n5444 & n22600 ) | ( n5444 & n22601 ) | ( n22600 & n22601 ) ;
  assign n22603 = ( ~n10624 & n22599 ) | ( ~n10624 & n22602 ) | ( n22599 & n22602 ) ;
  assign n22604 = n22597 & ~n22603 ;
  assign n22605 = ( ~n12637 & n13476 ) | ( ~n12637 & n22604 ) | ( n13476 & n22604 ) ;
  assign n22606 = n22596 & ~n22605 ;
  assign n22607 = n22606 ^ n3759 ^ 1'b0 ;
  assign n22608 = n14861 | n15336 ;
  assign n22609 = ( n4149 & n4757 ) | ( n4149 & n16675 ) | ( n4757 & n16675 ) ;
  assign n22610 = ( n16748 & n19294 ) | ( n16748 & n22609 ) | ( n19294 & n22609 ) ;
  assign n22611 = ~n676 & n2529 ;
  assign n22612 = n8924 & n22611 ;
  assign n22613 = n22612 ^ n11194 ^ n8244 ;
  assign n22614 = ( n406 & n15961 ) | ( n406 & n22613 ) | ( n15961 & n22613 ) ;
  assign n22620 = n13187 ^ n2366 ^ n1124 ;
  assign n22617 = n11907 ^ n10370 ^ n4244 ;
  assign n22618 = n22617 ^ n10404 ^ 1'b0 ;
  assign n22619 = ( ~n1560 & n3050 ) | ( ~n1560 & n22618 ) | ( n3050 & n22618 ) ;
  assign n22621 = n22620 ^ n22619 ^ n8235 ;
  assign n22622 = ~n684 & n22621 ;
  assign n22615 = ( n3469 & ~n6251 ) | ( n3469 & n8978 ) | ( ~n6251 & n8978 ) ;
  assign n22616 = n16443 & ~n22615 ;
  assign n22623 = n22622 ^ n22616 ^ 1'b0 ;
  assign n22624 = ( n5101 & n19591 ) | ( n5101 & n21583 ) | ( n19591 & n21583 ) ;
  assign n22626 = n8113 ^ n7680 ^ n4595 ;
  assign n22627 = ( n1491 & ~n6686 ) | ( n1491 & n8735 ) | ( ~n6686 & n8735 ) ;
  assign n22628 = ~n12411 & n22627 ;
  assign n22629 = n22626 & n22628 ;
  assign n22625 = n12822 ^ n12486 ^ n6526 ;
  assign n22630 = n22629 ^ n22625 ^ n4050 ;
  assign n22631 = n7849 | n16164 ;
  assign n22632 = n22630 & ~n22631 ;
  assign n22633 = ( n8554 & n19361 ) | ( n8554 & n22632 ) | ( n19361 & n22632 ) ;
  assign n22634 = ( n1565 & n3188 ) | ( n1565 & ~n7925 ) | ( n3188 & ~n7925 ) ;
  assign n22635 = ( ~x194 & n22633 ) | ( ~x194 & n22634 ) | ( n22633 & n22634 ) ;
  assign n22636 = x74 & ~n3753 ;
  assign n22637 = ( n4670 & n13851 ) | ( n4670 & n22636 ) | ( n13851 & n22636 ) ;
  assign n22638 = n17632 ^ n9883 ^ n9261 ;
  assign n22639 = ( n16190 & n22637 ) | ( n16190 & n22638 ) | ( n22637 & n22638 ) ;
  assign n22640 = n6430 & n9283 ;
  assign n22641 = n22640 ^ n2306 ^ 1'b0 ;
  assign n22642 = n22641 ^ n13229 ^ n3059 ;
  assign n22644 = n7966 ^ n5824 ^ n5082 ;
  assign n22645 = ( ~n962 & n1795 ) | ( ~n962 & n12713 ) | ( n1795 & n12713 ) ;
  assign n22646 = n22645 ^ n1155 ^ 1'b0 ;
  assign n22647 = n22644 | n22646 ;
  assign n22643 = n14175 ^ n8392 ^ n6480 ;
  assign n22648 = n22647 ^ n22643 ^ 1'b0 ;
  assign n22649 = ( n1324 & ~n3891 ) | ( n1324 & n16806 ) | ( ~n3891 & n16806 ) ;
  assign n22650 = n22649 ^ n4867 ^ 1'b0 ;
  assign n22655 = n14336 ^ n13162 ^ n12226 ;
  assign n22656 = ( n1130 & n2504 ) | ( n1130 & n22655 ) | ( n2504 & n22655 ) ;
  assign n22657 = n22656 ^ n7181 ^ n4746 ;
  assign n22651 = n2542 ^ n2424 ^ 1'b0 ;
  assign n22652 = ( n937 & n6428 ) | ( n937 & n22651 ) | ( n6428 & n22651 ) ;
  assign n22653 = ( n8793 & n21388 ) | ( n8793 & ~n22652 ) | ( n21388 & ~n22652 ) ;
  assign n22654 = n4795 | n22653 ;
  assign n22658 = n22657 ^ n22654 ^ 1'b0 ;
  assign n22659 = n22658 ^ n9941 ^ 1'b0 ;
  assign n22660 = n22104 & n22659 ;
  assign n22662 = n19419 ^ n15871 ^ n7123 ;
  assign n22661 = n19794 ^ n1543 ^ 1'b0 ;
  assign n22663 = n22662 ^ n22661 ^ n5543 ;
  assign n22670 = n13790 ^ n7965 ^ n1540 ;
  assign n22664 = n6160 & ~n11054 ;
  assign n22665 = ( ~n6144 & n12491 ) | ( ~n6144 & n13545 ) | ( n12491 & n13545 ) ;
  assign n22666 = ( n10509 & n22664 ) | ( n10509 & n22665 ) | ( n22664 & n22665 ) ;
  assign n22667 = ( n6168 & n21034 ) | ( n6168 & ~n22666 ) | ( n21034 & ~n22666 ) ;
  assign n22668 = n20048 & n22667 ;
  assign n22669 = n22668 ^ n5219 ^ 1'b0 ;
  assign n22671 = n22670 ^ n22669 ^ n2762 ;
  assign n22672 = ( n2302 & ~n9969 ) | ( n2302 & n22671 ) | ( ~n9969 & n22671 ) ;
  assign n22673 = n22672 ^ n16047 ^ n2439 ;
  assign n22674 = ( n903 & n15848 ) | ( n903 & n22673 ) | ( n15848 & n22673 ) ;
  assign n22675 = ( n6233 & n14767 ) | ( n6233 & n19670 ) | ( n14767 & n19670 ) ;
  assign n22683 = n12161 ^ n6586 ^ n4520 ;
  assign n22684 = n5135 & n22683 ;
  assign n22685 = n22684 ^ n18046 ^ 1'b0 ;
  assign n22682 = n8741 ^ n4115 ^ n3012 ;
  assign n22680 = n4643 & ~n5677 ;
  assign n22681 = ( n7557 & ~n15093 ) | ( n7557 & n22680 ) | ( ~n15093 & n22680 ) ;
  assign n22686 = n22685 ^ n22682 ^ n22681 ;
  assign n22676 = ( x189 & ~n3085 ) | ( x189 & n8945 ) | ( ~n3085 & n8945 ) ;
  assign n22677 = ~n1428 & n22676 ;
  assign n22678 = n22677 ^ n5523 ^ 1'b0 ;
  assign n22679 = n19668 & n22678 ;
  assign n22687 = n22686 ^ n22679 ^ 1'b0 ;
  assign n22700 = n7812 ^ n7028 ^ 1'b0 ;
  assign n22701 = ~n6408 & n22700 ;
  assign n22702 = n22701 ^ n17153 ^ n1515 ;
  assign n22703 = n22702 ^ n16743 ^ n7722 ;
  assign n22689 = ( ~n5926 & n9424 ) | ( ~n5926 & n17401 ) | ( n9424 & n17401 ) ;
  assign n22690 = n10576 & ~n19942 ;
  assign n22691 = n22690 ^ n19623 ^ 1'b0 ;
  assign n22696 = ( n5360 & n11577 ) | ( n5360 & ~n14905 ) | ( n11577 & ~n14905 ) ;
  assign n22693 = ( n661 & n770 ) | ( n661 & n8890 ) | ( n770 & n8890 ) ;
  assign n22694 = ( n12036 & n20857 ) | ( n12036 & ~n22693 ) | ( n20857 & ~n22693 ) ;
  assign n22695 = ( n12333 & n14400 ) | ( n12333 & ~n22694 ) | ( n14400 & ~n22694 ) ;
  assign n22692 = n17828 ^ n14974 ^ n11918 ;
  assign n22697 = n22696 ^ n22695 ^ n22692 ;
  assign n22698 = ( n22689 & ~n22691 ) | ( n22689 & n22697 ) | ( ~n22691 & n22697 ) ;
  assign n22699 = n22698 ^ n14171 ^ n7286 ;
  assign n22688 = n11682 ^ n5294 ^ 1'b0 ;
  assign n22704 = n22703 ^ n22699 ^ n22688 ;
  assign n22705 = ( n8418 & n18009 ) | ( n8418 & n20235 ) | ( n18009 & n20235 ) ;
  assign n22706 = ( n1416 & n3158 ) | ( n1416 & n11086 ) | ( n3158 & n11086 ) ;
  assign n22707 = ( n1203 & n1661 ) | ( n1203 & ~n22706 ) | ( n1661 & ~n22706 ) ;
  assign n22708 = n6519 ^ n4867 ^ n4672 ;
  assign n22709 = n22708 ^ n11636 ^ n6983 ;
  assign n22710 = ~n10653 & n20768 ;
  assign n22711 = n22710 ^ n15316 ^ n3995 ;
  assign n22712 = n15637 ^ n13236 ^ 1'b0 ;
  assign n22713 = n19251 ^ n1283 ^ n1055 ;
  assign n22714 = n14335 ^ n6623 ^ 1'b0 ;
  assign n22715 = ( n12338 & ~n22713 ) | ( n12338 & n22714 ) | ( ~n22713 & n22714 ) ;
  assign n22716 = ( n1598 & n9066 ) | ( n1598 & n22715 ) | ( n9066 & n22715 ) ;
  assign n22721 = ( n7714 & ~n11252 ) | ( n7714 & n12952 ) | ( ~n11252 & n12952 ) ;
  assign n22722 = n22721 ^ n7021 ^ n5518 ;
  assign n22723 = n22722 ^ n17456 ^ 1'b0 ;
  assign n22719 = ~n1350 & n5564 ;
  assign n22720 = ( n6821 & n8699 ) | ( n6821 & n22719 ) | ( n8699 & n22719 ) ;
  assign n22717 = n5343 ^ n3705 ^ n1980 ;
  assign n22718 = n22717 ^ n18296 ^ n3636 ;
  assign n22724 = n22723 ^ n22720 ^ n22718 ;
  assign n22725 = n22724 ^ n22717 ^ n7833 ;
  assign n22726 = n22725 ^ n19500 ^ n12587 ;
  assign n22728 = ( n6316 & n10111 ) | ( n6316 & ~n20293 ) | ( n10111 & ~n20293 ) ;
  assign n22727 = n15875 ^ n15065 ^ n2268 ;
  assign n22729 = n22728 ^ n22727 ^ n9847 ;
  assign n22730 = ( n6317 & n17054 ) | ( n6317 & ~n18090 ) | ( n17054 & ~n18090 ) ;
  assign n22731 = ( n10555 & n13768 ) | ( n10555 & ~n22730 ) | ( n13768 & ~n22730 ) ;
  assign n22732 = n22731 ^ n17058 ^ 1'b0 ;
  assign n22733 = ( n11075 & n22729 ) | ( n11075 & n22732 ) | ( n22729 & n22732 ) ;
  assign n22734 = ( ~n5087 & n13814 ) | ( ~n5087 & n19204 ) | ( n13814 & n19204 ) ;
  assign n22735 = ( n4235 & ~n12290 ) | ( n4235 & n22734 ) | ( ~n12290 & n22734 ) ;
  assign n22736 = n9730 ^ n9040 ^ n4882 ;
  assign n22737 = ( n5498 & n19829 ) | ( n5498 & n22736 ) | ( n19829 & n22736 ) ;
  assign n22738 = ~n454 & n9497 ;
  assign n22743 = n19121 ^ n6315 ^ n709 ;
  assign n22739 = ( n286 & ~n17438 ) | ( n286 & n18078 ) | ( ~n17438 & n18078 ) ;
  assign n22740 = n11051 ^ n10304 ^ n5662 ;
  assign n22741 = ( n16872 & n22739 ) | ( n16872 & ~n22740 ) | ( n22739 & ~n22740 ) ;
  assign n22742 = ( ~n15826 & n15892 ) | ( ~n15826 & n22741 ) | ( n15892 & n22741 ) ;
  assign n22744 = n22743 ^ n22742 ^ n11733 ;
  assign n22745 = n12117 ^ n11653 ^ n9066 ;
  assign n22746 = n15601 ^ n13900 ^ n5226 ;
  assign n22747 = n22746 ^ n1694 ^ 1'b0 ;
  assign n22748 = n20812 ^ n13570 ^ n8269 ;
  assign n22749 = n7901 ^ n7588 ^ n4540 ;
  assign n22750 = n22749 ^ n10009 ^ 1'b0 ;
  assign n22751 = n22750 ^ n15856 ^ n9788 ;
  assign n22757 = ( ~n5847 & n7646 ) | ( ~n5847 & n21424 ) | ( n7646 & n21424 ) ;
  assign n22758 = ( n9771 & ~n15219 ) | ( n9771 & n22757 ) | ( ~n15219 & n22757 ) ;
  assign n22752 = n17418 ^ n1249 ^ 1'b0 ;
  assign n22753 = n4851 & ~n22752 ;
  assign n22754 = n22753 ^ n21839 ^ n11354 ;
  assign n22755 = ( n7780 & n19112 ) | ( n7780 & n22754 ) | ( n19112 & n22754 ) ;
  assign n22756 = n22755 ^ n15433 ^ n11288 ;
  assign n22759 = n22758 ^ n22756 ^ n2105 ;
  assign n22760 = ( n5240 & ~n7260 ) | ( n5240 & n13047 ) | ( ~n7260 & n13047 ) ;
  assign n22761 = n1155 & ~n13051 ;
  assign n22762 = n22761 ^ n10620 ^ 1'b0 ;
  assign n22763 = n22762 ^ n16095 ^ n5994 ;
  assign n22764 = n20495 ^ n19812 ^ 1'b0 ;
  assign n22765 = ( ~n4665 & n20117 ) | ( ~n4665 & n22764 ) | ( n20117 & n22764 ) ;
  assign n22766 = n13822 ^ n11671 ^ n5427 ;
  assign n22767 = ( n2268 & n21111 ) | ( n2268 & ~n22766 ) | ( n21111 & ~n22766 ) ;
  assign n22769 = n5718 ^ n3019 ^ x227 ;
  assign n22768 = n11007 ^ n3164 ^ 1'b0 ;
  assign n22770 = n22769 ^ n22768 ^ n11588 ;
  assign n22771 = ( n849 & ~n1894 ) | ( n849 & n22770 ) | ( ~n1894 & n22770 ) ;
  assign n22772 = n9390 ^ n1262 ^ n382 ;
  assign n22773 = n22772 ^ n19585 ^ n1000 ;
  assign n22774 = n22773 ^ n17268 ^ 1'b0 ;
  assign n22775 = n1309 & ~n22774 ;
  assign n22776 = n11712 ^ n6521 ^ n3462 ;
  assign n22777 = n14843 ^ n13632 ^ n5116 ;
  assign n22778 = n22777 ^ n15154 ^ n13743 ;
  assign n22779 = n14436 ^ n4442 ^ 1'b0 ;
  assign n22780 = n16428 & ~n22779 ;
  assign n22781 = ( n8473 & n11237 ) | ( n8473 & ~n16959 ) | ( n11237 & ~n16959 ) ;
  assign n22782 = ( ~n9174 & n22780 ) | ( ~n9174 & n22781 ) | ( n22780 & n22781 ) ;
  assign n22783 = ( ~n13009 & n15581 ) | ( ~n13009 & n17482 ) | ( n15581 & n17482 ) ;
  assign n22784 = n22783 ^ n15792 ^ n11633 ;
  assign n22785 = n15477 ^ n9986 ^ n7088 ;
  assign n22786 = ( x0 & ~n8142 ) | ( x0 & n12472 ) | ( ~n8142 & n12472 ) ;
  assign n22787 = n22785 | n22786 ;
  assign n22788 = n12344 ^ n7468 ^ n5849 ;
  assign n22789 = ( n1248 & n7613 ) | ( n1248 & ~n13352 ) | ( n7613 & ~n13352 ) ;
  assign n22790 = n7365 ^ n5855 ^ n5271 ;
  assign n22791 = n22790 ^ n2055 ^ 1'b0 ;
  assign n22792 = ( n12102 & n22789 ) | ( n12102 & n22791 ) | ( n22789 & n22791 ) ;
  assign n22793 = n22788 & n22792 ;
  assign n22794 = n14704 ^ n3962 ^ n2784 ;
  assign n22795 = n22794 ^ n18962 ^ n3232 ;
  assign n22803 = n9585 & ~n15818 ;
  assign n22800 = n14501 ^ n4945 ^ n3065 ;
  assign n22799 = ( n6515 & ~n8207 ) | ( n6515 & n8376 ) | ( ~n8207 & n8376 ) ;
  assign n22801 = n22800 ^ n22799 ^ n5462 ;
  assign n22797 = n19313 ^ n16068 ^ n4145 ;
  assign n22796 = ( ~n1133 & n11342 ) | ( ~n1133 & n18974 ) | ( n11342 & n18974 ) ;
  assign n22798 = n22797 ^ n22796 ^ n2744 ;
  assign n22802 = n22801 ^ n22798 ^ n10815 ;
  assign n22804 = n22803 ^ n22802 ^ n11468 ;
  assign n22805 = n9942 ^ n499 ^ x120 ;
  assign n22806 = n22805 ^ n12007 ^ n2217 ;
  assign n22807 = n22806 ^ n21983 ^ n14843 ;
  assign n22808 = ( n1541 & n16049 ) | ( n1541 & n20816 ) | ( n16049 & n20816 ) ;
  assign n22809 = ( n762 & ~n2140 ) | ( n762 & n13260 ) | ( ~n2140 & n13260 ) ;
  assign n22810 = ( ~n13461 & n22808 ) | ( ~n13461 & n22809 ) | ( n22808 & n22809 ) ;
  assign n22811 = n14459 ^ n13567 ^ n4989 ;
  assign n22812 = ( n1395 & n2173 ) | ( n1395 & ~n9867 ) | ( n2173 & ~n9867 ) ;
  assign n22813 = ( n18038 & n21541 ) | ( n18038 & ~n22812 ) | ( n21541 & ~n22812 ) ;
  assign n22814 = ( n4923 & n17571 ) | ( n4923 & n22813 ) | ( n17571 & n22813 ) ;
  assign n22815 = n22814 ^ n19149 ^ n15197 ;
  assign n22816 = n15394 ^ n6008 ^ n3541 ;
  assign n22817 = n8469 ^ n5736 ^ n563 ;
  assign n22818 = ( n959 & ~n6232 ) | ( n959 & n16204 ) | ( ~n6232 & n16204 ) ;
  assign n22819 = ( n4740 & ~n22817 ) | ( n4740 & n22818 ) | ( ~n22817 & n22818 ) ;
  assign n22820 = ( ~n2751 & n22816 ) | ( ~n2751 & n22819 ) | ( n22816 & n22819 ) ;
  assign n22821 = n20916 ^ n14715 ^ n4229 ;
  assign n22822 = n21981 ^ n18066 ^ 1'b0 ;
  assign n22823 = x27 & ~n22822 ;
  assign n22824 = n12362 ^ n2097 ^ 1'b0 ;
  assign n22825 = ( n284 & n13697 ) | ( n284 & n22824 ) | ( n13697 & n22824 ) ;
  assign n22827 = ( n6068 & ~n7989 ) | ( n6068 & n9289 ) | ( ~n7989 & n9289 ) ;
  assign n22828 = ( ~n582 & n19921 ) | ( ~n582 & n22827 ) | ( n19921 & n22827 ) ;
  assign n22826 = ( x247 & n13907 ) | ( x247 & n16454 ) | ( n13907 & n16454 ) ;
  assign n22829 = n22828 ^ n22826 ^ n8716 ;
  assign n22830 = n3194 | n9524 ;
  assign n22831 = ( n3265 & n7228 ) | ( n3265 & ~n14612 ) | ( n7228 & ~n14612 ) ;
  assign n22832 = n13322 & n22831 ;
  assign n22833 = ~n22830 & n22832 ;
  assign n22834 = n9795 ^ n8084 ^ n4615 ;
  assign n22835 = ( ~n11744 & n22568 ) | ( ~n11744 & n22834 ) | ( n22568 & n22834 ) ;
  assign n22836 = ( n9721 & ~n10828 ) | ( n9721 & n22835 ) | ( ~n10828 & n22835 ) ;
  assign n22837 = ( n1879 & n2480 ) | ( n1879 & n6971 ) | ( n2480 & n6971 ) ;
  assign n22838 = ~n6723 & n22837 ;
  assign n22839 = n22838 ^ n20047 ^ n18686 ;
  assign n22840 = ~n6269 & n18397 ;
  assign n22841 = n13092 ^ n8269 ^ x40 ;
  assign n22842 = n22841 ^ n14076 ^ 1'b0 ;
  assign n22843 = ~n22840 & n22842 ;
  assign n22844 = n19181 ^ n6738 ^ n3390 ;
  assign n22845 = ( n2481 & n16933 ) | ( n2481 & n22844 ) | ( n16933 & n22844 ) ;
  assign n22846 = n4819 ^ n400 ^ 1'b0 ;
  assign n22847 = n3149 & ~n22846 ;
  assign n22848 = n12801 & n22847 ;
  assign n22849 = n9697 ^ n7482 ^ 1'b0 ;
  assign n22850 = n7032 | n22849 ;
  assign n22851 = n10880 & ~n22850 ;
  assign n22852 = n22851 ^ n12607 ^ 1'b0 ;
  assign n22853 = n22852 ^ n9986 ^ n9279 ;
  assign n22854 = ~n3240 & n20460 ;
  assign n22855 = ( n5680 & n7296 ) | ( n5680 & ~n11576 ) | ( n7296 & ~n11576 ) ;
  assign n22856 = n4471 & n6347 ;
  assign n22857 = n22856 ^ x5 ^ 1'b0 ;
  assign n22860 = n13386 ^ n12127 ^ n5235 ;
  assign n22861 = n22860 ^ n13337 ^ n10403 ;
  assign n22862 = n5621 | n14201 ;
  assign n22863 = n22861 | n22862 ;
  assign n22858 = n4033 ^ n2333 ^ 1'b0 ;
  assign n22859 = ~n6664 & n22858 ;
  assign n22864 = n22863 ^ n22859 ^ n17363 ;
  assign n22865 = ~n22235 & n22864 ;
  assign n22866 = ~n4577 & n11963 ;
  assign n22867 = n11625 & n22866 ;
  assign n22868 = n3225 | n22867 ;
  assign n22869 = n22868 ^ n15065 ^ n13240 ;
  assign n22870 = n22869 ^ n9143 ^ n8222 ;
  assign n22871 = n19692 ^ n15000 ^ n4406 ;
  assign n22872 = ( ~n20770 & n22870 ) | ( ~n20770 & n22871 ) | ( n22870 & n22871 ) ;
  assign n22873 = n18018 ^ n10073 ^ n7118 ;
  assign n22874 = n21687 ^ n21119 ^ n4735 ;
  assign n22875 = n19294 | n22874 ;
  assign n22876 = n22875 ^ n8394 ^ 1'b0 ;
  assign n22877 = ~n11671 & n22876 ;
  assign n22878 = n22877 ^ n11231 ^ 1'b0 ;
  assign n22879 = ( n3277 & n6665 ) | ( n3277 & ~n15463 ) | ( n6665 & ~n15463 ) ;
  assign n22880 = n17375 ^ n10286 ^ n10165 ;
  assign n22881 = ( n8743 & ~n16847 ) | ( n8743 & n22880 ) | ( ~n16847 & n22880 ) ;
  assign n22882 = n22881 ^ n8494 ^ 1'b0 ;
  assign n22888 = n14352 ^ n6497 ^ x45 ;
  assign n22886 = n4210 ^ n3798 ^ 1'b0 ;
  assign n22887 = n7499 & n22886 ;
  assign n22883 = n2881 ^ x70 ^ x44 ;
  assign n22884 = ( n3139 & n4839 ) | ( n3139 & ~n22883 ) | ( n4839 & ~n22883 ) ;
  assign n22885 = ( ~n5532 & n21537 ) | ( ~n5532 & n22884 ) | ( n21537 & n22884 ) ;
  assign n22889 = n22888 ^ n22887 ^ n22885 ;
  assign n22890 = n22275 ^ n7142 ^ n4245 ;
  assign n22891 = n17496 ^ n8413 ^ n8032 ;
  assign n22892 = ( n10986 & ~n14397 ) | ( n10986 & n22891 ) | ( ~n14397 & n22891 ) ;
  assign n22893 = n21961 ^ n13348 ^ n10547 ;
  assign n22894 = ( n4953 & n5330 ) | ( n4953 & ~n18313 ) | ( n5330 & ~n18313 ) ;
  assign n22895 = ( n1502 & n16335 ) | ( n1502 & n22548 ) | ( n16335 & n22548 ) ;
  assign n22896 = n22895 ^ n11538 ^ n3806 ;
  assign n22897 = ( n7556 & n11437 ) | ( n7556 & n22896 ) | ( n11437 & n22896 ) ;
  assign n22898 = ( n3491 & n5070 ) | ( n3491 & n8855 ) | ( n5070 & n8855 ) ;
  assign n22899 = n22898 ^ n15638 ^ 1'b0 ;
  assign n22900 = n6648 & n22899 ;
  assign n22901 = ( n890 & n10195 ) | ( n890 & n12929 ) | ( n10195 & n12929 ) ;
  assign n22902 = ( n17845 & n18012 ) | ( n17845 & ~n21963 ) | ( n18012 & ~n21963 ) ;
  assign n22903 = ( ~n6621 & n13726 ) | ( ~n6621 & n22902 ) | ( n13726 & n22902 ) ;
  assign n22904 = ( n10941 & ~n22901 ) | ( n10941 & n22903 ) | ( ~n22901 & n22903 ) ;
  assign n22905 = ( n7892 & n22900 ) | ( n7892 & n22904 ) | ( n22900 & n22904 ) ;
  assign n22906 = n16404 ^ n14367 ^ n12787 ;
  assign n22907 = ( n6249 & ~n11385 ) | ( n6249 & n18563 ) | ( ~n11385 & n18563 ) ;
  assign n22908 = n22907 ^ n645 ^ 1'b0 ;
  assign n22910 = n5656 ^ n256 ^ 1'b0 ;
  assign n22911 = n1884 | n22910 ;
  assign n22909 = n11159 ^ n9410 ^ n7733 ;
  assign n22912 = n22911 ^ n22909 ^ n13807 ;
  assign n22913 = ( ~n15894 & n22908 ) | ( ~n15894 & n22912 ) | ( n22908 & n22912 ) ;
  assign n22914 = n6783 ^ n5580 ^ 1'b0 ;
  assign n22915 = ( n9033 & ~n22798 ) | ( n9033 & n22914 ) | ( ~n22798 & n22914 ) ;
  assign n22916 = n22915 ^ n18506 ^ n7494 ;
  assign n22917 = ( n3518 & ~n14198 ) | ( n3518 & n21474 ) | ( ~n14198 & n21474 ) ;
  assign n22918 = n5849 & ~n11674 ;
  assign n22919 = n22918 ^ n7535 ^ 1'b0 ;
  assign n22920 = n17539 ^ n8413 ^ n4984 ;
  assign n22921 = n22920 ^ n6614 ^ 1'b0 ;
  assign n22922 = ( n22917 & n22919 ) | ( n22917 & ~n22921 ) | ( n22919 & ~n22921 ) ;
  assign n22923 = n14985 ^ n9109 ^ n3326 ;
  assign n22924 = n13882 ^ n1828 ^ 1'b0 ;
  assign n22925 = ( ~n5004 & n17916 ) | ( ~n5004 & n22924 ) | ( n17916 & n22924 ) ;
  assign n22926 = ~n3066 & n7621 ;
  assign n22928 = n20826 ^ n14784 ^ n6136 ;
  assign n22927 = ( n7635 & n11198 ) | ( n7635 & ~n20547 ) | ( n11198 & ~n20547 ) ;
  assign n22929 = n22928 ^ n22927 ^ n15826 ;
  assign n22930 = n22929 ^ n15063 ^ n607 ;
  assign n22932 = ( n1828 & ~n7682 ) | ( n1828 & n21752 ) | ( ~n7682 & n21752 ) ;
  assign n22931 = n12665 ^ n4490 ^ x111 ;
  assign n22933 = n22932 ^ n22931 ^ 1'b0 ;
  assign n22934 = ~n22930 & n22933 ;
  assign n22935 = n1705 & ~n3051 ;
  assign n22936 = n10829 & n22935 ;
  assign n22937 = ( x202 & n4883 ) | ( x202 & n17531 ) | ( n4883 & n17531 ) ;
  assign n22938 = ( ~n3734 & n22936 ) | ( ~n3734 & n22937 ) | ( n22936 & n22937 ) ;
  assign n22939 = ( n7117 & n9357 ) | ( n7117 & n17612 ) | ( n9357 & n17612 ) ;
  assign n22940 = n22939 ^ n14072 ^ n11348 ;
  assign n22941 = ( n859 & ~n3541 ) | ( n859 & n22940 ) | ( ~n3541 & n22940 ) ;
  assign n22942 = n20940 ^ n715 ^ 1'b0 ;
  assign n22943 = n22941 | n22942 ;
  assign n22944 = n22943 ^ n2551 ^ n2183 ;
  assign n22945 = n19074 ^ n7547 ^ n1191 ;
  assign n22946 = ( n4135 & n18707 ) | ( n4135 & ~n22945 ) | ( n18707 & ~n22945 ) ;
  assign n22947 = n19306 ^ n15747 ^ n15247 ;
  assign n22948 = ( ~n2478 & n12892 ) | ( ~n2478 & n19436 ) | ( n12892 & n19436 ) ;
  assign n22949 = n16742 ^ n16297 ^ n6167 ;
  assign n22950 = ( ~x254 & n5931 ) | ( ~x254 & n6093 ) | ( n5931 & n6093 ) ;
  assign n22951 = n2491 & ~n20223 ;
  assign n22952 = n22951 ^ n4794 ^ 1'b0 ;
  assign n22953 = ( n8067 & ~n22950 ) | ( n8067 & n22952 ) | ( ~n22950 & n22952 ) ;
  assign n22954 = ( ~n3417 & n5595 ) | ( ~n3417 & n7823 ) | ( n5595 & n7823 ) ;
  assign n22955 = ( ~n5764 & n6023 ) | ( ~n5764 & n22954 ) | ( n6023 & n22954 ) ;
  assign n22956 = ( n9854 & ~n10069 ) | ( n9854 & n22955 ) | ( ~n10069 & n22955 ) ;
  assign n22957 = n22953 & ~n22956 ;
  assign n22958 = ( n12936 & ~n22273 ) | ( n12936 & n22957 ) | ( ~n22273 & n22957 ) ;
  assign n22959 = ( ~n2962 & n7037 ) | ( ~n2962 & n9665 ) | ( n7037 & n9665 ) ;
  assign n22960 = n16595 ^ n15969 ^ 1'b0 ;
  assign n22961 = n3763 | n22960 ;
  assign n22962 = n11808 | n22961 ;
  assign n22964 = n12167 ^ n2093 ^ 1'b0 ;
  assign n22965 = n2773 | n9647 ;
  assign n22966 = ( ~n7870 & n22964 ) | ( ~n7870 & n22965 ) | ( n22964 & n22965 ) ;
  assign n22967 = n17724 & n22966 ;
  assign n22968 = n22967 ^ n5130 ^ 1'b0 ;
  assign n22963 = ( n5753 & n13192 ) | ( n5753 & n14098 ) | ( n13192 & n14098 ) ;
  assign n22969 = n22968 ^ n22963 ^ n8860 ;
  assign n22970 = ( n3097 & n4936 ) | ( n3097 & n22969 ) | ( n4936 & n22969 ) ;
  assign n22971 = n18375 ^ n8015 ^ n4768 ;
  assign n22972 = n22971 ^ n13894 ^ n8337 ;
  assign n22974 = ~x166 & n3266 ;
  assign n22973 = n17667 ^ n4844 ^ n297 ;
  assign n22975 = n22974 ^ n22973 ^ n21780 ;
  assign n22976 = ( n18618 & ~n22972 ) | ( n18618 & n22975 ) | ( ~n22972 & n22975 ) ;
  assign n22978 = n2374 | n8679 ;
  assign n22977 = n13110 ^ n8811 ^ 1'b0 ;
  assign n22979 = n22978 ^ n22977 ^ n10119 ;
  assign n22980 = n22042 ^ n808 ^ 1'b0 ;
  assign n22981 = ( n3027 & ~n5328 ) | ( n3027 & n22980 ) | ( ~n5328 & n22980 ) ;
  assign n22982 = ( n14936 & ~n22979 ) | ( n14936 & n22981 ) | ( ~n22979 & n22981 ) ;
  assign n22983 = ~n7207 & n16742 ;
  assign n22984 = n20252 & n22983 ;
  assign n22988 = n21630 & ~n22868 ;
  assign n22989 = ( n3938 & n5961 ) | ( n3938 & ~n22988 ) | ( n5961 & ~n22988 ) ;
  assign n22985 = ( ~n1276 & n4129 ) | ( ~n1276 & n5374 ) | ( n4129 & n5374 ) ;
  assign n22986 = n5763 & ~n22985 ;
  assign n22987 = n22986 ^ n2801 ^ 1'b0 ;
  assign n22990 = n22989 ^ n22987 ^ 1'b0 ;
  assign n22991 = n11709 | n14786 ;
  assign n22992 = ( n8541 & n10056 ) | ( n8541 & n15815 ) | ( n10056 & n15815 ) ;
  assign n22993 = ( ~n18948 & n21640 ) | ( ~n18948 & n22992 ) | ( n21640 & n22992 ) ;
  assign n22994 = n22993 ^ n13679 ^ n10380 ;
  assign n22995 = n22991 & ~n22994 ;
  assign n23004 = n7588 ^ n4347 ^ n3712 ;
  assign n23005 = ( n8603 & ~n14296 ) | ( n8603 & n23004 ) | ( ~n14296 & n23004 ) ;
  assign n23006 = ( ~n5057 & n8228 ) | ( ~n5057 & n23005 ) | ( n8228 & n23005 ) ;
  assign n22999 = n8333 ^ n7178 ^ n5434 ;
  assign n23000 = n15811 ^ n9937 ^ n3912 ;
  assign n23001 = n23000 ^ n15574 ^ n7948 ;
  assign n23002 = n23001 ^ n7323 ^ n899 ;
  assign n23003 = ( ~n1735 & n22999 ) | ( ~n1735 & n23002 ) | ( n22999 & n23002 ) ;
  assign n23007 = n23006 ^ n23003 ^ n18948 ;
  assign n22997 = ( n9621 & ~n13999 ) | ( n9621 & n22504 ) | ( ~n13999 & n22504 ) ;
  assign n22996 = n19917 ^ n11958 ^ n4570 ;
  assign n22998 = n22997 ^ n22996 ^ n16770 ;
  assign n23008 = n23007 ^ n22998 ^ n17567 ;
  assign n23010 = n14913 ^ n3683 ^ n1200 ;
  assign n23009 = n2578 & n10419 ;
  assign n23011 = n23010 ^ n23009 ^ n967 ;
  assign n23012 = ( n631 & n15197 ) | ( n631 & n20343 ) | ( n15197 & n20343 ) ;
  assign n23013 = ( n2469 & ~n3451 ) | ( n2469 & n6173 ) | ( ~n3451 & n6173 ) ;
  assign n23014 = n19846 ^ n18707 ^ n1109 ;
  assign n23015 = n23014 ^ n5192 ^ n1513 ;
  assign n23016 = n16898 ^ n12837 ^ n8059 ;
  assign n23017 = ( n7648 & n8191 ) | ( n7648 & n17837 ) | ( n8191 & n17837 ) ;
  assign n23018 = n23017 ^ n20814 ^ n5474 ;
  assign n23019 = n1866 & ~n6768 ;
  assign n23020 = n23019 ^ n13817 ^ n11982 ;
  assign n23021 = ( n2324 & n5687 ) | ( n2324 & n18531 ) | ( n5687 & n18531 ) ;
  assign n23022 = ( n22121 & n23020 ) | ( n22121 & n23021 ) | ( n23020 & n23021 ) ;
  assign n23023 = n23022 ^ n20437 ^ n510 ;
  assign n23024 = n23018 | n23023 ;
  assign n23025 = n23016 | n23024 ;
  assign n23026 = ( n12524 & ~n13763 ) | ( n12524 & n15049 ) | ( ~n13763 & n15049 ) ;
  assign n23027 = ( n10874 & ~n14491 ) | ( n10874 & n23026 ) | ( ~n14491 & n23026 ) ;
  assign n23028 = n19272 ^ n13742 ^ n1758 ;
  assign n23029 = ( ~n1000 & n3114 ) | ( ~n1000 & n23028 ) | ( n3114 & n23028 ) ;
  assign n23030 = n9459 ^ n7288 ^ n3098 ;
  assign n23031 = n10838 & ~n23030 ;
  assign n23032 = n23031 ^ n4968 ^ 1'b0 ;
  assign n23033 = n5803 ^ n5168 ^ 1'b0 ;
  assign n23034 = n23032 & n23033 ;
  assign n23035 = n20666 ^ n13748 ^ n2341 ;
  assign n23036 = ( ~n18825 & n19863 ) | ( ~n18825 & n23035 ) | ( n19863 & n23035 ) ;
  assign n23037 = ( n515 & n5491 ) | ( n515 & n18117 ) | ( n5491 & n18117 ) ;
  assign n23038 = n23037 ^ n17732 ^ n4422 ;
  assign n23039 = n14615 ^ n6976 ^ n1881 ;
  assign n23040 = n15478 ^ n4484 ^ 1'b0 ;
  assign n23041 = ~n23039 & n23040 ;
  assign n23042 = n6553 ^ n2473 ^ x223 ;
  assign n23043 = n17236 ^ n9477 ^ n1821 ;
  assign n23044 = ( n12329 & ~n23042 ) | ( n12329 & n23043 ) | ( ~n23042 & n23043 ) ;
  assign n23046 = ( n575 & n3213 ) | ( n575 & n8665 ) | ( n3213 & n8665 ) ;
  assign n23045 = ( n7698 & ~n14968 ) | ( n7698 & n20722 ) | ( ~n14968 & n20722 ) ;
  assign n23047 = n23046 ^ n23045 ^ n7599 ;
  assign n23048 = ( n5840 & ~n20633 ) | ( n5840 & n23047 ) | ( ~n20633 & n23047 ) ;
  assign n23049 = ( n15585 & ~n19975 ) | ( n15585 & n23048 ) | ( ~n19975 & n23048 ) ;
  assign n23050 = ( n885 & ~n23044 ) | ( n885 & n23049 ) | ( ~n23044 & n23049 ) ;
  assign n23060 = n18260 ^ n6293 ^ n2282 ;
  assign n23051 = ( n6509 & n8937 ) | ( n6509 & n20823 ) | ( n8937 & n20823 ) ;
  assign n23052 = ( n9909 & ~n11899 ) | ( n9909 & n16290 ) | ( ~n11899 & n16290 ) ;
  assign n23053 = ( n12496 & n17253 ) | ( n12496 & ~n19506 ) | ( n17253 & ~n19506 ) ;
  assign n23054 = n6468 ^ n6218 ^ n6041 ;
  assign n23055 = n23054 ^ n2255 ^ 1'b0 ;
  assign n23056 = n20478 & ~n23055 ;
  assign n23057 = n23056 ^ n15651 ^ 1'b0 ;
  assign n23058 = ( n23052 & n23053 ) | ( n23052 & ~n23057 ) | ( n23053 & ~n23057 ) ;
  assign n23059 = ( n10062 & n23051 ) | ( n10062 & n23058 ) | ( n23051 & n23058 ) ;
  assign n23061 = n23060 ^ n23059 ^ n7481 ;
  assign n23062 = ~n7375 & n15064 ;
  assign n23063 = ~n23061 & n23062 ;
  assign n23064 = ( n6600 & n7293 ) | ( n6600 & n12519 ) | ( n7293 & n12519 ) ;
  assign n23065 = ( x246 & n7602 ) | ( x246 & n8549 ) | ( n7602 & n8549 ) ;
  assign n23066 = n23065 ^ n22425 ^ n8256 ;
  assign n23067 = ( ~n15397 & n23064 ) | ( ~n15397 & n23066 ) | ( n23064 & n23066 ) ;
  assign n23068 = n1870 | n6029 ;
  assign n23069 = n6918 & ~n23068 ;
  assign n23070 = n23069 ^ n4144 ^ n2661 ;
  assign n23071 = ( n9889 & n20575 ) | ( n9889 & n22588 ) | ( n20575 & n22588 ) ;
  assign n23072 = ( n5624 & n23070 ) | ( n5624 & n23071 ) | ( n23070 & n23071 ) ;
  assign n23089 = ( n966 & n5155 ) | ( n966 & n7672 ) | ( n5155 & n7672 ) ;
  assign n23090 = ( n3081 & ~n4510 ) | ( n3081 & n23089 ) | ( ~n4510 & n23089 ) ;
  assign n23091 = n23090 ^ n568 ^ n379 ;
  assign n23092 = ~n21222 & n23091 ;
  assign n23093 = n23092 ^ n8741 ^ 1'b0 ;
  assign n23083 = ( ~n318 & n6595 ) | ( ~n318 & n17265 ) | ( n6595 & n17265 ) ;
  assign n23084 = n20743 ^ n1371 ^ 1'b0 ;
  assign n23085 = n19166 & n23084 ;
  assign n23086 = n23085 ^ n10927 ^ 1'b0 ;
  assign n23087 = n23086 ^ n13384 ^ n9869 ;
  assign n23088 = ( n17571 & n23083 ) | ( n17571 & n23087 ) | ( n23083 & n23087 ) ;
  assign n23073 = ( n3888 & ~n8118 ) | ( n3888 & n17180 ) | ( ~n8118 & n17180 ) ;
  assign n23074 = ~n1059 & n5021 ;
  assign n23075 = ( n17301 & n23073 ) | ( n17301 & ~n23074 ) | ( n23073 & ~n23074 ) ;
  assign n23076 = n23075 ^ n18106 ^ n1224 ;
  assign n23077 = n1588 & n5107 ;
  assign n23078 = n2087 & n23077 ;
  assign n23079 = ~n8191 & n23078 ;
  assign n23080 = ( ~n1276 & n5346 ) | ( ~n1276 & n23079 ) | ( n5346 & n23079 ) ;
  assign n23081 = n23080 ^ n20663 ^ n7078 ;
  assign n23082 = ( ~n18321 & n23076 ) | ( ~n18321 & n23081 ) | ( n23076 & n23081 ) ;
  assign n23094 = n23093 ^ n23088 ^ n23082 ;
  assign n23095 = ( n1210 & ~n6398 ) | ( n1210 & n7896 ) | ( ~n6398 & n7896 ) ;
  assign n23097 = ( n767 & ~n10044 ) | ( n767 & n19527 ) | ( ~n10044 & n19527 ) ;
  assign n23096 = ~n7296 & n12229 ;
  assign n23098 = n23097 ^ n23096 ^ 1'b0 ;
  assign n23099 = ( n6784 & n7936 ) | ( n6784 & n13599 ) | ( n7936 & n13599 ) ;
  assign n23100 = n10146 ^ n4374 ^ 1'b0 ;
  assign n23101 = ( ~n1136 & n4488 ) | ( ~n1136 & n23100 ) | ( n4488 & n23100 ) ;
  assign n23102 = ( n9833 & n17875 ) | ( n9833 & n23101 ) | ( n17875 & n23101 ) ;
  assign n23103 = ( ~n487 & n20459 ) | ( ~n487 & n23102 ) | ( n20459 & n23102 ) ;
  assign n23104 = ( ~n10838 & n23099 ) | ( ~n10838 & n23103 ) | ( n23099 & n23103 ) ;
  assign n23109 = n14152 ^ n11095 ^ n5852 ;
  assign n23107 = n11065 ^ n5968 ^ n3125 ;
  assign n23105 = n6876 ^ n3648 ^ 1'b0 ;
  assign n23106 = ~n5140 & n23105 ;
  assign n23108 = n23107 ^ n23106 ^ n2025 ;
  assign n23110 = n23109 ^ n23108 ^ n2857 ;
  assign n23111 = ( n4834 & n5822 ) | ( n4834 & n13717 ) | ( n5822 & n13717 ) ;
  assign n23112 = n18741 ^ n9101 ^ n8615 ;
  assign n23113 = ( n10238 & ~n12317 ) | ( n10238 & n23112 ) | ( ~n12317 & n23112 ) ;
  assign n23114 = n16006 & ~n23113 ;
  assign n23115 = n20744 ^ n18336 ^ n7981 ;
  assign n23116 = ( n7446 & ~n21541 ) | ( n7446 & n23115 ) | ( ~n21541 & n23115 ) ;
  assign n23117 = n21630 ^ n11216 ^ n2669 ;
  assign n23118 = n23117 ^ n11428 ^ n2552 ;
  assign n23119 = ( n8693 & n13627 ) | ( n8693 & ~n23118 ) | ( n13627 & ~n23118 ) ;
  assign n23120 = ( n6101 & n15673 ) | ( n6101 & ~n20339 ) | ( n15673 & ~n20339 ) ;
  assign n23121 = ( n3856 & n12331 ) | ( n3856 & ~n19962 ) | ( n12331 & ~n19962 ) ;
  assign n23122 = ( ~n8592 & n21531 ) | ( ~n8592 & n23121 ) | ( n21531 & n23121 ) ;
  assign n23123 = n23122 ^ n19831 ^ 1'b0 ;
  assign n23124 = n6848 ^ n5078 ^ 1'b0 ;
  assign n23125 = n8158 ^ n1656 ^ 1'b0 ;
  assign n23126 = n23124 & n23125 ;
  assign n23127 = n13048 ^ n7610 ^ 1'b0 ;
  assign n23128 = ~n17204 & n23127 ;
  assign n23129 = ( n1479 & n23126 ) | ( n1479 & n23128 ) | ( n23126 & n23128 ) ;
  assign n23130 = ( n6502 & ~n9044 ) | ( n6502 & n23129 ) | ( ~n9044 & n23129 ) ;
  assign n23131 = ( ~n18224 & n20481 ) | ( ~n18224 & n23130 ) | ( n20481 & n23130 ) ;
  assign n23132 = ( n5240 & n10367 ) | ( n5240 & ~n11468 ) | ( n10367 & ~n11468 ) ;
  assign n23133 = ~n9171 & n23132 ;
  assign n23134 = n23133 ^ n20715 ^ 1'b0 ;
  assign n23135 = n23134 ^ n18107 ^ 1'b0 ;
  assign n23136 = n8065 | n23135 ;
  assign n23137 = ( n2153 & n5814 ) | ( n2153 & n16814 ) | ( n5814 & n16814 ) ;
  assign n23138 = ( n3160 & n9067 ) | ( n3160 & n9920 ) | ( n9067 & n9920 ) ;
  assign n23139 = n23138 ^ n2747 ^ 1'b0 ;
  assign n23140 = n18259 & n23139 ;
  assign n23141 = ( n5938 & ~n23137 ) | ( n5938 & n23140 ) | ( ~n23137 & n23140 ) ;
  assign n23142 = ( ~n2537 & n15602 ) | ( ~n2537 & n22758 ) | ( n15602 & n22758 ) ;
  assign n23143 = n6289 ^ n4088 ^ n688 ;
  assign n23144 = ( n5490 & n16418 ) | ( n5490 & n23143 ) | ( n16418 & n23143 ) ;
  assign n23145 = n23144 ^ n17569 ^ n588 ;
  assign n23146 = n23145 ^ n11699 ^ n388 ;
  assign n23147 = x215 | n12507 ;
  assign n23148 = n22246 ^ n10515 ^ n7443 ;
  assign n23149 = n16614 ^ n1490 ^ 1'b0 ;
  assign n23150 = ( n8688 & n15034 ) | ( n8688 & ~n23149 ) | ( n15034 & ~n23149 ) ;
  assign n23151 = n1053 & ~n21580 ;
  assign n23152 = ( n12407 & ~n18442 ) | ( n12407 & n19445 ) | ( ~n18442 & n19445 ) ;
  assign n23153 = ~n6755 & n9726 ;
  assign n23154 = n23153 ^ n2625 ^ 1'b0 ;
  assign n23155 = ( n4329 & n7250 ) | ( n4329 & ~n23154 ) | ( n7250 & ~n23154 ) ;
  assign n23156 = n10784 ^ n8489 ^ 1'b0 ;
  assign n23157 = n23156 ^ n15152 ^ n410 ;
  assign n23158 = ( ~n4847 & n14091 ) | ( ~n4847 & n14712 ) | ( n14091 & n14712 ) ;
  assign n23159 = ( x110 & ~n2629 ) | ( x110 & n17077 ) | ( ~n2629 & n17077 ) ;
  assign n23160 = n23159 ^ n10306 ^ n3690 ;
  assign n23161 = ( ~n438 & n923 ) | ( ~n438 & n23160 ) | ( n923 & n23160 ) ;
  assign n23162 = ( n13884 & ~n15019 ) | ( n13884 & n23161 ) | ( ~n15019 & n23161 ) ;
  assign n23163 = n10670 | n14819 ;
  assign n23164 = n21728 | n23163 ;
  assign n23165 = ( n5877 & ~n19977 ) | ( n5877 & n23164 ) | ( ~n19977 & n23164 ) ;
  assign n23166 = n20293 ^ n19987 ^ n7674 ;
  assign n23167 = n21131 ^ n18834 ^ n11101 ;
  assign n23168 = ( n7607 & ~n23166 ) | ( n7607 & n23167 ) | ( ~n23166 & n23167 ) ;
  assign n23169 = ( n4787 & n6008 ) | ( n4787 & n17350 ) | ( n6008 & n17350 ) ;
  assign n23170 = ( n2853 & ~n4329 ) | ( n2853 & n7891 ) | ( ~n4329 & n7891 ) ;
  assign n23171 = ( n23168 & ~n23169 ) | ( n23168 & n23170 ) | ( ~n23169 & n23170 ) ;
  assign n23179 = n12514 ^ n1665 ^ n1159 ;
  assign n23176 = n5233 ^ n2997 ^ n840 ;
  assign n23173 = n3729 ^ n1404 ^ n904 ;
  assign n23172 = n1541 & ~n4862 ;
  assign n23174 = n23173 ^ n23172 ^ 1'b0 ;
  assign n23175 = n23174 ^ n8941 ^ n5280 ;
  assign n23177 = n23176 ^ n23175 ^ 1'b0 ;
  assign n23178 = n5414 | n23177 ;
  assign n23180 = n23179 ^ n23178 ^ n3174 ;
  assign n23181 = n13244 ^ n5040 ^ 1'b0 ;
  assign n23182 = n15316 ^ n8782 ^ n8550 ;
  assign n23183 = n14519 ^ n4067 ^ n2862 ;
  assign n23187 = n8237 ^ n6915 ^ n265 ;
  assign n23188 = ( x89 & n4700 ) | ( x89 & n23187 ) | ( n4700 & n23187 ) ;
  assign n23184 = n6845 ^ n6387 ^ n4871 ;
  assign n23185 = ( n6586 & n10072 ) | ( n6586 & n23184 ) | ( n10072 & n23184 ) ;
  assign n23186 = ( n11611 & n14147 ) | ( n11611 & n23185 ) | ( n14147 & n23185 ) ;
  assign n23189 = n23188 ^ n23186 ^ 1'b0 ;
  assign n23190 = n23183 & ~n23189 ;
  assign n23191 = ( ~n23181 & n23182 ) | ( ~n23181 & n23190 ) | ( n23182 & n23190 ) ;
  assign n23192 = ( ~n13314 & n23180 ) | ( ~n13314 & n23191 ) | ( n23180 & n23191 ) ;
  assign n23193 = n23192 ^ n21844 ^ n2362 ;
  assign n23196 = n8590 ^ n3677 ^ n760 ;
  assign n23197 = n23196 ^ n19655 ^ n7320 ;
  assign n23198 = ( x195 & ~n8020 ) | ( x195 & n23197 ) | ( ~n8020 & n23197 ) ;
  assign n23194 = ( n2697 & n4863 ) | ( n2697 & ~n13845 ) | ( n4863 & ~n13845 ) ;
  assign n23195 = n23194 ^ n20263 ^ x183 ;
  assign n23199 = n23198 ^ n23195 ^ n16184 ;
  assign n23200 = n8994 ^ n3305 ^ 1'b0 ;
  assign n23201 = n12474 ^ n7764 ^ n2013 ;
  assign n23202 = n23201 ^ n11120 ^ n3914 ;
  assign n23203 = n9455 & n19198 ;
  assign n23204 = ~n23202 & n23203 ;
  assign n23205 = ~n23200 & n23204 ;
  assign n23206 = ( ~n4460 & n4734 ) | ( ~n4460 & n20280 ) | ( n4734 & n20280 ) ;
  assign n23207 = ( n5027 & ~n17611 ) | ( n5027 & n18305 ) | ( ~n17611 & n18305 ) ;
  assign n23208 = ( n14927 & n23206 ) | ( n14927 & ~n23207 ) | ( n23206 & ~n23207 ) ;
  assign n23209 = n12525 ^ n7363 ^ n6276 ;
  assign n23210 = n23209 ^ n9541 ^ n7911 ;
  assign n23211 = n19656 ^ n13867 ^ n10944 ;
  assign n23216 = n20272 ^ n16980 ^ n7170 ;
  assign n23214 = n6170 ^ n3328 ^ x219 ;
  assign n23212 = n5621 ^ n430 ^ n308 ;
  assign n23213 = ( n12429 & n23070 ) | ( n12429 & ~n23212 ) | ( n23070 & ~n23212 ) ;
  assign n23215 = n23214 ^ n23213 ^ 1'b0 ;
  assign n23217 = n23216 ^ n23215 ^ n2804 ;
  assign n23218 = n6997 ^ n5438 ^ n2682 ;
  assign n23219 = ( n5281 & n21022 ) | ( n5281 & ~n23218 ) | ( n21022 & ~n23218 ) ;
  assign n23220 = n21072 ^ n13317 ^ n8268 ;
  assign n23221 = ( n1028 & n23219 ) | ( n1028 & n23220 ) | ( n23219 & n23220 ) ;
  assign n23222 = n6902 & n7320 ;
  assign n23223 = n23222 ^ n7833 ^ 1'b0 ;
  assign n23224 = n3802 | n23223 ;
  assign n23225 = n4427 & ~n23224 ;
  assign n23226 = n13274 ^ n10554 ^ n2835 ;
  assign n23227 = n4481 & n23226 ;
  assign n23228 = n23225 & n23227 ;
  assign n23229 = n23228 ^ n22554 ^ n14699 ;
  assign n23230 = ( ~n275 & n12267 ) | ( ~n275 & n19003 ) | ( n12267 & n19003 ) ;
  assign n23231 = ( n5474 & ~n11923 ) | ( n5474 & n23230 ) | ( ~n11923 & n23230 ) ;
  assign n23232 = n23231 ^ n2012 ^ n1528 ;
  assign n23233 = ( n7020 & n11549 ) | ( n7020 & n23232 ) | ( n11549 & n23232 ) ;
  assign n23234 = n5794 ^ n3027 ^ n982 ;
  assign n23235 = ( n6560 & ~n9080 ) | ( n6560 & n23234 ) | ( ~n9080 & n23234 ) ;
  assign n23237 = n18016 ^ n6886 ^ n485 ;
  assign n23238 = ~n4217 & n14235 ;
  assign n23239 = n23238 ^ n14356 ^ n6774 ;
  assign n23240 = ( n23107 & ~n23237 ) | ( n23107 & n23239 ) | ( ~n23237 & n23239 ) ;
  assign n23236 = n20818 ^ n5494 ^ n3862 ;
  assign n23241 = n23240 ^ n23236 ^ n18519 ;
  assign n23245 = n22063 ^ n8313 ^ n1361 ;
  assign n23242 = ( n4506 & n11057 ) | ( n4506 & ~n21986 ) | ( n11057 & ~n21986 ) ;
  assign n23243 = n23242 ^ n10759 ^ n5944 ;
  assign n23244 = n17244 | n23243 ;
  assign n23246 = n23245 ^ n23244 ^ n20876 ;
  assign n23247 = n22723 ^ n21200 ^ n3694 ;
  assign n23248 = n1716 | n2686 ;
  assign n23249 = n23248 ^ n1297 ^ 1'b0 ;
  assign n23250 = ( n7206 & n8718 ) | ( n7206 & n23249 ) | ( n8718 & n23249 ) ;
  assign n23251 = n6091 ^ n2910 ^ n1727 ;
  assign n23252 = ( n10163 & n23250 ) | ( n10163 & n23251 ) | ( n23250 & n23251 ) ;
  assign n23253 = ( ~n13219 & n15310 ) | ( ~n13219 & n19238 ) | ( n15310 & n19238 ) ;
  assign n23254 = ( ~n4042 & n21326 ) | ( ~n4042 & n23253 ) | ( n21326 & n23253 ) ;
  assign n23255 = n2711 & ~n23254 ;
  assign n23256 = n605 & n23255 ;
  assign n23259 = ( n1009 & n4117 ) | ( n1009 & ~n8392 ) | ( n4117 & ~n8392 ) ;
  assign n23257 = n13734 | n16966 ;
  assign n23258 = n21474 & ~n23257 ;
  assign n23260 = n23259 ^ n23258 ^ n23161 ;
  assign n23261 = n9047 ^ n6392 ^ n5860 ;
  assign n23262 = n16993 ^ n13223 ^ n1354 ;
  assign n23263 = n21171 ^ n20162 ^ n12841 ;
  assign n23264 = n14513 ^ x83 ^ 1'b0 ;
  assign n23265 = n18448 ^ n3549 ^ n3499 ;
  assign n23266 = ( ~n23263 & n23264 ) | ( ~n23263 & n23265 ) | ( n23264 & n23265 ) ;
  assign n23271 = n17474 ^ n15050 ^ n3012 ;
  assign n23267 = n3250 & ~n3261 ;
  assign n23268 = n3217 & n23267 ;
  assign n23269 = n23268 ^ n12021 ^ 1'b0 ;
  assign n23270 = n9892 & n23269 ;
  assign n23272 = n23271 ^ n23270 ^ n9071 ;
  assign n23273 = ( n3700 & n3760 ) | ( n3700 & ~n4204 ) | ( n3760 & ~n4204 ) ;
  assign n23274 = ( n8103 & n11614 ) | ( n8103 & ~n23273 ) | ( n11614 & ~n23273 ) ;
  assign n23275 = ( n10056 & ~n19814 ) | ( n10056 & n23274 ) | ( ~n19814 & n23274 ) ;
  assign n23276 = ( n3317 & n13016 ) | ( n3317 & ~n13840 ) | ( n13016 & ~n13840 ) ;
  assign n23277 = ( ~n1242 & n18077 ) | ( ~n1242 & n23276 ) | ( n18077 & n23276 ) ;
  assign n23278 = n23277 ^ n17849 ^ n1296 ;
  assign n23279 = ( n1957 & n2968 ) | ( n1957 & n4745 ) | ( n2968 & n4745 ) ;
  assign n23280 = ( n11228 & n17802 ) | ( n11228 & ~n23279 ) | ( n17802 & ~n23279 ) ;
  assign n23281 = ( ~n10079 & n15852 ) | ( ~n10079 & n23280 ) | ( n15852 & n23280 ) ;
  assign n23282 = ( n801 & n4833 ) | ( n801 & ~n22914 ) | ( n4833 & ~n22914 ) ;
  assign n23283 = n23282 ^ n14687 ^ n2530 ;
  assign n23284 = n15468 ^ n6139 ^ n3309 ;
  assign n23285 = ( ~n3826 & n6957 ) | ( ~n3826 & n10407 ) | ( n6957 & n10407 ) ;
  assign n23286 = n3000 & n23285 ;
  assign n23287 = ( x247 & n7209 ) | ( x247 & n23286 ) | ( n7209 & n23286 ) ;
  assign n23288 = ( ~n13179 & n23284 ) | ( ~n13179 & n23287 ) | ( n23284 & n23287 ) ;
  assign n23289 = ( n14127 & n23283 ) | ( n14127 & n23288 ) | ( n23283 & n23288 ) ;
  assign n23290 = ( n3564 & ~n9799 ) | ( n3564 & n10816 ) | ( ~n9799 & n10816 ) ;
  assign n23291 = ( n9364 & ~n13133 ) | ( n9364 & n23276 ) | ( ~n13133 & n23276 ) ;
  assign n23292 = n13757 ^ n7390 ^ n493 ;
  assign n23293 = n4015 & n23292 ;
  assign n23294 = n23293 ^ n1418 ^ 1'b0 ;
  assign n23295 = ( n13312 & n23291 ) | ( n13312 & n23294 ) | ( n23291 & n23294 ) ;
  assign n23296 = n4736 & n15647 ;
  assign n23297 = ~n9160 & n23296 ;
  assign n23298 = ( n9577 & ~n23295 ) | ( n9577 & n23297 ) | ( ~n23295 & n23297 ) ;
  assign n23301 = n12322 ^ n3726 ^ 1'b0 ;
  assign n23302 = n23301 ^ n8122 ^ n5064 ;
  assign n23299 = n18390 ^ n6452 ^ 1'b0 ;
  assign n23300 = n10825 & ~n23299 ;
  assign n23303 = n23302 ^ n23300 ^ n11979 ;
  assign n23305 = n12218 ^ n5979 ^ n2570 ;
  assign n23304 = n6231 ^ n4989 ^ n4493 ;
  assign n23306 = n23305 ^ n23304 ^ n7055 ;
  assign n23307 = ( n10269 & n11708 ) | ( n10269 & ~n19219 ) | ( n11708 & ~n19219 ) ;
  assign n23308 = ~n4482 & n23307 ;
  assign n23309 = ~n6106 & n10364 ;
  assign n23310 = n23309 ^ n21755 ^ n11962 ;
  assign n23311 = ( n6594 & n17482 ) | ( n6594 & ~n23310 ) | ( n17482 & ~n23310 ) ;
  assign n23321 = n16460 ^ n4765 ^ n988 ;
  assign n23317 = n12733 ^ n1092 ^ 1'b0 ;
  assign n23318 = n7606 & ~n23317 ;
  assign n23319 = n23318 ^ n22649 ^ n16338 ;
  assign n23315 = ( n3407 & n11148 ) | ( n3407 & n12484 ) | ( n11148 & n12484 ) ;
  assign n23312 = n5502 ^ n507 ^ 1'b0 ;
  assign n23313 = n15125 & n23312 ;
  assign n23314 = ( n5074 & n14296 ) | ( n5074 & n23313 ) | ( n14296 & n23313 ) ;
  assign n23316 = n23315 ^ n23314 ^ n12471 ;
  assign n23320 = n23319 ^ n23316 ^ n5546 ;
  assign n23322 = n23321 ^ n23320 ^ x95 ;
  assign n23323 = n2893 & ~n6201 ;
  assign n23324 = n1002 & n23323 ;
  assign n23325 = n23324 ^ n10416 ^ n5970 ;
  assign n23326 = n12812 ^ n7137 ^ n1220 ;
  assign n23327 = n16030 ^ n6875 ^ n1696 ;
  assign n23328 = ( n5014 & n23326 ) | ( n5014 & n23327 ) | ( n23326 & n23327 ) ;
  assign n23329 = ( ~n3031 & n3547 ) | ( ~n3031 & n23328 ) | ( n3547 & n23328 ) ;
  assign n23330 = ~n20358 & n23329 ;
  assign n23331 = n23325 & n23330 ;
  assign n23332 = ~n4997 & n8385 ;
  assign n23333 = n8668 ^ n2509 ^ n1465 ;
  assign n23334 = ( ~n14844 & n17987 ) | ( ~n14844 & n23333 ) | ( n17987 & n23333 ) ;
  assign n23335 = ( n3469 & ~n14937 ) | ( n3469 & n23334 ) | ( ~n14937 & n23334 ) ;
  assign n23336 = n12038 ^ n10773 ^ n7655 ;
  assign n23337 = n20401 ^ n12556 ^ n4922 ;
  assign n23338 = ~n17660 & n23337 ;
  assign n23343 = n17231 ^ n16263 ^ n4616 ;
  assign n23344 = n3181 & ~n3451 ;
  assign n23345 = ( n10277 & ~n23343 ) | ( n10277 & n23344 ) | ( ~n23343 & n23344 ) ;
  assign n23341 = n17644 ^ n11483 ^ n1581 ;
  assign n23342 = n23341 ^ n294 ^ 1'b0 ;
  assign n23339 = n365 & n11879 ;
  assign n23340 = n16997 & n23339 ;
  assign n23346 = n23345 ^ n23342 ^ n23340 ;
  assign n23351 = ( n5522 & ~n12484 ) | ( n5522 & n16595 ) | ( ~n12484 & n16595 ) ;
  assign n23347 = ( x175 & n1959 ) | ( x175 & ~n3579 ) | ( n1959 & ~n3579 ) ;
  assign n23348 = ( n6428 & n18831 ) | ( n6428 & ~n23347 ) | ( n18831 & ~n23347 ) ;
  assign n23349 = ( ~n7997 & n9197 ) | ( ~n7997 & n23348 ) | ( n9197 & n23348 ) ;
  assign n23350 = n23349 ^ n13020 ^ 1'b0 ;
  assign n23352 = n23351 ^ n23350 ^ n4132 ;
  assign n23356 = n9519 ^ n4344 ^ n1150 ;
  assign n23357 = n7208 | n23356 ;
  assign n23358 = n23357 ^ n6186 ^ 1'b0 ;
  assign n23353 = ( ~n4714 & n16986 ) | ( ~n4714 & n21419 ) | ( n16986 & n21419 ) ;
  assign n23354 = n23353 ^ n15164 ^ 1'b0 ;
  assign n23355 = ~n10504 & n23354 ;
  assign n23359 = n23358 ^ n23355 ^ n13169 ;
  assign n23360 = n14829 ^ n11872 ^ x61 ;
  assign n23361 = n23360 ^ n22072 ^ n4969 ;
  assign n23362 = ( x55 & n19420 ) | ( x55 & ~n23361 ) | ( n19420 & ~n23361 ) ;
  assign n23363 = ( n3806 & ~n15095 ) | ( n3806 & n23362 ) | ( ~n15095 & n23362 ) ;
  assign n23364 = n17758 ^ n1228 ^ n280 ;
  assign n23365 = ( ~n5053 & n16323 ) | ( ~n5053 & n23364 ) | ( n16323 & n23364 ) ;
  assign n23366 = n23365 ^ n15425 ^ n7250 ;
  assign n23367 = n23366 ^ n20530 ^ n9748 ;
  assign n23368 = n17468 ^ n14029 ^ n9496 ;
  assign n23369 = x80 & ~n22568 ;
  assign n23370 = n23369 ^ n10927 ^ 1'b0 ;
  assign n23371 = n10480 ^ n2108 ^ n762 ;
  assign n23372 = n23371 ^ n12405 ^ 1'b0 ;
  assign n23373 = ( n23368 & n23370 ) | ( n23368 & ~n23372 ) | ( n23370 & ~n23372 ) ;
  assign n23374 = ( n3402 & n4289 ) | ( n3402 & n19848 ) | ( n4289 & n19848 ) ;
  assign n23375 = n23374 ^ n6235 ^ n1010 ;
  assign n23379 = n4571 & ~n10904 ;
  assign n23380 = n4893 & n23379 ;
  assign n23381 = n13615 | n23380 ;
  assign n23376 = ( ~n686 & n3771 ) | ( ~n686 & n11084 ) | ( n3771 & n11084 ) ;
  assign n23377 = n10640 & ~n22796 ;
  assign n23378 = ( ~n3708 & n23376 ) | ( ~n3708 & n23377 ) | ( n23376 & n23377 ) ;
  assign n23382 = n23381 ^ n23378 ^ n11983 ;
  assign n23383 = n8901 ^ n1572 ^ n1002 ;
  assign n23384 = ~n520 & n7771 ;
  assign n23385 = ( n4754 & n7476 ) | ( n4754 & n23384 ) | ( n7476 & n23384 ) ;
  assign n23386 = ( n369 & n23383 ) | ( n369 & n23385 ) | ( n23383 & n23385 ) ;
  assign n23387 = n7633 & n14802 ;
  assign n23389 = n3643 ^ n843 ^ n450 ;
  assign n23388 = n5271 ^ n4297 ^ n4037 ;
  assign n23390 = n23389 ^ n23388 ^ 1'b0 ;
  assign n23391 = ~n21952 & n23390 ;
  assign n23392 = ( n11712 & n23387 ) | ( n11712 & n23391 ) | ( n23387 & n23391 ) ;
  assign n23393 = ( n1538 & ~n3659 ) | ( n1538 & n15068 ) | ( ~n3659 & n15068 ) ;
  assign n23394 = n17489 ^ n1436 ^ 1'b0 ;
  assign n23395 = n23394 ^ n14462 ^ n6976 ;
  assign n23396 = ~n5669 & n23395 ;
  assign n23397 = ~n23393 & n23396 ;
  assign n23398 = ( n6039 & n9950 ) | ( n6039 & n22988 ) | ( n9950 & n22988 ) ;
  assign n23399 = n15188 ^ n3401 ^ n2575 ;
  assign n23400 = ( ~n14687 & n16244 ) | ( ~n14687 & n23399 ) | ( n16244 & n23399 ) ;
  assign n23401 = ( ~n8228 & n11689 ) | ( ~n8228 & n19674 ) | ( n11689 & n19674 ) ;
  assign n23402 = ( n5038 & ~n14799 ) | ( n5038 & n23401 ) | ( ~n14799 & n23401 ) ;
  assign n23403 = ( n1615 & n8983 ) | ( n1615 & ~n17489 ) | ( n8983 & ~n17489 ) ;
  assign n23404 = ( n6999 & n12215 ) | ( n6999 & ~n23403 ) | ( n12215 & ~n23403 ) ;
  assign n23405 = ( ~n1924 & n4521 ) | ( ~n1924 & n23404 ) | ( n4521 & n23404 ) ;
  assign n23406 = ( n7236 & n10123 ) | ( n7236 & n17562 ) | ( n10123 & n17562 ) ;
  assign n23407 = ~n16271 & n23406 ;
  assign n23408 = n23405 & n23407 ;
  assign n23414 = n12413 ^ n11764 ^ n6525 ;
  assign n23413 = n2359 & n14321 ;
  assign n23411 = ( n5035 & ~n12724 ) | ( n5035 & n20442 ) | ( ~n12724 & n20442 ) ;
  assign n23409 = ( n3834 & n8897 ) | ( n3834 & n16288 ) | ( n8897 & n16288 ) ;
  assign n23410 = n14873 & ~n23409 ;
  assign n23412 = n23411 ^ n23410 ^ 1'b0 ;
  assign n23415 = n23414 ^ n23413 ^ n23412 ;
  assign n23419 = n4422 ^ n1993 ^ n645 ;
  assign n23420 = n23419 ^ n7369 ^ n1558 ;
  assign n23417 = n12799 ^ n8402 ^ n1958 ;
  assign n23416 = n14725 & n22137 ;
  assign n23418 = n23417 ^ n23416 ^ 1'b0 ;
  assign n23421 = n23420 ^ n23418 ^ n1561 ;
  assign n23422 = n2864 | n13837 ;
  assign n23423 = n5575 & n5852 ;
  assign n23424 = ~n7897 & n23423 ;
  assign n23425 = n2381 & ~n4772 ;
  assign n23426 = n23425 ^ n838 ^ 1'b0 ;
  assign n23427 = n15489 & n23426 ;
  assign n23428 = ( n4111 & n5700 ) | ( n4111 & n8796 ) | ( n5700 & n8796 ) ;
  assign n23429 = n14306 ^ n13885 ^ 1'b0 ;
  assign n23430 = n23429 ^ n17735 ^ n3851 ;
  assign n23431 = ( ~n3481 & n17533 ) | ( ~n3481 & n23430 ) | ( n17533 & n23430 ) ;
  assign n23432 = ( n23427 & ~n23428 ) | ( n23427 & n23431 ) | ( ~n23428 & n23431 ) ;
  assign n23433 = n9924 ^ n8025 ^ n854 ;
  assign n23434 = n23433 ^ n2065 ^ 1'b0 ;
  assign n23435 = ( n13204 & n18376 ) | ( n13204 & n21540 ) | ( n18376 & n21540 ) ;
  assign n23436 = n2536 & ~n4269 ;
  assign n23437 = ~n5758 & n23436 ;
  assign n23438 = ~n22225 & n23437 ;
  assign n23439 = n10135 | n18767 ;
  assign n23440 = n2843 & ~n23439 ;
  assign n23446 = ( n7149 & ~n8257 ) | ( n7149 & n11605 ) | ( ~n8257 & n11605 ) ;
  assign n23447 = ( n4508 & n15501 ) | ( n4508 & n23446 ) | ( n15501 & n23446 ) ;
  assign n23441 = ( n1104 & ~n4264 ) | ( n1104 & n8146 ) | ( ~n4264 & n8146 ) ;
  assign n23442 = n9287 ^ n6490 ^ n552 ;
  assign n23443 = ( n7029 & ~n8777 ) | ( n7029 & n23442 ) | ( ~n8777 & n23442 ) ;
  assign n23444 = n23443 ^ n828 ^ 1'b0 ;
  assign n23445 = ( n22780 & n23441 ) | ( n22780 & ~n23444 ) | ( n23441 & ~n23444 ) ;
  assign n23448 = n23447 ^ n23445 ^ n7696 ;
  assign n23449 = n14575 ^ n9525 ^ 1'b0 ;
  assign n23450 = ( n2767 & ~n13824 ) | ( n2767 & n23449 ) | ( ~n13824 & n23449 ) ;
  assign n23451 = ~n302 & n14248 ;
  assign n23452 = ~n20575 & n23451 ;
  assign n23453 = n23452 ^ n6851 ^ n1343 ;
  assign n23454 = n23453 ^ n10932 ^ n2312 ;
  assign n23457 = n16488 ^ n13351 ^ n3741 ;
  assign n23455 = ~n5242 & n15199 ;
  assign n23456 = n23455 ^ n7738 ^ 1'b0 ;
  assign n23458 = n23457 ^ n23456 ^ n14592 ;
  assign n23459 = n3071 & n23458 ;
  assign n23460 = n5566 & n23459 ;
  assign n23461 = ( n11335 & n23454 ) | ( n11335 & n23460 ) | ( n23454 & n23460 ) ;
  assign n23462 = n2428 ^ n271 ^ 1'b0 ;
  assign n23463 = n7598 | n23462 ;
  assign n23464 = ( n2658 & n19954 ) | ( n2658 & ~n20937 ) | ( n19954 & ~n20937 ) ;
  assign n23465 = ( n8782 & n23463 ) | ( n8782 & ~n23464 ) | ( n23463 & ~n23464 ) ;
  assign n23466 = ( ~n3326 & n14598 ) | ( ~n3326 & n23465 ) | ( n14598 & n23465 ) ;
  assign n23467 = ( ~n3286 & n4061 ) | ( ~n3286 & n5816 ) | ( n4061 & n5816 ) ;
  assign n23468 = n6185 & ~n23467 ;
  assign n23469 = n11269 ^ n8014 ^ n1131 ;
  assign n23470 = ( n9477 & ~n23468 ) | ( n9477 & n23469 ) | ( ~n23468 & n23469 ) ;
  assign n23471 = ( n2541 & n23466 ) | ( n2541 & n23470 ) | ( n23466 & n23470 ) ;
  assign n23472 = ( n18147 & ~n22168 ) | ( n18147 & n23107 ) | ( ~n22168 & n23107 ) ;
  assign n23473 = ( n5185 & n7244 ) | ( n5185 & n11119 ) | ( n7244 & n11119 ) ;
  assign n23474 = n11513 ^ n9569 ^ 1'b0 ;
  assign n23475 = ~n5519 & n23474 ;
  assign n23476 = ( n2375 & ~n4205 ) | ( n2375 & n23475 ) | ( ~n4205 & n23475 ) ;
  assign n23481 = n10178 & n12541 ;
  assign n23482 = n23481 ^ n14712 ^ 1'b0 ;
  assign n23477 = ~n8926 & n15048 ;
  assign n23478 = n23477 ^ n8335 ^ n7804 ;
  assign n23479 = ( ~n6371 & n10671 ) | ( ~n6371 & n23478 ) | ( n10671 & n23478 ) ;
  assign n23480 = ( ~n710 & n11529 ) | ( ~n710 & n23479 ) | ( n11529 & n23479 ) ;
  assign n23483 = n23482 ^ n23480 ^ n21024 ;
  assign n23484 = ( ~n21028 & n23476 ) | ( ~n21028 & n23483 ) | ( n23476 & n23483 ) ;
  assign n23485 = ( ~n365 & n23473 ) | ( ~n365 & n23484 ) | ( n23473 & n23484 ) ;
  assign n23486 = n1063 & n5730 ;
  assign n23487 = n23486 ^ n22092 ^ n17788 ;
  assign n23488 = n23487 ^ n3130 ^ n2669 ;
  assign n23489 = n8876 ^ n8318 ^ 1'b0 ;
  assign n23490 = ( n866 & ~n20009 ) | ( n866 & n23489 ) | ( ~n20009 & n23489 ) ;
  assign n23491 = n23490 ^ n7793 ^ n2958 ;
  assign n23492 = ~n23488 & n23491 ;
  assign n23493 = ~n23485 & n23492 ;
  assign n23494 = n9332 ^ n6348 ^ n4307 ;
  assign n23495 = n23494 ^ n9324 ^ n1746 ;
  assign n23496 = n17221 & ~n18877 ;
  assign n23497 = ( n1451 & n9182 ) | ( n1451 & n19829 ) | ( n9182 & n19829 ) ;
  assign n23498 = n3984 & n23497 ;
  assign n23499 = ~x32 & n23498 ;
  assign n23500 = n23499 ^ n22993 ^ n3705 ;
  assign n23501 = n23500 ^ n12809 ^ n6008 ;
  assign n23502 = ~n3768 & n15401 ;
  assign n23503 = n23502 ^ n19794 ^ 1'b0 ;
  assign n23504 = x107 & n2027 ;
  assign n23505 = ~n3476 & n23504 ;
  assign n23506 = n11159 ^ n1673 ^ n885 ;
  assign n23507 = n15179 ^ n12925 ^ 1'b0 ;
  assign n23508 = ~n23506 & n23507 ;
  assign n23509 = n23508 ^ n16309 ^ n4341 ;
  assign n23510 = ( n23503 & n23505 ) | ( n23503 & n23509 ) | ( n23505 & n23509 ) ;
  assign n23511 = ~n1031 & n14989 ;
  assign n23512 = ~n6521 & n23511 ;
  assign n23513 = n23512 ^ n22218 ^ n4036 ;
  assign n23514 = n17135 ^ n13980 ^ n9766 ;
  assign n23515 = ( n654 & n12493 ) | ( n654 & n23514 ) | ( n12493 & n23514 ) ;
  assign n23524 = n23039 ^ n19726 ^ n355 ;
  assign n23525 = x194 & ~n13287 ;
  assign n23526 = n23525 ^ n9780 ^ 1'b0 ;
  assign n23527 = n5875 ^ n2362 ^ n2061 ;
  assign n23528 = ( ~n15852 & n23526 ) | ( ~n15852 & n23527 ) | ( n23526 & n23527 ) ;
  assign n23529 = ~n23524 & n23528 ;
  assign n23521 = ( n4761 & ~n5726 ) | ( n4761 & n7128 ) | ( ~n5726 & n7128 ) ;
  assign n23522 = n23521 ^ n14634 ^ 1'b0 ;
  assign n23523 = ( n11001 & n20263 ) | ( n11001 & n23522 ) | ( n20263 & n23522 ) ;
  assign n23519 = n10835 | n20101 ;
  assign n23517 = n1291 ^ n985 ^ n969 ;
  assign n23516 = n1809 ^ n1309 ^ n1026 ;
  assign n23518 = n23517 ^ n23516 ^ n1823 ;
  assign n23520 = n23519 ^ n23518 ^ n10396 ;
  assign n23530 = n23529 ^ n23523 ^ n23520 ;
  assign n23531 = ( x13 & n17047 ) | ( x13 & ~n20772 ) | ( n17047 & ~n20772 ) ;
  assign n23532 = n22282 ^ n18822 ^ n2107 ;
  assign n23533 = n8240 & ~n12583 ;
  assign n23534 = n23533 ^ n17828 ^ 1'b0 ;
  assign n23535 = ( n9336 & n14283 ) | ( n9336 & n23534 ) | ( n14283 & n23534 ) ;
  assign n23536 = n15368 ^ n1742 ^ 1'b0 ;
  assign n23537 = n19600 ^ n17097 ^ n6932 ;
  assign n23538 = n23537 ^ n21159 ^ n15973 ;
  assign n23539 = ( ~n12354 & n23536 ) | ( ~n12354 & n23538 ) | ( n23536 & n23538 ) ;
  assign n23540 = n18328 ^ n1843 ^ 1'b0 ;
  assign n23541 = n23540 ^ n13623 ^ n2718 ;
  assign n23542 = n23138 ^ n15350 ^ n13938 ;
  assign n23543 = n23542 ^ n5787 ^ n915 ;
  assign n23544 = ( n9573 & ~n11970 ) | ( n9573 & n15169 ) | ( ~n11970 & n15169 ) ;
  assign n23545 = n23544 ^ n9033 ^ 1'b0 ;
  assign n23546 = n14710 ^ n10355 ^ n3092 ;
  assign n23549 = ( ~n1644 & n3890 ) | ( ~n1644 & n10637 ) | ( n3890 & n10637 ) ;
  assign n23547 = ( n704 & n1585 ) | ( n704 & n17715 ) | ( n1585 & n17715 ) ;
  assign n23548 = n23547 ^ n3479 ^ n2902 ;
  assign n23550 = n23549 ^ n23548 ^ 1'b0 ;
  assign n23551 = n23546 & ~n23550 ;
  assign n23558 = n18929 ^ n9522 ^ n8588 ;
  assign n23559 = n23558 ^ n18526 ^ n10933 ;
  assign n23560 = n23559 ^ n18747 ^ n1398 ;
  assign n23552 = n20198 ^ n8307 ^ n2654 ;
  assign n23553 = n753 | n14680 ;
  assign n23554 = ( n19500 & ~n23552 ) | ( n19500 & n23553 ) | ( ~n23552 & n23553 ) ;
  assign n23555 = n4861 | n6421 ;
  assign n23556 = n23555 ^ n2408 ^ 1'b0 ;
  assign n23557 = n23554 | n23556 ;
  assign n23561 = n23560 ^ n23557 ^ 1'b0 ;
  assign n23568 = n6503 | n10145 ;
  assign n23569 = n3714 & ~n23568 ;
  assign n23566 = n3573 | n9917 ;
  assign n23567 = n23566 ^ n15135 ^ 1'b0 ;
  assign n23562 = n13893 ^ n10502 ^ x179 ;
  assign n23563 = ( x98 & n7910 ) | ( x98 & n23562 ) | ( n7910 & n23562 ) ;
  assign n23564 = ( ~n12579 & n15377 ) | ( ~n12579 & n23563 ) | ( n15377 & n23563 ) ;
  assign n23565 = n23564 ^ n14957 ^ n312 ;
  assign n23570 = n23569 ^ n23567 ^ n23565 ;
  assign n23571 = n21949 ^ n18588 ^ n17641 ;
  assign n23572 = n2937 & n23357 ;
  assign n23573 = n23571 & n23572 ;
  assign n23575 = n18821 ^ n15735 ^ n14876 ;
  assign n23576 = n23575 ^ n7475 ^ n6931 ;
  assign n23574 = n7112 & n9385 ;
  assign n23577 = n23576 ^ n23574 ^ 1'b0 ;
  assign n23578 = ~n8148 & n18485 ;
  assign n23579 = n23578 ^ n21856 ^ 1'b0 ;
  assign n23580 = ~n13023 & n18691 ;
  assign n23581 = ~n22601 & n23580 ;
  assign n23582 = ( n20485 & n23579 ) | ( n20485 & n23581 ) | ( n23579 & n23581 ) ;
  assign n23583 = ( n6930 & n20924 ) | ( n6930 & n22091 ) | ( n20924 & n22091 ) ;
  assign n23584 = ~n13887 & n23583 ;
  assign n23590 = n5028 | n8810 ;
  assign n23587 = n10857 & ~n14189 ;
  assign n23586 = n1790 & ~n20656 ;
  assign n23588 = n23587 ^ n23586 ^ 1'b0 ;
  assign n23589 = ( n5666 & n7898 ) | ( n5666 & ~n23588 ) | ( n7898 & ~n23588 ) ;
  assign n23585 = ( n5828 & n11252 ) | ( n5828 & ~n23376 ) | ( n11252 & ~n23376 ) ;
  assign n23591 = n23590 ^ n23589 ^ n23585 ;
  assign n23592 = ( n3336 & n15016 ) | ( n3336 & n15357 ) | ( n15016 & n15357 ) ;
  assign n23593 = n23592 ^ n7334 ^ n2967 ;
  assign n23594 = n19785 ^ n19066 ^ n15104 ;
  assign n23595 = n23594 ^ n11228 ^ n7706 ;
  assign n23596 = n15368 ^ n12167 ^ n1638 ;
  assign n23597 = ( n3452 & ~n17005 ) | ( n3452 & n23506 ) | ( ~n17005 & n23506 ) ;
  assign n23598 = n23597 ^ n4703 ^ n3349 ;
  assign n23599 = n23598 ^ n18903 ^ n13792 ;
  assign n23600 = ( n5403 & n9283 ) | ( n5403 & n12222 ) | ( n9283 & n12222 ) ;
  assign n23601 = x10 & ~n23263 ;
  assign n23602 = ~n9125 & n23601 ;
  assign n23603 = n7690 & ~n22183 ;
  assign n23604 = ( n2372 & n5572 ) | ( n2372 & n11326 ) | ( n5572 & n11326 ) ;
  assign n23605 = n15125 & n23604 ;
  assign n23606 = n19062 ^ n15632 ^ n10087 ;
  assign n23607 = ( n16020 & n23605 ) | ( n16020 & n23606 ) | ( n23605 & n23606 ) ;
  assign n23608 = ( n1002 & n11122 ) | ( n1002 & ~n20251 ) | ( n11122 & ~n20251 ) ;
  assign n23609 = n23608 ^ n6211 ^ n3597 ;
  assign n23610 = n9647 ^ n8642 ^ n2826 ;
  assign n23611 = n23610 ^ n5505 ^ n3833 ;
  assign n23612 = n7246 & ~n7262 ;
  assign n23613 = ( n2349 & ~n23611 ) | ( n2349 & n23612 ) | ( ~n23611 & n23612 ) ;
  assign n23614 = n12588 ^ n10401 ^ 1'b0 ;
  assign n23615 = n3384 | n23614 ;
  assign n23616 = n23615 ^ n10445 ^ n3475 ;
  assign n23617 = n23616 ^ n21775 ^ n17535 ;
  assign n23618 = ( n8396 & n9654 ) | ( n8396 & n23617 ) | ( n9654 & n23617 ) ;
  assign n23619 = n17874 ^ n8536 ^ n3830 ;
  assign n23620 = ( n887 & n14294 ) | ( n887 & n23619 ) | ( n14294 & n23619 ) ;
  assign n23621 = n23620 ^ n20547 ^ n9230 ;
  assign n23622 = ( ~n20568 & n20795 ) | ( ~n20568 & n22510 ) | ( n20795 & n22510 ) ;
  assign n23624 = n21142 ^ n15549 ^ n1130 ;
  assign n23623 = n18226 | n18492 ;
  assign n23625 = n23624 ^ n23623 ^ 1'b0 ;
  assign n23626 = ( ~n971 & n2767 ) | ( ~n971 & n3814 ) | ( n2767 & n3814 ) ;
  assign n23627 = n12685 ^ n12445 ^ n401 ;
  assign n23628 = ( ~n22847 & n23626 ) | ( ~n22847 & n23627 ) | ( n23626 & n23627 ) ;
  assign n23629 = n18800 ^ n15200 ^ n4738 ;
  assign n23630 = n22334 ^ n3472 ^ n2620 ;
  assign n23631 = n2915 | n21419 ;
  assign n23632 = n23631 ^ n12086 ^ n8288 ;
  assign n23633 = n16789 ^ n9129 ^ n3723 ;
  assign n23634 = n19619 ^ n13368 ^ n11666 ;
  assign n23635 = n23634 ^ n16978 ^ n3680 ;
  assign n23636 = n11222 ^ n1547 ^ 1'b0 ;
  assign n23637 = n20401 & n23636 ;
  assign n23638 = ( n23633 & n23635 ) | ( n23633 & ~n23637 ) | ( n23635 & ~n23637 ) ;
  assign n23639 = n14764 ^ n13869 ^ n3356 ;
  assign n23640 = ( ~n834 & n19735 ) | ( ~n834 & n23639 ) | ( n19735 & n23639 ) ;
  assign n23641 = n7127 ^ n3306 ^ 1'b0 ;
  assign n23642 = x104 & ~n23641 ;
  assign n23643 = n23642 ^ n19249 ^ n6004 ;
  assign n23644 = ( n3619 & ~n7483 ) | ( n3619 & n8378 ) | ( ~n7483 & n8378 ) ;
  assign n23645 = n23644 ^ n16531 ^ n14371 ;
  assign n23646 = n18738 ^ n3834 ^ n2643 ;
  assign n23647 = ( ~n2480 & n23645 ) | ( ~n2480 & n23646 ) | ( n23645 & n23646 ) ;
  assign n23648 = n23643 | n23647 ;
  assign n23662 = ( ~n3426 & n4504 ) | ( ~n3426 & n19325 ) | ( n4504 & n19325 ) ;
  assign n23663 = ( n2223 & ~n7888 ) | ( n2223 & n23662 ) | ( ~n7888 & n23662 ) ;
  assign n23651 = n6177 ^ n3197 ^ x184 ;
  assign n23649 = ~n1956 & n9296 ;
  assign n23650 = n23649 ^ n1469 ^ 1'b0 ;
  assign n23652 = n23651 ^ n23650 ^ n11315 ;
  assign n23653 = n23652 ^ n19184 ^ n5142 ;
  assign n23658 = n3282 & ~n4741 ;
  assign n23659 = n23658 ^ n544 ^ 1'b0 ;
  assign n23656 = ( ~n1204 & n3487 ) | ( ~n1204 & n5235 ) | ( n3487 & n5235 ) ;
  assign n23654 = ( n4681 & n6830 ) | ( n4681 & n11530 ) | ( n6830 & n11530 ) ;
  assign n23655 = n23654 ^ n17233 ^ n9599 ;
  assign n23657 = n23656 ^ n23655 ^ n12107 ;
  assign n23660 = n23659 ^ n23657 ^ n23443 ;
  assign n23661 = n23653 & ~n23660 ;
  assign n23664 = n23663 ^ n23661 ^ 1'b0 ;
  assign n23665 = ( ~n2963 & n11010 ) | ( ~n2963 & n19418 ) | ( n11010 & n19418 ) ;
  assign n23666 = n23665 ^ n18406 ^ n16542 ;
  assign n23667 = ( n8476 & n9341 ) | ( n8476 & n22269 ) | ( n9341 & n22269 ) ;
  assign n23668 = ( n1600 & n4127 ) | ( n1600 & n5481 ) | ( n4127 & n5481 ) ;
  assign n23669 = n23668 ^ n14356 ^ n9566 ;
  assign n23670 = ( n8357 & n11172 ) | ( n8357 & n23669 ) | ( n11172 & n23669 ) ;
  assign n23671 = n23670 ^ n6844 ^ 1'b0 ;
  assign n23672 = n7370 & ~n23671 ;
  assign n23673 = n23672 ^ n17439 ^ n7746 ;
  assign n23674 = n13367 ^ n3239 ^ x161 ;
  assign n23675 = ( ~n1985 & n2099 ) | ( ~n1985 & n23674 ) | ( n2099 & n23674 ) ;
  assign n23676 = ~n14747 & n19064 ;
  assign n23677 = ( n9425 & ~n21122 ) | ( n9425 & n23676 ) | ( ~n21122 & n23676 ) ;
  assign n23678 = n16040 & n18085 ;
  assign n23679 = n23678 ^ n12296 ^ 1'b0 ;
  assign n23682 = ( n6969 & n7657 ) | ( n6969 & n12582 ) | ( n7657 & n12582 ) ;
  assign n23680 = n22596 ^ n22027 ^ n15711 ;
  assign n23681 = n23680 ^ n9555 ^ 1'b0 ;
  assign n23683 = n23682 ^ n23681 ^ n7528 ;
  assign n23684 = n7658 ^ n3138 ^ n1868 ;
  assign n23685 = n20601 ^ n19273 ^ n19004 ;
  assign n23686 = ( n15516 & n23684 ) | ( n15516 & ~n23685 ) | ( n23684 & ~n23685 ) ;
  assign n23687 = n19943 & n23686 ;
  assign n23688 = ~n23683 & n23687 ;
  assign n23690 = ( n7528 & n11165 ) | ( n7528 & ~n21958 ) | ( n11165 & ~n21958 ) ;
  assign n23689 = ~n12029 & n16926 ;
  assign n23691 = n23690 ^ n23689 ^ 1'b0 ;
  assign n23692 = n17542 & n23691 ;
  assign n23693 = n23692 ^ n20093 ^ n1189 ;
  assign n23694 = ( n717 & n9573 ) | ( n717 & ~n11853 ) | ( n9573 & ~n11853 ) ;
  assign n23695 = n23694 ^ n11816 ^ n1048 ;
  assign n23696 = ( n11902 & n12110 ) | ( n11902 & n21470 ) | ( n12110 & n21470 ) ;
  assign n23697 = ( n7744 & ~n13567 ) | ( n7744 & n23696 ) | ( ~n13567 & n23696 ) ;
  assign n23698 = ( n7460 & n15349 ) | ( n7460 & ~n23697 ) | ( n15349 & ~n23697 ) ;
  assign n23700 = n4473 & ~n15501 ;
  assign n23701 = n23700 ^ n8009 ^ 1'b0 ;
  assign n23702 = n23701 ^ n3903 ^ n582 ;
  assign n23699 = n10390 ^ n3869 ^ n3595 ;
  assign n23703 = n23702 ^ n23699 ^ n7923 ;
  assign n23704 = n23703 ^ n846 ^ 1'b0 ;
  assign n23705 = n23704 ^ n21426 ^ n14136 ;
  assign n23706 = ( ~n4938 & n9619 ) | ( ~n4938 & n17882 ) | ( n9619 & n17882 ) ;
  assign n23707 = n23706 ^ n8307 ^ n1985 ;
  assign n23708 = ( ~n7154 & n7501 ) | ( ~n7154 & n23707 ) | ( n7501 & n23707 ) ;
  assign n23709 = n18493 ^ n12254 ^ n1864 ;
  assign n23710 = ( ~n8025 & n23708 ) | ( ~n8025 & n23709 ) | ( n23708 & n23709 ) ;
  assign n23711 = n10735 ^ n8680 ^ n4167 ;
  assign n23712 = n12451 | n23711 ;
  assign n23713 = n23712 ^ n4747 ^ 1'b0 ;
  assign n23714 = n19907 ^ n16062 ^ n4307 ;
  assign n23715 = n23475 & n23714 ;
  assign n23716 = n23713 & n23715 ;
  assign n23722 = ( n597 & n3134 ) | ( n597 & n3395 ) | ( n3134 & n3395 ) ;
  assign n23723 = n20293 ^ n2656 ^ 1'b0 ;
  assign n23724 = n23722 & ~n23723 ;
  assign n23717 = n17182 ^ n5106 ^ 1'b0 ;
  assign n23718 = n6864 | n23717 ;
  assign n23719 = n12235 ^ n7539 ^ n4643 ;
  assign n23720 = ( n6403 & ~n11481 ) | ( n6403 & n23719 ) | ( ~n11481 & n23719 ) ;
  assign n23721 = ~n23718 & n23720 ;
  assign n23725 = n23724 ^ n23721 ^ n22010 ;
  assign n23726 = ( n2457 & n13119 ) | ( n2457 & n23725 ) | ( n13119 & n23725 ) ;
  assign n23727 = ~n2417 & n3008 ;
  assign n23728 = ( n9218 & ~n14112 ) | ( n9218 & n23727 ) | ( ~n14112 & n23727 ) ;
  assign n23729 = ( n3735 & ~n6446 ) | ( n3735 & n19475 ) | ( ~n6446 & n19475 ) ;
  assign n23730 = ( n2564 & n2727 ) | ( n2564 & n18414 ) | ( n2727 & n18414 ) ;
  assign n23731 = ( n615 & n13014 ) | ( n615 & ~n23730 ) | ( n13014 & ~n23730 ) ;
  assign n23732 = ( n20088 & n23729 ) | ( n20088 & n23731 ) | ( n23729 & n23731 ) ;
  assign n23733 = n18564 ^ n2565 ^ 1'b0 ;
  assign n23734 = n20754 ^ n3126 ^ n1750 ;
  assign n23735 = n1705 & ~n11015 ;
  assign n23736 = ( n8732 & ~n23734 ) | ( n8732 & n23735 ) | ( ~n23734 & n23735 ) ;
  assign n23737 = n11030 & n14234 ;
  assign n23738 = n23737 ^ n16775 ^ 1'b0 ;
  assign n23739 = n18330 & ~n23738 ;
  assign n23740 = n16087 ^ n9163 ^ 1'b0 ;
  assign n23741 = n23740 ^ n9939 ^ n4852 ;
  assign n23742 = n1417 | n11907 ;
  assign n23743 = n23741 | n23742 ;
  assign n23744 = n8617 & ~n20786 ;
  assign n23745 = ( n1250 & n7507 ) | ( n1250 & ~n23182 ) | ( n7507 & ~n23182 ) ;
  assign n23746 = ~n14349 & n15577 ;
  assign n23747 = n18868 ^ n15395 ^ n15097 ;
  assign n23748 = n21289 ^ n16743 ^ x181 ;
  assign n23749 = n7715 | n21108 ;
  assign n23750 = n14252 & ~n23749 ;
  assign n23751 = ( ~n23747 & n23748 ) | ( ~n23747 & n23750 ) | ( n23748 & n23750 ) ;
  assign n23752 = n16907 ^ n5224 ^ n5028 ;
  assign n23753 = n23752 ^ n6011 ^ n3921 ;
  assign n23754 = n23753 ^ n19980 ^ n16025 ;
  assign n23755 = ( ~n2349 & n16816 ) | ( ~n2349 & n21636 ) | ( n16816 & n21636 ) ;
  assign n23756 = ( x125 & ~n9509 ) | ( x125 & n9960 ) | ( ~n9509 & n9960 ) ;
  assign n23757 = x97 & n10600 ;
  assign n23758 = ~n20031 & n23757 ;
  assign n23759 = ( n1271 & n3218 ) | ( n1271 & ~n10335 ) | ( n3218 & ~n10335 ) ;
  assign n23760 = n23759 ^ n16545 ^ n4085 ;
  assign n23761 = n23760 ^ n8695 ^ x146 ;
  assign n23762 = n23758 | n23761 ;
  assign n23763 = n23756 & ~n23762 ;
  assign n23767 = ( ~n6068 & n12264 ) | ( ~n6068 & n21154 ) | ( n12264 & n21154 ) ;
  assign n23765 = n10357 & n20222 ;
  assign n23764 = ~n1859 & n15717 ;
  assign n23766 = n23765 ^ n23764 ^ 1'b0 ;
  assign n23768 = n23767 ^ n23766 ^ 1'b0 ;
  assign n23769 = n23394 ^ n17172 ^ n9119 ;
  assign n23777 = n20288 ^ n5291 ^ n2640 ;
  assign n23776 = n17405 ^ n5354 ^ 1'b0 ;
  assign n23771 = ( n10418 & ~n21132 ) | ( n10418 & n23477 ) | ( ~n21132 & n23477 ) ;
  assign n23772 = n23771 ^ n18059 ^ n15093 ;
  assign n23773 = ( n907 & n20099 ) | ( n907 & ~n23772 ) | ( n20099 & ~n23772 ) ;
  assign n23770 = n688 & ~n4166 ;
  assign n23774 = n23773 ^ n23770 ^ n6397 ;
  assign n23775 = n23774 ^ n566 ^ 1'b0 ;
  assign n23778 = n23777 ^ n23776 ^ n23775 ;
  assign n23779 = ~n10409 & n18785 ;
  assign n23783 = ( n909 & n4350 ) | ( n909 & n7115 ) | ( n4350 & n7115 ) ;
  assign n23784 = n23783 ^ n14181 ^ n4770 ;
  assign n23780 = n10065 ^ n7911 ^ n3562 ;
  assign n23781 = n23780 ^ n17738 ^ 1'b0 ;
  assign n23782 = n10937 | n23781 ;
  assign n23785 = n23784 ^ n23782 ^ n17476 ;
  assign n23786 = ( n3665 & n5780 ) | ( n3665 & n23785 ) | ( n5780 & n23785 ) ;
  assign n23787 = ( n23778 & ~n23779 ) | ( n23778 & n23786 ) | ( ~n23779 & n23786 ) ;
  assign n23788 = n7659 ^ n6056 ^ 1'b0 ;
  assign n23789 = n2045 & n23788 ;
  assign n23790 = n23789 ^ n21952 ^ n4668 ;
  assign n23791 = ( n5063 & n5257 ) | ( n5063 & n11098 ) | ( n5257 & n11098 ) ;
  assign n23792 = n4850 & ~n23791 ;
  assign n23795 = n14136 ^ n11758 ^ n10563 ;
  assign n23793 = ( n309 & n7059 ) | ( n309 & ~n14961 ) | ( n7059 & ~n14961 ) ;
  assign n23794 = n13274 | n23793 ;
  assign n23796 = n23795 ^ n23794 ^ 1'b0 ;
  assign n23797 = n3559 | n14353 ;
  assign n23798 = ( n9693 & n20599 ) | ( n9693 & n23797 ) | ( n20599 & n23797 ) ;
  assign n23805 = n13843 ^ n8098 ^ n5930 ;
  assign n23802 = n4884 & ~n5240 ;
  assign n23803 = ~n12693 & n23802 ;
  assign n23801 = n21353 ^ n11632 ^ n5778 ;
  assign n23804 = n23803 ^ n23801 ^ n23534 ;
  assign n23799 = n12390 ^ n11983 ^ n8852 ;
  assign n23800 = n23799 ^ n426 ^ 1'b0 ;
  assign n23806 = n23805 ^ n23804 ^ n23800 ;
  assign n23807 = ( n836 & n1567 ) | ( n836 & ~n6427 ) | ( n1567 & ~n6427 ) ;
  assign n23808 = n3124 & n23807 ;
  assign n23811 = n23249 ^ n13715 ^ 1'b0 ;
  assign n23809 = ( n16452 & ~n16772 ) | ( n16452 & n19540 ) | ( ~n16772 & n19540 ) ;
  assign n23810 = ( n937 & n14298 ) | ( n937 & n23809 ) | ( n14298 & n23809 ) ;
  assign n23812 = n23811 ^ n23810 ^ n6175 ;
  assign n23815 = n5160 & ~n11673 ;
  assign n23816 = n23815 ^ n13647 ^ 1'b0 ;
  assign n23817 = ( n4915 & n5023 ) | ( n4915 & n23816 ) | ( n5023 & n23816 ) ;
  assign n23813 = n11252 ^ n8223 ^ n579 ;
  assign n23814 = n5090 | n23813 ;
  assign n23818 = n23817 ^ n23814 ^ 1'b0 ;
  assign n23819 = n23818 ^ n22671 ^ n22233 ;
  assign n23820 = n13617 ^ n11141 ^ n9364 ;
  assign n23821 = n16775 ^ n8830 ^ n7397 ;
  assign n23822 = ( n4959 & ~n23820 ) | ( n4959 & n23821 ) | ( ~n23820 & n23821 ) ;
  assign n23824 = ( ~x93 & n9874 ) | ( ~x93 & n16148 ) | ( n9874 & n16148 ) ;
  assign n23823 = ( ~n2299 & n6064 ) | ( ~n2299 & n6174 ) | ( n6064 & n6174 ) ;
  assign n23825 = n23824 ^ n23823 ^ n1521 ;
  assign n23826 = n6908 & ~n23825 ;
  assign n23827 = ~n8106 & n23826 ;
  assign n23828 = ( ~n9416 & n10999 ) | ( ~n9416 & n18816 ) | ( n10999 & n18816 ) ;
  assign n23829 = n14191 ^ n12582 ^ n11443 ;
  assign n23830 = n23829 ^ n17723 ^ n9344 ;
  assign n23831 = n7861 ^ n5598 ^ 1'b0 ;
  assign n23832 = n11535 ^ n3164 ^ 1'b0 ;
  assign n23833 = n15140 & n23832 ;
  assign n23834 = ~n21728 & n23833 ;
  assign n23835 = ( n19111 & n23831 ) | ( n19111 & n23834 ) | ( n23831 & n23834 ) ;
  assign n23836 = n23835 ^ n11873 ^ n3711 ;
  assign n23837 = ~n12889 & n22101 ;
  assign n23838 = ~n20975 & n23837 ;
  assign n23846 = n11720 ^ n6679 ^ x60 ;
  assign n23845 = ( n4112 & ~n8062 ) | ( n4112 & n12548 ) | ( ~n8062 & n12548 ) ;
  assign n23847 = n23846 ^ n23845 ^ n19025 ;
  assign n23843 = n11482 ^ n9801 ^ n3782 ;
  assign n23839 = ( n9254 & ~n9507 ) | ( n9254 & n11577 ) | ( ~n9507 & n11577 ) ;
  assign n23840 = n23839 ^ n11168 ^ n1166 ;
  assign n23841 = n23019 ^ n12537 ^ n2814 ;
  assign n23842 = n23840 & n23841 ;
  assign n23844 = n23843 ^ n23842 ^ 1'b0 ;
  assign n23848 = n23847 ^ n23844 ^ n11659 ;
  assign n23849 = n12441 ^ n5763 ^ n2784 ;
  assign n23850 = ~n8985 & n14853 ;
  assign n23851 = ~n785 & n9805 ;
  assign n23852 = ( n23725 & ~n23850 ) | ( n23725 & n23851 ) | ( ~n23850 & n23851 ) ;
  assign n23855 = n11872 ^ n2397 ^ n510 ;
  assign n23856 = ( n8138 & n9931 ) | ( n8138 & ~n23855 ) | ( n9931 & ~n23855 ) ;
  assign n23857 = ( n1779 & n1810 ) | ( n1779 & ~n23856 ) | ( n1810 & ~n23856 ) ;
  assign n23853 = n20768 ^ n7037 ^ 1'b0 ;
  assign n23854 = ~n20099 & n23853 ;
  assign n23858 = n23857 ^ n23854 ^ n14695 ;
  assign n23859 = ( n1869 & n7073 ) | ( n1869 & ~n14306 ) | ( n7073 & ~n14306 ) ;
  assign n23860 = n15613 ^ n8740 ^ n5660 ;
  assign n23861 = ( x171 & n23859 ) | ( x171 & n23860 ) | ( n23859 & n23860 ) ;
  assign n23862 = ( n2390 & ~n4419 ) | ( n2390 & n18939 ) | ( ~n4419 & n18939 ) ;
  assign n23863 = n8841 ^ n5351 ^ 1'b0 ;
  assign n23864 = n23862 & n23863 ;
  assign n23865 = n23864 ^ n10635 ^ 1'b0 ;
  assign n23866 = ( n16700 & n18954 ) | ( n16700 & n23865 ) | ( n18954 & n23865 ) ;
  assign n23867 = n13828 & ~n23866 ;
  assign n23868 = n19982 & n23867 ;
  assign n23869 = n8346 & ~n21313 ;
  assign n23870 = ( n10600 & n15878 ) | ( n10600 & n16793 ) | ( n15878 & n16793 ) ;
  assign n23871 = ( n16091 & n23869 ) | ( n16091 & ~n23870 ) | ( n23869 & ~n23870 ) ;
  assign n23887 = n2118 & ~n16520 ;
  assign n23888 = n318 & n23887 ;
  assign n23881 = n23756 ^ n23519 ^ n11034 ;
  assign n23882 = ( n2941 & n4306 ) | ( n2941 & ~n13233 ) | ( n4306 & ~n13233 ) ;
  assign n23883 = n14748 ^ n12245 ^ 1'b0 ;
  assign n23884 = n7629 & n23883 ;
  assign n23885 = ( n4122 & ~n23882 ) | ( n4122 & n23884 ) | ( ~n23882 & n23884 ) ;
  assign n23886 = ( n10294 & ~n23881 ) | ( n10294 & n23885 ) | ( ~n23881 & n23885 ) ;
  assign n23879 = ( ~n1101 & n1676 ) | ( ~n1101 & n9726 ) | ( n1676 & n9726 ) ;
  assign n23877 = ( n3598 & ~n4073 ) | ( n3598 & n5901 ) | ( ~n4073 & n5901 ) ;
  assign n23878 = n23877 ^ n18088 ^ n12964 ;
  assign n23873 = n6845 ^ n6207 ^ 1'b0 ;
  assign n23874 = n23873 ^ n19952 ^ n14363 ;
  assign n23875 = ( ~n16268 & n19367 ) | ( ~n16268 & n23874 ) | ( n19367 & n23874 ) ;
  assign n23872 = ( ~n2084 & n22717 ) | ( ~n2084 & n23759 ) | ( n22717 & n23759 ) ;
  assign n23876 = n23875 ^ n23872 ^ n19640 ;
  assign n23880 = n23879 ^ n23878 ^ n23876 ;
  assign n23889 = n23888 ^ n23886 ^ n23880 ;
  assign n23890 = n5263 ^ n4418 ^ 1'b0 ;
  assign n23891 = n21207 | n23890 ;
  assign n23892 = n14730 | n16512 ;
  assign n23893 = ( n7057 & n10515 ) | ( n7057 & n12849 ) | ( n10515 & n12849 ) ;
  assign n23894 = n23893 ^ n6735 ^ 1'b0 ;
  assign n23895 = n23894 ^ n11047 ^ n5267 ;
  assign n23900 = n6202 | n22898 ;
  assign n23901 = n5575 | n23900 ;
  assign n23896 = n19457 ^ n16544 ^ n8876 ;
  assign n23897 = n5879 & ~n23896 ;
  assign n23898 = n4333 & n23897 ;
  assign n23899 = ( n6177 & ~n16156 ) | ( n6177 & n23898 ) | ( ~n16156 & n23898 ) ;
  assign n23902 = n23901 ^ n23899 ^ n8815 ;
  assign n23903 = n23902 ^ n1213 ^ 1'b0 ;
  assign n23904 = n22145 | n23903 ;
  assign n23905 = n10163 ^ n1992 ^ n507 ;
  assign n23906 = n23905 ^ n22599 ^ n6963 ;
  assign n23907 = n21954 ^ n2021 ^ n1381 ;
  assign n23916 = n13309 ^ n5576 ^ n5425 ;
  assign n23914 = n18904 ^ n16419 ^ 1'b0 ;
  assign n23908 = n17421 ^ n3793 ^ n1663 ;
  assign n23909 = n23347 ^ n7901 ^ n2504 ;
  assign n23910 = ( n725 & n3112 ) | ( n725 & ~n13063 ) | ( n3112 & ~n13063 ) ;
  assign n23911 = n23910 ^ n15720 ^ 1'b0 ;
  assign n23912 = n23909 & ~n23911 ;
  assign n23913 = ( n11066 & ~n23908 ) | ( n11066 & n23912 ) | ( ~n23908 & n23912 ) ;
  assign n23915 = n23914 ^ n23913 ^ n9121 ;
  assign n23917 = n23916 ^ n23915 ^ n21488 ;
  assign n23919 = n2701 & n15980 ;
  assign n23918 = ( n2962 & ~n19631 ) | ( n2962 & n22095 ) | ( ~n19631 & n22095 ) ;
  assign n23920 = n23919 ^ n23918 ^ n22426 ;
  assign n23921 = n2386 & n2827 ;
  assign n23922 = n18181 ^ n13429 ^ n7312 ;
  assign n23923 = n6189 ^ n3959 ^ n1886 ;
  assign n23924 = ( n3894 & n14838 ) | ( n3894 & ~n23923 ) | ( n14838 & ~n23923 ) ;
  assign n23925 = ( n23921 & n23922 ) | ( n23921 & ~n23924 ) | ( n23922 & ~n23924 ) ;
  assign n23926 = n16545 ^ n11945 ^ 1'b0 ;
  assign n23927 = n23926 ^ n13808 ^ 1'b0 ;
  assign n23928 = n10883 | n23927 ;
  assign n23933 = n16927 ^ n4077 ^ n999 ;
  assign n23934 = ( n9864 & n13987 ) | ( n9864 & ~n23933 ) | ( n13987 & ~n23933 ) ;
  assign n23929 = n4743 ^ n3564 ^ n420 ;
  assign n23930 = ( n6073 & n21846 ) | ( n6073 & ~n23929 ) | ( n21846 & ~n23929 ) ;
  assign n23931 = n23930 ^ n16475 ^ n9141 ;
  assign n23932 = n23931 ^ n8894 ^ n4223 ;
  assign n23935 = n23934 ^ n23932 ^ n7819 ;
  assign n23936 = ( n2880 & n4933 ) | ( n2880 & ~n19179 ) | ( n4933 & ~n19179 ) ;
  assign n23937 = n23936 ^ n13606 ^ 1'b0 ;
  assign n23938 = ( ~n6045 & n10307 ) | ( ~n6045 & n20841 ) | ( n10307 & n20841 ) ;
  assign n23939 = n23938 ^ n2991 ^ x185 ;
  assign n23940 = ( n5196 & n12485 ) | ( n5196 & ~n12861 ) | ( n12485 & ~n12861 ) ;
  assign n23941 = ( n2771 & n22651 ) | ( n2771 & ~n23940 ) | ( n22651 & ~n23940 ) ;
  assign n23942 = n23356 ^ n10788 ^ n5467 ;
  assign n23943 = ( n5468 & n22018 ) | ( n5468 & n23942 ) | ( n22018 & n23942 ) ;
  assign n23944 = n20989 ^ n10575 ^ 1'b0 ;
  assign n23945 = n17601 | n23944 ;
  assign n23946 = n7354 ^ n5187 ^ x68 ;
  assign n23947 = n6716 | n9081 ;
  assign n23948 = n14190 ^ n12122 ^ x252 ;
  assign n23949 = n13735 ^ n7082 ^ n1196 ;
  assign n23950 = ( n17809 & n23948 ) | ( n17809 & n23949 ) | ( n23948 & n23949 ) ;
  assign n23951 = n14663 ^ n8078 ^ 1'b0 ;
  assign n23952 = ~n14166 & n23951 ;
  assign n23953 = ( ~n2780 & n12627 ) | ( ~n2780 & n21770 ) | ( n12627 & n21770 ) ;
  assign n23954 = ( n14653 & n23952 ) | ( n14653 & ~n23953 ) | ( n23952 & ~n23953 ) ;
  assign n23955 = n18278 | n22429 ;
  assign n23956 = ( n3236 & n8009 ) | ( n3236 & ~n23955 ) | ( n8009 & ~n23955 ) ;
  assign n23960 = n16075 ^ n11756 ^ n7518 ;
  assign n23959 = ( n8745 & ~n11746 ) | ( n8745 & n19119 ) | ( ~n11746 & n19119 ) ;
  assign n23957 = n13430 & ~n23320 ;
  assign n23958 = n7217 & n23957 ;
  assign n23961 = n23960 ^ n23959 ^ n23958 ;
  assign n23962 = n19288 ^ n17469 ^ n4258 ;
  assign n23963 = n23962 ^ n12831 ^ 1'b0 ;
  assign n23964 = n23963 ^ n17746 ^ n10599 ;
  assign n23965 = n23964 ^ n5476 ^ n357 ;
  assign n23969 = ( n3811 & ~n10879 ) | ( n3811 & n17423 ) | ( ~n10879 & n17423 ) ;
  assign n23967 = x221 & ~n2727 ;
  assign n23968 = n23967 ^ n7456 ^ 1'b0 ;
  assign n23970 = n23969 ^ n23968 ^ n9167 ;
  assign n23966 = n3749 & ~n14786 ;
  assign n23971 = n23970 ^ n23966 ^ 1'b0 ;
  assign n23972 = n23971 ^ n17541 ^ n6451 ;
  assign n23973 = ( n12243 & n23965 ) | ( n12243 & ~n23972 ) | ( n23965 & ~n23972 ) ;
  assign n23974 = n4467 | n10729 ;
  assign n23975 = ( n7149 & n7528 ) | ( n7149 & n14200 ) | ( n7528 & n14200 ) ;
  assign n23976 = ( n14978 & n23974 ) | ( n14978 & n23975 ) | ( n23974 & n23975 ) ;
  assign n23977 = ( n7655 & n12642 ) | ( n7655 & n23976 ) | ( n12642 & n23976 ) ;
  assign n23978 = n23977 ^ x236 ^ 1'b0 ;
  assign n23979 = n23978 ^ n21681 ^ n5960 ;
  assign n23980 = n22662 ^ n19308 ^ n5368 ;
  assign n23981 = ( n7473 & n12951 ) | ( n7473 & n13105 ) | ( n12951 & n13105 ) ;
  assign n23982 = n17737 ^ n11196 ^ n4631 ;
  assign n23983 = ~n13010 & n23183 ;
  assign n23984 = n23983 ^ n17708 ^ 1'b0 ;
  assign n23985 = ( n10271 & ~n23982 ) | ( n10271 & n23984 ) | ( ~n23982 & n23984 ) ;
  assign n23986 = ( x167 & n12625 ) | ( x167 & ~n23985 ) | ( n12625 & ~n23985 ) ;
  assign n23987 = ( ~n2619 & n23981 ) | ( ~n2619 & n23986 ) | ( n23981 & n23986 ) ;
  assign n23988 = ( n15989 & n17542 ) | ( n15989 & ~n22751 ) | ( n17542 & ~n22751 ) ;
  assign n23990 = n3924 & ~n5935 ;
  assign n23991 = n23990 ^ n1213 ^ 1'b0 ;
  assign n23989 = n3039 & n13661 ;
  assign n23992 = n23991 ^ n23989 ^ 1'b0 ;
  assign n23993 = n23992 ^ n13031 ^ n12167 ;
  assign n24000 = ( x27 & n3693 ) | ( x27 & n17323 ) | ( n3693 & n17323 ) ;
  assign n23994 = n12297 ^ n1115 ^ 1'b0 ;
  assign n23995 = n13391 & ~n23994 ;
  assign n23996 = n23995 ^ n18531 ^ n2391 ;
  assign n23997 = ( x3 & n2809 ) | ( x3 & ~n23996 ) | ( n2809 & ~n23996 ) ;
  assign n23998 = n23997 ^ n20234 ^ x70 ;
  assign n23999 = ( n2099 & n10758 ) | ( n2099 & ~n23998 ) | ( n10758 & ~n23998 ) ;
  assign n24001 = n24000 ^ n23999 ^ n9592 ;
  assign n24002 = n10836 ^ n3527 ^ n3229 ;
  assign n24003 = n1643 | n2814 ;
  assign n24004 = n4655 & ~n24003 ;
  assign n24005 = n24004 ^ n21345 ^ n300 ;
  assign n24006 = ( n1540 & n5792 ) | ( n1540 & n24005 ) | ( n5792 & n24005 ) ;
  assign n24007 = ( n17934 & n24002 ) | ( n17934 & n24006 ) | ( n24002 & n24006 ) ;
  assign n24008 = ( n3988 & n4158 ) | ( n3988 & n6452 ) | ( n4158 & n6452 ) ;
  assign n24009 = ( n859 & n1745 ) | ( n859 & ~n14977 ) | ( n1745 & ~n14977 ) ;
  assign n24010 = ( n20157 & n24008 ) | ( n20157 & ~n24009 ) | ( n24008 & ~n24009 ) ;
  assign n24011 = n8848 & ~n18939 ;
  assign n24012 = n2413 & n24011 ;
  assign n24013 = n24012 ^ n15983 ^ n12323 ;
  assign n24014 = n24013 ^ n23023 ^ n14283 ;
  assign n24022 = ( n5199 & n6748 ) | ( n5199 & n20051 ) | ( n6748 & n20051 ) ;
  assign n24015 = n21111 ^ n9008 ^ n2959 ;
  assign n24018 = ~n3897 & n5867 ;
  assign n24019 = ( n1835 & ~n5560 ) | ( n1835 & n24018 ) | ( ~n5560 & n24018 ) ;
  assign n24016 = n12960 ^ n11710 ^ 1'b0 ;
  assign n24017 = ( n12893 & n14077 ) | ( n12893 & n24016 ) | ( n14077 & n24016 ) ;
  assign n24020 = n24019 ^ n24017 ^ 1'b0 ;
  assign n24021 = n24015 & n24020 ;
  assign n24023 = n24022 ^ n24021 ^ n3501 ;
  assign n24024 = ( n2247 & n11319 ) | ( n2247 & ~n15376 ) | ( n11319 & ~n15376 ) ;
  assign n24025 = n24024 ^ n6694 ^ 1'b0 ;
  assign n24026 = n20278 ^ n15837 ^ n4361 ;
  assign n24027 = n24026 ^ n12651 ^ n10519 ;
  assign n24028 = n15492 ^ n4659 ^ n522 ;
  assign n24029 = ( n12273 & ~n19583 ) | ( n12273 & n24028 ) | ( ~n19583 & n24028 ) ;
  assign n24034 = n18362 ^ n4937 ^ 1'b0 ;
  assign n24035 = n18493 | n24034 ;
  assign n24033 = n15135 ^ n12245 ^ n3873 ;
  assign n24030 = n9346 ^ n8326 ^ n1629 ;
  assign n24031 = ( n10690 & n15351 ) | ( n10690 & n18432 ) | ( n15351 & n18432 ) ;
  assign n24032 = ( n1494 & ~n24030 ) | ( n1494 & n24031 ) | ( ~n24030 & n24031 ) ;
  assign n24036 = n24035 ^ n24033 ^ n24032 ;
  assign n24037 = ( ~n9599 & n13755 ) | ( ~n9599 & n24036 ) | ( n13755 & n24036 ) ;
  assign n24040 = n20670 ^ n8582 ^ 1'b0 ;
  assign n24041 = n5187 & ~n24040 ;
  assign n24038 = n15197 ^ n11929 ^ n4194 ;
  assign n24039 = n11906 | n24038 ;
  assign n24042 = n24041 ^ n24039 ^ 1'b0 ;
  assign n24043 = n24042 ^ n7832 ^ n4431 ;
  assign n24044 = ( n8478 & ~n21508 ) | ( n8478 & n24043 ) | ( ~n21508 & n24043 ) ;
  assign n24047 = n21607 ^ n17100 ^ n2535 ;
  assign n24045 = n22057 ^ n7178 ^ n2360 ;
  assign n24046 = n16103 & n24045 ;
  assign n24048 = n24047 ^ n24046 ^ 1'b0 ;
  assign n24049 = ( x112 & ~n3881 ) | ( x112 & n24048 ) | ( ~n3881 & n24048 ) ;
  assign n24050 = ( n364 & ~n507 ) | ( n364 & n12684 ) | ( ~n507 & n12684 ) ;
  assign n24051 = ( n10906 & n23075 ) | ( n10906 & n24050 ) | ( n23075 & n24050 ) ;
  assign n24052 = n11711 & n12964 ;
  assign n24053 = n24052 ^ n2046 ^ n901 ;
  assign n24054 = ( n1286 & n18349 ) | ( n1286 & ~n21761 ) | ( n18349 & ~n21761 ) ;
  assign n24055 = n6816 ^ n6665 ^ 1'b0 ;
  assign n24058 = n15471 ^ n10395 ^ n1122 ;
  assign n24056 = n4879 ^ n4651 ^ n3760 ;
  assign n24057 = n24056 ^ n1523 ^ 1'b0 ;
  assign n24059 = n24058 ^ n24057 ^ n9528 ;
  assign n24060 = n11898 ^ n9106 ^ n2019 ;
  assign n24061 = ( n7454 & n13666 ) | ( n7454 & n19606 ) | ( n13666 & n19606 ) ;
  assign n24062 = ( n16365 & ~n24060 ) | ( n16365 & n24061 ) | ( ~n24060 & n24061 ) ;
  assign n24063 = n24062 ^ n2553 ^ 1'b0 ;
  assign n24064 = n4968 | n24063 ;
  assign n24065 = n2230 & ~n16757 ;
  assign n24066 = n1760 & ~n4331 ;
  assign n24067 = ( ~n8415 & n14572 ) | ( ~n8415 & n24066 ) | ( n14572 & n24066 ) ;
  assign n24068 = n24067 ^ n4235 ^ 1'b0 ;
  assign n24069 = n4769 & n24068 ;
  assign n24070 = n14164 & ~n18230 ;
  assign n24071 = ~n20851 & n24070 ;
  assign n24072 = n14919 ^ n9275 ^ n6253 ;
  assign n24073 = ( n4264 & n19789 ) | ( n4264 & ~n24072 ) | ( n19789 & ~n24072 ) ;
  assign n24074 = n4827 ^ n3528 ^ n978 ;
  assign n24075 = n24074 ^ n7990 ^ n654 ;
  assign n24076 = ( x192 & ~n10262 ) | ( x192 & n12359 ) | ( ~n10262 & n12359 ) ;
  assign n24077 = n9165 ^ n3167 ^ 1'b0 ;
  assign n24078 = n20400 & n24077 ;
  assign n24079 = n9863 | n24078 ;
  assign n24082 = n8232 ^ n269 ^ x10 ;
  assign n24083 = ( n4370 & ~n12220 ) | ( n4370 & n24082 ) | ( ~n12220 & n24082 ) ;
  assign n24080 = n3391 ^ n3186 ^ 1'b0 ;
  assign n24081 = n21903 & n24080 ;
  assign n24084 = n24083 ^ n24081 ^ 1'b0 ;
  assign n24085 = ( n2766 & n8234 ) | ( n2766 & ~n13307 ) | ( n8234 & ~n13307 ) ;
  assign n24086 = n9479 ^ n1770 ^ n427 ;
  assign n24087 = n12326 ^ n2847 ^ 1'b0 ;
  assign n24088 = ( n1967 & ~n24086 ) | ( n1967 & n24087 ) | ( ~n24086 & n24087 ) ;
  assign n24089 = ( n1898 & n4310 ) | ( n1898 & n10396 ) | ( n4310 & n10396 ) ;
  assign n24090 = n11661 ^ n9344 ^ n8267 ;
  assign n24091 = n24090 ^ n13387 ^ n2351 ;
  assign n24092 = n24089 | n24091 ;
  assign n24093 = n24092 ^ n21045 ^ n17893 ;
  assign n24094 = n24093 ^ n21370 ^ n12329 ;
  assign n24095 = n4333 | n21434 ;
  assign n24096 = ( n5884 & n24094 ) | ( n5884 & ~n24095 ) | ( n24094 & ~n24095 ) ;
  assign n24097 = ( n459 & ~n7031 ) | ( n459 & n10874 ) | ( ~n7031 & n10874 ) ;
  assign n24099 = n17947 ^ n9767 ^ n3489 ;
  assign n24100 = ( ~n1266 & n2351 ) | ( ~n1266 & n21595 ) | ( n2351 & n21595 ) ;
  assign n24101 = ( n23309 & n24099 ) | ( n23309 & n24100 ) | ( n24099 & n24100 ) ;
  assign n24098 = n16577 ^ n10720 ^ n5281 ;
  assign n24102 = n24101 ^ n24098 ^ n16448 ;
  assign n24103 = n24102 ^ n22596 ^ n8878 ;
  assign n24104 = n5865 ^ n2516 ^ n364 ;
  assign n24105 = ( ~n3057 & n4810 ) | ( ~n3057 & n19025 ) | ( n4810 & n19025 ) ;
  assign n24106 = ( ~n21938 & n24104 ) | ( ~n21938 & n24105 ) | ( n24104 & n24105 ) ;
  assign n24107 = n6808 ^ n4316 ^ 1'b0 ;
  assign n24109 = ( ~n835 & n7923 ) | ( ~n835 & n21567 ) | ( n7923 & n21567 ) ;
  assign n24110 = n24109 ^ n9494 ^ n9029 ;
  assign n24108 = n11791 ^ n10651 ^ n10227 ;
  assign n24111 = n24110 ^ n24108 ^ n8653 ;
  assign n24112 = ( n1974 & n18741 ) | ( n1974 & n24111 ) | ( n18741 & n24111 ) ;
  assign n24113 = n20165 ^ n18108 ^ n14436 ;
  assign n24119 = ( ~n4301 & n5397 ) | ( ~n4301 & n7451 ) | ( n5397 & n7451 ) ;
  assign n24120 = n24119 ^ n4939 ^ n1709 ;
  assign n24114 = n15589 | n17108 ;
  assign n24115 = n4884 ^ n2667 ^ 1'b0 ;
  assign n24116 = ( n2853 & n24114 ) | ( n2853 & n24115 ) | ( n24114 & n24115 ) ;
  assign n24117 = ( n2117 & n3624 ) | ( n2117 & n21829 ) | ( n3624 & n21829 ) ;
  assign n24118 = ( n18945 & n24116 ) | ( n18945 & n24117 ) | ( n24116 & n24117 ) ;
  assign n24121 = n24120 ^ n24118 ^ n9982 ;
  assign n24122 = n17722 ^ n2752 ^ n2625 ;
  assign n24123 = n1583 & ~n11599 ;
  assign n24124 = ( n12998 & n21860 ) | ( n12998 & ~n24123 ) | ( n21860 & ~n24123 ) ;
  assign n24125 = n21138 & ~n21213 ;
  assign n24126 = ( ~n5281 & n8473 ) | ( ~n5281 & n24125 ) | ( n8473 & n24125 ) ;
  assign n24127 = ( n10096 & n24124 ) | ( n10096 & ~n24126 ) | ( n24124 & ~n24126 ) ;
  assign n24128 = ( n18023 & n19119 ) | ( n18023 & ~n24127 ) | ( n19119 & ~n24127 ) ;
  assign n24129 = ( n21881 & ~n24122 ) | ( n21881 & n24128 ) | ( ~n24122 & n24128 ) ;
  assign n24130 = ( ~n7727 & n19251 ) | ( ~n7727 & n21231 ) | ( n19251 & n21231 ) ;
  assign n24131 = n18871 ^ n10330 ^ n1194 ;
  assign n24132 = n5959 ^ n3592 ^ x42 ;
  assign n24133 = ( n1732 & n20633 ) | ( n1732 & ~n24132 ) | ( n20633 & ~n24132 ) ;
  assign n24134 = ( ~n3849 & n8641 ) | ( ~n3849 & n24133 ) | ( n8641 & n24133 ) ;
  assign n24135 = ( n24130 & n24131 ) | ( n24130 & n24134 ) | ( n24131 & n24134 ) ;
  assign n24136 = n24135 ^ n24024 ^ n18300 ;
  assign n24137 = ( n8346 & n8450 ) | ( n8346 & n9073 ) | ( n8450 & n9073 ) ;
  assign n24138 = n24137 ^ n13783 ^ n6855 ;
  assign n24139 = n7439 ^ n5575 ^ n2892 ;
  assign n24140 = ~n3989 & n16496 ;
  assign n24141 = n24140 ^ n7647 ^ 1'b0 ;
  assign n24142 = n24141 ^ n3147 ^ 1'b0 ;
  assign n24143 = n24142 ^ n10899 ^ n6344 ;
  assign n24144 = ~n21076 & n23132 ;
  assign n24145 = n24144 ^ n10937 ^ n2881 ;
  assign n24151 = n9466 & ~n15846 ;
  assign n24152 = n24151 ^ n14017 ^ 1'b0 ;
  assign n24153 = n4527 ^ n4002 ^ n1389 ;
  assign n24154 = ( n1946 & n24152 ) | ( n1946 & ~n24153 ) | ( n24152 & ~n24153 ) ;
  assign n24146 = n19718 ^ n8042 ^ n6962 ;
  assign n24148 = n4575 ^ n4191 ^ n3804 ;
  assign n24147 = n4310 & ~n17280 ;
  assign n24149 = n24148 ^ n24147 ^ 1'b0 ;
  assign n24150 = ( n11269 & ~n24146 ) | ( n11269 & n24149 ) | ( ~n24146 & n24149 ) ;
  assign n24155 = n24154 ^ n24150 ^ n12392 ;
  assign n24156 = ( n4113 & ~n24145 ) | ( n4113 & n24155 ) | ( ~n24145 & n24155 ) ;
  assign n24157 = ( n24139 & n24143 ) | ( n24139 & n24156 ) | ( n24143 & n24156 ) ;
  assign n24158 = n593 | n13443 ;
  assign n24159 = ( ~n1445 & n4218 ) | ( ~n1445 & n11892 ) | ( n4218 & n11892 ) ;
  assign n24160 = n24159 ^ n14463 ^ n11492 ;
  assign n24161 = ( n18964 & ~n24158 ) | ( n18964 & n24160 ) | ( ~n24158 & n24160 ) ;
  assign n24162 = n19250 ^ n17504 ^ x116 ;
  assign n24163 = n24162 ^ n7590 ^ n2050 ;
  assign n24164 = n24163 ^ n8552 ^ n4702 ;
  assign n24173 = ( n516 & n16769 ) | ( n516 & n18586 ) | ( n16769 & n18586 ) ;
  assign n24174 = ( ~n453 & n3393 ) | ( ~n453 & n24173 ) | ( n3393 & n24173 ) ;
  assign n24167 = n5698 ^ n4036 ^ n3450 ;
  assign n24165 = n7745 ^ n7526 ^ n4874 ;
  assign n24166 = n6883 & n24165 ;
  assign n24168 = n24167 ^ n24166 ^ 1'b0 ;
  assign n24169 = n19055 ^ n12079 ^ n2183 ;
  assign n24170 = ( n2761 & n24168 ) | ( n2761 & ~n24169 ) | ( n24168 & ~n24169 ) ;
  assign n24171 = ( n2710 & n11520 ) | ( n2710 & ~n24170 ) | ( n11520 & ~n24170 ) ;
  assign n24172 = n16190 & ~n24171 ;
  assign n24175 = n24174 ^ n24172 ^ 1'b0 ;
  assign n24176 = n14280 ^ n14139 ^ n9677 ;
  assign n24177 = n4497 ^ n4344 ^ n787 ;
  assign n24178 = ( n4098 & ~n11420 ) | ( n4098 & n24177 ) | ( ~n11420 & n24177 ) ;
  assign n24179 = n7098 ^ n588 ^ 1'b0 ;
  assign n24180 = ( ~n2756 & n6908 ) | ( ~n2756 & n24179 ) | ( n6908 & n24179 ) ;
  assign n24181 = n24180 ^ n3451 ^ 1'b0 ;
  assign n24182 = n1898 & n24181 ;
  assign n24183 = n14650 & n24182 ;
  assign n24184 = n9667 & n24183 ;
  assign n24185 = ( n12079 & n24178 ) | ( n12079 & n24184 ) | ( n24178 & n24184 ) ;
  assign n24186 = ( ~n14551 & n24176 ) | ( ~n14551 & n24185 ) | ( n24176 & n24185 ) ;
  assign n24187 = n18961 ^ n13425 ^ n11948 ;
  assign n24188 = n23304 ^ n17133 ^ n10269 ;
  assign n24190 = ( n14344 & n15388 ) | ( n14344 & ~n19326 ) | ( n15388 & ~n19326 ) ;
  assign n24189 = ( n497 & n4103 ) | ( n497 & n13522 ) | ( n4103 & n13522 ) ;
  assign n24191 = n24190 ^ n24189 ^ n22406 ;
  assign n24195 = n22095 ^ n14749 ^ 1'b0 ;
  assign n24196 = n14541 & n24195 ;
  assign n24192 = ( n2695 & ~n4096 ) | ( n2695 & n10441 ) | ( ~n4096 & n10441 ) ;
  assign n24193 = n24192 ^ n5800 ^ n692 ;
  assign n24194 = ( ~n4743 & n5909 ) | ( ~n4743 & n24193 ) | ( n5909 & n24193 ) ;
  assign n24197 = n24196 ^ n24194 ^ n10815 ;
  assign n24198 = ( n3093 & ~n14544 ) | ( n3093 & n24197 ) | ( ~n14544 & n24197 ) ;
  assign n24199 = ( n4775 & n5761 ) | ( n4775 & ~n9406 ) | ( n5761 & ~n9406 ) ;
  assign n24200 = n12654 ^ n802 ^ 1'b0 ;
  assign n24201 = ( n2124 & n24199 ) | ( n2124 & ~n24200 ) | ( n24199 & ~n24200 ) ;
  assign n24202 = n6349 ^ n3555 ^ 1'b0 ;
  assign n24203 = n17440 & n24202 ;
  assign n24204 = ( ~n10922 & n13065 ) | ( ~n10922 & n24203 ) | ( n13065 & n24203 ) ;
  assign n24205 = n3180 & ~n8849 ;
  assign n24206 = n24205 ^ n12158 ^ 1'b0 ;
  assign n24207 = n24206 ^ n17901 ^ 1'b0 ;
  assign n24208 = n21182 ^ n16656 ^ n9536 ;
  assign n24209 = ( n2122 & ~n5887 ) | ( n2122 & n22358 ) | ( ~n5887 & n22358 ) ;
  assign n24210 = n22098 ^ n13680 ^ n11078 ;
  assign n24216 = n9742 ^ n5525 ^ n3865 ;
  assign n24217 = ~n13773 & n24216 ;
  assign n24211 = ( n1407 & ~n6840 ) | ( n1407 & n15492 ) | ( ~n6840 & n15492 ) ;
  assign n24212 = ( x5 & n2580 ) | ( x5 & ~n24211 ) | ( n2580 & ~n24211 ) ;
  assign n24213 = ( n10790 & n17743 ) | ( n10790 & n24212 ) | ( n17743 & n24212 ) ;
  assign n24214 = ~n2869 & n24213 ;
  assign n24215 = n24214 ^ n15324 ^ n1776 ;
  assign n24218 = n24217 ^ n24215 ^ n15173 ;
  assign n24223 = ( n2682 & ~n3733 ) | ( n2682 & n13438 ) | ( ~n3733 & n13438 ) ;
  assign n24224 = ( ~n9522 & n16652 ) | ( ~n9522 & n24223 ) | ( n16652 & n24223 ) ;
  assign n24222 = ( n7355 & n19960 ) | ( n7355 & n21166 ) | ( n19960 & n21166 ) ;
  assign n24219 = ( n1175 & ~n5763 ) | ( n1175 & n5768 ) | ( ~n5763 & n5768 ) ;
  assign n24220 = n24219 ^ n19180 ^ n978 ;
  assign n24221 = ( n2930 & n12942 ) | ( n2930 & ~n24220 ) | ( n12942 & ~n24220 ) ;
  assign n24225 = n24224 ^ n24222 ^ n24221 ;
  assign n24226 = n15390 ^ n4240 ^ n2271 ;
  assign n24227 = n24226 ^ n20006 ^ n6119 ;
  assign n24228 = ( n4289 & ~n18586 ) | ( n4289 & n19320 ) | ( ~n18586 & n19320 ) ;
  assign n24229 = ( ~n14604 & n24227 ) | ( ~n14604 & n24228 ) | ( n24227 & n24228 ) ;
  assign n24230 = ( n478 & ~n24225 ) | ( n478 & n24229 ) | ( ~n24225 & n24229 ) ;
  assign n24231 = n10788 ^ n9325 ^ n9064 ;
  assign n24232 = n10480 ^ n5818 ^ n4110 ;
  assign n24233 = n24232 ^ n20978 ^ n2698 ;
  assign n24234 = n24072 ^ n5272 ^ n2394 ;
  assign n24235 = n24234 ^ n6405 ^ n3218 ;
  assign n24236 = n24235 ^ n15826 ^ n693 ;
  assign n24237 = n24236 ^ n11426 ^ n7189 ;
  assign n24238 = ( x1 & n1813 ) | ( x1 & n11660 ) | ( n1813 & n11660 ) ;
  assign n24239 = n3600 ^ n1308 ^ n467 ;
  assign n24240 = ( n1904 & n3579 ) | ( n1904 & ~n24239 ) | ( n3579 & ~n24239 ) ;
  assign n24241 = ( ~n2805 & n4048 ) | ( ~n2805 & n24240 ) | ( n4048 & n24240 ) ;
  assign n24242 = ( ~n21096 & n22691 ) | ( ~n21096 & n24241 ) | ( n22691 & n24241 ) ;
  assign n24243 = n24242 ^ n1411 ^ 1'b0 ;
  assign n24244 = n16806 ^ n10354 ^ n5749 ;
  assign n24245 = ( n868 & n20142 ) | ( n868 & ~n24244 ) | ( n20142 & ~n24244 ) ;
  assign n24246 = n19265 ^ n11209 ^ x94 ;
  assign n24247 = n18892 ^ n9576 ^ n9560 ;
  assign n24248 = ( n18131 & n24246 ) | ( n18131 & n24247 ) | ( n24246 & n24247 ) ;
  assign n24249 = n24248 ^ n8554 ^ n3763 ;
  assign n24250 = n4989 | n6962 ;
  assign n24251 = n24250 ^ n3637 ^ 1'b0 ;
  assign n24252 = ( n7872 & n11124 ) | ( n7872 & n24251 ) | ( n11124 & n24251 ) ;
  assign n24253 = ( n1384 & ~n9813 ) | ( n1384 & n21184 ) | ( ~n9813 & n21184 ) ;
  assign n24254 = n7103 ^ n2020 ^ 1'b0 ;
  assign n24255 = ( n24252 & n24253 ) | ( n24252 & ~n24254 ) | ( n24253 & ~n24254 ) ;
  assign n24256 = n19913 ^ n19492 ^ n14936 ;
  assign n24257 = n24256 ^ n8536 ^ n6676 ;
  assign n24258 = n24257 ^ n17133 ^ n6529 ;
  assign n24259 = n20988 ^ n20606 ^ n6763 ;
  assign n24263 = ( n5616 & n10579 ) | ( n5616 & ~n22310 ) | ( n10579 & ~n22310 ) ;
  assign n24264 = n24263 ^ n5369 ^ n3962 ;
  assign n24261 = ( n3347 & n16300 ) | ( n3347 & n17420 ) | ( n16300 & n17420 ) ;
  assign n24262 = n24261 ^ n483 ^ 1'b0 ;
  assign n24260 = n5780 & ~n22490 ;
  assign n24265 = n24264 ^ n24262 ^ n24260 ;
  assign n24266 = ( n10244 & n10525 ) | ( n10244 & ~n13341 ) | ( n10525 & ~n13341 ) ;
  assign n24267 = n24266 ^ n19101 ^ n3175 ;
  assign n24268 = n14617 ^ n12647 ^ n10227 ;
  assign n24269 = ( n7864 & n10121 ) | ( n7864 & ~n18436 ) | ( n10121 & ~n18436 ) ;
  assign n24270 = n11652 ^ n3263 ^ x210 ;
  assign n24271 = n8327 & n17802 ;
  assign n24272 = ~n24270 & n24271 ;
  assign n24273 = ( ~n7560 & n23318 ) | ( ~n7560 & n24272 ) | ( n23318 & n24272 ) ;
  assign n24274 = ( n7246 & n24269 ) | ( n7246 & n24273 ) | ( n24269 & n24273 ) ;
  assign n24275 = n13671 ^ n13645 ^ n5138 ;
  assign n24276 = ( n2762 & n10158 ) | ( n2762 & ~n24275 ) | ( n10158 & ~n24275 ) ;
  assign n24277 = ( n2857 & ~n19570 ) | ( n2857 & n21224 ) | ( ~n19570 & n21224 ) ;
  assign n24278 = ~n11899 & n24277 ;
  assign n24279 = n24276 & n24278 ;
  assign n24280 = n3575 & n10247 ;
  assign n24281 = ( n13610 & n22583 ) | ( n13610 & n24280 ) | ( n22583 & n24280 ) ;
  assign n24282 = ( n5489 & n17499 ) | ( n5489 & ~n23617 ) | ( n17499 & ~n23617 ) ;
  assign n24283 = n24282 ^ n17678 ^ n7626 ;
  assign n24284 = ( x198 & n7012 ) | ( x198 & n11299 ) | ( n7012 & n11299 ) ;
  assign n24285 = ( n6472 & n7968 ) | ( n6472 & n24284 ) | ( n7968 & n24284 ) ;
  assign n24286 = n24285 ^ n7505 ^ 1'b0 ;
  assign n24287 = ( n4134 & ~n6717 ) | ( n4134 & n24286 ) | ( ~n6717 & n24286 ) ;
  assign n24288 = n17957 ^ n14495 ^ n10932 ;
  assign n24289 = n24288 ^ n18272 ^ n5274 ;
  assign n24290 = ( ~n10807 & n13316 ) | ( ~n10807 & n14768 ) | ( n13316 & n14768 ) ;
  assign n24291 = n22121 ^ n7089 ^ 1'b0 ;
  assign n24292 = ( n10191 & n18273 ) | ( n10191 & n24291 ) | ( n18273 & n24291 ) ;
  assign n24293 = n4076 | n19921 ;
  assign n24294 = ( n19228 & n23984 ) | ( n19228 & n24293 ) | ( n23984 & n24293 ) ;
  assign n24295 = ( ~n4703 & n7887 ) | ( ~n4703 & n11169 ) | ( n7887 & n11169 ) ;
  assign n24296 = n23286 ^ n6167 ^ n899 ;
  assign n24297 = ( ~n19975 & n24295 ) | ( ~n19975 & n24296 ) | ( n24295 & n24296 ) ;
  assign n24298 = ~n1582 & n6206 ;
  assign n24299 = ~n5330 & n24298 ;
  assign n24300 = ( ~n9710 & n11847 ) | ( ~n9710 & n24299 ) | ( n11847 & n24299 ) ;
  assign n24301 = n24300 ^ n23594 ^ n4127 ;
  assign n24302 = ( n3639 & n5191 ) | ( n3639 & ~n24301 ) | ( n5191 & ~n24301 ) ;
  assign n24303 = ~n9511 & n14387 ;
  assign n24304 = n24303 ^ n15996 ^ 1'b0 ;
  assign n24305 = n3589 & ~n19971 ;
  assign n24306 = n10083 ^ n10082 ^ n651 ;
  assign n24307 = n24306 ^ n6828 ^ n1621 ;
  assign n24308 = n24307 ^ n14429 ^ n1729 ;
  assign n24309 = n10683 | n20559 ;
  assign n24310 = n24309 ^ n23519 ^ 1'b0 ;
  assign n24311 = ( x238 & n681 ) | ( x238 & n4922 ) | ( n681 & n4922 ) ;
  assign n24312 = ( n1787 & n15817 ) | ( n1787 & ~n19490 ) | ( n15817 & ~n19490 ) ;
  assign n24313 = n24311 & ~n24312 ;
  assign n24314 = n24313 ^ n13182 ^ n8703 ;
  assign n24319 = ( ~n2412 & n12182 ) | ( ~n2412 & n15236 ) | ( n12182 & n15236 ) ;
  assign n24320 = ( x210 & n6769 ) | ( x210 & n24319 ) | ( n6769 & n24319 ) ;
  assign n24321 = n24320 ^ n23181 ^ n16888 ;
  assign n24317 = n22757 ^ n15387 ^ n4662 ;
  assign n24315 = n3032 & ~n15532 ;
  assign n24316 = ( n6960 & n16624 ) | ( n6960 & n24315 ) | ( n16624 & n24315 ) ;
  assign n24318 = n24317 ^ n24316 ^ n21770 ;
  assign n24322 = n24321 ^ n24318 ^ n12888 ;
  assign n24323 = ( n2932 & n4386 ) | ( n2932 & n23909 ) | ( n4386 & n23909 ) ;
  assign n24324 = ( n1503 & ~n3407 ) | ( n1503 & n10233 ) | ( ~n3407 & n10233 ) ;
  assign n24325 = ( n12116 & n23784 ) | ( n12116 & ~n24324 ) | ( n23784 & ~n24324 ) ;
  assign n24326 = ( ~n466 & n24323 ) | ( ~n466 & n24325 ) | ( n24323 & n24325 ) ;
  assign n24332 = ( ~n1653 & n9182 ) | ( ~n1653 & n11733 ) | ( n9182 & n11733 ) ;
  assign n24327 = n18679 ^ n14355 ^ n5402 ;
  assign n24328 = n24327 ^ n10772 ^ x175 ;
  assign n24329 = n24328 ^ n10779 ^ n2552 ;
  assign n24330 = n24329 ^ n20930 ^ n18001 ;
  assign n24331 = ( n7387 & n15555 ) | ( n7387 & ~n24330 ) | ( n15555 & ~n24330 ) ;
  assign n24333 = n24332 ^ n24331 ^ n4623 ;
  assign n24334 = ( n8871 & n11479 ) | ( n8871 & ~n18360 ) | ( n11479 & ~n18360 ) ;
  assign n24335 = n24334 ^ n5780 ^ n3064 ;
  assign n24336 = ( n1328 & n7830 ) | ( n1328 & n24335 ) | ( n7830 & n24335 ) ;
  assign n24337 = n2237 | n7349 ;
  assign n24338 = n3109 | n24337 ;
  assign n24339 = ( n875 & n1499 ) | ( n875 & ~n24338 ) | ( n1499 & ~n24338 ) ;
  assign n24342 = n8032 ^ x39 ^ 1'b0 ;
  assign n24343 = ( n5006 & n7602 ) | ( n5006 & n24342 ) | ( n7602 & n24342 ) ;
  assign n24340 = ( n1226 & n1795 ) | ( n1226 & n18318 ) | ( n1795 & n18318 ) ;
  assign n24341 = ( ~n6266 & n8944 ) | ( ~n6266 & n24340 ) | ( n8944 & n24340 ) ;
  assign n24344 = n24343 ^ n24341 ^ n8384 ;
  assign n24345 = n24344 ^ n17460 ^ n13403 ;
  assign n24346 = n22664 ^ n10361 ^ n5862 ;
  assign n24347 = ( n575 & ~n4357 ) | ( n575 & n15984 ) | ( ~n4357 & n15984 ) ;
  assign n24348 = ( n3917 & n24346 ) | ( n3917 & ~n24347 ) | ( n24346 & ~n24347 ) ;
  assign n24349 = n17622 ^ n12375 ^ n770 ;
  assign n24350 = ( n21908 & n23259 ) | ( n21908 & n24349 ) | ( n23259 & n24349 ) ;
  assign n24351 = ( n14613 & n24348 ) | ( n14613 & ~n24350 ) | ( n24348 & ~n24350 ) ;
  assign n24357 = n11659 ^ n8018 ^ 1'b0 ;
  assign n24358 = ~n6238 & n24357 ;
  assign n24355 = n14697 ^ n7371 ^ n2469 ;
  assign n24356 = n24355 ^ n647 ^ n633 ;
  assign n24359 = n24358 ^ n24356 ^ n18526 ;
  assign n24360 = ( ~n13760 & n23748 ) | ( ~n13760 & n24359 ) | ( n23748 & n24359 ) ;
  assign n24352 = ( n2121 & n11208 ) | ( n2121 & n13713 ) | ( n11208 & n13713 ) ;
  assign n24353 = n11411 & n24352 ;
  assign n24354 = n20853 & n24353 ;
  assign n24361 = n24360 ^ n24354 ^ n15513 ;
  assign n24362 = ( n2918 & n11612 ) | ( n2918 & ~n15781 ) | ( n11612 & ~n15781 ) ;
  assign n24373 = n1762 & ~n6085 ;
  assign n24371 = n2724 | n4990 ;
  assign n24367 = n13311 ^ n7400 ^ n3224 ;
  assign n24368 = n24367 ^ n2020 ^ 1'b0 ;
  assign n24369 = ~n6834 & n24368 ;
  assign n24370 = ( n2324 & n3140 ) | ( n2324 & n24369 ) | ( n3140 & n24369 ) ;
  assign n24372 = n24371 ^ n24370 ^ n3199 ;
  assign n24364 = n10119 & ~n12373 ;
  assign n24365 = ~n261 & n24364 ;
  assign n24363 = ( n1903 & n4226 ) | ( n1903 & ~n5605 ) | ( n4226 & ~n5605 ) ;
  assign n24366 = n24365 ^ n24363 ^ n16831 ;
  assign n24374 = n24373 ^ n24372 ^ n24366 ;
  assign n24375 = n24374 ^ n10310 ^ n3703 ;
  assign n24376 = n6250 ^ n4180 ^ n967 ;
  assign n24377 = ( n9416 & n14699 ) | ( n9416 & ~n24235 ) | ( n14699 & ~n24235 ) ;
  assign n24378 = n15256 ^ n5041 ^ n1214 ;
  assign n24379 = n24378 ^ n11045 ^ 1'b0 ;
  assign n24380 = n1350 & n24379 ;
  assign n24381 = ( ~n6399 & n19017 ) | ( ~n6399 & n24380 ) | ( n19017 & n24380 ) ;
  assign n24384 = n16624 ^ n3991 ^ 1'b0 ;
  assign n24383 = ( ~n2790 & n8622 ) | ( ~n2790 & n18419 ) | ( n8622 & n18419 ) ;
  assign n24382 = n11248 ^ n2477 ^ 1'b0 ;
  assign n24385 = n24384 ^ n24383 ^ n24382 ;
  assign n24386 = n14672 ^ n8023 ^ n4074 ;
  assign n24387 = n24386 ^ n21218 ^ n15232 ;
  assign n24388 = ( ~n5220 & n6318 ) | ( ~n5220 & n12052 ) | ( n6318 & n12052 ) ;
  assign n24389 = ( n3526 & n8485 ) | ( n3526 & n20551 ) | ( n8485 & n20551 ) ;
  assign n24390 = ~n1943 & n10902 ;
  assign n24391 = n24390 ^ x94 ^ 1'b0 ;
  assign n24392 = ( n24388 & ~n24389 ) | ( n24388 & n24391 ) | ( ~n24389 & n24391 ) ;
  assign n24393 = n4985 ^ n2684 ^ 1'b0 ;
  assign n24394 = n23467 | n24393 ;
  assign n24395 = ( x78 & n4915 ) | ( x78 & n24394 ) | ( n4915 & n24394 ) ;
  assign n24396 = n24395 ^ n17392 ^ n2838 ;
  assign n24397 = ( n4958 & ~n6935 ) | ( n4958 & n24396 ) | ( ~n6935 & n24396 ) ;
  assign n24398 = ( n19284 & n24392 ) | ( n19284 & n24397 ) | ( n24392 & n24397 ) ;
  assign n24399 = n14263 ^ n1267 ^ n650 ;
  assign n24400 = ~n4935 & n20761 ;
  assign n24401 = ~n22478 & n24400 ;
  assign n24402 = n22065 ^ n5455 ^ n2162 ;
  assign n24410 = ( n1537 & ~n3239 ) | ( n1537 & n15702 ) | ( ~n3239 & n15702 ) ;
  assign n24411 = n10810 & ~n24410 ;
  assign n24403 = ( n1360 & ~n5682 ) | ( n1360 & n12455 ) | ( ~n5682 & n12455 ) ;
  assign n24404 = ( n3492 & ~n15501 ) | ( n3492 & n18925 ) | ( ~n15501 & n18925 ) ;
  assign n24405 = ( ~n8751 & n24403 ) | ( ~n8751 & n24404 ) | ( n24403 & n24404 ) ;
  assign n24406 = n24405 ^ n20743 ^ n8587 ;
  assign n24407 = n24406 ^ n14846 ^ n11847 ;
  assign n24408 = n24407 ^ n9932 ^ n6340 ;
  assign n24409 = n24408 ^ n9707 ^ x194 ;
  assign n24412 = n24411 ^ n24409 ^ n3044 ;
  assign n24413 = n10094 ^ n2106 ^ n837 ;
  assign n24414 = ~n6995 & n12489 ;
  assign n24415 = n24414 ^ n4942 ^ 1'b0 ;
  assign n24416 = n24415 ^ n19192 ^ n11555 ;
  assign n24417 = n24416 ^ n23349 ^ n14926 ;
  assign n24418 = ( n10148 & n11464 ) | ( n10148 & n23069 ) | ( n11464 & n23069 ) ;
  assign n24419 = n4314 & n24418 ;
  assign n24420 = n24419 ^ n13223 ^ 1'b0 ;
  assign n24421 = ( n6646 & n16846 ) | ( n6646 & n24420 ) | ( n16846 & n24420 ) ;
  assign n24422 = ( n1964 & n2121 ) | ( n1964 & ~n4220 ) | ( n2121 & ~n4220 ) ;
  assign n24423 = n14527 ^ n13233 ^ n5234 ;
  assign n24424 = n16079 & ~n24423 ;
  assign n24425 = n15765 | n24424 ;
  assign n24426 = n24422 & ~n24425 ;
  assign n24427 = n4444 & ~n24426 ;
  assign n24428 = n24427 ^ n1461 ^ 1'b0 ;
  assign n24429 = ( n1915 & ~n7767 ) | ( n1915 & n12212 ) | ( ~n7767 & n12212 ) ;
  assign n24430 = ( n5393 & n16660 ) | ( n5393 & n24429 ) | ( n16660 & n24429 ) ;
  assign n24431 = ( n5996 & n18827 ) | ( n5996 & ~n19292 ) | ( n18827 & ~n19292 ) ;
  assign n24432 = ( n21681 & n24430 ) | ( n21681 & ~n24431 ) | ( n24430 & ~n24431 ) ;
  assign n24433 = ( x199 & n20808 ) | ( x199 & n24432 ) | ( n20808 & n24432 ) ;
  assign n24434 = ( ~n477 & n2451 ) | ( ~n477 & n10614 ) | ( n2451 & n10614 ) ;
  assign n24435 = n24434 ^ n8692 ^ n3619 ;
  assign n24436 = n24435 ^ n14899 ^ n13185 ;
  assign n24437 = ( n7175 & n10226 ) | ( n7175 & ~n24436 ) | ( n10226 & ~n24436 ) ;
  assign n24439 = ( n2877 & n6918 ) | ( n2877 & ~n16786 ) | ( n6918 & ~n16786 ) ;
  assign n24438 = ( x55 & ~n17770 ) | ( x55 & n21579 ) | ( ~n17770 & n21579 ) ;
  assign n24440 = n24439 ^ n24438 ^ x158 ;
  assign n24441 = ( n3871 & n4285 ) | ( n3871 & n8226 ) | ( n4285 & n8226 ) ;
  assign n24442 = ( n1448 & ~n1557 ) | ( n1448 & n24441 ) | ( ~n1557 & n24441 ) ;
  assign n24443 = ( ~n16101 & n19484 ) | ( ~n16101 & n24442 ) | ( n19484 & n24442 ) ;
  assign n24444 = ( n3105 & n11340 ) | ( n3105 & n24443 ) | ( n11340 & n24443 ) ;
  assign n24447 = n23590 ^ n10186 ^ n5501 ;
  assign n24448 = ( n16164 & ~n24384 ) | ( n16164 & n24447 ) | ( ~n24384 & n24447 ) ;
  assign n24445 = ~n5033 & n6473 ;
  assign n24446 = n24445 ^ n11269 ^ 1'b0 ;
  assign n24449 = n24448 ^ n24446 ^ n12348 ;
  assign n24450 = ( ~n1178 & n12651 ) | ( ~n1178 & n19849 ) | ( n12651 & n19849 ) ;
  assign n24451 = n24450 ^ n11104 ^ 1'b0 ;
  assign n24452 = ( n3432 & n14677 ) | ( n3432 & n21436 ) | ( n14677 & n21436 ) ;
  assign n24453 = n24452 ^ n5121 ^ n3971 ;
  assign n24454 = ( n883 & ~n6229 ) | ( n883 & n7814 ) | ( ~n6229 & n7814 ) ;
  assign n24455 = n17046 ^ n8882 ^ n2786 ;
  assign n24456 = n24455 ^ n23780 ^ n4916 ;
  assign n24457 = n24456 ^ n22114 ^ n16408 ;
  assign n24458 = ( ~n6615 & n6950 ) | ( ~n6615 & n24457 ) | ( n6950 & n24457 ) ;
  assign n24459 = ( n8484 & n9199 ) | ( n8484 & n11141 ) | ( n9199 & n11141 ) ;
  assign n24460 = n20841 ^ n3278 ^ n2659 ;
  assign n24461 = n24460 ^ n19804 ^ n11946 ;
  assign n24462 = ( n5196 & ~n24459 ) | ( n5196 & n24461 ) | ( ~n24459 & n24461 ) ;
  assign n24463 = ( n473 & n24458 ) | ( n473 & ~n24462 ) | ( n24458 & ~n24462 ) ;
  assign n24464 = ( n20707 & ~n24454 ) | ( n20707 & n24463 ) | ( ~n24454 & n24463 ) ;
  assign n24465 = n941 & n2691 ;
  assign n24466 = n24465 ^ n1187 ^ 1'b0 ;
  assign n24467 = n18753 ^ n1522 ^ 1'b0 ;
  assign n24468 = ( n7054 & n13190 ) | ( n7054 & n24467 ) | ( n13190 & n24467 ) ;
  assign n24469 = ( n1746 & n6947 ) | ( n1746 & ~n24468 ) | ( n6947 & ~n24468 ) ;
  assign n24470 = n24469 ^ n18251 ^ n6044 ;
  assign n24471 = ( n13173 & ~n24466 ) | ( n13173 & n24470 ) | ( ~n24466 & n24470 ) ;
  assign n24473 = n22461 ^ n2330 ^ 1'b0 ;
  assign n24472 = ~n6063 & n22109 ;
  assign n24474 = n24473 ^ n24472 ^ 1'b0 ;
  assign n24475 = ( n19164 & ~n20995 ) | ( n19164 & n24474 ) | ( ~n20995 & n24474 ) ;
  assign n24476 = ( n2261 & ~n20923 ) | ( n2261 & n24475 ) | ( ~n20923 & n24475 ) ;
  assign n24477 = ( n1968 & ~n5618 ) | ( n1968 & n24476 ) | ( ~n5618 & n24476 ) ;
  assign n24478 = n8725 ^ x157 ^ 1'b0 ;
  assign n24479 = ( ~n7446 & n12494 ) | ( ~n7446 & n24478 ) | ( n12494 & n24478 ) ;
  assign n24480 = ( n7800 & ~n8877 ) | ( n7800 & n14205 ) | ( ~n8877 & n14205 ) ;
  assign n24481 = n1863 ^ n1420 ^ 1'b0 ;
  assign n24482 = n10228 ^ n5913 ^ n4129 ;
  assign n24483 = n24482 ^ n21426 ^ n851 ;
  assign n24484 = n23341 ^ n14949 ^ 1'b0 ;
  assign n24485 = ~n3883 & n5968 ;
  assign n24486 = ~n24484 & n24485 ;
  assign n24487 = n11306 ^ n6626 ^ n387 ;
  assign n24488 = ( ~n3346 & n18361 ) | ( ~n3346 & n24487 ) | ( n18361 & n24487 ) ;
  assign n24489 = ( ~n5723 & n20594 ) | ( ~n5723 & n24488 ) | ( n20594 & n24488 ) ;
  assign n24490 = n24489 ^ n6251 ^ 1'b0 ;
  assign n24491 = n6378 | n24490 ;
  assign n24495 = n3610 ^ n3047 ^ n1576 ;
  assign n24496 = ( ~n5901 & n9888 ) | ( ~n5901 & n24495 ) | ( n9888 & n24495 ) ;
  assign n24492 = n16653 ^ n11201 ^ n4741 ;
  assign n24493 = n16300 ^ n14628 ^ n4493 ;
  assign n24494 = n24492 & n24493 ;
  assign n24497 = n24496 ^ n24494 ^ 1'b0 ;
  assign n24498 = ( ~n1355 & n11101 ) | ( ~n1355 & n18389 ) | ( n11101 & n18389 ) ;
  assign n24499 = ( n7502 & n20101 ) | ( n7502 & n24498 ) | ( n20101 & n24498 ) ;
  assign n24500 = ( n4958 & n8603 ) | ( n4958 & ~n24499 ) | ( n8603 & ~n24499 ) ;
  assign n24501 = ( n6772 & n8121 ) | ( n6772 & ~n24500 ) | ( n8121 & ~n24500 ) ;
  assign n24502 = n24501 ^ n21025 ^ n8033 ;
  assign n24503 = ( n11538 & ~n24384 ) | ( n11538 & n24502 ) | ( ~n24384 & n24502 ) ;
  assign n24504 = n22772 & n24503 ;
  assign n24505 = n24497 & n24504 ;
  assign n24506 = ( n5148 & n5332 ) | ( n5148 & ~n14101 ) | ( n5332 & ~n14101 ) ;
  assign n24507 = n20933 ^ n16998 ^ n2934 ;
  assign n24508 = ( ~n8066 & n24506 ) | ( ~n8066 & n24507 ) | ( n24506 & n24507 ) ;
  assign n24509 = ( ~n12418 & n14204 ) | ( ~n12418 & n24508 ) | ( n14204 & n24508 ) ;
  assign n24510 = ( ~n17088 & n21402 ) | ( ~n17088 & n23101 ) | ( n21402 & n23101 ) ;
  assign n24511 = ( n386 & ~n7066 ) | ( n386 & n15897 ) | ( ~n7066 & n15897 ) ;
  assign n24512 = n24511 ^ n22313 ^ n19194 ;
  assign n24516 = n17015 ^ n16814 ^ n4525 ;
  assign n24514 = n13353 ^ n12210 ^ n6324 ;
  assign n24515 = ~n5449 & n24514 ;
  assign n24517 = n24516 ^ n24515 ^ 1'b0 ;
  assign n24513 = ( n6422 & n12489 ) | ( n6422 & n21624 ) | ( n12489 & n21624 ) ;
  assign n24518 = n24517 ^ n24513 ^ n13648 ;
  assign n24528 = ( n10772 & ~n11757 ) | ( n10772 & n13822 ) | ( ~n11757 & n13822 ) ;
  assign n24526 = n21801 ^ n493 ^ 1'b0 ;
  assign n24527 = n21784 & ~n24526 ;
  assign n24519 = n8588 | n21640 ;
  assign n24522 = n21871 ^ n13874 ^ x239 ;
  assign n24520 = n9730 & ~n13936 ;
  assign n24521 = n2355 & n24520 ;
  assign n24523 = n24522 ^ n24521 ^ n9988 ;
  assign n24524 = n24523 ^ n11045 ^ n9095 ;
  assign n24525 = ( ~n13729 & n24519 ) | ( ~n13729 & n24524 ) | ( n24519 & n24524 ) ;
  assign n24529 = n24528 ^ n24527 ^ n24525 ;
  assign n24530 = n20650 ^ n9640 ^ n2893 ;
  assign n24539 = n5929 ^ n4715 ^ n3553 ;
  assign n24538 = n7775 ^ n2498 ^ n484 ;
  assign n24540 = n24539 ^ n24538 ^ n15356 ;
  assign n24541 = ( n9032 & ~n15430 ) | ( n9032 & n24540 ) | ( ~n15430 & n24540 ) ;
  assign n24531 = n12327 ^ n9854 ^ n7150 ;
  assign n24532 = n18237 ^ n8188 ^ 1'b0 ;
  assign n24533 = n21834 | n24532 ;
  assign n24534 = ( n3833 & n6067 ) | ( n3833 & n24533 ) | ( n6067 & n24533 ) ;
  assign n24535 = n11765 | n19577 ;
  assign n24536 = n24534 & ~n24535 ;
  assign n24537 = ( n13643 & ~n24531 ) | ( n13643 & n24536 ) | ( ~n24531 & n24536 ) ;
  assign n24542 = n24541 ^ n24537 ^ 1'b0 ;
  assign n24543 = n17996 ^ n12466 ^ n7173 ;
  assign n24544 = n17431 ^ n14680 ^ n5297 ;
  assign n24545 = ( n297 & n24543 ) | ( n297 & ~n24544 ) | ( n24543 & ~n24544 ) ;
  assign n24546 = n1345 ^ n989 ^ 1'b0 ;
  assign n24547 = ~n870 & n24546 ;
  assign n24548 = ( n1726 & n19272 ) | ( n1726 & n24547 ) | ( n19272 & n24547 ) ;
  assign n24549 = n13983 ^ n11077 ^ n6018 ;
  assign n24550 = n24549 ^ n8033 ^ n6736 ;
  assign n24551 = n9924 ^ n967 ^ 1'b0 ;
  assign n24552 = ( n24548 & ~n24550 ) | ( n24548 & n24551 ) | ( ~n24550 & n24551 ) ;
  assign n24563 = n11553 ^ n2157 ^ x50 ;
  assign n24560 = n1063 & n1314 ;
  assign n24561 = n24560 ^ n857 ^ 1'b0 ;
  assign n24562 = n24561 ^ n19274 ^ n3912 ;
  assign n24553 = ~n1439 & n1989 ;
  assign n24554 = n24553 ^ n883 ^ 1'b0 ;
  assign n24555 = ( n12840 & ~n15373 ) | ( n12840 & n24554 ) | ( ~n15373 & n24554 ) ;
  assign n24556 = n12338 & ~n24555 ;
  assign n24557 = n21300 & n24556 ;
  assign n24558 = ( n1402 & ~n15122 ) | ( n1402 & n17967 ) | ( ~n15122 & n17967 ) ;
  assign n24559 = ( n9860 & n24557 ) | ( n9860 & ~n24558 ) | ( n24557 & ~n24558 ) ;
  assign n24564 = n24563 ^ n24562 ^ n24559 ;
  assign n24565 = n13141 ^ n8660 ^ n1119 ;
  assign n24566 = ( n893 & n7556 ) | ( n893 & n24565 ) | ( n7556 & n24565 ) ;
  assign n24567 = n13718 ^ n8702 ^ n5347 ;
  assign n24568 = n24567 ^ n10033 ^ n9311 ;
  assign n24569 = n11006 ^ n10181 ^ n1145 ;
  assign n24570 = ( n5132 & n20843 ) | ( n5132 & ~n24569 ) | ( n20843 & ~n24569 ) ;
  assign n24571 = ( n24566 & n24568 ) | ( n24566 & ~n24570 ) | ( n24568 & ~n24570 ) ;
  assign n24574 = ( n4694 & ~n4852 ) | ( n4694 & n14541 ) | ( ~n4852 & n14541 ) ;
  assign n24572 = n11726 ^ n10663 ^ 1'b0 ;
  assign n24573 = ~n1319 & n24572 ;
  assign n24575 = n24574 ^ n24573 ^ n8853 ;
  assign n24576 = n24575 ^ n20249 ^ n11217 ;
  assign n24577 = ( n16076 & ~n24571 ) | ( n16076 & n24576 ) | ( ~n24571 & n24576 ) ;
  assign n24578 = ( ~n20488 & n20490 ) | ( ~n20488 & n24577 ) | ( n20490 & n24577 ) ;
  assign n24582 = n13054 & ~n14430 ;
  assign n24579 = n1522 ^ x169 ^ x149 ;
  assign n24580 = n19281 ^ n9258 ^ n2302 ;
  assign n24581 = n24579 | n24580 ;
  assign n24583 = n24582 ^ n24581 ^ 1'b0 ;
  assign n24592 = n10464 ^ n8818 ^ n903 ;
  assign n24589 = ( n13152 & n13493 ) | ( n13152 & n21260 ) | ( n13493 & n21260 ) ;
  assign n24590 = n24589 ^ n21365 ^ n9384 ;
  assign n24591 = ( ~n2712 & n12366 ) | ( ~n2712 & n24590 ) | ( n12366 & n24590 ) ;
  assign n24593 = n24592 ^ n24591 ^ n22978 ;
  assign n24594 = n24593 ^ n7508 ^ n3712 ;
  assign n24584 = n16866 & ~n17931 ;
  assign n24585 = ~n18799 & n24584 ;
  assign n24586 = ( n4529 & n22515 ) | ( n4529 & ~n24585 ) | ( n22515 & ~n24585 ) ;
  assign n24587 = n23615 ^ n8616 ^ n2323 ;
  assign n24588 = n24586 & ~n24587 ;
  assign n24595 = n24594 ^ n24588 ^ 1'b0 ;
  assign n24596 = ( ~n6733 & n10975 ) | ( ~n6733 & n20823 ) | ( n10975 & n20823 ) ;
  assign n24597 = ( n15582 & ~n17405 ) | ( n15582 & n24596 ) | ( ~n17405 & n24596 ) ;
  assign n24598 = n9066 ^ n7625 ^ n4307 ;
  assign n24599 = ~n4189 & n14689 ;
  assign n24605 = n8550 ^ n3371 ^ n806 ;
  assign n24600 = n5780 & ~n13906 ;
  assign n24601 = n24600 ^ n1449 ^ 1'b0 ;
  assign n24602 = ( n1856 & n5918 ) | ( n1856 & ~n24601 ) | ( n5918 & ~n24601 ) ;
  assign n24603 = n23057 & ~n24602 ;
  assign n24604 = n21265 & n24603 ;
  assign n24606 = n24605 ^ n24604 ^ n7897 ;
  assign n24607 = n24606 ^ n11078 ^ n2021 ;
  assign n24608 = ~n9949 & n17253 ;
  assign n24609 = n4154 & n6435 ;
  assign n24610 = n24609 ^ n9232 ^ 1'b0 ;
  assign n24611 = ( n4428 & n12483 ) | ( n4428 & ~n19483 ) | ( n12483 & ~n19483 ) ;
  assign n24612 = n12159 | n21471 ;
  assign n24613 = ( n15522 & ~n24611 ) | ( n15522 & n24612 ) | ( ~n24611 & n24612 ) ;
  assign n24614 = ( ~n7205 & n24610 ) | ( ~n7205 & n24613 ) | ( n24610 & n24613 ) ;
  assign n24615 = n14997 ^ n631 ^ 1'b0 ;
  assign n24616 = n24615 ^ n11048 ^ n5256 ;
  assign n24617 = ( n10494 & n16571 ) | ( n10494 & n24616 ) | ( n16571 & n24616 ) ;
  assign n24618 = n8396 ^ n7754 ^ 1'b0 ;
  assign n24619 = n21550 ^ n18913 ^ n16168 ;
  assign n24620 = n16932 | n24455 ;
  assign n24621 = n24620 ^ n14113 ^ n13955 ;
  assign n24622 = n2403 ^ n1030 ^ 1'b0 ;
  assign n24623 = n15326 | n24622 ;
  assign n24624 = n3896 & n15974 ;
  assign n24625 = n24624 ^ n16104 ^ 1'b0 ;
  assign n24626 = ~n9750 & n24625 ;
  assign n24627 = ( n3641 & ~n17849 ) | ( n3641 & n18096 ) | ( ~n17849 & n18096 ) ;
  assign n24628 = n12001 | n24627 ;
  assign n24629 = ( n2160 & ~n13999 ) | ( n2160 & n24628 ) | ( ~n13999 & n24628 ) ;
  assign n24630 = ( n19565 & n24626 ) | ( n19565 & n24629 ) | ( n24626 & n24629 ) ;
  assign n24631 = n8058 ^ n1536 ^ 1'b0 ;
  assign n24632 = n24631 ^ n13182 ^ 1'b0 ;
  assign n24633 = ( n444 & n6396 ) | ( n444 & ~n11750 ) | ( n6396 & ~n11750 ) ;
  assign n24635 = n17651 ^ n14835 ^ n2017 ;
  assign n24634 = ( ~n13740 & n14765 ) | ( ~n13740 & n17371 ) | ( n14765 & n17371 ) ;
  assign n24636 = n24635 ^ n24634 ^ n11914 ;
  assign n24637 = ( n4339 & ~n22955 ) | ( n4339 & n24636 ) | ( ~n22955 & n24636 ) ;
  assign n24638 = ( n9133 & n24633 ) | ( n9133 & n24637 ) | ( n24633 & n24637 ) ;
  assign n24639 = n19486 ^ n17948 ^ n6355 ;
  assign n24640 = n24435 ^ n21428 ^ n11429 ;
  assign n24641 = n20401 ^ n5458 ^ n529 ;
  assign n24642 = n24641 ^ n17282 ^ n6106 ;
  assign n24643 = ( n19062 & ~n23020 ) | ( n19062 & n24642 ) | ( ~n23020 & n24642 ) ;
  assign n24644 = ( n10712 & ~n24640 ) | ( n10712 & n24643 ) | ( ~n24640 & n24643 ) ;
  assign n24645 = n1482 & ~n2336 ;
  assign n24646 = ~n4665 & n24645 ;
  assign n24647 = n10076 ^ n9336 ^ n5741 ;
  assign n24648 = ( n5655 & n22994 ) | ( n5655 & ~n24647 ) | ( n22994 & ~n24647 ) ;
  assign n24655 = n16960 ^ n4640 ^ n2489 ;
  assign n24649 = n14089 ^ n6078 ^ n1760 ;
  assign n24650 = n21206 & n24649 ;
  assign n24651 = n24650 ^ n11128 ^ 1'b0 ;
  assign n24652 = n15271 & n24651 ;
  assign n24653 = n24652 ^ n10913 ^ 1'b0 ;
  assign n24654 = n24653 ^ n7039 ^ n6947 ;
  assign n24656 = n24655 ^ n24654 ^ n11020 ;
  assign n24660 = ( ~n691 & n3141 ) | ( ~n691 & n3217 ) | ( n3141 & n3217 ) ;
  assign n24661 = n24660 ^ n11149 ^ n10508 ;
  assign n24657 = n11052 ^ n2290 ^ n899 ;
  assign n24658 = ( ~n3683 & n11353 ) | ( ~n3683 & n24657 ) | ( n11353 & n24657 ) ;
  assign n24659 = n24658 ^ n8899 ^ 1'b0 ;
  assign n24662 = n24661 ^ n24659 ^ n21323 ;
  assign n24663 = n23962 ^ n22452 ^ n10899 ;
  assign n24664 = n24663 ^ n9339 ^ 1'b0 ;
  assign n24665 = n9786 | n21035 ;
  assign n24666 = n24665 ^ n5905 ^ 1'b0 ;
  assign n24667 = ( ~n18139 & n18230 ) | ( ~n18139 & n24666 ) | ( n18230 & n24666 ) ;
  assign n24668 = n24667 ^ n17348 ^ 1'b0 ;
  assign n24669 = n24668 ^ n21183 ^ 1'b0 ;
  assign n24670 = n16577 ^ n13201 ^ n5533 ;
  assign n24671 = ( n1246 & n1936 ) | ( n1246 & ~n14243 ) | ( n1936 & ~n14243 ) ;
  assign n24675 = n11204 ^ n7945 ^ n7381 ;
  assign n24676 = n951 | n1756 ;
  assign n24677 = n409 & ~n24676 ;
  assign n24678 = n24675 & ~n24677 ;
  assign n24679 = n13906 & n24678 ;
  assign n24672 = n14502 ^ n3886 ^ n1538 ;
  assign n24673 = n4915 | n17967 ;
  assign n24674 = ( n5279 & n24672 ) | ( n5279 & ~n24673 ) | ( n24672 & ~n24673 ) ;
  assign n24680 = n24679 ^ n24674 ^ n1081 ;
  assign n24681 = n15602 & n24680 ;
  assign n24682 = n24681 ^ n22248 ^ 1'b0 ;
  assign n24683 = ( ~n1906 & n24671 ) | ( ~n1906 & n24682 ) | ( n24671 & n24682 ) ;
  assign n24684 = ( ~n5584 & n12665 ) | ( ~n5584 & n17313 ) | ( n12665 & n17313 ) ;
  assign n24685 = n24684 ^ n15854 ^ n9579 ;
  assign n24686 = ( ~x97 & n9420 ) | ( ~x97 & n13907 ) | ( n9420 & n13907 ) ;
  assign n24687 = ~n1868 & n5742 ;
  assign n24688 = n24687 ^ n1009 ^ 1'b0 ;
  assign n24689 = n24005 & n24688 ;
  assign n24690 = n23017 ^ n8674 ^ 1'b0 ;
  assign n24691 = n20451 ^ n14506 ^ n2098 ;
  assign n24692 = n24691 ^ n19086 ^ n1620 ;
  assign n24693 = ( n1663 & ~n13427 ) | ( n1663 & n16001 ) | ( ~n13427 & n16001 ) ;
  assign n24694 = n24693 ^ n15573 ^ 1'b0 ;
  assign n24695 = ( n318 & n6716 ) | ( n318 & n24694 ) | ( n6716 & n24694 ) ;
  assign n24697 = n5689 ^ n1680 ^ n865 ;
  assign n24698 = ( n1383 & ~n5082 ) | ( n1383 & n24697 ) | ( ~n5082 & n24697 ) ;
  assign n24699 = ( x5 & ~n21266 ) | ( x5 & n24698 ) | ( ~n21266 & n24698 ) ;
  assign n24696 = ( n1246 & n4640 ) | ( n1246 & n13394 ) | ( n4640 & n13394 ) ;
  assign n24700 = n24699 ^ n24696 ^ 1'b0 ;
  assign n24701 = ( n14061 & n16714 ) | ( n14061 & n21180 ) | ( n16714 & n21180 ) ;
  assign n24702 = n24701 ^ n13020 ^ 1'b0 ;
  assign n24703 = n24700 | n24702 ;
  assign n24704 = ( ~n8421 & n15506 ) | ( ~n8421 & n21082 ) | ( n15506 & n21082 ) ;
  assign n24705 = ( ~n1490 & n1808 ) | ( ~n1490 & n5987 ) | ( n1808 & n5987 ) ;
  assign n24713 = ( ~n6205 & n8119 ) | ( ~n6205 & n20650 ) | ( n8119 & n20650 ) ;
  assign n24711 = n4905 | n8850 ;
  assign n24712 = ( ~n17657 & n18538 ) | ( ~n17657 & n24711 ) | ( n18538 & n24711 ) ;
  assign n24709 = ( n6741 & ~n11322 ) | ( n6741 & n19286 ) | ( ~n11322 & n19286 ) ;
  assign n24706 = n6922 ^ n5214 ^ n1859 ;
  assign n24707 = n19092 ^ n3807 ^ 1'b0 ;
  assign n24708 = n24706 & n24707 ;
  assign n24710 = n24709 ^ n24708 ^ n23190 ;
  assign n24714 = n24713 ^ n24712 ^ n24710 ;
  assign n24715 = ( n15447 & ~n24705 ) | ( n15447 & n24714 ) | ( ~n24705 & n24714 ) ;
  assign n24716 = ( n14150 & n24704 ) | ( n14150 & ~n24715 ) | ( n24704 & ~n24715 ) ;
  assign n24717 = ( n335 & n342 ) | ( n335 & n4260 ) | ( n342 & n4260 ) ;
  assign n24718 = ( ~n556 & n8998 ) | ( ~n556 & n10403 ) | ( n8998 & n10403 ) ;
  assign n24719 = ( n1529 & n24717 ) | ( n1529 & ~n24718 ) | ( n24717 & ~n24718 ) ;
  assign n24722 = n7563 ^ n5647 ^ n5098 ;
  assign n24720 = ~n9180 & n22651 ;
  assign n24721 = n24720 ^ n13473 ^ n2041 ;
  assign n24723 = n24722 ^ n24721 ^ n21635 ;
  assign n24724 = n18904 & n24723 ;
  assign n24726 = n18158 ^ n14764 ^ n2432 ;
  assign n24727 = ( n8116 & n20770 ) | ( n8116 & ~n24726 ) | ( n20770 & ~n24726 ) ;
  assign n24725 = ~n8969 & n22063 ;
  assign n24728 = n24727 ^ n24725 ^ n2885 ;
  assign n24729 = n24728 ^ n2879 ^ n796 ;
  assign n24730 = ( n384 & ~n1904 ) | ( n384 & n18690 ) | ( ~n1904 & n18690 ) ;
  assign n24731 = ( n8899 & n9498 ) | ( n8899 & ~n24730 ) | ( n9498 & ~n24730 ) ;
  assign n24732 = n21265 & ~n24731 ;
  assign n24733 = ( n1056 & ~n6551 ) | ( n1056 & n14954 ) | ( ~n6551 & n14954 ) ;
  assign n24734 = n24733 ^ n13300 ^ n4696 ;
  assign n24735 = ( ~n3666 & n19532 ) | ( ~n3666 & n24734 ) | ( n19532 & n24734 ) ;
  assign n24736 = ( n7635 & ~n24732 ) | ( n7635 & n24735 ) | ( ~n24732 & n24735 ) ;
  assign n24737 = n24736 ^ n15876 ^ n10142 ;
  assign n24738 = n20302 ^ n11338 ^ n550 ;
  assign n24739 = ( n4156 & n6939 ) | ( n4156 & n19054 ) | ( n6939 & n19054 ) ;
  assign n24740 = n24739 ^ n24723 ^ n13954 ;
  assign n24741 = ( ~n720 & n24738 ) | ( ~n720 & n24740 ) | ( n24738 & n24740 ) ;
  assign n24742 = n12098 ^ n5037 ^ n3025 ;
  assign n24743 = ( n5308 & ~n7154 ) | ( n5308 & n20084 ) | ( ~n7154 & n20084 ) ;
  assign n24744 = ( n20506 & n24742 ) | ( n20506 & ~n24743 ) | ( n24742 & ~n24743 ) ;
  assign n24745 = n6631 ^ n1407 ^ 1'b0 ;
  assign n24746 = n24744 & ~n24745 ;
  assign n24747 = ( n8574 & ~n14939 ) | ( n8574 & n24746 ) | ( ~n14939 & n24746 ) ;
  assign n24748 = n5456 & ~n17019 ;
  assign n24749 = n24748 ^ n4722 ^ 1'b0 ;
  assign n24750 = n24749 ^ n18280 ^ n4656 ;
  assign n24751 = n1671 & ~n10949 ;
  assign n24752 = n24751 ^ n17503 ^ n4890 ;
  assign n24753 = n24752 ^ n21482 ^ n16636 ;
  assign n24754 = n1577 | n24753 ;
  assign n24755 = n24754 ^ n22847 ^ 1'b0 ;
  assign n24756 = n9479 ^ n9105 ^ n7470 ;
  assign n24757 = n24756 ^ n20047 ^ n2183 ;
  assign n24758 = n10345 & ~n20661 ;
  assign n24759 = n24758 ^ n11700 ^ 1'b0 ;
  assign n24760 = n24759 ^ n11010 ^ n5816 ;
  assign n24761 = n24760 ^ n6493 ^ n4714 ;
  assign n24762 = ( n13043 & n16021 ) | ( n13043 & ~n21511 ) | ( n16021 & ~n21511 ) ;
  assign n24763 = ( n3894 & n4011 ) | ( n3894 & n24762 ) | ( n4011 & n24762 ) ;
  assign n24764 = n19683 ^ n12456 ^ x108 ;
  assign n24767 = ( n1180 & n7430 ) | ( n1180 & n12633 ) | ( n7430 & n12633 ) ;
  assign n24765 = n22435 ^ n16991 ^ n8237 ;
  assign n24766 = ~n21702 & n24765 ;
  assign n24768 = n24767 ^ n24766 ^ 1'b0 ;
  assign n24769 = ~n22751 & n24768 ;
  assign n24770 = n24764 & n24769 ;
  assign n24773 = ( n3457 & ~n11029 ) | ( n3457 & n20002 ) | ( ~n11029 & n20002 ) ;
  assign n24771 = n23273 ^ n21547 ^ n10712 ;
  assign n24772 = ( n736 & n6803 ) | ( n736 & n24771 ) | ( n6803 & n24771 ) ;
  assign n24774 = n24773 ^ n24772 ^ n299 ;
  assign n24777 = n6453 & n18115 ;
  assign n24778 = n24777 ^ n1357 ^ 1'b0 ;
  assign n24775 = n7952 ^ n4086 ^ 1'b0 ;
  assign n24776 = n22641 & ~n24775 ;
  assign n24779 = n24778 ^ n24776 ^ n1722 ;
  assign n24780 = n24779 ^ n18746 ^ 1'b0 ;
  assign n24781 = n12274 ^ n1166 ^ 1'b0 ;
  assign n24782 = n24781 ^ n17830 ^ n5460 ;
  assign n24783 = ( n1729 & n7513 ) | ( n1729 & ~n8534 ) | ( n7513 & ~n8534 ) ;
  assign n24784 = ( ~n12837 & n15341 ) | ( ~n12837 & n24783 ) | ( n15341 & n24783 ) ;
  assign n24785 = n24782 & n24784 ;
  assign n24786 = ~n1464 & n24785 ;
  assign n24787 = n12383 ^ n10885 ^ n8554 ;
  assign n24788 = n8616 ^ n1741 ^ n1148 ;
  assign n24792 = ~n1072 & n2252 ;
  assign n24793 = ~n10152 & n24792 ;
  assign n24794 = n24793 ^ n3914 ^ n2957 ;
  assign n24789 = ( n9713 & ~n15557 ) | ( n9713 & n19618 ) | ( ~n15557 & n19618 ) ;
  assign n24790 = ( n5760 & n10839 ) | ( n5760 & n24789 ) | ( n10839 & n24789 ) ;
  assign n24791 = n24790 ^ x40 ^ 1'b0 ;
  assign n24795 = n24794 ^ n24791 ^ n9652 ;
  assign n24796 = n21032 ^ n1421 ^ 1'b0 ;
  assign n24797 = n6470 & ~n24796 ;
  assign n24798 = ( n995 & n2725 ) | ( n995 & ~n9951 ) | ( n2725 & ~n9951 ) ;
  assign n24799 = n1795 & n11223 ;
  assign n24800 = ( n12041 & n16060 ) | ( n12041 & n24799 ) | ( n16060 & n24799 ) ;
  assign n24801 = n24798 & n24800 ;
  assign n24802 = n24797 & ~n24801 ;
  assign n24803 = ( x241 & ~n12804 ) | ( x241 & n16518 ) | ( ~n12804 & n16518 ) ;
  assign n24804 = ( ~n8750 & n20939 ) | ( ~n8750 & n24803 ) | ( n20939 & n24803 ) ;
  assign n24805 = n24804 ^ n5310 ^ n4367 ;
  assign n24806 = ( n4861 & n13933 ) | ( n4861 & n23132 ) | ( n13933 & n23132 ) ;
  assign n24807 = n16481 ^ n15937 ^ n6202 ;
  assign n24808 = ( n8685 & n13360 ) | ( n8685 & n24807 ) | ( n13360 & n24807 ) ;
  assign n24809 = ( n3223 & ~n17069 ) | ( n3223 & n24701 ) | ( ~n17069 & n24701 ) ;
  assign n24810 = n24809 ^ n16245 ^ n2943 ;
  assign n24811 = ( ~n5317 & n8821 ) | ( ~n5317 & n24810 ) | ( n8821 & n24810 ) ;
  assign n24812 = ( ~n3040 & n5000 ) | ( ~n3040 & n13390 ) | ( n5000 & n13390 ) ;
  assign n24813 = n24812 ^ n18436 ^ n7651 ;
  assign n24815 = n19320 ^ n2508 ^ 1'b0 ;
  assign n24816 = ( n6801 & n10286 ) | ( n6801 & n24815 ) | ( n10286 & n24815 ) ;
  assign n24814 = ( n477 & n1265 ) | ( n477 & ~n2118 ) | ( n1265 & ~n2118 ) ;
  assign n24817 = n24816 ^ n24814 ^ n9419 ;
  assign n24818 = n5515 ^ n534 ^ n287 ;
  assign n24819 = ( n1745 & n6758 ) | ( n1745 & n20961 ) | ( n6758 & n20961 ) ;
  assign n24820 = ( n1326 & ~n18902 ) | ( n1326 & n24819 ) | ( ~n18902 & n24819 ) ;
  assign n24821 = ( ~n24649 & n24818 ) | ( ~n24649 & n24820 ) | ( n24818 & n24820 ) ;
  assign n24822 = ( n12655 & ~n24817 ) | ( n12655 & n24821 ) | ( ~n24817 & n24821 ) ;
  assign n24823 = n23583 ^ n18544 ^ 1'b0 ;
  assign n24824 = n18707 & n24823 ;
  assign n24825 = n7757 ^ n3727 ^ n2098 ;
  assign n24830 = ( n692 & n14503 ) | ( n692 & n24165 ) | ( n14503 & n24165 ) ;
  assign n24826 = n12994 ^ n5402 ^ n4118 ;
  assign n24827 = ~n11221 & n24826 ;
  assign n24828 = ( n13141 & n13808 ) | ( n13141 & ~n24827 ) | ( n13808 & ~n24827 ) ;
  assign n24829 = ( n4077 & n17535 ) | ( n4077 & ~n24828 ) | ( n17535 & ~n24828 ) ;
  assign n24831 = n24830 ^ n24829 ^ n8989 ;
  assign n24832 = n23840 ^ n9121 ^ n5145 ;
  assign n24833 = ( n757 & ~n1122 ) | ( n757 & n11850 ) | ( ~n1122 & n11850 ) ;
  assign n24834 = ( n20585 & ~n24832 ) | ( n20585 & n24833 ) | ( ~n24832 & n24833 ) ;
  assign n24835 = ( n16142 & n20627 ) | ( n16142 & ~n24834 ) | ( n20627 & ~n24834 ) ;
  assign n24836 = n2140 | n24835 ;
  assign n24837 = ( n485 & ~n2869 ) | ( n485 & n14748 ) | ( ~n2869 & n14748 ) ;
  assign n24838 = n24837 ^ n14854 ^ 1'b0 ;
  assign n24839 = n16995 ^ n16827 ^ n11016 ;
  assign n24840 = n19122 ^ n14716 ^ 1'b0 ;
  assign n24841 = n24839 & ~n24840 ;
  assign n24842 = n21466 ^ n15736 ^ n3075 ;
  assign n24843 = n8597 ^ n2840 ^ n577 ;
  assign n24844 = n10932 | n24843 ;
  assign n24845 = n7018 | n24844 ;
  assign n24846 = ( n4061 & n5316 ) | ( n4061 & n24845 ) | ( n5316 & n24845 ) ;
  assign n24849 = n16653 ^ n4374 ^ 1'b0 ;
  assign n24850 = ( ~n1960 & n5285 ) | ( ~n1960 & n14436 ) | ( n5285 & n14436 ) ;
  assign n24851 = ( ~n1992 & n5277 ) | ( ~n1992 & n24850 ) | ( n5277 & n24850 ) ;
  assign n24852 = ~n24849 & n24851 ;
  assign n24847 = n14692 ^ n3530 ^ n2372 ;
  assign n24848 = ( n8590 & n14874 ) | ( n8590 & ~n24847 ) | ( n14874 & ~n24847 ) ;
  assign n24853 = n24852 ^ n24848 ^ n17604 ;
  assign n24854 = n24853 ^ n9964 ^ n1344 ;
  assign n24855 = ( ~n12542 & n15151 ) | ( ~n12542 & n24854 ) | ( n15151 & n24854 ) ;
  assign n24856 = n24108 ^ n8320 ^ n5716 ;
  assign n24857 = n20744 ^ n12717 ^ n7123 ;
  assign n24858 = ( n13539 & n24856 ) | ( n13539 & n24857 ) | ( n24856 & n24857 ) ;
  assign n24859 = ( n11408 & ~n16466 ) | ( n11408 & n24858 ) | ( ~n16466 & n24858 ) ;
  assign n24860 = ( ~n9414 & n11056 ) | ( ~n9414 & n14853 ) | ( n11056 & n14853 ) ;
  assign n24861 = ( ~n11465 & n24506 ) | ( ~n11465 & n24860 ) | ( n24506 & n24860 ) ;
  assign n24862 = ( ~n6309 & n6861 ) | ( ~n6309 & n24861 ) | ( n6861 & n24861 ) ;
  assign n24863 = ( n14031 & n19295 ) | ( n14031 & n24862 ) | ( n19295 & n24862 ) ;
  assign n24864 = n5754 ^ n3307 ^ 1'b0 ;
  assign n24865 = n7623 ^ n1552 ^ n636 ;
  assign n24866 = ( n12942 & n24864 ) | ( n12942 & n24865 ) | ( n24864 & n24865 ) ;
  assign n24869 = n3826 ^ n1322 ^ n747 ;
  assign n24867 = n21554 ^ n19068 ^ n4849 ;
  assign n24868 = ( x99 & n6691 ) | ( x99 & n24867 ) | ( n6691 & n24867 ) ;
  assign n24870 = n24869 ^ n24868 ^ n11958 ;
  assign n24871 = n24845 ^ n16296 ^ n8035 ;
  assign n24872 = ( n1653 & ~n3809 ) | ( n1653 & n4165 ) | ( ~n3809 & n4165 ) ;
  assign n24873 = ( ~n16168 & n17458 ) | ( ~n16168 & n24872 ) | ( n17458 & n24872 ) ;
  assign n24874 = ( n16369 & n24871 ) | ( n16369 & n24873 ) | ( n24871 & n24873 ) ;
  assign n24875 = ( n1104 & n14699 ) | ( n1104 & ~n21132 ) | ( n14699 & ~n21132 ) ;
  assign n24876 = ( ~n4294 & n16441 ) | ( ~n4294 & n24565 ) | ( n16441 & n24565 ) ;
  assign n24877 = n24876 ^ n17460 ^ n15570 ;
  assign n24878 = ( n309 & n866 ) | ( n309 & n5662 ) | ( n866 & n5662 ) ;
  assign n24879 = ( n9618 & ~n18818 ) | ( n9618 & n24878 ) | ( ~n18818 & n24878 ) ;
  assign n24880 = n15141 ^ n14905 ^ 1'b0 ;
  assign n24881 = n19354 | n24880 ;
  assign n24882 = n24881 ^ n21424 ^ 1'b0 ;
  assign n24883 = n24882 ^ n15028 ^ n11695 ;
  assign n24884 = n7442 & ~n18960 ;
  assign n24885 = n9370 & n24884 ;
  assign n24886 = ( n11646 & ~n23360 ) | ( n11646 & n24885 ) | ( ~n23360 & n24885 ) ;
  assign n24887 = ( n8577 & n9504 ) | ( n8577 & ~n9539 ) | ( n9504 & ~n9539 ) ;
  assign n24888 = ( ~n8812 & n19887 ) | ( ~n8812 & n24887 ) | ( n19887 & n24887 ) ;
  assign n24889 = n24888 ^ n22924 ^ n9070 ;
  assign n24890 = ( n1628 & n7641 ) | ( n1628 & n16874 ) | ( n7641 & n16874 ) ;
  assign n24891 = ( x240 & ~n2484 ) | ( x240 & n17740 ) | ( ~n2484 & n17740 ) ;
  assign n24892 = ( n6987 & ~n11795 ) | ( n6987 & n15150 ) | ( ~n11795 & n15150 ) ;
  assign n24893 = ( n20598 & n24891 ) | ( n20598 & ~n24892 ) | ( n24891 & ~n24892 ) ;
  assign n24894 = ~n21531 & n24893 ;
  assign n24895 = n13581 ^ n9692 ^ n263 ;
  assign n24896 = n24895 ^ n11030 ^ n5730 ;
  assign n24897 = n14972 ^ n8040 ^ n5746 ;
  assign n24898 = ( ~n13388 & n14288 ) | ( ~n13388 & n20200 ) | ( n14288 & n20200 ) ;
  assign n24899 = n24898 ^ n24142 ^ n7552 ;
  assign n24900 = ( n8199 & ~n24897 ) | ( n8199 & n24899 ) | ( ~n24897 & n24899 ) ;
  assign n24901 = ( n3723 & n12764 ) | ( n3723 & ~n13526 ) | ( n12764 & ~n13526 ) ;
  assign n24902 = n21707 ^ n15840 ^ n6352 ;
  assign n24903 = ~n9359 & n12790 ;
  assign n24904 = n5434 ^ n5058 ^ 1'b0 ;
  assign n24905 = ( n4660 & ~n10616 ) | ( n4660 & n24904 ) | ( ~n10616 & n24904 ) ;
  assign n24906 = n9060 ^ n3695 ^ n2888 ;
  assign n24907 = ( n8563 & n21972 ) | ( n8563 & ~n24605 ) | ( n21972 & ~n24605 ) ;
  assign n24908 = n24907 ^ n14417 ^ n13441 ;
  assign n24909 = ( n3234 & ~n21894 ) | ( n3234 & n24908 ) | ( ~n21894 & n24908 ) ;
  assign n24910 = n17043 ^ n10702 ^ n1925 ;
  assign n24911 = ( n10166 & n11285 ) | ( n10166 & ~n24042 ) | ( n11285 & ~n24042 ) ;
  assign n24912 = n24911 ^ n12859 ^ n6073 ;
  assign n24913 = ( n11390 & ~n24910 ) | ( n11390 & n24912 ) | ( ~n24910 & n24912 ) ;
  assign n24914 = ( ~n12332 & n19397 ) | ( ~n12332 & n24913 ) | ( n19397 & n24913 ) ;
  assign n24916 = ( n3300 & n12359 ) | ( n3300 & n15406 ) | ( n12359 & n15406 ) ;
  assign n24915 = n11274 ^ n7660 ^ n3986 ;
  assign n24917 = n24916 ^ n24915 ^ 1'b0 ;
  assign n24918 = n14006 ^ n6244 ^ n2523 ;
  assign n24919 = n15430 ^ n5460 ^ 1'b0 ;
  assign n24920 = n2262 | n10148 ;
  assign n24921 = n9016 | n24920 ;
  assign n24922 = n24921 ^ n7409 ^ 1'b0 ;
  assign n24923 = ( ~n12420 & n24919 ) | ( ~n12420 & n24922 ) | ( n24919 & n24922 ) ;
  assign n24924 = ( ~n3288 & n10073 ) | ( ~n3288 & n24752 ) | ( n10073 & n24752 ) ;
  assign n24925 = n16874 | n24924 ;
  assign n24926 = n1229 | n10129 ;
  assign n24927 = n24926 ^ n8277 ^ 1'b0 ;
  assign n24928 = ( n809 & ~n10801 ) | ( n809 & n14200 ) | ( ~n10801 & n14200 ) ;
  assign n24929 = ( ~n2265 & n2549 ) | ( ~n2265 & n24928 ) | ( n2549 & n24928 ) ;
  assign n24930 = ( n10182 & n20236 ) | ( n10182 & ~n24929 ) | ( n20236 & ~n24929 ) ;
  assign n24931 = ( ~n1943 & n5268 ) | ( ~n1943 & n6223 ) | ( n5268 & n6223 ) ;
  assign n24932 = n24931 ^ n20341 ^ n11746 ;
  assign n24933 = n4171 & ~n24932 ;
  assign n24934 = n24933 ^ n12231 ^ 1'b0 ;
  assign n24935 = n24934 ^ n16428 ^ n12564 ;
  assign n24936 = ( ~n604 & n10257 ) | ( ~n604 & n15151 ) | ( n10257 & n15151 ) ;
  assign n24937 = ( n9131 & ~n12123 ) | ( n9131 & n12318 ) | ( ~n12123 & n12318 ) ;
  assign n24938 = ( n15413 & n24936 ) | ( n15413 & ~n24937 ) | ( n24936 & ~n24937 ) ;
  assign n24939 = n965 | n17563 ;
  assign n24940 = ( n6871 & n19415 ) | ( n6871 & n24939 ) | ( n19415 & n24939 ) ;
  assign n24941 = n21357 ^ n5172 ^ x17 ;
  assign n24942 = n14196 ^ n6991 ^ n4529 ;
  assign n24944 = n16084 ^ n8055 ^ 1'b0 ;
  assign n24945 = n24944 ^ n17486 ^ n16598 ;
  assign n24943 = n21472 ^ n15634 ^ n3445 ;
  assign n24946 = n24945 ^ n24943 ^ n3887 ;
  assign n24947 = ( n9469 & ~n11625 ) | ( n9469 & n17348 ) | ( ~n11625 & n17348 ) ;
  assign n24948 = n9953 & n24947 ;
  assign n24949 = n24948 ^ n22609 ^ n5968 ;
  assign n24959 = n3234 & ~n9026 ;
  assign n24958 = n18958 ^ n2063 ^ 1'b0 ;
  assign n24960 = n24959 ^ n24958 ^ n358 ;
  assign n24961 = ( n9124 & n11155 ) | ( n9124 & ~n24960 ) | ( n11155 & ~n24960 ) ;
  assign n24957 = n15983 ^ n13491 ^ n13407 ;
  assign n24950 = n18487 ^ n5539 ^ n1801 ;
  assign n24951 = n24950 ^ n3751 ^ n1121 ;
  assign n24952 = ( n3230 & n15790 ) | ( n3230 & n24951 ) | ( n15790 & n24951 ) ;
  assign n24953 = n11375 ^ x232 ^ 1'b0 ;
  assign n24954 = n5661 ^ n3795 ^ n1570 ;
  assign n24955 = n24953 & ~n24954 ;
  assign n24956 = ( n17958 & n24952 ) | ( n17958 & ~n24955 ) | ( n24952 & ~n24955 ) ;
  assign n24962 = n24961 ^ n24957 ^ n24956 ;
  assign n24963 = n12904 ^ n12896 ^ n4163 ;
  assign n24964 = n22630 ^ n16242 ^ n1601 ;
  assign n24965 = n6775 ^ n3847 ^ n3086 ;
  assign n24966 = ( n3980 & n20843 ) | ( n3980 & ~n24965 ) | ( n20843 & ~n24965 ) ;
  assign n24967 = ( ~n11713 & n24964 ) | ( ~n11713 & n24966 ) | ( n24964 & n24966 ) ;
  assign n24968 = ( n16170 & n24963 ) | ( n16170 & n24967 ) | ( n24963 & n24967 ) ;
  assign n24969 = n8450 ^ n6187 ^ n1288 ;
  assign n24970 = n24969 ^ n24932 ^ n8995 ;
  assign n24971 = n15076 ^ n11009 ^ n5394 ;
  assign n24972 = n19003 ^ n4691 ^ n719 ;
  assign n24973 = ~n6376 & n24972 ;
  assign n24974 = n9725 & n24973 ;
  assign n24975 = ( n17199 & ~n17999 ) | ( n17199 & n19295 ) | ( ~n17999 & n19295 ) ;
  assign n24976 = ~n6506 & n24975 ;
  assign n24977 = ( n15585 & ~n21545 ) | ( n15585 & n24976 ) | ( ~n21545 & n24976 ) ;
  assign n24979 = ( ~n7234 & n7887 ) | ( ~n7234 & n14445 ) | ( n7887 & n14445 ) ;
  assign n24978 = n5595 ^ n1618 ^ 1'b0 ;
  assign n24980 = n24979 ^ n24978 ^ n23149 ;
  assign n24981 = n20059 ^ n2575 ^ x131 ;
  assign n24982 = n24981 ^ n20217 ^ n901 ;
  assign n24983 = ( ~n1448 & n24610 ) | ( ~n1448 & n24982 ) | ( n24610 & n24982 ) ;
  assign n24984 = ( n12455 & n15212 ) | ( n12455 & ~n16881 ) | ( n15212 & ~n16881 ) ;
  assign n24985 = ( ~n721 & n13500 ) | ( ~n721 & n24984 ) | ( n13500 & n24984 ) ;
  assign n24986 = n20027 ^ n10028 ^ n3708 ;
  assign n24987 = ( n15147 & n19781 ) | ( n15147 & n24986 ) | ( n19781 & n24986 ) ;
  assign n24988 = ( n2781 & n9652 ) | ( n2781 & n24987 ) | ( n9652 & n24987 ) ;
  assign n24989 = ( n24983 & n24985 ) | ( n24983 & n24988 ) | ( n24985 & n24988 ) ;
  assign n24990 = ( ~n2351 & n8946 ) | ( ~n2351 & n15493 ) | ( n8946 & n15493 ) ;
  assign n24991 = ( n6178 & n20559 ) | ( n6178 & n24990 ) | ( n20559 & n24990 ) ;
  assign n24992 = n24991 ^ n24047 ^ n15741 ;
  assign n24993 = ( ~n9114 & n11604 ) | ( ~n9114 & n12215 ) | ( n11604 & n12215 ) ;
  assign n24994 = n24993 ^ n19974 ^ n6199 ;
  assign n24995 = ( n4036 & ~n9336 ) | ( n4036 & n24994 ) | ( ~n9336 & n24994 ) ;
  assign n24996 = n14491 ^ n5286 ^ 1'b0 ;
  assign n24997 = n24996 ^ n24928 ^ n14675 ;
  assign n24998 = ( ~n7256 & n14668 ) | ( ~n7256 & n20424 ) | ( n14668 & n20424 ) ;
  assign n24999 = n16789 & n24998 ;
  assign n25000 = n24999 ^ n15452 ^ n8113 ;
  assign n25001 = n10831 ^ n8634 ^ n3864 ;
  assign n25002 = n3638 & n6407 ;
  assign n25003 = n25002 ^ n10955 ^ 1'b0 ;
  assign n25004 = n25003 ^ n12380 ^ n536 ;
  assign n25005 = ( ~n1700 & n10195 ) | ( ~n1700 & n25004 ) | ( n10195 & n25004 ) ;
  assign n25006 = n21394 ^ n10442 ^ n4744 ;
  assign n25007 = ( ~n20828 & n23042 ) | ( ~n20828 & n25006 ) | ( n23042 & n25006 ) ;
  assign n25008 = n25007 ^ n12593 ^ n9897 ;
  assign n25009 = ( n25001 & n25005 ) | ( n25001 & ~n25008 ) | ( n25005 & ~n25008 ) ;
  assign n25010 = n9898 & ~n13535 ;
  assign n25011 = n20552 | n25010 ;
  assign n25012 = n4213 | n25011 ;
  assign n25013 = ~n21540 & n24233 ;
  assign n25014 = ( n2657 & ~n9855 ) | ( n2657 & n17371 ) | ( ~n9855 & n17371 ) ;
  assign n25015 = ( ~n3262 & n4789 ) | ( ~n3262 & n19665 ) | ( n4789 & n19665 ) ;
  assign n25016 = ( ~n7087 & n24009 ) | ( ~n7087 & n25015 ) | ( n24009 & n25015 ) ;
  assign n25017 = n20722 ^ n18565 ^ 1'b0 ;
  assign n25018 = n1880 & ~n25017 ;
  assign n25019 = ( ~n25014 & n25016 ) | ( ~n25014 & n25018 ) | ( n25016 & n25018 ) ;
  assign n25025 = ( n8707 & n12684 ) | ( n8707 & n18983 ) | ( n12684 & n18983 ) ;
  assign n25026 = n25025 ^ n14009 ^ n4564 ;
  assign n25024 = n10385 ^ n9983 ^ n1464 ;
  assign n25020 = n11126 ^ n7624 ^ n3456 ;
  assign n25021 = n536 | n25020 ;
  assign n25022 = n25021 ^ n3988 ^ 1'b0 ;
  assign n25023 = n25022 ^ n16736 ^ n9964 ;
  assign n25027 = n25026 ^ n25024 ^ n25023 ;
  assign n25028 = n5984 ^ n5725 ^ n382 ;
  assign n25029 = n25028 ^ n24587 ^ n7545 ;
  assign n25030 = n11588 ^ n7195 ^ 1'b0 ;
  assign n25031 = n25030 ^ n18909 ^ n13790 ;
  assign n25032 = n25031 ^ n3845 ^ 1'b0 ;
  assign n25033 = n7493 & ~n25032 ;
  assign n25034 = ( n12331 & ~n12702 ) | ( n12331 & n21636 ) | ( ~n12702 & n21636 ) ;
  assign n25035 = ( ~n7092 & n10570 ) | ( ~n7092 & n25034 ) | ( n10570 & n25034 ) ;
  assign n25036 = ( n2098 & n17940 ) | ( n2098 & n18001 ) | ( n17940 & n18001 ) ;
  assign n25037 = ( n8488 & ~n12056 ) | ( n8488 & n21190 ) | ( ~n12056 & n21190 ) ;
  assign n25038 = n25037 ^ n14590 ^ n3153 ;
  assign n25039 = ( n7060 & ~n11514 ) | ( n7060 & n14014 ) | ( ~n11514 & n14014 ) ;
  assign n25040 = n20281 & n25039 ;
  assign n25041 = n9086 & n25040 ;
  assign n25042 = ( n2403 & n21351 ) | ( n2403 & n25041 ) | ( n21351 & n25041 ) ;
  assign n25043 = ( n11122 & ~n16631 ) | ( n11122 & n25042 ) | ( ~n16631 & n25042 ) ;
  assign n25044 = n25043 ^ n7425 ^ n5595 ;
  assign n25045 = n13110 ^ n1424 ^ 1'b0 ;
  assign n25046 = n25045 ^ n12994 ^ n9192 ;
  assign n25047 = ( n25038 & n25044 ) | ( n25038 & ~n25046 ) | ( n25044 & ~n25046 ) ;
  assign n25048 = n8350 ^ n7628 ^ n953 ;
  assign n25049 = ( n2373 & n19328 ) | ( n2373 & ~n25048 ) | ( n19328 & ~n25048 ) ;
  assign n25050 = n25049 ^ n10401 ^ n4568 ;
  assign n25051 = n25050 ^ n20576 ^ n4735 ;
  assign n25052 = ( n5989 & n11994 ) | ( n5989 & n19332 ) | ( n11994 & n19332 ) ;
  assign n25053 = n1945 & n12594 ;
  assign n25054 = n23327 ^ n11380 ^ n5131 ;
  assign n25055 = ( n2481 & n4403 ) | ( n2481 & ~n16568 ) | ( n4403 & ~n16568 ) ;
  assign n25056 = ( n14384 & ~n25054 ) | ( n14384 & n25055 ) | ( ~n25054 & n25055 ) ;
  assign n25057 = ( n5061 & n5458 ) | ( n5061 & n11074 ) | ( n5458 & n11074 ) ;
  assign n25058 = n18723 ^ n17839 ^ n17025 ;
  assign n25059 = ( n734 & n25057 ) | ( n734 & ~n25058 ) | ( n25057 & ~n25058 ) ;
  assign n25060 = ( n25053 & ~n25056 ) | ( n25053 & n25059 ) | ( ~n25056 & n25059 ) ;
  assign n25061 = n2776 & ~n22027 ;
  assign n25062 = n23183 ^ n13423 ^ n947 ;
  assign n25063 = n25062 ^ n4494 ^ 1'b0 ;
  assign n25064 = n4334 | n22941 ;
  assign n25065 = n25063 & ~n25064 ;
  assign n25066 = ( n17787 & ~n25061 ) | ( n17787 & n25065 ) | ( ~n25061 & n25065 ) ;
  assign n25067 = ~n15576 & n19364 ;
  assign n25068 = n25067 ^ n20521 ^ 1'b0 ;
  assign n25069 = ( ~n6546 & n7216 ) | ( ~n6546 & n7281 ) | ( n7216 & n7281 ) ;
  assign n25070 = ( ~n3828 & n7596 ) | ( ~n3828 & n18606 ) | ( n7596 & n18606 ) ;
  assign n25071 = ( n4922 & n18738 ) | ( n4922 & ~n21019 ) | ( n18738 & ~n21019 ) ;
  assign n25072 = ~n4277 & n17578 ;
  assign n25073 = n25072 ^ n17949 ^ 1'b0 ;
  assign n25074 = ( n2293 & ~n8059 ) | ( n2293 & n10298 ) | ( ~n8059 & n10298 ) ;
  assign n25075 = ( ~n1361 & n3453 ) | ( ~n1361 & n5930 ) | ( n3453 & n5930 ) ;
  assign n25078 = n3768 | n4879 ;
  assign n25079 = n25078 ^ n13615 ^ n4620 ;
  assign n25076 = ( n7187 & n11264 ) | ( n7187 & ~n19239 ) | ( n11264 & ~n19239 ) ;
  assign n25077 = n25076 ^ n18975 ^ n6940 ;
  assign n25080 = n25079 ^ n25077 ^ n12207 ;
  assign n25083 = n10864 ^ n8380 ^ n7737 ;
  assign n25082 = ( n18132 & ~n22363 ) | ( n18132 & n23090 ) | ( ~n22363 & n23090 ) ;
  assign n25081 = n15095 ^ n12855 ^ n506 ;
  assign n25084 = n25083 ^ n25082 ^ n25081 ;
  assign n25085 = n7038 ^ n1120 ^ 1'b0 ;
  assign n25086 = ~n2570 & n25085 ;
  assign n25087 = n10185 & ~n19921 ;
  assign n25088 = ( n4727 & ~n12781 ) | ( n4727 & n25087 ) | ( ~n12781 & n25087 ) ;
  assign n25089 = n25088 ^ n6381 ^ n3836 ;
  assign n25090 = ( n3104 & n3267 ) | ( n3104 & n20549 ) | ( n3267 & n20549 ) ;
  assign n25091 = n971 | n25090 ;
  assign n25092 = n11094 | n25091 ;
  assign n25093 = ( ~n10287 & n25089 ) | ( ~n10287 & n25092 ) | ( n25089 & n25092 ) ;
  assign n25094 = ( n6188 & ~n6292 ) | ( n6188 & n22196 ) | ( ~n6292 & n22196 ) ;
  assign n25095 = n25094 ^ n14304 ^ n4049 ;
  assign n25096 = n25095 ^ n4659 ^ n1081 ;
  assign n25097 = ( n308 & n23646 ) | ( n308 & ~n25096 ) | ( n23646 & ~n25096 ) ;
  assign n25098 = ( ~n8777 & n14227 ) | ( ~n8777 & n25097 ) | ( n14227 & n25097 ) ;
  assign n25099 = ( n2523 & n8707 ) | ( n2523 & n13999 ) | ( n8707 & n13999 ) ;
  assign n25100 = ( n8293 & n15075 ) | ( n8293 & n25099 ) | ( n15075 & n25099 ) ;
  assign n25101 = n14739 ^ n5494 ^ x33 ;
  assign n25102 = ( n7692 & n12326 ) | ( n7692 & ~n13804 ) | ( n12326 & ~n13804 ) ;
  assign n25103 = ~n25101 & n25102 ;
  assign n25104 = n25103 ^ n4825 ^ 1'b0 ;
  assign n25105 = n21115 ^ n14180 ^ n10939 ;
  assign n25106 = n25105 ^ n10279 ^ n8438 ;
  assign n25107 = n25106 ^ n16308 ^ n7747 ;
  assign n25108 = n9776 ^ n3491 ^ n909 ;
  assign n25109 = n25108 ^ n18270 ^ n14778 ;
  assign n25110 = n17668 ^ n17392 ^ n4928 ;
  assign n25111 = n25110 ^ n6183 ^ n2254 ;
  assign n25112 = ( ~n10379 & n25109 ) | ( ~n10379 & n25111 ) | ( n25109 & n25111 ) ;
  assign n25114 = n21559 ^ n17762 ^ n12472 ;
  assign n25113 = ( n14768 & ~n18547 ) | ( n14768 & n22961 ) | ( ~n18547 & n22961 ) ;
  assign n25115 = n25114 ^ n25113 ^ n13361 ;
  assign n25116 = ( ~x253 & n6737 ) | ( ~x253 & n21559 ) | ( n6737 & n21559 ) ;
  assign n25117 = ( ~x51 & n14784 ) | ( ~x51 & n25116 ) | ( n14784 & n25116 ) ;
  assign n25118 = ( ~n4069 & n9412 ) | ( ~n4069 & n10784 ) | ( n9412 & n10784 ) ;
  assign n25119 = ( x26 & n278 ) | ( x26 & ~n3375 ) | ( n278 & ~n3375 ) ;
  assign n25120 = ( n15691 & ~n20220 ) | ( n15691 & n25119 ) | ( ~n20220 & n25119 ) ;
  assign n25121 = n25120 ^ n11744 ^ 1'b0 ;
  assign n25122 = n17613 ^ n13628 ^ n7902 ;
  assign n25123 = n15058 ^ n4518 ^ n3035 ;
  assign n25124 = n25123 ^ n15876 ^ n5027 ;
  assign n25125 = n21024 ^ n6913 ^ n6267 ;
  assign n25126 = ( n22538 & n25124 ) | ( n22538 & ~n25125 ) | ( n25124 & ~n25125 ) ;
  assign n25131 = ( x59 & n4621 ) | ( x59 & n22714 ) | ( n4621 & n22714 ) ;
  assign n25128 = n5427 ^ n4661 ^ 1'b0 ;
  assign n25129 = n10825 & n25128 ;
  assign n25127 = ( n1230 & ~n3500 ) | ( n1230 & n9717 ) | ( ~n3500 & n9717 ) ;
  assign n25130 = n25129 ^ n25127 ^ n20547 ;
  assign n25132 = n25131 ^ n25130 ^ n13684 ;
  assign n25133 = ( n3714 & n16676 ) | ( n3714 & n25132 ) | ( n16676 & n25132 ) ;
  assign n25138 = n8573 ^ n7845 ^ n5614 ;
  assign n25134 = ( n2398 & ~n5081 ) | ( n2398 & n7873 ) | ( ~n5081 & n7873 ) ;
  assign n25135 = ( ~n1790 & n3579 ) | ( ~n1790 & n25134 ) | ( n3579 & n25134 ) ;
  assign n25136 = n13583 & ~n25135 ;
  assign n25137 = ( ~n12815 & n15376 ) | ( ~n12815 & n25136 ) | ( n15376 & n25136 ) ;
  assign n25139 = n25138 ^ n25137 ^ n13824 ;
  assign n25141 = n23230 ^ n2439 ^ n371 ;
  assign n25140 = n11543 & ~n16097 ;
  assign n25142 = n25141 ^ n25140 ^ n18745 ;
  assign n25143 = n11965 ^ n5120 ^ 1'b0 ;
  assign n25144 = ~n25142 & n25143 ;
  assign n25145 = ( n1886 & n3904 ) | ( n1886 & n6548 ) | ( n3904 & n6548 ) ;
  assign n25146 = n13902 ^ n11801 ^ n10790 ;
  assign n25147 = ( n8465 & ~n25145 ) | ( n8465 & n25146 ) | ( ~n25145 & n25146 ) ;
  assign n25148 = ( n1358 & n3737 ) | ( n1358 & ~n14181 ) | ( n3737 & ~n14181 ) ;
  assign n25149 = ~n7926 & n25148 ;
  assign n25150 = n25149 ^ n17994 ^ 1'b0 ;
  assign n25151 = n25150 ^ n2346 ^ n1410 ;
  assign n25157 = ( ~n10094 & n11897 ) | ( ~n10094 & n14613 ) | ( n11897 & n14613 ) ;
  assign n25152 = n3194 ^ x96 ^ 1'b0 ;
  assign n25153 = x249 & ~n25152 ;
  assign n25154 = n14985 ^ n1015 ^ 1'b0 ;
  assign n25155 = ( n802 & ~n6194 ) | ( n802 & n10741 ) | ( ~n6194 & n10741 ) ;
  assign n25156 = ( n25153 & n25154 ) | ( n25153 & n25155 ) | ( n25154 & n25155 ) ;
  assign n25158 = n25157 ^ n25156 ^ n9283 ;
  assign n25159 = ( n2351 & n25151 ) | ( n2351 & n25158 ) | ( n25151 & n25158 ) ;
  assign n25162 = ( ~n8741 & n10142 ) | ( ~n8741 & n14242 ) | ( n10142 & n14242 ) ;
  assign n25160 = n14724 ^ n3119 ^ n703 ;
  assign n25161 = n25160 ^ n9281 ^ n5944 ;
  assign n25163 = n25162 ^ n25161 ^ 1'b0 ;
  assign n25166 = n21209 ^ n12512 ^ n5809 ;
  assign n25167 = ( n2326 & n12529 ) | ( n2326 & n25166 ) | ( n12529 & n25166 ) ;
  assign n25164 = ( n2031 & n11876 ) | ( n2031 & ~n23230 ) | ( n11876 & ~n23230 ) ;
  assign n25165 = n15678 & ~n25164 ;
  assign n25168 = n25167 ^ n25165 ^ n21447 ;
  assign n25170 = ( n1759 & n2874 ) | ( n1759 & n16670 ) | ( n2874 & n16670 ) ;
  assign n25169 = n23590 ^ n22422 ^ n11112 ;
  assign n25171 = n25170 ^ n25169 ^ n3488 ;
  assign n25172 = n25171 ^ n2405 ^ n1503 ;
  assign n25173 = n9488 ^ n1252 ^ 1'b0 ;
  assign n25174 = n6093 | n21373 ;
  assign n25175 = n25174 ^ n13795 ^ 1'b0 ;
  assign n25176 = ( n370 & n14132 ) | ( n370 & n25175 ) | ( n14132 & n25175 ) ;
  assign n25177 = ( n449 & n25173 ) | ( n449 & n25176 ) | ( n25173 & n25176 ) ;
  assign n25178 = ( n5739 & n16693 ) | ( n5739 & ~n25177 ) | ( n16693 & ~n25177 ) ;
  assign n25179 = n21820 ^ n19769 ^ n2652 ;
  assign n25180 = ( n1430 & ~n11667 ) | ( n1430 & n25179 ) | ( ~n11667 & n25179 ) ;
  assign n25181 = n8244 & ~n25180 ;
  assign n25182 = ~n1418 & n25181 ;
  assign n25183 = ( ~n22525 & n24824 ) | ( ~n22525 & n25182 ) | ( n24824 & n25182 ) ;
  assign n25184 = n18654 ^ n7685 ^ n1648 ;
  assign n25185 = ( n2643 & n24293 ) | ( n2643 & n25184 ) | ( n24293 & n25184 ) ;
  assign n25186 = n14132 & ~n18825 ;
  assign n25187 = n25186 ^ n9555 ^ n8022 ;
  assign n25188 = n14618 ^ n9799 ^ n6940 ;
  assign n25189 = ( n6444 & n11590 ) | ( n6444 & ~n25188 ) | ( n11590 & ~n25188 ) ;
  assign n25190 = n25189 ^ n21633 ^ n4191 ;
  assign n25191 = n11993 ^ n5568 ^ n3962 ;
  assign n25192 = ( ~n3303 & n10033 ) | ( ~n3303 & n19315 ) | ( n10033 & n19315 ) ;
  assign n25193 = ( n5792 & n25191 ) | ( n5792 & n25192 ) | ( n25191 & n25192 ) ;
  assign n25194 = ( n7577 & n11474 ) | ( n7577 & ~n15748 ) | ( n11474 & ~n15748 ) ;
  assign n25195 = ( n2080 & ~n4897 ) | ( n2080 & n13291 ) | ( ~n4897 & n13291 ) ;
  assign n25196 = ( n9850 & n25194 ) | ( n9850 & n25195 ) | ( n25194 & n25195 ) ;
  assign n25197 = ( n9390 & n25193 ) | ( n9390 & ~n25196 ) | ( n25193 & ~n25196 ) ;
  assign n25198 = n11521 ^ n4789 ^ n285 ;
  assign n25199 = ( n2104 & n10555 ) | ( n2104 & ~n16130 ) | ( n10555 & ~n16130 ) ;
  assign n25200 = n1262 | n6156 ;
  assign n25201 = n25199 & ~n25200 ;
  assign n25202 = n25201 ^ n12687 ^ n3481 ;
  assign n25203 = n25202 ^ n7219 ^ n3343 ;
  assign n25204 = ( n9190 & n25198 ) | ( n9190 & n25203 ) | ( n25198 & n25203 ) ;
  assign n25205 = n25204 ^ n21034 ^ n17572 ;
  assign n25206 = ( ~n676 & n1591 ) | ( ~n676 & n6413 ) | ( n1591 & n6413 ) ;
  assign n25207 = ( n2336 & n7840 ) | ( n2336 & n25206 ) | ( n7840 & n25206 ) ;
  assign n25208 = n21082 ^ n16609 ^ n2116 ;
  assign n25209 = n25208 ^ n8813 ^ n2069 ;
  assign n25210 = n25207 | n25209 ;
  assign n25211 = n25205 & ~n25210 ;
  assign n25216 = ( n6403 & ~n16542 ) | ( n6403 & n23899 ) | ( ~n16542 & n23899 ) ;
  assign n25213 = n1686 | n1843 ;
  assign n25214 = n1346 & ~n25213 ;
  assign n25212 = ( n1215 & n2457 ) | ( n1215 & n10492 ) | ( n2457 & n10492 ) ;
  assign n25215 = n25214 ^ n25212 ^ n442 ;
  assign n25217 = n25216 ^ n25215 ^ n8628 ;
  assign n25218 = n25217 ^ n1530 ^ n1377 ;
  assign n25220 = n13500 ^ n7190 ^ n336 ;
  assign n25219 = n7932 ^ n2493 ^ n1903 ;
  assign n25221 = n25220 ^ n25219 ^ 1'b0 ;
  assign n25222 = n6776 ^ n5984 ^ n4687 ;
  assign n25223 = n8496 ^ n1695 ^ x204 ;
  assign n25224 = ( n8524 & n25222 ) | ( n8524 & ~n25223 ) | ( n25222 & ~n25223 ) ;
  assign n25225 = n25224 ^ n8387 ^ n323 ;
  assign n25226 = ( n5981 & ~n6455 ) | ( n5981 & n9986 ) | ( ~n6455 & n9986 ) ;
  assign n25227 = ( n2231 & ~n25225 ) | ( n2231 & n25226 ) | ( ~n25225 & n25226 ) ;
  assign n25234 = ~n1472 & n13351 ;
  assign n25233 = ( n1593 & n4759 ) | ( n1593 & n6792 ) | ( n4759 & n6792 ) ;
  assign n25235 = n25234 ^ n25233 ^ n7640 ;
  assign n25232 = ~n8012 & n17939 ;
  assign n25236 = n25235 ^ n25232 ^ n10520 ;
  assign n25228 = ( n1880 & ~n2828 ) | ( n1880 & n10674 ) | ( ~n2828 & n10674 ) ;
  assign n25229 = ( n9209 & n21695 ) | ( n9209 & ~n25228 ) | ( n21695 & ~n25228 ) ;
  assign n25230 = n7635 ^ x8 ^ 1'b0 ;
  assign n25231 = ( ~n7270 & n25229 ) | ( ~n7270 & n25230 ) | ( n25229 & n25230 ) ;
  assign n25237 = n25236 ^ n25231 ^ n20594 ;
  assign n25238 = ( n678 & n829 ) | ( n678 & ~n2209 ) | ( n829 & ~n2209 ) ;
  assign n25239 = n25238 ^ n17927 ^ n322 ;
  assign n25240 = ( n11444 & ~n25237 ) | ( n11444 & n25239 ) | ( ~n25237 & n25239 ) ;
  assign n25241 = n5951 ^ n4911 ^ n1990 ;
  assign n25242 = ( n18480 & n19315 ) | ( n18480 & n22963 ) | ( n19315 & n22963 ) ;
  assign n25243 = ( n4481 & n5450 ) | ( n4481 & n6056 ) | ( n5450 & n6056 ) ;
  assign n25244 = n25243 ^ n8293 ^ n2800 ;
  assign n25245 = n11688 ^ n5136 ^ 1'b0 ;
  assign n25246 = ( n23467 & ~n25244 ) | ( n23467 & n25245 ) | ( ~n25244 & n25245 ) ;
  assign n25247 = n15010 ^ n8437 ^ n873 ;
  assign n25248 = n4963 & ~n15245 ;
  assign n25249 = n25248 ^ n22827 ^ 1'b0 ;
  assign n25250 = n25249 ^ n13799 ^ n5292 ;
  assign n25261 = ( n4589 & n15872 ) | ( n4589 & ~n23604 ) | ( n15872 & ~n23604 ) ;
  assign n25251 = n8736 ^ n4945 ^ n2280 ;
  assign n25252 = n5964 ^ x98 ^ 1'b0 ;
  assign n25253 = n11208 & ~n25252 ;
  assign n25254 = n11337 ^ n6589 ^ n2091 ;
  assign n25255 = ( x113 & n4141 ) | ( x113 & ~n10395 ) | ( n4141 & ~n10395 ) ;
  assign n25256 = n25255 ^ n4367 ^ 1'b0 ;
  assign n25257 = n1392 & n25256 ;
  assign n25258 = ( n11468 & n25254 ) | ( n11468 & n25257 ) | ( n25254 & n25257 ) ;
  assign n25259 = ( n18932 & n25253 ) | ( n18932 & ~n25258 ) | ( n25253 & ~n25258 ) ;
  assign n25260 = ( n7691 & n25251 ) | ( n7691 & n25259 ) | ( n25251 & n25259 ) ;
  assign n25262 = n25261 ^ n25260 ^ n6022 ;
  assign n25263 = n21965 ^ n9511 ^ n4978 ;
  assign n25264 = n25263 ^ n16050 ^ n1561 ;
  assign n25271 = n20865 ^ n18711 ^ n7521 ;
  assign n25265 = ( n3739 & ~n4147 ) | ( n3739 & n20707 ) | ( ~n4147 & n20707 ) ;
  assign n25266 = n11057 ^ n8312 ^ 1'b0 ;
  assign n25267 = ~n2677 & n25266 ;
  assign n25268 = n25267 ^ n20995 ^ 1'b0 ;
  assign n25269 = ~n25111 & n25268 ;
  assign n25270 = ( n7717 & n25265 ) | ( n7717 & ~n25269 ) | ( n25265 & ~n25269 ) ;
  assign n25272 = n25271 ^ n25270 ^ x151 ;
  assign n25275 = ( ~n1464 & n7535 ) | ( ~n1464 & n21091 ) | ( n7535 & n21091 ) ;
  assign n25273 = n24869 ^ n18324 ^ n13842 ;
  assign n25274 = n8802 | n25273 ;
  assign n25276 = n25275 ^ n25274 ^ n17407 ;
  assign n25282 = n15974 ^ n13932 ^ n536 ;
  assign n25283 = n25282 ^ n6141 ^ n2254 ;
  assign n25280 = n1787 & n19545 ;
  assign n25279 = ( n3570 & ~n8134 ) | ( n3570 & n13133 ) | ( ~n8134 & n13133 ) ;
  assign n25281 = n25280 ^ n25279 ^ 1'b0 ;
  assign n25277 = n6959 ^ n4347 ^ 1'b0 ;
  assign n25278 = n25277 ^ n17464 ^ n7953 ;
  assign n25284 = n25283 ^ n25281 ^ n25278 ;
  assign n25285 = ~n16719 & n20551 ;
  assign n25286 = ~n7173 & n25285 ;
  assign n25287 = n22978 ^ n1249 ^ 1'b0 ;
  assign n25288 = n25287 ^ n23355 ^ n6057 ;
  assign n25290 = ( ~n1243 & n4834 ) | ( ~n1243 & n12780 ) | ( n4834 & n12780 ) ;
  assign n25289 = n16489 ^ n16475 ^ 1'b0 ;
  assign n25291 = n25290 ^ n25289 ^ n18805 ;
  assign n25292 = n5609 ^ n3248 ^ n2944 ;
  assign n25293 = n25292 ^ n4970 ^ 1'b0 ;
  assign n25294 = ( ~n6927 & n14197 ) | ( ~n6927 & n25293 ) | ( n14197 & n25293 ) ;
  assign n25295 = ~n5041 & n25294 ;
  assign n25296 = ( n2192 & ~n13786 ) | ( n2192 & n20837 ) | ( ~n13786 & n20837 ) ;
  assign n25297 = n25296 ^ n15118 ^ n12279 ;
  assign n25305 = n17022 ^ n8371 ^ n5608 ;
  assign n25298 = ( n3224 & ~n7341 ) | ( n3224 & n13030 ) | ( ~n7341 & n13030 ) ;
  assign n25299 = ( n5374 & n13492 ) | ( n5374 & ~n25298 ) | ( n13492 & ~n25298 ) ;
  assign n25300 = ( ~n9479 & n19727 ) | ( ~n9479 & n22898 ) | ( n19727 & n22898 ) ;
  assign n25301 = n25300 ^ n18906 ^ n4028 ;
  assign n25302 = n25299 & ~n25301 ;
  assign n25303 = n25302 ^ n8590 ^ 1'b0 ;
  assign n25304 = ( n11087 & n12937 ) | ( n11087 & n25303 ) | ( n12937 & n25303 ) ;
  assign n25306 = n25305 ^ n25304 ^ n6538 ;
  assign n25307 = ( ~n2097 & n11782 ) | ( ~n2097 & n16021 ) | ( n11782 & n16021 ) ;
  assign n25310 = n6302 ^ n2335 ^ n983 ;
  assign n25309 = ( x26 & ~n9622 ) | ( x26 & n22530 ) | ( ~n9622 & n22530 ) ;
  assign n25308 = ( ~n2150 & n8654 ) | ( ~n2150 & n10338 ) | ( n8654 & n10338 ) ;
  assign n25311 = n25310 ^ n25309 ^ n25308 ;
  assign n25312 = n15620 | n25311 ;
  assign n25313 = n25312 ^ n21888 ^ n17837 ;
  assign n25314 = ( n2389 & n8981 ) | ( n2389 & ~n11614 ) | ( n8981 & ~n11614 ) ;
  assign n25315 = n25314 ^ n22121 ^ n3740 ;
  assign n25322 = n22617 ^ n6871 ^ n276 ;
  assign n25316 = n12335 ^ n1542 ^ 1'b0 ;
  assign n25317 = ( n9708 & ~n10579 ) | ( n9708 & n25316 ) | ( ~n10579 & n25316 ) ;
  assign n25318 = ( x62 & n24276 ) | ( x62 & n25317 ) | ( n24276 & n25317 ) ;
  assign n25319 = n25318 ^ n13411 ^ n4563 ;
  assign n25320 = n25319 ^ n18064 ^ n9619 ;
  assign n25321 = ( n3948 & n18469 ) | ( n3948 & n25320 ) | ( n18469 & n25320 ) ;
  assign n25323 = n25322 ^ n25321 ^ n21574 ;
  assign n25324 = n25323 ^ n18232 ^ n6439 ;
  assign n25325 = n5495 ^ n4961 ^ 1'b0 ;
  assign n25326 = ~n5082 & n25325 ;
  assign n25327 = n1833 & n25326 ;
  assign n25328 = n25327 ^ n13583 ^ 1'b0 ;
  assign n25329 = n25328 ^ n24242 ^ n7948 ;
  assign n25330 = n17876 ^ n16851 ^ x86 ;
  assign n25333 = n6995 ^ n3243 ^ n360 ;
  assign n25334 = n5960 & ~n25333 ;
  assign n25335 = n19201 & n25334 ;
  assign n25331 = ~n1079 & n4593 ;
  assign n25332 = ( n2852 & n17412 ) | ( n2852 & ~n25331 ) | ( n17412 & ~n25331 ) ;
  assign n25336 = n25335 ^ n25332 ^ n14654 ;
  assign n25337 = ( n7216 & ~n7903 ) | ( n7216 & n13559 ) | ( ~n7903 & n13559 ) ;
  assign n25338 = n7818 & n17376 ;
  assign n25339 = ~n25337 & n25338 ;
  assign n25340 = n25151 ^ n19239 ^ n3752 ;
  assign n25341 = ( n273 & n12028 ) | ( n273 & n25340 ) | ( n12028 & n25340 ) ;
  assign n25342 = n6161 & n13578 ;
  assign n25343 = n21782 ^ n12628 ^ n5588 ;
  assign n25344 = n25343 ^ n22342 ^ n13351 ;
  assign n25345 = n7094 & ~n25344 ;
  assign n25346 = n8809 ^ n8736 ^ n3620 ;
  assign n25347 = ( n7120 & n10304 ) | ( n7120 & ~n24130 ) | ( n10304 & ~n24130 ) ;
  assign n25348 = n25347 ^ n19453 ^ n5877 ;
  assign n25349 = ( n7810 & n12367 ) | ( n7810 & n18318 ) | ( n12367 & n18318 ) ;
  assign n25350 = n18803 ^ n18501 ^ 1'b0 ;
  assign n25351 = ~n3494 & n25350 ;
  assign n25352 = n6244 ^ n6058 ^ n1489 ;
  assign n25353 = ( n3895 & n10940 ) | ( n3895 & n25352 ) | ( n10940 & n25352 ) ;
  assign n25354 = ( ~n9430 & n25351 ) | ( ~n9430 & n25353 ) | ( n25351 & n25353 ) ;
  assign n25355 = n16965 ^ n7378 ^ n6581 ;
  assign n25356 = n25355 ^ n19875 ^ n19827 ;
  assign n25362 = n10557 ^ n9844 ^ n7028 ;
  assign n25357 = n17636 ^ n11483 ^ n7913 ;
  assign n25358 = n25357 ^ n3204 ^ n607 ;
  assign n25359 = n22033 ^ n5383 ^ n4698 ;
  assign n25360 = n25359 ^ n10077 ^ n661 ;
  assign n25361 = ( ~n4142 & n25358 ) | ( ~n4142 & n25360 ) | ( n25358 & n25360 ) ;
  assign n25363 = n25362 ^ n25361 ^ n5269 ;
  assign n25364 = n22699 ^ n2291 ^ n1783 ;
  assign n25365 = n15330 ^ n11017 ^ n1961 ;
  assign n25366 = ( ~n1424 & n2133 ) | ( ~n1424 & n4604 ) | ( n2133 & n4604 ) ;
  assign n25367 = n25366 ^ n4417 ^ n3132 ;
  assign n25368 = n25367 ^ n16978 ^ n16730 ;
  assign n25369 = ( n9725 & n25365 ) | ( n9725 & ~n25368 ) | ( n25365 & ~n25368 ) ;
  assign n25370 = ( n2464 & n6415 ) | ( n2464 & n13595 ) | ( n6415 & n13595 ) ;
  assign n25371 = ( ~n4754 & n5039 ) | ( ~n4754 & n6530 ) | ( n5039 & n6530 ) ;
  assign n25372 = ( n13975 & n24082 ) | ( n13975 & n25371 ) | ( n24082 & n25371 ) ;
  assign n25373 = n25372 ^ n18473 ^ n18434 ;
  assign n25374 = n25373 ^ n20223 ^ 1'b0 ;
  assign n25376 = n766 & n22424 ;
  assign n25377 = ~n16721 & n25376 ;
  assign n25378 = ( ~n548 & n22397 ) | ( ~n548 & n25377 ) | ( n22397 & n25377 ) ;
  assign n25379 = ( n7054 & ~n9277 ) | ( n7054 & n25378 ) | ( ~n9277 & n25378 ) ;
  assign n25375 = n20663 ^ n3922 ^ 1'b0 ;
  assign n25380 = n25379 ^ n25375 ^ n7558 ;
  assign n25381 = n9689 ^ n3045 ^ 1'b0 ;
  assign n25382 = n19876 ^ n12638 ^ n8348 ;
  assign n25383 = n25381 & ~n25382 ;
  assign n25384 = ~n25380 & n25383 ;
  assign n25389 = n10751 ^ n6633 ^ 1'b0 ;
  assign n25388 = n1160 & n4209 ;
  assign n25390 = n25389 ^ n25388 ^ 1'b0 ;
  assign n25385 = n7119 ^ x90 ^ 1'b0 ;
  assign n25386 = n25385 ^ n16894 ^ 1'b0 ;
  assign n25387 = n25386 ^ n12700 ^ 1'b0 ;
  assign n25391 = n25390 ^ n25387 ^ n512 ;
  assign n25392 = n14194 ^ n1548 ^ 1'b0 ;
  assign n25393 = ~n2998 & n25392 ;
  assign n25394 = ( ~x10 & n3514 ) | ( ~x10 & n25393 ) | ( n3514 & n25393 ) ;
  assign n25395 = ( ~n1539 & n7043 ) | ( ~n1539 & n20143 ) | ( n7043 & n20143 ) ;
  assign n25396 = ( ~n6281 & n8660 ) | ( ~n6281 & n25395 ) | ( n8660 & n25395 ) ;
  assign n25401 = ( n6583 & n19320 ) | ( n6583 & n23283 ) | ( n19320 & n23283 ) ;
  assign n25399 = ( n1124 & n3871 ) | ( n1124 & ~n4502 ) | ( n3871 & ~n4502 ) ;
  assign n25397 = n8523 & ~n24286 ;
  assign n25398 = ~n23785 & n25397 ;
  assign n25400 = n25399 ^ n25398 ^ 1'b0 ;
  assign n25402 = n25401 ^ n25400 ^ 1'b0 ;
  assign n25403 = ~n14201 & n25402 ;
  assign n25404 = n15316 ^ n11354 ^ n2711 ;
  assign n25405 = n25404 ^ n19614 ^ n4587 ;
  assign n25406 = n25405 ^ n10212 ^ 1'b0 ;
  assign n25407 = ( n6634 & ~n13302 ) | ( n6634 & n13547 ) | ( ~n13302 & n13547 ) ;
  assign n25408 = ( ~n1986 & n7789 ) | ( ~n1986 & n25407 ) | ( n7789 & n25407 ) ;
  assign n25409 = n25408 ^ n10431 ^ 1'b0 ;
  assign n25410 = ( n3959 & ~n9616 ) | ( n3959 & n14666 ) | ( ~n9616 & n14666 ) ;
  assign n25411 = n13135 ^ n9044 ^ n8081 ;
  assign n25412 = ( n16687 & n25410 ) | ( n16687 & n25411 ) | ( n25410 & n25411 ) ;
  assign n25413 = n13108 ^ n5587 ^ 1'b0 ;
  assign n25414 = n9280 & n25413 ;
  assign n25415 = ( n25409 & ~n25412 ) | ( n25409 & n25414 ) | ( ~n25412 & n25414 ) ;
  assign n25416 = ( n943 & n8782 ) | ( n943 & ~n12925 ) | ( n8782 & ~n12925 ) ;
  assign n25417 = n25416 ^ n21221 ^ n17924 ;
  assign n25418 = n25417 ^ n11706 ^ n544 ;
  assign n25419 = n14099 ^ n7158 ^ n590 ;
  assign n25420 = ~n4780 & n25419 ;
  assign n25421 = ~n25418 & n25420 ;
  assign n25422 = n25421 ^ n20075 ^ n8244 ;
  assign n25427 = n14692 ^ n13219 ^ n2918 ;
  assign n25425 = ( ~n1009 & n2767 ) | ( ~n1009 & n8739 ) | ( n2767 & n8739 ) ;
  assign n25426 = ( ~n9688 & n21053 ) | ( ~n9688 & n25425 ) | ( n21053 & n25425 ) ;
  assign n25423 = ( n9502 & ~n15255 ) | ( n9502 & n15880 ) | ( ~n15255 & n15880 ) ;
  assign n25424 = n25423 ^ n21393 ^ n10152 ;
  assign n25428 = n25427 ^ n25426 ^ n25424 ;
  assign n25429 = n2684 & ~n19429 ;
  assign n25430 = ~n25428 & n25429 ;
  assign n25434 = ( n12971 & ~n17711 ) | ( n12971 & n18917 ) | ( ~n17711 & n18917 ) ;
  assign n25431 = ( n4292 & ~n7031 ) | ( n4292 & n7574 ) | ( ~n7031 & n7574 ) ;
  assign n25432 = ( n8057 & ~n8299 ) | ( n8057 & n25431 ) | ( ~n8299 & n25431 ) ;
  assign n25433 = n11010 | n25432 ;
  assign n25435 = n25434 ^ n25433 ^ 1'b0 ;
  assign n25436 = n5030 & ~n6308 ;
  assign n25437 = n25436 ^ n22572 ^ n12305 ;
  assign n25438 = ( n11385 & ~n23660 ) | ( n11385 & n25437 ) | ( ~n23660 & n25437 ) ;
  assign n25439 = n14567 ^ n11002 ^ n6289 ;
  assign n25440 = ~n14735 & n21218 ;
  assign n25441 = ( n8181 & ~n16034 ) | ( n8181 & n20802 ) | ( ~n16034 & n20802 ) ;
  assign n25442 = n17075 ^ n6795 ^ 1'b0 ;
  assign n25443 = n25442 ^ n700 ^ 1'b0 ;
  assign n25444 = n4528 & ~n25443 ;
  assign n25446 = ( n6546 & n19153 ) | ( n6546 & n23212 ) | ( n19153 & n23212 ) ;
  assign n25445 = n13281 ^ n8645 ^ n921 ;
  assign n25447 = n25446 ^ n25445 ^ n19325 ;
  assign n25448 = n21407 ^ n5690 ^ n2471 ;
  assign n25449 = ( ~n3592 & n7704 ) | ( ~n3592 & n25448 ) | ( n7704 & n25448 ) ;
  assign n25450 = n25449 ^ n20901 ^ n6086 ;
  assign n25461 = ( n407 & n2171 ) | ( n407 & n8749 ) | ( n2171 & n8749 ) ;
  assign n25460 = ( n18325 & n22155 ) | ( n18325 & n22600 ) | ( n22155 & n22600 ) ;
  assign n25459 = n9539 ^ n4586 ^ n1735 ;
  assign n25462 = n25461 ^ n25460 ^ n25459 ;
  assign n25455 = n9458 ^ n2661 ^ n1379 ;
  assign n25456 = n17732 ^ n10194 ^ 1'b0 ;
  assign n25457 = n25455 & ~n25456 ;
  assign n25454 = ( n8686 & ~n14269 ) | ( n8686 & n15269 ) | ( ~n14269 & n15269 ) ;
  assign n25458 = n25457 ^ n25454 ^ n24216 ;
  assign n25451 = ( n1026 & n6672 ) | ( n1026 & ~n9180 ) | ( n6672 & ~n9180 ) ;
  assign n25452 = ( n2478 & n5014 ) | ( n2478 & ~n25451 ) | ( n5014 & ~n25451 ) ;
  assign n25453 = n25452 ^ n25150 ^ n19484 ;
  assign n25463 = n25462 ^ n25458 ^ n25453 ;
  assign n25464 = ( ~n4362 & n19459 ) | ( ~n4362 & n24854 ) | ( n19459 & n24854 ) ;
  assign n25467 = ( n1091 & n10252 ) | ( n1091 & ~n22834 ) | ( n10252 & ~n22834 ) ;
  assign n25465 = ( n1207 & n8198 ) | ( n1207 & n22156 ) | ( n8198 & n22156 ) ;
  assign n25466 = ( ~n1766 & n15655 ) | ( ~n1766 & n25465 ) | ( n15655 & n25465 ) ;
  assign n25468 = n25467 ^ n25466 ^ n10721 ;
  assign n25469 = n22577 & ~n25468 ;
  assign n25470 = n25469 ^ n17453 ^ 1'b0 ;
  assign n25471 = ( n1775 & n2716 ) | ( n1775 & n17590 ) | ( n2716 & n17590 ) ;
  assign n25472 = ( n1698 & n3014 ) | ( n1698 & ~n25471 ) | ( n3014 & ~n25471 ) ;
  assign n25473 = n1399 ^ n1146 ^ 1'b0 ;
  assign n25474 = ~n544 & n25473 ;
  assign n25475 = ~n11883 & n25474 ;
  assign n25476 = ~n25472 & n25475 ;
  assign n25477 = ( n4371 & n15145 ) | ( n4371 & ~n20223 ) | ( n15145 & ~n20223 ) ;
  assign n25478 = ( n14571 & n16082 ) | ( n14571 & ~n25477 ) | ( n16082 & ~n25477 ) ;
  assign n25482 = ( n2408 & n9153 ) | ( n2408 & ~n17266 ) | ( n9153 & ~n17266 ) ;
  assign n25479 = x21 & n1799 ;
  assign n25480 = n25479 ^ n14967 ^ 1'b0 ;
  assign n25481 = n25480 ^ n8341 ^ n6744 ;
  assign n25483 = n25482 ^ n25481 ^ n3032 ;
  assign n25484 = n18519 ^ n15748 ^ n5637 ;
  assign n25485 = ( n8678 & n24752 ) | ( n8678 & n25484 ) | ( n24752 & n25484 ) ;
  assign n25486 = ( n3759 & ~n5944 ) | ( n3759 & n11183 ) | ( ~n5944 & n11183 ) ;
  assign n25487 = n8900 ^ n2846 ^ 1'b0 ;
  assign n25488 = n25487 ^ n17623 ^ n12060 ;
  assign n25489 = ( n16640 & n25486 ) | ( n16640 & ~n25488 ) | ( n25486 & ~n25488 ) ;
  assign n25490 = n23642 ^ n20252 ^ n5141 ;
  assign n25491 = ( n18826 & n24982 ) | ( n18826 & ~n25490 ) | ( n24982 & ~n25490 ) ;
  assign n25492 = n17173 ^ n12510 ^ n5615 ;
  assign n25493 = n10820 ^ n9444 ^ 1'b0 ;
  assign n25497 = n5931 ^ n982 ^ n552 ;
  assign n25498 = n25497 ^ n5317 ^ n4302 ;
  assign n25494 = ( ~n1777 & n17866 ) | ( ~n1777 & n22764 ) | ( n17866 & n22764 ) ;
  assign n25495 = n25494 ^ n17992 ^ 1'b0 ;
  assign n25496 = n5746 & n25495 ;
  assign n25499 = n25498 ^ n25496 ^ n9012 ;
  assign n25500 = n8254 ^ n6843 ^ n3174 ;
  assign n25501 = n25500 ^ n17612 ^ n9354 ;
  assign n25502 = ( ~n4745 & n7913 ) | ( ~n4745 & n25501 ) | ( n7913 & n25501 ) ;
  assign n25503 = n25502 ^ n423 ^ 1'b0 ;
  assign n25504 = n6079 & n25503 ;
  assign n25505 = n23740 ^ n7750 ^ n6108 ;
  assign n25506 = n25505 ^ n22484 ^ 1'b0 ;
  assign n25507 = n20278 ^ n10674 ^ n6227 ;
  assign n25508 = n6935 | n13613 ;
  assign n25509 = n23173 | n25508 ;
  assign n25510 = n20952 ^ n19683 ^ n10643 ;
  assign n25511 = n25510 ^ n20746 ^ n16049 ;
  assign n25512 = ( ~n8269 & n20463 ) | ( ~n8269 & n21011 ) | ( n20463 & n21011 ) ;
  assign n25516 = n15385 ^ n4036 ^ 1'b0 ;
  assign n25517 = n19483 | n25516 ;
  assign n25518 = n25517 ^ n13919 ^ n8674 ;
  assign n25514 = n20133 ^ n11164 ^ n3214 ;
  assign n25513 = ( ~n1326 & n21011 ) | ( ~n1326 & n21917 ) | ( n21011 & n21917 ) ;
  assign n25515 = n25514 ^ n25513 ^ n19153 ;
  assign n25519 = n25518 ^ n25515 ^ n12305 ;
  assign n25520 = n8531 & n16982 ;
  assign n25521 = n5700 & n25520 ;
  assign n25522 = ( n19036 & n21112 ) | ( n19036 & ~n25521 ) | ( n21112 & ~n25521 ) ;
  assign n25523 = n13405 ^ n6407 ^ n946 ;
  assign n25524 = ~n2345 & n13927 ;
  assign n25525 = n25523 & n25524 ;
  assign n25529 = n5131 & ~n5817 ;
  assign n25530 = n20061 & n25529 ;
  assign n25526 = ( n622 & n3976 ) | ( n622 & ~n11711 ) | ( n3976 & ~n11711 ) ;
  assign n25527 = n675 & ~n25526 ;
  assign n25528 = n23697 & n25527 ;
  assign n25531 = n25530 ^ n25528 ^ n25514 ;
  assign n25532 = ( n3028 & ~n5693 ) | ( n3028 & n12760 ) | ( ~n5693 & n12760 ) ;
  assign n25536 = n13006 ^ n4088 ^ n2373 ;
  assign n25533 = n10553 & ~n20360 ;
  assign n25534 = ~n800 & n25533 ;
  assign n25535 = n15118 & ~n25534 ;
  assign n25537 = n25536 ^ n25535 ^ 1'b0 ;
  assign n25538 = ( n25167 & n25532 ) | ( n25167 & n25537 ) | ( n25532 & n25537 ) ;
  assign n25539 = n13110 ^ n9703 ^ n1434 ;
  assign n25540 = n11528 ^ n4907 ^ n1457 ;
  assign n25541 = ~n17916 & n25540 ;
  assign n25542 = ( ~n13852 & n14973 ) | ( ~n13852 & n25541 ) | ( n14973 & n25541 ) ;
  assign n25543 = n25542 ^ n16304 ^ x38 ;
  assign n25544 = ( n20351 & n25539 ) | ( n20351 & ~n25543 ) | ( n25539 & ~n25543 ) ;
  assign n25545 = n18744 ^ n16252 ^ n5591 ;
  assign n25546 = n22096 ^ n11583 ^ n8041 ;
  assign n25547 = ( ~n675 & n10350 ) | ( ~n675 & n11841 ) | ( n10350 & n11841 ) ;
  assign n25548 = n25547 ^ n23357 ^ n15572 ;
  assign n25549 = n25546 | n25548 ;
  assign n25550 = n25549 ^ n13943 ^ x202 ;
  assign n25551 = ~n12911 & n20295 ;
  assign n25552 = ( n12039 & n12492 ) | ( n12039 & ~n16491 ) | ( n12492 & ~n16491 ) ;
  assign n25553 = ( ~n10541 & n16449 ) | ( ~n10541 & n25552 ) | ( n16449 & n25552 ) ;
  assign n25554 = ( ~n7927 & n11516 ) | ( ~n7927 & n25553 ) | ( n11516 & n25553 ) ;
  assign n25555 = n25112 ^ n1813 ^ 1'b0 ;
  assign n25556 = n25554 & ~n25555 ;
  assign n25557 = n11815 ^ n6082 ^ 1'b0 ;
  assign n25558 = ~n1033 & n25557 ;
  assign n25559 = ( n9898 & ~n17174 ) | ( n9898 & n25558 ) | ( ~n17174 & n25558 ) ;
  assign n25560 = n25559 ^ n20514 ^ n12649 ;
  assign n25561 = n13427 ^ n2489 ^ 1'b0 ;
  assign n25562 = n25561 ^ n10776 ^ n7477 ;
  assign n25563 = n18588 ^ n12985 ^ n904 ;
  assign n25564 = ( n4121 & ~n25562 ) | ( n4121 & n25563 ) | ( ~n25562 & n25563 ) ;
  assign n25565 = n1009 | n19181 ;
  assign n25566 = n25565 ^ n13894 ^ n3325 ;
  assign n25567 = n25566 ^ n25534 ^ n8513 ;
  assign n25574 = n20781 ^ n14993 ^ n5752 ;
  assign n25573 = n23479 ^ n5395 ^ n4336 ;
  assign n25575 = n25574 ^ n25573 ^ n11735 ;
  assign n25576 = ( n12312 & n12617 ) | ( n12312 & ~n25575 ) | ( n12617 & ~n25575 ) ;
  assign n25570 = n20982 ^ n11164 ^ n6299 ;
  assign n25571 = ( ~n4509 & n8323 ) | ( ~n4509 & n12544 ) | ( n8323 & n12544 ) ;
  assign n25572 = ( n7820 & n25570 ) | ( n7820 & ~n25571 ) | ( n25570 & ~n25571 ) ;
  assign n25568 = n23223 ^ n1552 ^ 1'b0 ;
  assign n25569 = ( ~n17871 & n18764 ) | ( ~n17871 & n25568 ) | ( n18764 & n25568 ) ;
  assign n25577 = n25576 ^ n25572 ^ n25569 ;
  assign n25578 = n13171 ^ n11244 ^ n10832 ;
  assign n25579 = ( x190 & n3211 ) | ( x190 & ~n23879 ) | ( n3211 & ~n23879 ) ;
  assign n25580 = n22090 ^ n11030 ^ n8396 ;
  assign n25581 = ( n1880 & ~n24406 ) | ( n1880 & n25580 ) | ( ~n24406 & n25580 ) ;
  assign n25582 = ( n14555 & n25579 ) | ( n14555 & ~n25581 ) | ( n25579 & ~n25581 ) ;
  assign n25583 = n16855 ^ n7848 ^ n1180 ;
  assign n25584 = n25583 ^ n9807 ^ n8056 ;
  assign n25585 = n25584 ^ n16193 ^ n7588 ;
  assign n25586 = n17323 ^ n15201 ^ n15179 ;
  assign n25587 = n23238 ^ n10046 ^ n7385 ;
  assign n25588 = ( n5169 & ~n8044 ) | ( n5169 & n25587 ) | ( ~n8044 & n25587 ) ;
  assign n25589 = n13577 ^ n1442 ^ 1'b0 ;
  assign n25590 = n799 & n25589 ;
  assign n25591 = n25590 ^ n24442 ^ n3945 ;
  assign n25592 = ( ~n7719 & n14155 ) | ( ~n7719 & n14289 ) | ( n14155 & n14289 ) ;
  assign n25593 = n13733 ^ n4355 ^ 1'b0 ;
  assign n25594 = n25593 ^ n18090 ^ 1'b0 ;
  assign n25595 = ( n25591 & n25592 ) | ( n25591 & ~n25594 ) | ( n25592 & ~n25594 ) ;
  assign n25596 = ( n2380 & ~n21431 ) | ( n2380 & n22753 ) | ( ~n21431 & n22753 ) ;
  assign n25597 = n25596 ^ n16916 ^ n13764 ;
  assign n25598 = ( n5462 & n9514 ) | ( n5462 & ~n23934 ) | ( n9514 & ~n23934 ) ;
  assign n25599 = ( n24858 & n25541 ) | ( n24858 & ~n25598 ) | ( n25541 & ~n25598 ) ;
  assign n25600 = n25597 & n25599 ;
  assign n25601 = n25600 ^ n19447 ^ 1'b0 ;
  assign n25602 = ( n1035 & n2952 ) | ( n1035 & n5849 ) | ( n2952 & n5849 ) ;
  assign n25603 = ( ~n20608 & n24531 ) | ( ~n20608 & n25602 ) | ( n24531 & n25602 ) ;
  assign n25604 = n6686 ^ n1448 ^ n1065 ;
  assign n25605 = n25604 ^ n18999 ^ n5150 ;
  assign n25606 = ( n24360 & n25603 ) | ( n24360 & n25605 ) | ( n25603 & n25605 ) ;
  assign n25607 = n18653 ^ n7465 ^ n3680 ;
  assign n25608 = ( n6142 & n13428 ) | ( n6142 & n25607 ) | ( n13428 & n25607 ) ;
  assign n25609 = n25608 ^ n24461 ^ n5395 ;
  assign n25612 = n7808 & ~n16291 ;
  assign n25610 = n8210 ^ n2325 ^ 1'b0 ;
  assign n25611 = ( n12915 & n15693 ) | ( n12915 & n25610 ) | ( n15693 & n25610 ) ;
  assign n25613 = n25612 ^ n25611 ^ n6273 ;
  assign n25624 = n22729 ^ n21690 ^ n10070 ;
  assign n25619 = n21447 ^ n11505 ^ n3470 ;
  assign n25620 = n4863 & n25619 ;
  assign n25621 = n25620 ^ n11767 ^ 1'b0 ;
  assign n25622 = n25621 ^ n10226 ^ n1566 ;
  assign n25623 = ( ~n4941 & n5460 ) | ( ~n4941 & n25622 ) | ( n5460 & n25622 ) ;
  assign n25614 = ( x22 & ~n7123 ) | ( x22 & n19253 ) | ( ~n7123 & n19253 ) ;
  assign n25615 = n6934 ^ n3105 ^ 1'b0 ;
  assign n25616 = n18876 | n25615 ;
  assign n25617 = ( ~n1716 & n11065 ) | ( ~n1716 & n25616 ) | ( n11065 & n25616 ) ;
  assign n25618 = ( n990 & ~n25614 ) | ( n990 & n25617 ) | ( ~n25614 & n25617 ) ;
  assign n25625 = n25624 ^ n25623 ^ n25618 ;
  assign n25626 = ( n5891 & ~n22218 ) | ( n5891 & n22593 ) | ( ~n22218 & n22593 ) ;
  assign n25627 = n25626 ^ n12974 ^ n2350 ;
  assign n25628 = ~n3228 & n7176 ;
  assign n25629 = n25628 ^ n6816 ^ 1'b0 ;
  assign n25630 = ( n20293 & n22655 ) | ( n20293 & n25629 ) | ( n22655 & n25629 ) ;
  assign n25631 = ( n5021 & n8232 ) | ( n5021 & n11397 ) | ( n8232 & n11397 ) ;
  assign n25632 = n25631 ^ n12922 ^ n1181 ;
  assign n25633 = n6945 & n25632 ;
  assign n25634 = n13365 ^ n10753 ^ 1'b0 ;
  assign n25635 = ( n25630 & n25633 ) | ( n25630 & n25634 ) | ( n25633 & n25634 ) ;
  assign n25639 = n9048 ^ x164 ^ 1'b0 ;
  assign n25640 = n25639 ^ n21792 ^ n1746 ;
  assign n25636 = n7306 ^ n5574 ^ n4569 ;
  assign n25637 = ( n5283 & n20736 ) | ( n5283 & n25636 ) | ( n20736 & n25636 ) ;
  assign n25638 = n25637 ^ n23479 ^ n13771 ;
  assign n25641 = n25640 ^ n25638 ^ n11752 ;
  assign n25642 = n3473 & ~n18205 ;
  assign n25643 = ~n8914 & n25642 ;
  assign n25644 = n6422 | n20106 ;
  assign n25645 = n25644 ^ n5058 ^ 1'b0 ;
  assign n25646 = n25645 ^ n16940 ^ n9044 ;
  assign n25647 = n3908 ^ n3401 ^ x163 ;
  assign n25648 = n25647 ^ n571 ^ 1'b0 ;
  assign n25649 = ( n5926 & ~n15275 ) | ( n5926 & n25648 ) | ( ~n15275 & n25648 ) ;
  assign n25650 = ( n4707 & n6233 ) | ( n4707 & ~n21547 ) | ( n6233 & ~n21547 ) ;
  assign n25652 = ( n1651 & n5733 ) | ( n1651 & n21748 ) | ( n5733 & n21748 ) ;
  assign n25651 = n18295 ^ n7652 ^ n413 ;
  assign n25653 = n25652 ^ n25651 ^ n9200 ;
  assign n25654 = ( n21488 & n25650 ) | ( n21488 & n25653 ) | ( n25650 & n25653 ) ;
  assign n25656 = ( n1547 & n9912 ) | ( n1547 & n13106 ) | ( n9912 & n13106 ) ;
  assign n25655 = n11059 | n17563 ;
  assign n25657 = n25656 ^ n25655 ^ 1'b0 ;
  assign n25658 = ~n13067 & n20345 ;
  assign n25659 = ( n2289 & n22852 ) | ( n2289 & ~n25658 ) | ( n22852 & ~n25658 ) ;
  assign n25660 = n15758 & n24110 ;
  assign n25661 = n21359 ^ n11776 ^ n7436 ;
  assign n25662 = n25661 ^ n24082 ^ 1'b0 ;
  assign n25663 = ( n7171 & n7313 ) | ( n7171 & ~n8429 ) | ( n7313 & ~n8429 ) ;
  assign n25664 = ( n6273 & ~n10145 ) | ( n6273 & n25663 ) | ( ~n10145 & n25663 ) ;
  assign n25665 = ~n17308 & n25664 ;
  assign n25666 = n18157 & n25665 ;
  assign n25667 = ( ~n1945 & n3523 ) | ( ~n1945 & n6174 ) | ( n3523 & n6174 ) ;
  assign n25668 = ( n1780 & ~n15460 ) | ( n1780 & n25667 ) | ( ~n15460 & n25667 ) ;
  assign n25669 = n25668 ^ n22218 ^ n6549 ;
  assign n25670 = n17893 & n25669 ;
  assign n25671 = ~n2220 & n25670 ;
  assign n25672 = n14478 & n25671 ;
  assign n25673 = n25672 ^ n16650 ^ n1011 ;
  assign n25674 = n25673 ^ n2738 ^ 1'b0 ;
  assign n25675 = ( ~n24608 & n25666 ) | ( ~n24608 & n25674 ) | ( n25666 & n25674 ) ;
  assign n25676 = ( ~n3216 & n6567 ) | ( ~n3216 & n16259 ) | ( n6567 & n16259 ) ;
  assign n25677 = n14330 ^ n3133 ^ 1'b0 ;
  assign n25678 = n4833 | n25677 ;
  assign n25679 = ( n24718 & n25676 ) | ( n24718 & n25678 ) | ( n25676 & n25678 ) ;
  assign n25680 = ( n11120 & ~n20645 ) | ( n11120 & n25679 ) | ( ~n20645 & n25679 ) ;
  assign n25681 = n18749 ^ n9803 ^ n1893 ;
  assign n25682 = n14136 & n25681 ;
  assign n25683 = n25682 ^ n9380 ^ 1'b0 ;
  assign n25684 = n25683 ^ n3140 ^ 1'b0 ;
  assign n25685 = n14878 & n23908 ;
  assign n25686 = n25684 & n25685 ;
  assign n25687 = n3639 & ~n8345 ;
  assign n25688 = ( n4215 & n10946 ) | ( n4215 & n25687 ) | ( n10946 & n25687 ) ;
  assign n25689 = n25688 ^ n20776 ^ n768 ;
  assign n25690 = n22583 ^ n11803 ^ n9681 ;
  assign n25691 = ( ~n2566 & n25689 ) | ( ~n2566 & n25690 ) | ( n25689 & n25690 ) ;
  assign n25692 = ( ~n10367 & n25686 ) | ( ~n10367 & n25691 ) | ( n25686 & n25691 ) ;
  assign n25693 = ( n11853 & ~n25680 ) | ( n11853 & n25692 ) | ( ~n25680 & n25692 ) ;
  assign n25696 = n19808 ^ n17740 ^ n4133 ;
  assign n25694 = ( n3981 & ~n6591 ) | ( n3981 & n6689 ) | ( ~n6591 & n6689 ) ;
  assign n25695 = ( n1471 & n2218 ) | ( n1471 & ~n25694 ) | ( n2218 & ~n25694 ) ;
  assign n25697 = n25696 ^ n25695 ^ x171 ;
  assign n25699 = n7012 ^ n3342 ^ n2350 ;
  assign n25698 = n23899 ^ n20653 ^ n10057 ;
  assign n25700 = n25699 ^ n25698 ^ n4510 ;
  assign n25701 = ( n8172 & ~n17284 ) | ( n8172 & n23608 ) | ( ~n17284 & n23608 ) ;
  assign n25702 = n25701 ^ n10099 ^ n6648 ;
  assign n25703 = n17519 ^ n13582 ^ n2006 ;
  assign n25704 = n3958 & ~n4363 ;
  assign n25705 = n18916 & ~n25704 ;
  assign n25706 = n25703 & n25705 ;
  assign n25707 = x14 | n25706 ;
  assign n25717 = n24848 ^ n21310 ^ n4215 ;
  assign n25713 = ( x188 & n5163 ) | ( x188 & ~n5165 ) | ( n5163 & ~n5165 ) ;
  assign n25714 = ( n3802 & ~n14919 ) | ( n3802 & n25713 ) | ( ~n14919 & n25713 ) ;
  assign n25711 = n14218 ^ n1330 ^ 1'b0 ;
  assign n25712 = ~n12331 & n25711 ;
  assign n25708 = n24148 ^ n10710 ^ n3705 ;
  assign n25709 = n25708 ^ n10224 ^ n6795 ;
  assign n25710 = ( n9391 & n14685 ) | ( n9391 & ~n25709 ) | ( n14685 & ~n25709 ) ;
  assign n25715 = n25714 ^ n25712 ^ n25710 ;
  assign n25716 = x79 & ~n25715 ;
  assign n25718 = n25717 ^ n25716 ^ 1'b0 ;
  assign n25720 = ~n5421 & n14192 ;
  assign n25721 = n13665 & n25720 ;
  assign n25719 = n10746 ^ n10111 ^ 1'b0 ;
  assign n25722 = n25721 ^ n25719 ^ n7018 ;
  assign n25723 = n25722 ^ n23556 ^ 1'b0 ;
  assign n25724 = n4948 & n25723 ;
  assign n25725 = ( ~n400 & n20403 ) | ( ~n400 & n25724 ) | ( n20403 & n25724 ) ;
  assign n25726 = n20272 ^ n19991 ^ n4930 ;
  assign n25727 = ( n4390 & ~n25725 ) | ( n4390 & n25726 ) | ( ~n25725 & n25726 ) ;
  assign n25728 = n24506 ^ n13530 ^ n8772 ;
  assign n25729 = n12443 ^ n6097 ^ n2272 ;
  assign n25730 = n14964 ^ n3779 ^ n3530 ;
  assign n25731 = ( n3085 & n25729 ) | ( n3085 & ~n25730 ) | ( n25729 & ~n25730 ) ;
  assign n25732 = ( ~x238 & n19351 ) | ( ~x238 & n25731 ) | ( n19351 & n25731 ) ;
  assign n25735 = n15471 ^ n8441 ^ n565 ;
  assign n25733 = ( n2741 & ~n3035 ) | ( n2741 & n3267 ) | ( ~n3035 & n3267 ) ;
  assign n25734 = n2241 | n25733 ;
  assign n25736 = n25735 ^ n25734 ^ 1'b0 ;
  assign n25737 = ( n25728 & n25732 ) | ( n25728 & ~n25736 ) | ( n25732 & ~n25736 ) ;
  assign n25744 = n13982 ^ n7298 ^ n5239 ;
  assign n25745 = ( ~n473 & n8526 ) | ( ~n473 & n25744 ) | ( n8526 & n25744 ) ;
  assign n25740 = n2237 | n11014 ;
  assign n25741 = ( n5264 & n6001 ) | ( n5264 & n8627 ) | ( n6001 & n8627 ) ;
  assign n25742 = ( n10105 & n25740 ) | ( n10105 & ~n25741 ) | ( n25740 & ~n25741 ) ;
  assign n25739 = n6119 ^ n375 ^ 1'b0 ;
  assign n25738 = n24850 ^ n10505 ^ n7444 ;
  assign n25743 = n25742 ^ n25739 ^ n25738 ;
  assign n25746 = n25745 ^ n25743 ^ n687 ;
  assign n25747 = ( n1987 & ~n7046 ) | ( n1987 & n10421 ) | ( ~n7046 & n10421 ) ;
  assign n25748 = ( n5128 & n9465 ) | ( n5128 & ~n25747 ) | ( n9465 & ~n25747 ) ;
  assign n25749 = ( n2218 & ~n8487 ) | ( n2218 & n12545 ) | ( ~n8487 & n12545 ) ;
  assign n25750 = ( n3178 & n11885 ) | ( n3178 & ~n21606 ) | ( n11885 & ~n21606 ) ;
  assign n25751 = ( n25748 & n25749 ) | ( n25748 & ~n25750 ) | ( n25749 & ~n25750 ) ;
  assign n25752 = n20964 ^ n15215 ^ x55 ;
  assign n25754 = ( n3640 & n6849 ) | ( n3640 & ~n10187 ) | ( n6849 & ~n10187 ) ;
  assign n25753 = ( n793 & ~n3866 ) | ( n793 & n23226 ) | ( ~n3866 & n23226 ) ;
  assign n25755 = n25754 ^ n25753 ^ 1'b0 ;
  assign n25756 = n25752 & ~n25755 ;
  assign n25757 = n17449 ^ n5338 ^ 1'b0 ;
  assign n25763 = ( n1684 & n3224 ) | ( n1684 & ~n7396 ) | ( n3224 & ~n7396 ) ;
  assign n25762 = n14456 ^ n14397 ^ n5496 ;
  assign n25758 = n15669 ^ n647 ^ 1'b0 ;
  assign n25759 = ~n21207 & n25758 ;
  assign n25760 = n25759 ^ n19110 ^ n2226 ;
  assign n25761 = ( n1816 & n8078 ) | ( n1816 & n25760 ) | ( n8078 & n25760 ) ;
  assign n25764 = n25763 ^ n25762 ^ n25761 ;
  assign n25765 = n17734 ^ n15366 ^ n4508 ;
  assign n25766 = n20112 ^ n18872 ^ n8073 ;
  assign n25767 = n25766 ^ n14196 ^ n8901 ;
  assign n25768 = n8699 & ~n25767 ;
  assign n25769 = n24300 ^ n17777 ^ n12492 ;
  assign n25770 = ( x129 & n1696 ) | ( x129 & n7972 ) | ( n1696 & n7972 ) ;
  assign n25771 = n25770 ^ n17501 ^ n680 ;
  assign n25772 = n12994 ^ n4229 ^ n3200 ;
  assign n25773 = ( n5181 & ~n8163 ) | ( n5181 & n25772 ) | ( ~n8163 & n25772 ) ;
  assign n25774 = n23793 ^ n17513 ^ n816 ;
  assign n25782 = n15346 ^ n7030 ^ n3326 ;
  assign n25775 = n9766 & n24839 ;
  assign n25776 = ~n5921 & n25775 ;
  assign n25777 = ( ~n5248 & n8097 ) | ( ~n5248 & n9670 ) | ( n8097 & n9670 ) ;
  assign n25778 = ( n7202 & n25517 ) | ( n7202 & ~n25777 ) | ( n25517 & ~n25777 ) ;
  assign n25779 = n25778 ^ n23722 ^ n12415 ;
  assign n25780 = n25779 ^ n23934 ^ n13225 ;
  assign n25781 = ( ~n2094 & n25776 ) | ( ~n2094 & n25780 ) | ( n25776 & n25780 ) ;
  assign n25783 = n25782 ^ n25781 ^ n11139 ;
  assign n25784 = ( n11640 & n15150 ) | ( n11640 & n25783 ) | ( n15150 & n25783 ) ;
  assign n25785 = n14194 ^ n665 ^ 1'b0 ;
  assign n25786 = n25785 ^ n22151 ^ n11538 ;
  assign n25787 = ( n8947 & ~n10814 ) | ( n8947 & n25786 ) | ( ~n10814 & n25786 ) ;
  assign n25788 = ( n13762 & ~n18177 ) | ( n13762 & n24939 ) | ( ~n18177 & n24939 ) ;
  assign n25789 = ( n10422 & ~n18409 ) | ( n10422 & n25788 ) | ( ~n18409 & n25788 ) ;
  assign n25790 = n17334 ^ n14162 ^ n7003 ;
  assign n25792 = ( ~x223 & n5848 ) | ( ~x223 & n7780 ) | ( n5848 & n7780 ) ;
  assign n25791 = n20759 ^ n14675 ^ n2737 ;
  assign n25793 = n25792 ^ n25791 ^ n6690 ;
  assign n25794 = ( n14129 & ~n25790 ) | ( n14129 & n25793 ) | ( ~n25790 & n25793 ) ;
  assign n25795 = x185 & ~n4852 ;
  assign n25796 = n25795 ^ n7738 ^ 1'b0 ;
  assign n25797 = ( n5859 & ~n15708 ) | ( n5859 & n25796 ) | ( ~n15708 & n25796 ) ;
  assign n25798 = ( n8870 & ~n16134 ) | ( n8870 & n21367 ) | ( ~n16134 & n21367 ) ;
  assign n25799 = n25798 ^ n18634 ^ n2347 ;
  assign n25800 = n25799 ^ n21171 ^ n520 ;
  assign n25802 = n8699 ^ n8259 ^ n6960 ;
  assign n25801 = n873 | n8931 ;
  assign n25803 = n25802 ^ n25801 ^ 1'b0 ;
  assign n25804 = ( n8692 & n13592 ) | ( n8692 & n19398 ) | ( n13592 & n19398 ) ;
  assign n25805 = ( n15985 & n25803 ) | ( n15985 & n25804 ) | ( n25803 & n25804 ) ;
  assign n25806 = ( n760 & n6373 ) | ( n760 & n11963 ) | ( n6373 & n11963 ) ;
  assign n25807 = n25806 ^ n17097 ^ n1606 ;
  assign n25808 = n9857 ^ n9050 ^ x12 ;
  assign n25809 = n13352 ^ n12914 ^ n9266 ;
  assign n25810 = ( n8873 & n18487 ) | ( n8873 & ~n25809 ) | ( n18487 & ~n25809 ) ;
  assign n25811 = n19937 ^ n13738 ^ n7123 ;
  assign n25812 = n25811 ^ n10813 ^ 1'b0 ;
  assign n25813 = n17912 & ~n25812 ;
  assign n25814 = ( n6795 & n25810 ) | ( n6795 & n25813 ) | ( n25810 & n25813 ) ;
  assign n25818 = ( ~n11841 & n21862 ) | ( ~n11841 & n25722 ) | ( n21862 & n25722 ) ;
  assign n25815 = n18738 ^ n12960 ^ n9488 ;
  assign n25816 = n25815 ^ n25574 ^ n5882 ;
  assign n25817 = n25816 ^ n19806 ^ n1396 ;
  assign n25819 = n25818 ^ n25817 ^ 1'b0 ;
  assign n25822 = ( n4608 & n11363 ) | ( n4608 & n11795 ) | ( n11363 & n11795 ) ;
  assign n25823 = ( ~n1637 & n3232 ) | ( ~n1637 & n25822 ) | ( n3232 & n25822 ) ;
  assign n25824 = ( n837 & n12810 ) | ( n837 & n25823 ) | ( n12810 & n25823 ) ;
  assign n25820 = ( n810 & n1804 ) | ( n810 & ~n2567 ) | ( n1804 & ~n2567 ) ;
  assign n25821 = n25820 ^ n8401 ^ n416 ;
  assign n25825 = n25824 ^ n25821 ^ n1729 ;
  assign n25826 = n25825 ^ n21871 ^ n2905 ;
  assign n25827 = n13031 ^ n9650 ^ n6025 ;
  assign n25831 = ( n7274 & n11806 ) | ( n7274 & n20589 ) | ( n11806 & n20589 ) ;
  assign n25828 = ( x183 & n1711 ) | ( x183 & ~n7725 ) | ( n1711 & ~n7725 ) ;
  assign n25829 = ( n2695 & ~n3914 ) | ( n2695 & n4681 ) | ( ~n3914 & n4681 ) ;
  assign n25830 = ( n2134 & n25828 ) | ( n2134 & ~n25829 ) | ( n25828 & ~n25829 ) ;
  assign n25832 = n25831 ^ n25830 ^ n22136 ;
  assign n25833 = ( n5817 & ~n15057 ) | ( n5817 & n25832 ) | ( ~n15057 & n25832 ) ;
  assign n25836 = ( x8 & n5499 ) | ( x8 & ~n13090 ) | ( n5499 & ~n13090 ) ;
  assign n25834 = ( n6648 & ~n15674 ) | ( n6648 & n16337 ) | ( ~n15674 & n16337 ) ;
  assign n25835 = n22168 & n25834 ;
  assign n25837 = n25836 ^ n25835 ^ 1'b0 ;
  assign n25838 = ( ~n1991 & n12956 ) | ( ~n1991 & n21293 ) | ( n12956 & n21293 ) ;
  assign n25839 = ( ~n4322 & n4366 ) | ( ~n4322 & n20619 ) | ( n4366 & n20619 ) ;
  assign n25840 = n22163 & n25839 ;
  assign n25841 = ( n7010 & n14584 ) | ( n7010 & n25840 ) | ( n14584 & n25840 ) ;
  assign n25842 = n6090 ^ n3923 ^ n327 ;
  assign n25843 = n1575 | n25842 ;
  assign n25844 = n25843 ^ n20791 ^ n15265 ;
  assign n25845 = n25844 ^ n10554 ^ 1'b0 ;
  assign n25848 = ( ~n2841 & n4539 ) | ( ~n2841 & n15329 ) | ( n4539 & n15329 ) ;
  assign n25849 = n24182 & n25848 ;
  assign n25846 = n22164 ^ n11657 ^ n11635 ;
  assign n25847 = ~n6636 & n25846 ;
  assign n25850 = n25849 ^ n25847 ^ 1'b0 ;
  assign n25851 = n2771 ^ n2220 ^ n955 ;
  assign n25852 = n25851 ^ n16790 ^ n7967 ;
  assign n25853 = n25852 ^ n14917 ^ n8608 ;
  assign n25854 = ( n15996 & n20299 ) | ( n15996 & n25853 ) | ( n20299 & n25853 ) ;
  assign n25859 = n13740 ^ n3650 ^ 1'b0 ;
  assign n25860 = n25859 ^ n12468 ^ 1'b0 ;
  assign n25861 = n25860 ^ n8972 ^ n7015 ;
  assign n25857 = n15211 ^ n4258 ^ n4221 ;
  assign n25855 = ( n3576 & n5741 ) | ( n3576 & n10939 ) | ( n5741 & n10939 ) ;
  assign n25856 = n25855 ^ n23517 ^ 1'b0 ;
  assign n25858 = n25857 ^ n25856 ^ n11471 ;
  assign n25862 = n25861 ^ n25858 ^ n8269 ;
  assign n25863 = n21647 ^ n18946 ^ n11501 ;
  assign n25864 = n25863 ^ n2378 ^ 1'b0 ;
  assign n25865 = n10433 | n25864 ;
  assign n25866 = n1716 & ~n25865 ;
  assign n25867 = n22568 ^ n7891 ^ n2613 ;
  assign n25868 = ( ~n3294 & n10487 ) | ( ~n3294 & n25867 ) | ( n10487 & n25867 ) ;
  assign n25869 = n25868 ^ n24083 ^ n22615 ;
  assign n25870 = n25869 ^ n14851 ^ n384 ;
  assign n25871 = n23545 ^ n21970 ^ n8216 ;
  assign n25872 = ( n502 & n12176 ) | ( n502 & n25871 ) | ( n12176 & n25871 ) ;
  assign n25873 = ( n5822 & n6095 ) | ( n5822 & n16006 ) | ( n6095 & n16006 ) ;
  assign n25874 = ( n14625 & n19315 ) | ( n14625 & ~n24473 ) | ( n19315 & ~n24473 ) ;
  assign n25875 = ( ~n16542 & n24694 ) | ( ~n16542 & n25874 ) | ( n24694 & n25874 ) ;
  assign n25887 = ( ~n1111 & n1325 ) | ( ~n1111 & n11590 ) | ( n1325 & n11590 ) ;
  assign n25888 = ~n24349 & n25887 ;
  assign n25876 = n13401 ^ n9942 ^ x4 ;
  assign n25877 = n11192 | n25876 ;
  assign n25878 = n488 | n25877 ;
  assign n25879 = ( ~n585 & n4655 ) | ( ~n585 & n6115 ) | ( n4655 & n6115 ) ;
  assign n25880 = n11569 ^ n7418 ^ n831 ;
  assign n25881 = n4915 | n25880 ;
  assign n25882 = n25274 | n25881 ;
  assign n25883 = ( n19281 & n25879 ) | ( n19281 & ~n25882 ) | ( n25879 & ~n25882 ) ;
  assign n25884 = n25883 ^ n7881 ^ 1'b0 ;
  assign n25885 = n4261 & n25884 ;
  assign n25886 = ( n4640 & n25878 ) | ( n4640 & ~n25885 ) | ( n25878 & ~n25885 ) ;
  assign n25889 = n25888 ^ n25886 ^ n11194 ;
  assign n25896 = ( n5028 & n16435 ) | ( n5028 & ~n25749 ) | ( n16435 & ~n25749 ) ;
  assign n25890 = ~n2014 & n15215 ;
  assign n25891 = n25890 ^ n5169 ^ 1'b0 ;
  assign n25892 = n25891 ^ n13291 ^ n3265 ;
  assign n25893 = n25892 ^ n22468 ^ n6788 ;
  assign n25894 = ( n10546 & n17720 ) | ( n10546 & n20473 ) | ( n17720 & n20473 ) ;
  assign n25895 = ( ~n12045 & n25893 ) | ( ~n12045 & n25894 ) | ( n25893 & n25894 ) ;
  assign n25897 = n25896 ^ n25895 ^ n578 ;
  assign n25898 = ( ~n4669 & n23220 ) | ( ~n4669 & n25897 ) | ( n23220 & n25897 ) ;
  assign n25899 = n10339 & ~n11155 ;
  assign n25900 = n24566 & n25899 ;
  assign n25901 = n25900 ^ n6699 ^ n1154 ;
  assign n25902 = x77 & n25901 ;
  assign n25903 = n25902 ^ n8975 ^ 1'b0 ;
  assign n25904 = ~n868 & n2166 ;
  assign n25905 = n25904 ^ n3494 ^ 1'b0 ;
  assign n25906 = n25905 ^ n24442 ^ n4033 ;
  assign n25907 = n17184 ^ n14901 ^ n9616 ;
  assign n25908 = n1457 & n25907 ;
  assign n25909 = ~n25906 & n25908 ;
  assign n25910 = n6496 ^ n2204 ^ n1985 ;
  assign n25911 = n25910 ^ n2086 ^ 1'b0 ;
  assign n25912 = ( n13364 & n13734 ) | ( n13364 & ~n25911 ) | ( n13734 & ~n25911 ) ;
  assign n25913 = ( n5220 & ~n5751 ) | ( n5220 & n20869 ) | ( ~n5751 & n20869 ) ;
  assign n25914 = n9554 ^ n6878 ^ n4065 ;
  assign n25922 = ( n14898 & n20554 ) | ( n14898 & ~n22692 ) | ( n20554 & ~n22692 ) ;
  assign n25915 = ( ~n3121 & n10713 ) | ( ~n3121 & n13817 ) | ( n10713 & n13817 ) ;
  assign n25918 = n6182 ^ n4370 ^ 1'b0 ;
  assign n25919 = n25918 ^ n17365 ^ n13947 ;
  assign n25916 = n10159 ^ n5060 ^ n2045 ;
  assign n25917 = ( ~n4401 & n8724 ) | ( ~n4401 & n25916 ) | ( n8724 & n25916 ) ;
  assign n25920 = n25919 ^ n25917 ^ n16325 ;
  assign n25921 = ( n11924 & ~n25915 ) | ( n11924 & n25920 ) | ( ~n25915 & n25920 ) ;
  assign n25923 = n25922 ^ n25921 ^ n1056 ;
  assign n25924 = ( n16109 & n25914 ) | ( n16109 & n25923 ) | ( n25914 & n25923 ) ;
  assign n25925 = n21494 ^ n15219 ^ n1201 ;
  assign n25927 = n8799 ^ x46 ^ 1'b0 ;
  assign n25928 = n5767 | n25927 ;
  assign n25926 = n15888 ^ n14629 ^ n1905 ;
  assign n25929 = n25928 ^ n25926 ^ x72 ;
  assign n25930 = n15654 ^ n7842 ^ n7698 ;
  assign n25931 = n23078 ^ n20759 ^ n6690 ;
  assign n25932 = ( n2895 & n25930 ) | ( n2895 & ~n25931 ) | ( n25930 & ~n25931 ) ;
  assign n25933 = ( n1316 & n1349 ) | ( n1316 & ~n18016 ) | ( n1349 & ~n18016 ) ;
  assign n25934 = ~n7044 & n25933 ;
  assign n25935 = n25934 ^ n20605 ^ 1'b0 ;
  assign n25942 = ( n9748 & n18077 ) | ( n9748 & n20929 ) | ( n18077 & n20929 ) ;
  assign n25943 = n25942 ^ n16141 ^ 1'b0 ;
  assign n25944 = n3901 & n25943 ;
  assign n25938 = n13151 ^ n7319 ^ 1'b0 ;
  assign n25939 = n9790 | n25938 ;
  assign n25940 = n25939 ^ n2902 ^ n2305 ;
  assign n25936 = n6558 | n21687 ;
  assign n25937 = n18926 & ~n25936 ;
  assign n25941 = n25940 ^ n25937 ^ n25244 ;
  assign n25945 = n25944 ^ n25941 ^ n25667 ;
  assign n25946 = n23286 ^ n17411 ^ n6816 ;
  assign n25947 = n20152 ^ n17905 ^ n10764 ;
  assign n25948 = n23948 & n25947 ;
  assign n25949 = n23604 ^ n9323 ^ 1'b0 ;
  assign n25950 = n12943 & ~n25949 ;
  assign n25951 = ( n3756 & ~n4636 ) | ( n3756 & n25427 ) | ( ~n4636 & n25427 ) ;
  assign n25952 = n17334 ^ n12268 ^ n8607 ;
  assign n25953 = ( n10241 & n13481 ) | ( n10241 & n15290 ) | ( n13481 & n15290 ) ;
  assign n25954 = ( ~n2474 & n25952 ) | ( ~n2474 & n25953 ) | ( n25952 & n25953 ) ;
  assign n25955 = n12842 ^ n10379 ^ n6969 ;
  assign n25956 = n2428 & n8378 ;
  assign n25957 = n2306 | n25956 ;
  assign n25958 = n25957 ^ n22696 ^ n10054 ;
  assign n25959 = n25958 ^ n11164 ^ x0 ;
  assign n25960 = ( ~n5628 & n14295 ) | ( ~n5628 & n14653 ) | ( n14295 & n14653 ) ;
  assign n25961 = n25960 ^ n14565 ^ n10650 ;
  assign n25962 = ( ~n6433 & n10420 ) | ( ~n6433 & n16239 ) | ( n10420 & n16239 ) ;
  assign n25963 = ( ~n8220 & n10880 ) | ( ~n8220 & n25962 ) | ( n10880 & n25962 ) ;
  assign n25964 = ( n20420 & n22554 ) | ( n20420 & n25963 ) | ( n22554 & n25963 ) ;
  assign n25965 = n25729 ^ n23183 ^ n4005 ;
  assign n25966 = ( ~n9327 & n11490 ) | ( ~n9327 & n12396 ) | ( n11490 & n12396 ) ;
  assign n25967 = n6633 ^ n1545 ^ 1'b0 ;
  assign n25968 = n25966 | n25967 ;
  assign n25969 = n25968 ^ x142 ^ 1'b0 ;
  assign n25970 = n25969 ^ n21784 ^ n8789 ;
  assign n25971 = ( ~n13703 & n25965 ) | ( ~n13703 & n25970 ) | ( n25965 & n25970 ) ;
  assign n25972 = ( ~n10484 & n20493 ) | ( ~n10484 & n25971 ) | ( n20493 & n25971 ) ;
  assign n25973 = n25465 ^ n5141 ^ n2516 ;
  assign n25974 = ( n565 & n25048 ) | ( n565 & n25973 ) | ( n25048 & n25973 ) ;
  assign n25975 = ( n8096 & ~n17122 ) | ( n8096 & n19545 ) | ( ~n17122 & n19545 ) ;
  assign n25976 = n25975 ^ n18709 ^ n6858 ;
  assign n25977 = ( ~n11216 & n18057 ) | ( ~n11216 & n22263 ) | ( n18057 & n22263 ) ;
  assign n25978 = n10671 ^ n7287 ^ 1'b0 ;
  assign n25979 = n25977 | n25978 ;
  assign n25980 = n16522 ^ n2809 ^ 1'b0 ;
  assign n25981 = ( n10600 & n14320 ) | ( n10600 & n15313 ) | ( n14320 & n15313 ) ;
  assign n25982 = n25981 ^ n24193 ^ n3158 ;
  assign n25983 = n25982 ^ n22411 ^ n6227 ;
  assign n25984 = ( n8567 & n11368 ) | ( n8567 & n24102 ) | ( n11368 & n24102 ) ;
  assign n25985 = ( n9682 & n20491 ) | ( n9682 & ~n25984 ) | ( n20491 & ~n25984 ) ;
  assign n25986 = ( n3409 & n4308 ) | ( n3409 & n16094 ) | ( n4308 & n16094 ) ;
  assign n25987 = n25986 ^ n19582 ^ n2749 ;
  assign n25988 = n1051 & ~n5667 ;
  assign n25989 = ( n1527 & n14730 ) | ( n1527 & n25988 ) | ( n14730 & n25988 ) ;
  assign n25990 = ( n13807 & ~n20059 ) | ( n13807 & n23300 ) | ( ~n20059 & n23300 ) ;
  assign n25991 = n22725 ^ n18587 ^ n5057 ;
  assign n25992 = ( n1594 & ~n5116 ) | ( n1594 & n12974 ) | ( ~n5116 & n12974 ) ;
  assign n25993 = n25992 ^ n18004 ^ 1'b0 ;
  assign n25994 = n1969 & ~n25993 ;
  assign n25995 = ( n2254 & n3439 ) | ( n2254 & n3818 ) | ( n3439 & n3818 ) ;
  assign n25996 = ( n9575 & n9683 ) | ( n9575 & ~n22140 ) | ( n9683 & ~n22140 ) ;
  assign n25997 = n21981 ^ n10940 ^ 1'b0 ;
  assign n25998 = ( n25995 & n25996 ) | ( n25995 & ~n25997 ) | ( n25996 & ~n25997 ) ;
  assign n25999 = ( n3525 & n11431 ) | ( n3525 & n18719 ) | ( n11431 & n18719 ) ;
  assign n26000 = n8225 ^ n1053 ^ x101 ;
  assign n26001 = n26000 ^ n1522 ^ 1'b0 ;
  assign n26002 = n3717 | n26001 ;
  assign n26003 = n26002 ^ n18408 ^ n1276 ;
  assign n26004 = ( n3751 & n25490 ) | ( n3751 & ~n26003 ) | ( n25490 & ~n26003 ) ;
  assign n26005 = n4879 | n8065 ;
  assign n26006 = n26005 ^ n1232 ^ 1'b0 ;
  assign n26007 = n26006 ^ n2834 ^ n806 ;
  assign n26008 = n26007 ^ n18268 ^ 1'b0 ;
  assign n26009 = n20183 & ~n26008 ;
  assign n26010 = n17877 ^ n4958 ^ 1'b0 ;
  assign n26011 = ( ~n13970 & n16284 ) | ( ~n13970 & n26010 ) | ( n16284 & n26010 ) ;
  assign n26012 = n24857 ^ n19525 ^ n431 ;
  assign n26013 = ( ~n5042 & n26011 ) | ( ~n5042 & n26012 ) | ( n26011 & n26012 ) ;
  assign n26014 = n26013 ^ n19917 ^ n13981 ;
  assign n26015 = n1665 & n14304 ;
  assign n26016 = n26015 ^ n19763 ^ 1'b0 ;
  assign n26017 = n15758 ^ n10361 ^ 1'b0 ;
  assign n26018 = n8868 | n26017 ;
  assign n26019 = n3083 | n15976 ;
  assign n26020 = n23594 & ~n26019 ;
  assign n26021 = n6218 | n12929 ;
  assign n26022 = n26020 & ~n26021 ;
  assign n26023 = ( n6418 & n26018 ) | ( n6418 & ~n26022 ) | ( n26018 & ~n26022 ) ;
  assign n26024 = ( ~n4482 & n26016 ) | ( ~n4482 & n26023 ) | ( n26016 & n26023 ) ;
  assign n26025 = ( n3135 & n7943 ) | ( n3135 & n19380 ) | ( n7943 & n19380 ) ;
  assign n26026 = ( x123 & n20721 ) | ( x123 & ~n26025 ) | ( n20721 & ~n26025 ) ;
  assign n26027 = n13645 ^ n9352 ^ n3728 ;
  assign n26028 = ( ~n2649 & n16901 ) | ( ~n2649 & n20594 ) | ( n16901 & n20594 ) ;
  assign n26029 = n26027 & n26028 ;
  assign n26030 = ( ~n14787 & n26026 ) | ( ~n14787 & n26029 ) | ( n26026 & n26029 ) ;
  assign n26033 = n3305 & n16991 ;
  assign n26034 = n26033 ^ n2616 ^ 1'b0 ;
  assign n26035 = n24212 ^ n601 ^ 1'b0 ;
  assign n26036 = ( n3898 & n26034 ) | ( n3898 & n26035 ) | ( n26034 & n26035 ) ;
  assign n26037 = ( n14335 & n20222 ) | ( n14335 & ~n26036 ) | ( n20222 & ~n26036 ) ;
  assign n26031 = ( ~n6887 & n14632 ) | ( ~n6887 & n15212 ) | ( n14632 & n15212 ) ;
  assign n26032 = ~n7565 & n26031 ;
  assign n26038 = n26037 ^ n26032 ^ n13777 ;
  assign n26039 = n17475 ^ n15100 ^ n10584 ;
  assign n26040 = n26039 ^ n14113 ^ n3750 ;
  assign n26041 = ( n8255 & ~n9624 ) | ( n8255 & n16783 ) | ( ~n9624 & n16783 ) ;
  assign n26042 = ( n5079 & n10429 ) | ( n5079 & ~n22317 ) | ( n10429 & ~n22317 ) ;
  assign n26043 = ( n26040 & ~n26041 ) | ( n26040 & n26042 ) | ( ~n26041 & n26042 ) ;
  assign n26044 = n24193 ^ n1509 ^ 1'b0 ;
  assign n26045 = n15840 & n20919 ;
  assign n26046 = ~n26044 & n26045 ;
  assign n26047 = ( n8116 & ~n11425 ) | ( n8116 & n14811 ) | ( ~n11425 & n14811 ) ;
  assign n26048 = n17436 ^ n3090 ^ 1'b0 ;
  assign n26049 = ( n17056 & n23878 ) | ( n17056 & n26048 ) | ( n23878 & n26048 ) ;
  assign n26050 = n10458 ^ n3373 ^ 1'b0 ;
  assign n26055 = ~n14180 & n25709 ;
  assign n26056 = n26055 ^ n291 ^ 1'b0 ;
  assign n26051 = ( n605 & n13709 ) | ( n605 & n15479 ) | ( n13709 & n15479 ) ;
  assign n26052 = n24405 | n26051 ;
  assign n26053 = n26052 ^ n12427 ^ 1'b0 ;
  assign n26054 = n707 & ~n26053 ;
  assign n26057 = n26056 ^ n26054 ^ 1'b0 ;
  assign n26058 = ~n26050 & n26057 ;
  assign n26059 = n26058 ^ n18206 ^ n8756 ;
  assign n26060 = n26059 ^ n23010 ^ n17146 ;
  assign n26061 = ( n5409 & n17132 ) | ( n5409 & n17735 ) | ( n17132 & n17735 ) ;
  assign n26062 = ( n2555 & n9883 ) | ( n2555 & ~n14084 ) | ( n9883 & ~n14084 ) ;
  assign n26063 = n13078 ^ n10165 ^ n7675 ;
  assign n26064 = ( n5694 & n14411 ) | ( n5694 & ~n26063 ) | ( n14411 & ~n26063 ) ;
  assign n26065 = ( n5233 & n26062 ) | ( n5233 & n26064 ) | ( n26062 & n26064 ) ;
  assign n26066 = ( n4234 & n6068 ) | ( n4234 & n26065 ) | ( n6068 & n26065 ) ;
  assign n26068 = n19466 ^ n13322 ^ n269 ;
  assign n26067 = n10199 ^ n2264 ^ 1'b0 ;
  assign n26069 = n26068 ^ n26067 ^ n11347 ;
  assign n26070 = n1167 & ~n26069 ;
  assign n26071 = ( n26061 & n26066 ) | ( n26061 & ~n26070 ) | ( n26066 & ~n26070 ) ;
  assign n26072 = n18727 ^ n9131 ^ n8104 ;
  assign n26073 = n25261 ^ n22617 ^ n3389 ;
  assign n26074 = ( n5784 & ~n26072 ) | ( n5784 & n26073 ) | ( ~n26072 & n26073 ) ;
  assign n26075 = n26074 ^ n18519 ^ n477 ;
  assign n26076 = ~n7137 & n26075 ;
  assign n26077 = n19620 & n26076 ;
  assign n26078 = n26077 ^ n18825 ^ n2608 ;
  assign n26079 = ( ~n12653 & n14046 ) | ( ~n12653 & n23670 ) | ( n14046 & n23670 ) ;
  assign n26080 = n8613 ^ n7007 ^ n4174 ;
  assign n26081 = ( n2845 & n21116 ) | ( n2845 & ~n26080 ) | ( n21116 & ~n26080 ) ;
  assign n26082 = ( ~n15977 & n23846 ) | ( ~n15977 & n26081 ) | ( n23846 & n26081 ) ;
  assign n26083 = n20251 ^ n1449 ^ x253 ;
  assign n26084 = ( n1651 & n25839 ) | ( n1651 & ~n26083 ) | ( n25839 & ~n26083 ) ;
  assign n26085 = n26084 ^ n10069 ^ 1'b0 ;
  assign n26086 = n26082 & ~n26085 ;
  assign n26087 = ( n1416 & ~n1552 ) | ( n1416 & n6119 ) | ( ~n1552 & n6119 ) ;
  assign n26088 = n26087 ^ n17379 ^ n8808 ;
  assign n26089 = ( ~n615 & n10779 ) | ( ~n615 & n26088 ) | ( n10779 & n26088 ) ;
  assign n26090 = n20408 ^ n17606 ^ n17428 ;
  assign n26094 = ( n2927 & n6626 ) | ( n2927 & ~n14352 ) | ( n6626 & ~n14352 ) ;
  assign n26091 = ~n8640 & n16220 ;
  assign n26092 = ~n18318 & n26091 ;
  assign n26093 = n26092 ^ n13713 ^ n5395 ;
  assign n26095 = n26094 ^ n26093 ^ n5070 ;
  assign n26096 = ( n2374 & ~n4877 ) | ( n2374 & n13349 ) | ( ~n4877 & n13349 ) ;
  assign n26098 = n8071 ^ n7833 ^ n6143 ;
  assign n26097 = ( n4245 & ~n8112 ) | ( n4245 & n19163 ) | ( ~n8112 & n19163 ) ;
  assign n26099 = n26098 ^ n26097 ^ n5680 ;
  assign n26100 = ( n3202 & n8712 ) | ( n3202 & ~n26099 ) | ( n8712 & ~n26099 ) ;
  assign n26111 = n8311 ^ n6373 ^ n1662 ;
  assign n26109 = n21655 ^ n20445 ^ n13348 ;
  assign n26110 = n26109 ^ n6708 ^ n6409 ;
  assign n26101 = n18074 ^ n8699 ^ n3201 ;
  assign n26102 = n26101 ^ n17020 ^ n11764 ;
  assign n26105 = n7859 ^ n6189 ^ n2106 ;
  assign n26103 = n20507 ^ n10740 ^ n284 ;
  assign n26104 = n26103 ^ n10509 ^ n1159 ;
  assign n26106 = n26105 ^ n26104 ^ n8769 ;
  assign n26107 = ( n8437 & ~n10123 ) | ( n8437 & n26106 ) | ( ~n10123 & n26106 ) ;
  assign n26108 = ( n12283 & ~n26102 ) | ( n12283 & n26107 ) | ( ~n26102 & n26107 ) ;
  assign n26112 = n26111 ^ n26110 ^ n26108 ;
  assign n26115 = n22033 ^ n3261 ^ 1'b0 ;
  assign n26113 = n20497 ^ n14304 ^ n11619 ;
  assign n26114 = ( n11222 & n11270 ) | ( n11222 & ~n26113 ) | ( n11270 & ~n26113 ) ;
  assign n26116 = n26115 ^ n26114 ^ n18272 ;
  assign n26117 = n25043 ^ n4780 ^ n2004 ;
  assign n26118 = n26117 ^ n13845 ^ n1880 ;
  assign n26119 = ( n13412 & n23064 ) | ( n13412 & ~n25222 ) | ( n23064 & ~n25222 ) ;
  assign n26120 = n26119 ^ n9301 ^ 1'b0 ;
  assign n26121 = ~n26118 & n26120 ;
  assign n26122 = ( ~n11844 & n14843 ) | ( ~n11844 & n25199 ) | ( n14843 & n25199 ) ;
  assign n26123 = ( n6501 & n11503 ) | ( n6501 & n26122 ) | ( n11503 & n26122 ) ;
  assign n26124 = ( n4219 & n5555 ) | ( n4219 & n10879 ) | ( n5555 & n10879 ) ;
  assign n26125 = n26124 ^ n7734 ^ n7426 ;
  assign n26126 = n22221 ^ n19994 ^ n11275 ;
  assign n26127 = n24827 ^ n4758 ^ n4594 ;
  assign n26128 = ( n2096 & ~n23800 ) | ( n2096 & n26127 ) | ( ~n23800 & n26127 ) ;
  assign n26129 = ( ~x191 & n8071 ) | ( ~x191 & n20031 ) | ( n8071 & n20031 ) ;
  assign n26130 = n26129 ^ n1664 ^ 1'b0 ;
  assign n26131 = n5433 | n26130 ;
  assign n26132 = n11512 ^ n10710 ^ n3814 ;
  assign n26133 = ( ~n6346 & n20619 ) | ( ~n6346 & n23652 ) | ( n20619 & n23652 ) ;
  assign n26134 = n26133 ^ n24013 ^ n6748 ;
  assign n26135 = ( n3596 & n14592 ) | ( n3596 & ~n14660 ) | ( n14592 & ~n14660 ) ;
  assign n26136 = ( n659 & ~n6752 ) | ( n659 & n9703 ) | ( ~n6752 & n9703 ) ;
  assign n26137 = ( n8306 & n15883 ) | ( n8306 & ~n26136 ) | ( n15883 & ~n26136 ) ;
  assign n26138 = ( n2017 & n9384 ) | ( n2017 & n12159 ) | ( n9384 & n12159 ) ;
  assign n26139 = n11110 | n13232 ;
  assign n26140 = n26139 ^ n11904 ^ n933 ;
  assign n26146 = n10643 & ~n11808 ;
  assign n26147 = n26146 ^ n10794 ^ 1'b0 ;
  assign n26148 = n5026 | n6560 ;
  assign n26149 = n26148 ^ n22826 ^ n7546 ;
  assign n26150 = ( n3335 & ~n26147 ) | ( n3335 & n26149 ) | ( ~n26147 & n26149 ) ;
  assign n26143 = n9823 ^ n4119 ^ n611 ;
  assign n26144 = ( ~x154 & n13136 ) | ( ~x154 & n26143 ) | ( n13136 & n26143 ) ;
  assign n26141 = n17364 ^ n9215 ^ n7002 ;
  assign n26142 = n6792 & n26141 ;
  assign n26145 = n26144 ^ n26142 ^ 1'b0 ;
  assign n26151 = n26150 ^ n26145 ^ n1489 ;
  assign n26152 = n10183 ^ n4043 ^ n3680 ;
  assign n26153 = n26152 ^ n9056 ^ 1'b0 ;
  assign n26154 = n5460 | n26153 ;
  assign n26156 = n10348 ^ n6607 ^ n5495 ;
  assign n26155 = n9630 & n13659 ;
  assign n26157 = n26156 ^ n26155 ^ n18727 ;
  assign n26158 = n13899 ^ n12408 ^ n8010 ;
  assign n26159 = x50 & ~n26158 ;
  assign n26160 = n19722 ^ n8633 ^ n5816 ;
  assign n26161 = n26160 ^ n6686 ^ 1'b0 ;
  assign n26162 = n8153 | n26161 ;
  assign n26163 = ~n3706 & n24960 ;
  assign n26164 = n989 & n26163 ;
  assign n26165 = n26164 ^ n20518 ^ n3185 ;
  assign n26166 = ( n9831 & n18093 ) | ( n9831 & ~n26165 ) | ( n18093 & ~n26165 ) ;
  assign n26168 = n8645 & n19729 ;
  assign n26167 = n23198 ^ n14316 ^ n9290 ;
  assign n26169 = n26168 ^ n26167 ^ n18181 ;
  assign n26170 = ( ~n5189 & n6217 ) | ( ~n5189 & n6317 ) | ( n6217 & n6317 ) ;
  assign n26171 = ( ~n23592 & n24693 ) | ( ~n23592 & n26170 ) | ( n24693 & n26170 ) ;
  assign n26172 = ( ~n2268 & n13394 ) | ( ~n2268 & n20103 ) | ( n13394 & n20103 ) ;
  assign n26173 = ( n15208 & n19697 ) | ( n15208 & n26172 ) | ( n19697 & n26172 ) ;
  assign n26174 = ~n9841 & n14829 ;
  assign n26175 = ( n2613 & ~n9177 ) | ( n2613 & n10760 ) | ( ~n9177 & n10760 ) ;
  assign n26176 = n26175 ^ n14317 ^ n6031 ;
  assign n26177 = ( n18015 & ~n21324 ) | ( n18015 & n26176 ) | ( ~n21324 & n26176 ) ;
  assign n26178 = ( n1750 & ~n2463 ) | ( n1750 & n21898 ) | ( ~n2463 & n21898 ) ;
  assign n26179 = ( n20063 & n21377 ) | ( n20063 & n26178 ) | ( n21377 & n26178 ) ;
  assign n26190 = ( ~n4917 & n9214 ) | ( ~n4917 & n9700 ) | ( n9214 & n9700 ) ;
  assign n26188 = n16042 ^ n13833 ^ n5033 ;
  assign n26189 = ~n12992 & n26188 ;
  assign n26183 = ~n1034 & n17045 ;
  assign n26184 = n2453 & n26183 ;
  assign n26185 = n26184 ^ n12285 ^ n2997 ;
  assign n26180 = ~n2013 & n21209 ;
  assign n26181 = n26180 ^ n16128 ^ 1'b0 ;
  assign n26182 = ( n3465 & ~n4406 ) | ( n3465 & n26181 ) | ( ~n4406 & n26181 ) ;
  assign n26186 = n26185 ^ n26182 ^ n25224 ;
  assign n26187 = n26186 ^ n21571 ^ n14045 ;
  assign n26191 = n26190 ^ n26189 ^ n26187 ;
  assign n26192 = ~n1630 & n15310 ;
  assign n26193 = n26192 ^ n11579 ^ n10965 ;
  assign n26194 = n10861 ^ n6126 ^ n3382 ;
  assign n26195 = n6195 & ~n7157 ;
  assign n26196 = ~n26194 & n26195 ;
  assign n26197 = ( ~n7690 & n19111 ) | ( ~n7690 & n26196 ) | ( n19111 & n26196 ) ;
  assign n26198 = ( n12186 & n16066 ) | ( n12186 & n17939 ) | ( n16066 & n17939 ) ;
  assign n26199 = n23758 | n25633 ;
  assign n26200 = n23783 & ~n26199 ;
  assign n26201 = n6061 ^ n4153 ^ 1'b0 ;
  assign n26202 = ~n2115 & n26201 ;
  assign n26203 = ( n1033 & ~n26200 ) | ( n1033 & n26202 ) | ( ~n26200 & n26202 ) ;
  assign n26204 = n16385 ^ n12921 ^ 1'b0 ;
  assign n26205 = n5971 & n26204 ;
  assign n26208 = n9517 ^ n2641 ^ n772 ;
  assign n26209 = n2609 | n13152 ;
  assign n26210 = n26209 ^ n7890 ^ 1'b0 ;
  assign n26211 = ( n7368 & ~n26208 ) | ( n7368 & n26210 ) | ( ~n26208 & n26210 ) ;
  assign n26206 = n16316 & ~n16602 ;
  assign n26207 = ~n11650 & n26206 ;
  assign n26212 = n26211 ^ n26207 ^ n18205 ;
  assign n26213 = n14566 ^ n3464 ^ n1814 ;
  assign n26214 = n18976 ^ n15941 ^ 1'b0 ;
  assign n26215 = ~n14227 & n26214 ;
  assign n26216 = ~n519 & n15333 ;
  assign n26217 = n15468 & n26216 ;
  assign n26218 = n26217 ^ n15395 ^ n11097 ;
  assign n26219 = n18781 | n19233 ;
  assign n26220 = n1019 & ~n26219 ;
  assign n26221 = n26220 ^ n25090 ^ 1'b0 ;
  assign n26222 = n20917 ^ n18966 ^ n8348 ;
  assign n26223 = ( ~n5985 & n6567 ) | ( ~n5985 & n18648 ) | ( n6567 & n18648 ) ;
  assign n26224 = ( n13505 & n26222 ) | ( n13505 & ~n26223 ) | ( n26222 & ~n26223 ) ;
  assign n26225 = ( ~n1980 & n9052 ) | ( ~n1980 & n13283 ) | ( n9052 & n13283 ) ;
  assign n26226 = n4505 & n7553 ;
  assign n26227 = n24713 & n26226 ;
  assign n26228 = ( n8737 & ~n11043 ) | ( n8737 & n25741 ) | ( ~n11043 & n25741 ) ;
  assign n26229 = ( n19181 & ~n26227 ) | ( n19181 & n26228 ) | ( ~n26227 & n26228 ) ;
  assign n26230 = n26229 ^ n21433 ^ n8876 ;
  assign n26231 = ( ~n6137 & n26225 ) | ( ~n6137 & n26230 ) | ( n26225 & n26230 ) ;
  assign n26232 = n544 | n26231 ;
  assign n26233 = n26232 ^ n2725 ^ 1'b0 ;
  assign n26235 = n12037 ^ n5845 ^ n2198 ;
  assign n26236 = n26235 ^ n2513 ^ n1977 ;
  assign n26234 = n13494 ^ n5237 ^ n318 ;
  assign n26237 = n26236 ^ n26234 ^ 1'b0 ;
  assign n26238 = n4584 & n26237 ;
  assign n26239 = ( n6318 & n9703 ) | ( n6318 & ~n25591 ) | ( n9703 & ~n25591 ) ;
  assign n26240 = n14731 ^ n13063 ^ n3989 ;
  assign n26241 = n17656 ^ n10082 ^ n1838 ;
  assign n26242 = ( ~n26239 & n26240 ) | ( ~n26239 & n26241 ) | ( n26240 & n26241 ) ;
  assign n26243 = n19602 ^ n11074 ^ n5827 ;
  assign n26244 = ( n12129 & ~n19761 ) | ( n12129 & n26243 ) | ( ~n19761 & n26243 ) ;
  assign n26249 = ( n1492 & n6491 ) | ( n1492 & ~n13256 ) | ( n6491 & ~n13256 ) ;
  assign n26250 = ( n1290 & ~n3717 ) | ( n1290 & n19499 ) | ( ~n3717 & n19499 ) ;
  assign n26251 = n11298 ^ n2367 ^ 1'b0 ;
  assign n26252 = n10779 & ~n26251 ;
  assign n26253 = ( ~n26249 & n26250 ) | ( ~n26249 & n26252 ) | ( n26250 & n26252 ) ;
  assign n26247 = ( n1171 & n9718 ) | ( n1171 & ~n16198 ) | ( n9718 & ~n16198 ) ;
  assign n26245 = ( ~n7393 & n8590 ) | ( ~n7393 & n13436 ) | ( n8590 & n13436 ) ;
  assign n26246 = ( n11817 & ~n18218 ) | ( n11817 & n26245 ) | ( ~n18218 & n26245 ) ;
  assign n26248 = n26247 ^ n26246 ^ n10191 ;
  assign n26254 = n26253 ^ n26248 ^ n16283 ;
  assign n26255 = n1804 | n12078 ;
  assign n26256 = n26254 | n26255 ;
  assign n26257 = n5798 | n18936 ;
  assign n26258 = n12482 ^ n9136 ^ n8041 ;
  assign n26259 = x202 & ~n1349 ;
  assign n26260 = ( n4884 & n26258 ) | ( n4884 & n26259 ) | ( n26258 & n26259 ) ;
  assign n26261 = ( n4076 & ~n15034 ) | ( n4076 & n21448 ) | ( ~n15034 & n21448 ) ;
  assign n26262 = n8721 ^ x208 ^ 1'b0 ;
  assign n26263 = n26262 ^ n12667 ^ n7585 ;
  assign n26264 = n11738 & n26263 ;
  assign n26265 = ~n13537 & n26264 ;
  assign n26266 = ( n7276 & ~n11220 ) | ( n7276 & n26265 ) | ( ~n11220 & n26265 ) ;
  assign n26267 = n24487 ^ n11514 ^ n7042 ;
  assign n26268 = n383 | n16371 ;
  assign n26269 = n26267 | n26268 ;
  assign n26270 = n13581 ^ n9315 ^ n1174 ;
  assign n26271 = n20201 ^ n9293 ^ n5811 ;
  assign n26272 = n26270 | n26271 ;
  assign n26279 = ( n910 & n12471 ) | ( n910 & n15973 ) | ( n12471 & n15973 ) ;
  assign n26277 = n23054 ^ n11768 ^ 1'b0 ;
  assign n26278 = n26277 ^ n22814 ^ n17722 ;
  assign n26280 = n26279 ^ n26278 ^ n7417 ;
  assign n26274 = n1538 & ~n11265 ;
  assign n26275 = n24585 & n26274 ;
  assign n26273 = n14050 ^ n11359 ^ n8501 ;
  assign n26276 = n26275 ^ n26273 ^ n19877 ;
  assign n26281 = n26280 ^ n26276 ^ n9482 ;
  assign n26282 = ~n7214 & n18544 ;
  assign n26283 = n22297 & n26282 ;
  assign n26284 = ( n1409 & ~n1716 ) | ( n1409 & n2268 ) | ( ~n1716 & n2268 ) ;
  assign n26285 = n26284 ^ n17634 ^ n9725 ;
  assign n26286 = n17503 ^ n5346 ^ n4324 ;
  assign n26287 = ( n6379 & n6397 ) | ( n6379 & n11207 ) | ( n6397 & n11207 ) ;
  assign n26288 = ( n6876 & ~n14265 ) | ( n6876 & n26287 ) | ( ~n14265 & n26287 ) ;
  assign n26289 = n26288 ^ n5113 ^ 1'b0 ;
  assign n26290 = ( n2825 & n26286 ) | ( n2825 & n26289 ) | ( n26286 & n26289 ) ;
  assign n26291 = n2199 ^ n1691 ^ x90 ;
  assign n26292 = n26291 ^ n12880 ^ 1'b0 ;
  assign n26293 = ( n4642 & n5384 ) | ( n4642 & n15356 ) | ( n5384 & n15356 ) ;
  assign n26294 = n26293 ^ n7739 ^ n2883 ;
  assign n26295 = ( n11781 & ~n26292 ) | ( n11781 & n26294 ) | ( ~n26292 & n26294 ) ;
  assign n26296 = n12550 ^ n9328 ^ 1'b0 ;
  assign n26297 = ( n5940 & ~n18071 ) | ( n5940 & n26296 ) | ( ~n18071 & n26296 ) ;
  assign n26298 = n26297 ^ n11922 ^ 1'b0 ;
  assign n26299 = n26298 ^ n4888 ^ 1'b0 ;
  assign n26300 = n23627 ^ n20883 ^ n9608 ;
  assign n26301 = n22895 ^ n21351 ^ n14445 ;
  assign n26302 = ( ~n4195 & n11189 ) | ( ~n4195 & n13186 ) | ( n11189 & n13186 ) ;
  assign n26303 = n26302 ^ n24849 ^ n13633 ;
  assign n26304 = n18645 ^ n11481 ^ n8727 ;
  assign n26305 = ( n11617 & n18104 ) | ( n11617 & n26304 ) | ( n18104 & n26304 ) ;
  assign n26306 = ( ~n5750 & n10617 ) | ( ~n5750 & n14400 ) | ( n10617 & n14400 ) ;
  assign n26307 = n14001 ^ n8813 ^ n2769 ;
  assign n26308 = ~n3448 & n26307 ;
  assign n26309 = ~n2410 & n26308 ;
  assign n26310 = n26306 | n26309 ;
  assign n26311 = ( x148 & n26305 ) | ( x148 & n26310 ) | ( n26305 & n26310 ) ;
  assign n26312 = ~n26303 & n26311 ;
  assign n26313 = n1633 | n4824 ;
  assign n26314 = n9179 ^ n8071 ^ n7153 ;
  assign n26315 = n26314 ^ n18266 ^ n4965 ;
  assign n26316 = ( x17 & ~n14090 ) | ( x17 & n26315 ) | ( ~n14090 & n26315 ) ;
  assign n26317 = n17571 ^ n15457 ^ n7378 ;
  assign n26318 = n26317 ^ n7538 ^ 1'b0 ;
  assign n26319 = ~n13717 & n26318 ;
  assign n26320 = ( n20911 & n26316 ) | ( n20911 & ~n26319 ) | ( n26316 & ~n26319 ) ;
  assign n26321 = ( n3880 & n4141 ) | ( n3880 & n18901 ) | ( n4141 & n18901 ) ;
  assign n26322 = n19353 ^ n6628 ^ n5235 ;
  assign n26323 = n26322 ^ n16427 ^ 1'b0 ;
  assign n26324 = n23111 ^ n16263 ^ n8465 ;
  assign n26325 = ( n11549 & ~n17496 ) | ( n11549 & n18408 ) | ( ~n17496 & n18408 ) ;
  assign n26326 = n26325 ^ n20818 ^ n1074 ;
  assign n26327 = ( n3196 & n7744 ) | ( n3196 & n26326 ) | ( n7744 & n26326 ) ;
  assign n26328 = ( n800 & ~n22290 ) | ( n800 & n26327 ) | ( ~n22290 & n26327 ) ;
  assign n26329 = ( n4307 & n13761 ) | ( n4307 & ~n17517 ) | ( n13761 & ~n17517 ) ;
  assign n26330 = n26329 ^ n8005 ^ n742 ;
  assign n26331 = ( n7851 & n25471 ) | ( n7851 & ~n26330 ) | ( n25471 & ~n26330 ) ;
  assign n26332 = ( n4823 & n7028 ) | ( n4823 & n26331 ) | ( n7028 & n26331 ) ;
  assign n26333 = ~n8349 & n20910 ;
  assign n26334 = ( ~n1269 & n7631 ) | ( ~n1269 & n26333 ) | ( n7631 & n26333 ) ;
  assign n26341 = n7367 & ~n13121 ;
  assign n26342 = n26341 ^ n11636 ^ 1'b0 ;
  assign n26343 = n13966 ^ n13664 ^ n3212 ;
  assign n26344 = ( n8239 & n26342 ) | ( n8239 & ~n26343 ) | ( n26342 & ~n26343 ) ;
  assign n26345 = n21287 & n26344 ;
  assign n26336 = n25326 ^ n15515 ^ n774 ;
  assign n26335 = ( n893 & n3844 ) | ( n893 & ~n20950 ) | ( n3844 & ~n20950 ) ;
  assign n26337 = n26336 ^ n26335 ^ n4406 ;
  assign n26338 = n10942 ^ n4525 ^ 1'b0 ;
  assign n26339 = ~n26337 & n26338 ;
  assign n26340 = n26339 ^ n22369 ^ n4863 ;
  assign n26346 = n26345 ^ n26340 ^ 1'b0 ;
  assign n26347 = ( ~n12396 & n18460 ) | ( ~n12396 & n26346 ) | ( n18460 & n26346 ) ;
  assign n26348 = ~n705 & n8585 ;
  assign n26349 = n26348 ^ n1229 ^ 1'b0 ;
  assign n26350 = ~n4334 & n26349 ;
  assign n26351 = n26350 ^ n2495 ^ 1'b0 ;
  assign n26352 = n8433 ^ n6714 ^ n5502 ;
  assign n26353 = ( n4438 & n26351 ) | ( n4438 & n26352 ) | ( n26351 & n26352 ) ;
  assign n26354 = ( n1335 & n1887 ) | ( n1335 & n12667 ) | ( n1887 & n12667 ) ;
  assign n26355 = n26354 ^ n12574 ^ n1162 ;
  assign n26356 = ( n12946 & n15656 ) | ( n12946 & n22488 ) | ( n15656 & n22488 ) ;
  assign n26359 = n12694 ^ x197 ^ 1'b0 ;
  assign n26360 = ~n5434 & n26359 ;
  assign n26357 = n22028 ^ n8870 ^ n4667 ;
  assign n26358 = ( n1531 & n2061 ) | ( n1531 & n26357 ) | ( n2061 & n26357 ) ;
  assign n26361 = n26360 ^ n26358 ^ n10429 ;
  assign n26362 = ( n3410 & n26356 ) | ( n3410 & ~n26361 ) | ( n26356 & ~n26361 ) ;
  assign n26363 = ~n22388 & n26362 ;
  assign n26364 = ( n11673 & n22397 ) | ( n11673 & n23491 ) | ( n22397 & n23491 ) ;
  assign n26372 = ( ~n6318 & n8819 ) | ( ~n6318 & n13348 ) | ( n8819 & n13348 ) ;
  assign n26367 = n1151 ^ x114 ^ 1'b0 ;
  assign n26368 = n7746 & n26367 ;
  assign n26369 = ( n2510 & n12940 ) | ( n2510 & n26368 ) | ( n12940 & n26368 ) ;
  assign n26370 = n26369 ^ n25326 ^ 1'b0 ;
  assign n26365 = n17245 ^ n16106 ^ n9570 ;
  assign n26366 = n26365 ^ n3008 ^ 1'b0 ;
  assign n26371 = n26370 ^ n26366 ^ n6563 ;
  assign n26373 = n26372 ^ n26371 ^ n21314 ;
  assign n26374 = ( ~n423 & n3736 ) | ( ~n423 & n17585 ) | ( n3736 & n17585 ) ;
  assign n26375 = ( ~n8114 & n10470 ) | ( ~n8114 & n11817 ) | ( n10470 & n11817 ) ;
  assign n26376 = ( ~n2672 & n10103 ) | ( ~n2672 & n26375 ) | ( n10103 & n26375 ) ;
  assign n26377 = ( n4155 & ~n26374 ) | ( n4155 & n26376 ) | ( ~n26374 & n26376 ) ;
  assign n26378 = ( ~n2712 & n6683 ) | ( ~n2712 & n8918 ) | ( n6683 & n8918 ) ;
  assign n26379 = n26378 ^ n18070 ^ n459 ;
  assign n26380 = n20634 ^ n18695 ^ n16119 ;
  assign n26381 = ( n6048 & n6868 ) | ( n6048 & ~n22909 ) | ( n6868 & ~n22909 ) ;
  assign n26382 = ( n20823 & n24004 ) | ( n20823 & ~n26381 ) | ( n24004 & ~n26381 ) ;
  assign n26383 = n26382 ^ n25007 ^ n12891 ;
  assign n26385 = ~x104 & n1623 ;
  assign n26386 = ( n826 & n9415 ) | ( n826 & n26385 ) | ( n9415 & n26385 ) ;
  assign n26384 = ( ~n1113 & n6443 ) | ( ~n1113 & n13505 ) | ( n6443 & n13505 ) ;
  assign n26387 = n26386 ^ n26384 ^ n3514 ;
  assign n26388 = n11213 | n16285 ;
  assign n26389 = n26388 ^ n11220 ^ n7383 ;
  assign n26390 = ( ~n496 & n3328 ) | ( ~n496 & n9937 ) | ( n3328 & n9937 ) ;
  assign n26391 = n7460 | n7511 ;
  assign n26392 = n26390 | n26391 ;
  assign n26393 = n8407 & n13342 ;
  assign n26394 = ~n17090 & n26393 ;
  assign n26395 = n2372 & ~n6637 ;
  assign n26396 = n26395 ^ n25451 ^ 1'b0 ;
  assign n26397 = ( ~n4604 & n26394 ) | ( ~n4604 & n26396 ) | ( n26394 & n26396 ) ;
  assign n26399 = ( ~n2324 & n11289 ) | ( ~n2324 & n16732 ) | ( n11289 & n16732 ) ;
  assign n26398 = n1217 & ~n20582 ;
  assign n26400 = n26399 ^ n26398 ^ 1'b0 ;
  assign n26401 = n15150 ^ n2809 ^ 1'b0 ;
  assign n26402 = n26401 ^ n20234 ^ n11831 ;
  assign n26403 = ( n19494 & ~n26400 ) | ( n19494 & n26402 ) | ( ~n26400 & n26402 ) ;
  assign n26405 = n15429 ^ n11953 ^ n5126 ;
  assign n26404 = n23121 ^ n22590 ^ n8657 ;
  assign n26406 = n26405 ^ n26404 ^ n9460 ;
  assign n26407 = n24675 ^ n12619 ^ n2378 ;
  assign n26408 = n26407 ^ n7619 ^ n1666 ;
  assign n26411 = n13876 ^ n12226 ^ 1'b0 ;
  assign n26409 = ( n1583 & ~n7774 ) | ( n1583 & n12876 ) | ( ~n7774 & n12876 ) ;
  assign n26410 = n26409 ^ n9320 ^ n1795 ;
  assign n26412 = n26411 ^ n26410 ^ n11436 ;
  assign n26413 = n24082 ^ n6363 ^ n2112 ;
  assign n26414 = n22235 ^ n16927 ^ n5264 ;
  assign n26415 = ( n1422 & ~n19960 ) | ( n1422 & n26414 ) | ( ~n19960 & n26414 ) ;
  assign n26416 = ( ~n624 & n26413 ) | ( ~n624 & n26415 ) | ( n26413 & n26415 ) ;
  assign n26417 = ( n6511 & n18585 ) | ( n6511 & ~n26416 ) | ( n18585 & ~n26416 ) ;
  assign n26418 = ( n13163 & n19009 ) | ( n13163 & n23562 ) | ( n19009 & n23562 ) ;
  assign n26419 = ( n9738 & n10828 ) | ( n9738 & n26418 ) | ( n10828 & n26418 ) ;
  assign n26420 = ( ~n1467 & n2722 ) | ( ~n1467 & n26419 ) | ( n2722 & n26419 ) ;
  assign n26421 = n15403 ^ n7721 ^ n5601 ;
  assign n26424 = ( ~x102 & n7365 ) | ( ~x102 & n21777 ) | ( n7365 & n21777 ) ;
  assign n26425 = ( n4100 & n15196 ) | ( n4100 & ~n26424 ) | ( n15196 & ~n26424 ) ;
  assign n26422 = n9240 | n26199 ;
  assign n26423 = n26422 ^ n8084 ^ 1'b0 ;
  assign n26426 = n26425 ^ n26423 ^ n21193 ;
  assign n26427 = ( n18378 & ~n26421 ) | ( n18378 & n26426 ) | ( ~n26421 & n26426 ) ;
  assign n26428 = n18215 ^ n8752 ^ n2389 ;
  assign n26429 = n26428 ^ n23324 ^ n2614 ;
  assign n26431 = ( n1433 & n10990 ) | ( n1433 & n24994 ) | ( n10990 & n24994 ) ;
  assign n26432 = ( n2121 & n20217 ) | ( n2121 & ~n26431 ) | ( n20217 & ~n26431 ) ;
  assign n26430 = ( n2890 & ~n11990 ) | ( n2890 & n12011 ) | ( ~n11990 & n12011 ) ;
  assign n26433 = n26432 ^ n26430 ^ n19124 ;
  assign n26434 = n21769 ^ n7333 ^ n654 ;
  assign n26435 = n21953 & ~n26434 ;
  assign n26436 = n4128 & ~n8258 ;
  assign n26437 = ( n21053 & ~n24891 ) | ( n21053 & n26436 ) | ( ~n24891 & n26436 ) ;
  assign n26438 = ( n8897 & n26435 ) | ( n8897 & ~n26437 ) | ( n26435 & ~n26437 ) ;
  assign n26439 = ( n13432 & n17277 ) | ( n13432 & n24953 ) | ( n17277 & n24953 ) ;
  assign n26440 = ( n7059 & n12605 ) | ( n7059 & n19139 ) | ( n12605 & n19139 ) ;
  assign n26441 = ( n8134 & n26439 ) | ( n8134 & ~n26440 ) | ( n26439 & ~n26440 ) ;
  assign n26443 = n20144 ^ n16383 ^ n6988 ;
  assign n26442 = n2129 & n10251 ;
  assign n26444 = n26443 ^ n26442 ^ 1'b0 ;
  assign n26445 = n26444 ^ n11104 ^ n9991 ;
  assign n26446 = n3983 & ~n5473 ;
  assign n26447 = ( x189 & n15955 ) | ( x189 & ~n26446 ) | ( n15955 & ~n26446 ) ;
  assign n26448 = n26447 ^ n6320 ^ n2591 ;
  assign n26449 = n26448 ^ n8838 ^ n8578 ;
  assign n26451 = ~n9801 & n20828 ;
  assign n26452 = n26451 ^ n4110 ^ 1'b0 ;
  assign n26450 = ( ~n2959 & n3789 ) | ( ~n2959 & n17231 ) | ( n3789 & n17231 ) ;
  assign n26453 = n26452 ^ n26450 ^ n19289 ;
  assign n26454 = ( n9777 & ~n19152 ) | ( n9777 & n26453 ) | ( ~n19152 & n26453 ) ;
  assign n26455 = n8646 ^ n7486 ^ x252 ;
  assign n26456 = n9846 ^ n9022 ^ n6214 ;
  assign n26457 = ( n17471 & n21623 ) | ( n17471 & n26456 ) | ( n21623 & n26456 ) ;
  assign n26458 = ( n10430 & n26455 ) | ( n10430 & n26457 ) | ( n26455 & n26457 ) ;
  assign n26461 = ( ~n7067 & n10683 ) | ( ~n7067 & n16212 ) | ( n10683 & n16212 ) ;
  assign n26460 = n15926 ^ n14321 ^ n1757 ;
  assign n26462 = n26461 ^ n26460 ^ n2537 ;
  assign n26463 = ( ~n6742 & n8782 ) | ( ~n6742 & n26462 ) | ( n8782 & n26462 ) ;
  assign n26459 = n20399 & n24350 ;
  assign n26464 = n26463 ^ n26459 ^ 1'b0 ;
  assign n26465 = n16969 ^ n6263 ^ n6247 ;
  assign n26466 = n26465 ^ n12720 ^ 1'b0 ;
  assign n26467 = ~n11591 & n19255 ;
  assign n26468 = ~n7936 & n26467 ;
  assign n26469 = ( n7755 & ~n10648 ) | ( n7755 & n16353 ) | ( ~n10648 & n16353 ) ;
  assign n26473 = ( n9425 & n15089 ) | ( n9425 & ~n18547 ) | ( n15089 & ~n18547 ) ;
  assign n26470 = n12126 ^ n11919 ^ n7956 ;
  assign n26471 = n18535 ^ n15147 ^ n13844 ;
  assign n26472 = ( ~n4129 & n26470 ) | ( ~n4129 & n26471 ) | ( n26470 & n26471 ) ;
  assign n26474 = n26473 ^ n26472 ^ n5699 ;
  assign n26475 = n22625 ^ n10308 ^ n7487 ;
  assign n26476 = n26475 ^ n18162 ^ n13413 ;
  assign n26477 = n26476 ^ n1561 ^ 1'b0 ;
  assign n26478 = n26477 ^ n12688 ^ n4376 ;
  assign n26479 = ( n1873 & n2397 ) | ( n1873 & n11785 ) | ( n2397 & n11785 ) ;
  assign n26480 = n26479 ^ n19279 ^ n16636 ;
  assign n26481 = ( n1964 & n5038 ) | ( n1964 & n26480 ) | ( n5038 & n26480 ) ;
  assign n26485 = n8941 | n24444 ;
  assign n26486 = n21334 | n26485 ;
  assign n26482 = n8685 ^ n1170 ^ n919 ;
  assign n26483 = n26482 ^ n15001 ^ n13918 ;
  assign n26484 = x113 & n26483 ;
  assign n26487 = n26486 ^ n26484 ^ 1'b0 ;
  assign n26488 = ( n2025 & n5847 ) | ( n2025 & ~n7612 ) | ( n5847 & ~n7612 ) ;
  assign n26489 = n3518 ^ n1262 ^ n1031 ;
  assign n26490 = ( n18583 & n26488 ) | ( n18583 & ~n26489 ) | ( n26488 & ~n26489 ) ;
  assign n26491 = ( ~n20743 & n23117 ) | ( ~n20743 & n26490 ) | ( n23117 & n26490 ) ;
  assign n26492 = n7260 ^ n939 ^ 1'b0 ;
  assign n26493 = x233 & n26492 ;
  assign n26494 = n26493 ^ n12738 ^ n2204 ;
  assign n26495 = ( ~n4264 & n5322 ) | ( ~n4264 & n26494 ) | ( n5322 & n26494 ) ;
  assign n26498 = n16264 ^ n12938 ^ n11210 ;
  assign n26496 = ( ~n3890 & n7187 ) | ( ~n3890 & n16031 ) | ( n7187 & n16031 ) ;
  assign n26497 = n26496 ^ n19766 ^ n3974 ;
  assign n26499 = n26498 ^ n26497 ^ n8983 ;
  assign n26500 = n6906 | n26499 ;
  assign n26501 = ( n9155 & ~n18691 ) | ( n9155 & n25366 ) | ( ~n18691 & n25366 ) ;
  assign n26502 = ( n14708 & n19667 ) | ( n14708 & ~n26501 ) | ( n19667 & ~n26501 ) ;
  assign n26503 = n16805 ^ n7216 ^ 1'b0 ;
  assign n26504 = n26503 ^ n16517 ^ 1'b0 ;
  assign n26505 = ~n694 & n17863 ;
  assign n26506 = n26505 ^ n9847 ^ 1'b0 ;
  assign n26507 = ( x248 & n4371 ) | ( x248 & ~n17829 ) | ( n4371 & ~n17829 ) ;
  assign n26508 = n26507 ^ n21454 ^ n11785 ;
  assign n26509 = n21670 ^ n10671 ^ 1'b0 ;
  assign n26510 = n26508 & ~n26509 ;
  assign n26511 = ( ~n3342 & n10120 ) | ( ~n3342 & n14102 ) | ( n10120 & n14102 ) ;
  assign n26512 = ( n8696 & n9893 ) | ( n8696 & ~n12514 ) | ( n9893 & ~n12514 ) ;
  assign n26513 = ( n4772 & ~n7655 ) | ( n4772 & n16812 ) | ( ~n7655 & n16812 ) ;
  assign n26514 = ( x172 & ~x230 ) | ( x172 & n8273 ) | ( ~x230 & n8273 ) ;
  assign n26515 = n1564 & n26514 ;
  assign n26516 = n16305 ^ n5915 ^ n3492 ;
  assign n26517 = n15363 ^ n14204 ^ n8244 ;
  assign n26518 = n26517 ^ n18619 ^ n11451 ;
  assign n26519 = n7128 | n9641 ;
  assign n26520 = n26519 ^ n15024 ^ 1'b0 ;
  assign n26521 = ( ~n10494 & n18232 ) | ( ~n10494 & n26520 ) | ( n18232 & n26520 ) ;
  assign n26522 = n25207 ^ n24352 ^ n11448 ;
  assign n26523 = ( ~n2689 & n10492 ) | ( ~n2689 & n12295 ) | ( n10492 & n12295 ) ;
  assign n26527 = ( x168 & n5958 ) | ( x168 & ~n7603 ) | ( n5958 & ~n7603 ) ;
  assign n26524 = n25371 ^ n18033 ^ n6969 ;
  assign n26525 = n26524 ^ n22618 ^ n10354 ;
  assign n26526 = ~n17442 & n26525 ;
  assign n26528 = n26527 ^ n26526 ^ 1'b0 ;
  assign n26529 = ( n5701 & n17953 ) | ( n5701 & n26528 ) | ( n17953 & n26528 ) ;
  assign n26530 = ( n5026 & n26523 ) | ( n5026 & ~n26529 ) | ( n26523 & ~n26529 ) ;
  assign n26531 = ( n363 & n21045 ) | ( n363 & ~n26530 ) | ( n21045 & ~n26530 ) ;
  assign n26532 = ( n2415 & ~n3385 ) | ( n2415 & n20112 ) | ( ~n3385 & n20112 ) ;
  assign n26533 = n1243 | n26532 ;
  assign n26534 = n20916 & ~n26533 ;
  assign n26535 = n3413 | n26534 ;
  assign n26536 = n15552 ^ n11021 ^ n5262 ;
  assign n26537 = ~n14943 & n22246 ;
  assign n26538 = n23718 & n26537 ;
  assign n26539 = ( n2549 & n5769 ) | ( n2549 & ~n26538 ) | ( n5769 & ~n26538 ) ;
  assign n26540 = ( n2184 & n26536 ) | ( n2184 & n26539 ) | ( n26536 & n26539 ) ;
  assign n26541 = ( n16970 & n26535 ) | ( n16970 & n26540 ) | ( n26535 & n26540 ) ;
  assign n26543 = n10541 ^ n3081 ^ n1417 ;
  assign n26544 = n26543 ^ n19911 ^ n19341 ;
  assign n26542 = n22812 ^ n21567 ^ n2630 ;
  assign n26545 = n26544 ^ n26542 ^ n11741 ;
  assign n26552 = n13299 ^ n8760 ^ n4041 ;
  assign n26553 = n21871 ^ n14486 ^ n2220 ;
  assign n26554 = ( n19892 & ~n26552 ) | ( n19892 & n26553 ) | ( ~n26552 & n26553 ) ;
  assign n26550 = ( n1224 & ~n4807 ) | ( n1224 & n18722 ) | ( ~n4807 & n18722 ) ;
  assign n26548 = n13820 ^ n4037 ^ n3206 ;
  assign n26546 = ( n1006 & n3370 ) | ( n1006 & ~n18976 ) | ( n3370 & ~n18976 ) ;
  assign n26547 = ( ~n4909 & n17992 ) | ( ~n4909 & n26546 ) | ( n17992 & n26546 ) ;
  assign n26549 = n26548 ^ n26547 ^ n5143 ;
  assign n26551 = n26550 ^ n26549 ^ n17771 ;
  assign n26555 = n26554 ^ n26551 ^ n16834 ;
  assign n26556 = n19806 ^ n15072 ^ n4129 ;
  assign n26557 = n8296 ^ n5788 ^ n4791 ;
  assign n26558 = ( n7153 & n24948 ) | ( n7153 & n26557 ) | ( n24948 & n26557 ) ;
  assign n26559 = ( n8955 & n18033 ) | ( n8955 & ~n26558 ) | ( n18033 & ~n26558 ) ;
  assign n26560 = n4944 ^ n3361 ^ n3249 ;
  assign n26561 = ( ~n9409 & n10625 ) | ( ~n9409 & n26560 ) | ( n10625 & n26560 ) ;
  assign n26562 = ( n4393 & n13030 ) | ( n4393 & n24849 ) | ( n13030 & n24849 ) ;
  assign n26563 = n26562 ^ n9149 ^ n7359 ;
  assign n26564 = n1382 & ~n26563 ;
  assign n26565 = ( n9040 & n26561 ) | ( n9040 & n26564 ) | ( n26561 & n26564 ) ;
  assign n26566 = n18495 ^ n17561 ^ n1049 ;
  assign n26567 = n16380 ^ n9493 ^ n7234 ;
  assign n26568 = n15187 ^ n13016 ^ n10408 ;
  assign n26569 = n26568 ^ n17322 ^ n17162 ;
  assign n26570 = n20162 ^ n19023 ^ n17913 ;
  assign n26571 = n14559 ^ n3134 ^ 1'b0 ;
  assign n26572 = n10085 & ~n26571 ;
  assign n26573 = n26572 ^ n14443 ^ n6435 ;
  assign n26574 = ( n8511 & n9290 ) | ( n8511 & ~n13169 ) | ( n9290 & ~n13169 ) ;
  assign n26575 = n26574 ^ n10588 ^ n3298 ;
  assign n26576 = n8285 | n26575 ;
  assign n26577 = n26573 | n26576 ;
  assign n26578 = n26577 ^ n15792 ^ 1'b0 ;
  assign n26580 = n10583 ^ n5743 ^ n444 ;
  assign n26579 = n15729 ^ n12424 ^ n3100 ;
  assign n26581 = n26580 ^ n26579 ^ n24728 ;
  assign n26582 = x63 & ~n10976 ;
  assign n26583 = n7466 & n26582 ;
  assign n26584 = n21494 ^ n3856 ^ n1261 ;
  assign n26589 = n15450 ^ n9939 ^ n1044 ;
  assign n26588 = n4476 & ~n5561 ;
  assign n26585 = n6681 ^ n5267 ^ n4465 ;
  assign n26586 = n16001 | n26585 ;
  assign n26587 = n26586 ^ n23231 ^ 1'b0 ;
  assign n26590 = n26589 ^ n26588 ^ n26587 ;
  assign n26591 = n26590 ^ n10585 ^ n2545 ;
  assign n26592 = n9057 | n9581 ;
  assign n26593 = n26592 ^ n11582 ^ 1'b0 ;
  assign n26594 = ( n12052 & n14724 ) | ( n12052 & n26593 ) | ( n14724 & n26593 ) ;
  assign n26595 = n13989 | n22895 ;
  assign n26596 = ( ~n23302 & n26594 ) | ( ~n23302 & n26595 ) | ( n26594 & n26595 ) ;
  assign n26597 = n20989 ^ n12151 ^ 1'b0 ;
  assign n26598 = n24672 ^ n12345 ^ x103 ;
  assign n26599 = ( n14738 & n16101 ) | ( n14738 & n26598 ) | ( n16101 & n26598 ) ;
  assign n26600 = ( n22468 & n26597 ) | ( n22468 & n26599 ) | ( n26597 & n26599 ) ;
  assign n26603 = n10809 ^ n1281 ^ 1'b0 ;
  assign n26604 = n881 & ~n26603 ;
  assign n26601 = n6594 ^ n1737 ^ x225 ;
  assign n26602 = n26601 ^ n24699 ^ n13793 ;
  assign n26605 = n26604 ^ n26602 ^ n15401 ;
  assign n26606 = n26605 ^ n19030 ^ n5587 ;
  assign n26607 = ~n5188 & n13399 ;
  assign n26608 = n19484 & n26607 ;
  assign n26609 = ( n16139 & n20405 ) | ( n16139 & ~n26608 ) | ( n20405 & ~n26608 ) ;
  assign n26616 = n16948 ^ n12542 ^ n7431 ;
  assign n26610 = ~n4863 & n6119 ;
  assign n26611 = n26610 ^ n22172 ^ 1'b0 ;
  assign n26612 = n26611 ^ n13827 ^ 1'b0 ;
  assign n26613 = ~n2317 & n26612 ;
  assign n26614 = ( n9610 & n19794 ) | ( n9610 & n26613 ) | ( n19794 & n26613 ) ;
  assign n26615 = n26614 ^ n25653 ^ n11723 ;
  assign n26617 = n26616 ^ n26615 ^ 1'b0 ;
  assign n26618 = n13015 ^ n1932 ^ n1766 ;
  assign n26619 = ~n1507 & n4676 ;
  assign n26620 = ( ~n14310 & n26618 ) | ( ~n14310 & n26619 ) | ( n26618 & n26619 ) ;
  assign n26621 = n9317 ^ n4535 ^ 1'b0 ;
  assign n26622 = n12116 | n26621 ;
  assign n26623 = n17819 & ~n26622 ;
  assign n26624 = n26623 ^ n1549 ^ 1'b0 ;
  assign n26625 = n26139 ^ n22753 ^ n10512 ;
  assign n26626 = ( ~n6529 & n17220 ) | ( ~n6529 & n26354 ) | ( n17220 & n26354 ) ;
  assign n26627 = n26626 ^ n16884 ^ n9647 ;
  assign n26628 = ( ~n11029 & n14926 ) | ( ~n11029 & n16947 ) | ( n14926 & n16947 ) ;
  assign n26629 = ( ~n4277 & n7519 ) | ( ~n4277 & n22435 ) | ( n7519 & n22435 ) ;
  assign n26630 = n11434 ^ n7089 ^ n379 ;
  assign n26631 = ( ~n12293 & n17777 ) | ( ~n12293 & n26630 ) | ( n17777 & n26630 ) ;
  assign n26632 = n9550 & n26631 ;
  assign n26633 = n13596 & ~n26632 ;
  assign n26634 = ~n3795 & n26633 ;
  assign n26643 = ( ~n847 & n3790 ) | ( ~n847 & n16167 ) | ( n3790 & n16167 ) ;
  assign n26644 = n26643 ^ n13240 ^ n9650 ;
  assign n26635 = ( ~n4612 & n12475 ) | ( ~n4612 & n16156 ) | ( n12475 & n16156 ) ;
  assign n26637 = n5215 ^ n5107 ^ 1'b0 ;
  assign n26638 = n9950 & ~n26637 ;
  assign n26636 = ( ~n821 & n3281 ) | ( ~n821 & n7407 ) | ( n3281 & n7407 ) ;
  assign n26639 = n26638 ^ n26636 ^ n2513 ;
  assign n26640 = n26639 ^ n13301 ^ 1'b0 ;
  assign n26641 = n25083 & n26640 ;
  assign n26642 = n26635 & n26641 ;
  assign n26645 = n26644 ^ n26642 ^ 1'b0 ;
  assign n26646 = n12866 ^ n10503 ^ n8911 ;
  assign n26647 = n26646 ^ n16988 ^ n3711 ;
  assign n26648 = ~n19488 & n21744 ;
  assign n26649 = n5152 & n26648 ;
  assign n26650 = n1133 & ~n26649 ;
  assign n26651 = ~n2518 & n26650 ;
  assign n26652 = n26651 ^ n13601 ^ n12269 ;
  assign n26653 = ( n2955 & n3571 ) | ( n2955 & ~n5152 ) | ( n3571 & ~n5152 ) ;
  assign n26654 = ~n6788 & n14544 ;
  assign n26655 = ( n3515 & n13498 ) | ( n3515 & n26654 ) | ( n13498 & n26654 ) ;
  assign n26656 = n26655 ^ n8254 ^ n8007 ;
  assign n26657 = n10163 & n26153 ;
  assign n26658 = n14673 ^ n8103 ^ n7224 ;
  assign n26659 = ( ~n12338 & n21795 ) | ( ~n12338 & n26658 ) | ( n21795 & n26658 ) ;
  assign n26660 = n26659 ^ n21074 ^ n16207 ;
  assign n26661 = ( n2481 & ~n10788 ) | ( n2481 & n18433 ) | ( ~n10788 & n18433 ) ;
  assign n26662 = n26661 ^ n16523 ^ n12803 ;
  assign n26663 = n26662 ^ n23353 ^ n19680 ;
  assign n26664 = n25238 ^ n21790 ^ n5966 ;
  assign n26665 = n26664 ^ n5450 ^ n3990 ;
  assign n26666 = ( ~n493 & n9189 ) | ( ~n493 & n26665 ) | ( n9189 & n26665 ) ;
  assign n26667 = ( n2579 & ~n19863 ) | ( n2579 & n26666 ) | ( ~n19863 & n26666 ) ;
  assign n26668 = n7721 | n8894 ;
  assign n26669 = n26668 ^ n10306 ^ 1'b0 ;
  assign n26670 = ( n10257 & n22992 ) | ( n10257 & ~n26669 ) | ( n22992 & ~n26669 ) ;
  assign n26671 = n26670 ^ n6106 ^ n3706 ;
  assign n26672 = n26671 ^ n24290 ^ n21646 ;
  assign n26673 = ( n2011 & ~n17805 ) | ( n2011 & n23884 ) | ( ~n17805 & n23884 ) ;
  assign n26678 = n12390 ^ n7876 ^ n5734 ;
  assign n26674 = n1651 | n15002 ;
  assign n26675 = ( n1019 & ~n8235 ) | ( n1019 & n26674 ) | ( ~n8235 & n26674 ) ;
  assign n26676 = n26675 ^ n8346 ^ 1'b0 ;
  assign n26677 = n21106 | n26676 ;
  assign n26679 = n26678 ^ n26677 ^ n11235 ;
  assign n26680 = n26679 ^ n20826 ^ n3225 ;
  assign n26681 = n5683 | n26680 ;
  assign n26682 = n26673 | n26681 ;
  assign n26683 = ( n10062 & n11683 ) | ( n10062 & ~n26682 ) | ( n11683 & ~n26682 ) ;
  assign n26684 = n22664 ^ n16054 ^ n9681 ;
  assign n26685 = n26684 ^ n8977 ^ n2557 ;
  assign n26686 = n10006 ^ n8431 ^ 1'b0 ;
  assign n26687 = n9627 ^ n4020 ^ n2677 ;
  assign n26688 = ( n5134 & ~n9611 ) | ( n5134 & n14031 ) | ( ~n9611 & n14031 ) ;
  assign n26689 = ( ~n5169 & n26687 ) | ( ~n5169 & n26688 ) | ( n26687 & n26688 ) ;
  assign n26690 = n26689 ^ n6293 ^ n4819 ;
  assign n26691 = ( ~n5074 & n16249 ) | ( ~n5074 & n26690 ) | ( n16249 & n26690 ) ;
  assign n26701 = ( n2432 & n4748 ) | ( n2432 & ~n12834 ) | ( n4748 & ~n12834 ) ;
  assign n26702 = n26701 ^ n19667 ^ n13009 ;
  assign n26703 = ~n18291 & n26702 ;
  assign n26704 = n26703 ^ n1229 ^ 1'b0 ;
  assign n26705 = n23734 ^ n22288 ^ n15424 ;
  assign n26706 = ( n4000 & n26704 ) | ( n4000 & ~n26705 ) | ( n26704 & ~n26705 ) ;
  assign n26693 = ( n11339 & ~n11488 ) | ( n11339 & n25823 ) | ( ~n11488 & n25823 ) ;
  assign n26694 = n462 & ~n26693 ;
  assign n26698 = n25796 ^ n2974 ^ n1240 ;
  assign n26695 = ( n311 & n5124 ) | ( n311 & ~n7247 ) | ( n5124 & ~n7247 ) ;
  assign n26696 = ( n3052 & n4743 ) | ( n3052 & n26695 ) | ( n4743 & n26695 ) ;
  assign n26697 = n26696 ^ n16790 ^ n7477 ;
  assign n26699 = n26698 ^ n26697 ^ n548 ;
  assign n26700 = ( n4478 & n26694 ) | ( n4478 & n26699 ) | ( n26694 & n26699 ) ;
  assign n26692 = n9241 ^ n3999 ^ 1'b0 ;
  assign n26707 = n26706 ^ n26700 ^ n26692 ;
  assign n26708 = n11155 ^ n3507 ^ n2695 ;
  assign n26709 = ( n13884 & n18621 ) | ( n13884 & ~n25309 ) | ( n18621 & ~n25309 ) ;
  assign n26710 = ( ~n9633 & n26708 ) | ( ~n9633 & n26709 ) | ( n26708 & n26709 ) ;
  assign n26711 = n19786 ^ n15906 ^ n6303 ;
  assign n26712 = ~n410 & n26711 ;
  assign n26713 = n5729 & n26712 ;
  assign n26714 = n14716 ^ n14529 ^ 1'b0 ;
  assign n26715 = n26713 | n26714 ;
  assign n26716 = n16700 ^ n4801 ^ n2518 ;
  assign n26717 = ~n2112 & n8182 ;
  assign n26718 = n26717 ^ n13899 ^ n1717 ;
  assign n26719 = ( x66 & n5173 ) | ( x66 & ~n13755 ) | ( n5173 & ~n13755 ) ;
  assign n26720 = n3271 & ~n6859 ;
  assign n26721 = ~n21150 & n26720 ;
  assign n26722 = ( n18576 & n26719 ) | ( n18576 & ~n26721 ) | ( n26719 & ~n26721 ) ;
  assign n26723 = ( n11458 & n13645 ) | ( n11458 & ~n15945 ) | ( n13645 & ~n15945 ) ;
  assign n26731 = ( n2768 & ~n3919 ) | ( n2768 & n4510 ) | ( ~n3919 & n4510 ) ;
  assign n26728 = ( n2699 & n7240 ) | ( n2699 & ~n20207 ) | ( n7240 & ~n20207 ) ;
  assign n26727 = n569 & ~n11337 ;
  assign n26729 = n26728 ^ n26727 ^ 1'b0 ;
  assign n26724 = n1869 & n10256 ;
  assign n26725 = ( n16514 & n20540 ) | ( n16514 & ~n26724 ) | ( n20540 & ~n26724 ) ;
  assign n26726 = ( n4493 & n13478 ) | ( n4493 & ~n26725 ) | ( n13478 & ~n26725 ) ;
  assign n26730 = n26729 ^ n26726 ^ n14104 ;
  assign n26732 = n26731 ^ n26730 ^ 1'b0 ;
  assign n26733 = n10557 ^ n5426 ^ n3570 ;
  assign n26734 = n19153 | n26733 ;
  assign n26735 = n26734 ^ n17493 ^ 1'b0 ;
  assign n26736 = n20111 ^ n10790 ^ n3497 ;
  assign n26738 = n8448 ^ n6201 ^ n4793 ;
  assign n26739 = ( ~n3154 & n3303 ) | ( ~n3154 & n26738 ) | ( n3303 & n26738 ) ;
  assign n26740 = n3065 | n26739 ;
  assign n26741 = n6048 & ~n26740 ;
  assign n26742 = n26741 ^ n13257 ^ 1'b0 ;
  assign n26743 = n1151 & ~n11469 ;
  assign n26744 = n26743 ^ n5961 ^ 1'b0 ;
  assign n26745 = ( n1171 & n26742 ) | ( n1171 & n26744 ) | ( n26742 & n26744 ) ;
  assign n26737 = n25407 ^ n22802 ^ n16349 ;
  assign n26746 = n26745 ^ n26737 ^ n19712 ;
  assign n26747 = n11539 & n23313 ;
  assign n26748 = n11673 ^ n4230 ^ 1'b0 ;
  assign n26749 = ( ~n3201 & n12188 ) | ( ~n3201 & n20622 ) | ( n12188 & n20622 ) ;
  assign n26757 = ( n910 & ~n15401 ) | ( n910 & n24579 ) | ( ~n15401 & n24579 ) ;
  assign n26758 = n26757 ^ n22797 ^ n1741 ;
  assign n26759 = ( n10508 & n10643 ) | ( n10508 & n26758 ) | ( n10643 & n26758 ) ;
  assign n26756 = n16269 ^ n11996 ^ n7855 ;
  assign n26760 = n26759 ^ n26756 ^ n22168 ;
  assign n26752 = n3428 ^ n977 ^ 1'b0 ;
  assign n26753 = n5792 & ~n26752 ;
  assign n26750 = n5226 ^ n3636 ^ n2752 ;
  assign n26751 = n5287 & ~n26750 ;
  assign n26754 = n26753 ^ n26751 ^ n13472 ;
  assign n26755 = n26754 ^ n6934 ^ n465 ;
  assign n26761 = n26760 ^ n26755 ^ n14431 ;
  assign n26763 = n17015 ^ n15471 ^ 1'b0 ;
  assign n26762 = n6554 & ~n17799 ;
  assign n26764 = n26763 ^ n26762 ^ 1'b0 ;
  assign n26765 = ( ~n5274 & n12097 ) | ( ~n5274 & n26764 ) | ( n12097 & n26764 ) ;
  assign n26766 = ( ~n2118 & n8839 ) | ( ~n2118 & n16485 ) | ( n8839 & n16485 ) ;
  assign n26767 = n9866 ^ n5494 ^ n4690 ;
  assign n26768 = ( n9116 & ~n16221 ) | ( n9116 & n26767 ) | ( ~n16221 & n26767 ) ;
  assign n26773 = n3880 | n5733 ;
  assign n26774 = ( n2106 & n6735 ) | ( n2106 & n26773 ) | ( n6735 & n26773 ) ;
  assign n26775 = n26774 ^ n5686 ^ n3921 ;
  assign n26769 = ( ~n305 & n9183 ) | ( ~n305 & n13757 ) | ( n9183 & n13757 ) ;
  assign n26770 = n26769 ^ n13710 ^ n9394 ;
  assign n26771 = n26770 ^ n1859 ^ 1'b0 ;
  assign n26772 = ~n964 & n26771 ;
  assign n26776 = n26775 ^ n26772 ^ n25880 ;
  assign n26777 = n9547 ^ n6263 ^ n3846 ;
  assign n26778 = n26777 ^ n20192 ^ n5242 ;
  assign n26780 = n24454 ^ n5894 ^ n5096 ;
  assign n26779 = ( n433 & ~n3064 ) | ( n433 & n15246 ) | ( ~n3064 & n15246 ) ;
  assign n26781 = n26780 ^ n26779 ^ n22184 ;
  assign n26782 = n26781 ^ n16291 ^ n13003 ;
  assign n26785 = n5395 ^ n2681 ^ 1'b0 ;
  assign n26783 = n16203 ^ n8657 ^ n2044 ;
  assign n26784 = n26783 ^ n922 ^ x222 ;
  assign n26786 = n26785 ^ n26784 ^ n13143 ;
  assign n26787 = ( n7002 & n10512 ) | ( n7002 & n15091 ) | ( n10512 & n15091 ) ;
  assign n26788 = ( n9544 & ~n10277 ) | ( n9544 & n13031 ) | ( ~n10277 & n13031 ) ;
  assign n26789 = n1350 & n22551 ;
  assign n26790 = n26788 & n26789 ;
  assign n26791 = n26790 ^ n7601 ^ n4340 ;
  assign n26792 = ( n1917 & ~n3795 ) | ( n1917 & n9840 ) | ( ~n3795 & n9840 ) ;
  assign n26793 = n7154 & n26792 ;
  assign n26794 = ( ~n22985 & n24631 ) | ( ~n22985 & n26793 ) | ( n24631 & n26793 ) ;
  assign n26795 = n3073 & ~n6570 ;
  assign n26796 = ( n2039 & ~n6350 ) | ( n2039 & n21834 ) | ( ~n6350 & n21834 ) ;
  assign n26797 = ~n1646 & n1905 ;
  assign n26798 = ~n460 & n26797 ;
  assign n26799 = n4616 ^ n3951 ^ 1'b0 ;
  assign n26800 = n1391 & n26799 ;
  assign n26801 = ( n26796 & ~n26798 ) | ( n26796 & n26800 ) | ( ~n26798 & n26800 ) ;
  assign n26802 = ( ~n26794 & n26795 ) | ( ~n26794 & n26801 ) | ( n26795 & n26801 ) ;
  assign n26803 = n11158 ^ n9071 ^ n3279 ;
  assign n26804 = n26803 ^ n10979 ^ n2780 ;
  assign n26805 = ( n2394 & n15842 ) | ( n2394 & n23348 ) | ( n15842 & n23348 ) ;
  assign n26806 = ( n5445 & n15746 ) | ( n5445 & n19104 ) | ( n15746 & n19104 ) ;
  assign n26807 = n26806 ^ n22120 ^ n17564 ;
  assign n26808 = n4024 & n9432 ;
  assign n26809 = n12067 & n26808 ;
  assign n26810 = n19714 ^ n6494 ^ n4830 ;
  assign n26811 = ( n9520 & n14953 ) | ( n9520 & n26810 ) | ( n14953 & n26810 ) ;
  assign n26812 = n6498 & n6630 ;
  assign n26813 = n26812 ^ n1521 ^ 1'b0 ;
  assign n26814 = n13797 ^ n5788 ^ 1'b0 ;
  assign n26815 = ~n26813 & n26814 ;
  assign n26816 = n26815 ^ n5601 ^ n3912 ;
  assign n26817 = ( n1505 & ~n3420 ) | ( n1505 & n18947 ) | ( ~n3420 & n18947 ) ;
  assign n26818 = ( n23901 & n25090 ) | ( n23901 & n26817 ) | ( n25090 & n26817 ) ;
  assign n26819 = ( ~n2203 & n8706 ) | ( ~n2203 & n11641 ) | ( n8706 & n11641 ) ;
  assign n26820 = ( n11546 & n15144 ) | ( n11546 & n26819 ) | ( n15144 & n26819 ) ;
  assign n26821 = ( n12113 & n21981 ) | ( n12113 & n26820 ) | ( n21981 & n26820 ) ;
  assign n26822 = ( n11688 & ~n13940 ) | ( n11688 & n15778 ) | ( ~n13940 & n15778 ) ;
  assign n26823 = ( n18300 & ~n24593 ) | ( n18300 & n26822 ) | ( ~n24593 & n26822 ) ;
  assign n26824 = n26823 ^ n14707 ^ n4319 ;
  assign n26825 = ( ~n26818 & n26821 ) | ( ~n26818 & n26824 ) | ( n26821 & n26824 ) ;
  assign n26828 = ( n2528 & ~n7912 ) | ( n2528 & n13335 ) | ( ~n7912 & n13335 ) ;
  assign n26826 = ( ~n4746 & n6413 ) | ( ~n4746 & n10095 ) | ( n6413 & n10095 ) ;
  assign n26827 = n26826 ^ n8722 ^ n3197 ;
  assign n26829 = n26828 ^ n26827 ^ n16741 ;
  assign n26830 = ( n7748 & n8637 ) | ( n7748 & n26829 ) | ( n8637 & n26829 ) ;
  assign n26831 = ~n26694 & n26830 ;
  assign n26832 = n26831 ^ x227 ^ 1'b0 ;
  assign n26833 = n26832 ^ n24415 ^ n16755 ;
  assign n26834 = ( ~n7667 & n10753 ) | ( ~n7667 & n25154 ) | ( n10753 & n25154 ) ;
  assign n26835 = n25006 ^ n14034 ^ n12725 ;
  assign n26836 = ( n5425 & n7764 ) | ( n5425 & n17120 ) | ( n7764 & n17120 ) ;
  assign n26837 = ( n13829 & n26835 ) | ( n13829 & ~n26836 ) | ( n26835 & ~n26836 ) ;
  assign n26838 = ( n1954 & n5918 ) | ( n1954 & n6294 ) | ( n5918 & n6294 ) ;
  assign n26839 = ( n9308 & ~n17530 ) | ( n9308 & n26838 ) | ( ~n17530 & n26838 ) ;
  assign n26840 = n26839 ^ n13647 ^ n484 ;
  assign n26841 = n16920 ^ n16225 ^ n2235 ;
  assign n26842 = ( n5032 & n26840 ) | ( n5032 & ~n26841 ) | ( n26840 & ~n26841 ) ;
  assign n26847 = n14292 ^ n3517 ^ n2647 ;
  assign n26845 = n3100 | n11855 ;
  assign n26846 = n26845 ^ n23368 ^ n13953 ;
  assign n26843 = ( n1565 & ~n3542 ) | ( n1565 & n3668 ) | ( ~n3542 & n3668 ) ;
  assign n26844 = ( n5372 & n9010 ) | ( n5372 & ~n26843 ) | ( n9010 & ~n26843 ) ;
  assign n26848 = n26847 ^ n26846 ^ n26844 ;
  assign n26849 = n11405 ^ n6408 ^ n476 ;
  assign n26850 = n26849 ^ n18330 ^ n3275 ;
  assign n26851 = ( ~n8256 & n11516 ) | ( ~n8256 & n26850 ) | ( n11516 & n26850 ) ;
  assign n26852 = ( ~n13895 & n26848 ) | ( ~n13895 & n26851 ) | ( n26848 & n26851 ) ;
  assign n26853 = n5953 | n13660 ;
  assign n26854 = n26853 ^ n13035 ^ 1'b0 ;
  assign n26855 = n26854 ^ n10298 ^ n7552 ;
  assign n26858 = ( n2864 & n6279 ) | ( n2864 & n8854 ) | ( n6279 & n8854 ) ;
  assign n26859 = n26858 ^ n12489 ^ n4557 ;
  assign n26856 = n8784 ^ n5646 ^ x90 ;
  assign n26857 = n26856 ^ n17595 ^ n2407 ;
  assign n26860 = n26859 ^ n26857 ^ 1'b0 ;
  assign n26861 = ( n2850 & n3180 ) | ( n2850 & n4865 ) | ( n3180 & n4865 ) ;
  assign n26862 = n26861 ^ n26044 ^ n5507 ;
  assign n26863 = ( n364 & n12577 ) | ( n364 & ~n24550 ) | ( n12577 & ~n24550 ) ;
  assign n26864 = n19953 ^ n5848 ^ 1'b0 ;
  assign n26865 = ( n26862 & n26863 ) | ( n26862 & n26864 ) | ( n26863 & n26864 ) ;
  assign n26866 = n14347 ^ n12739 ^ n5876 ;
  assign n26867 = n26866 ^ n26856 ^ n9104 ;
  assign n26868 = n8171 ^ n5377 ^ n5338 ;
  assign n26869 = n3771 | n26868 ;
  assign n26870 = n26867 & ~n26869 ;
  assign n26871 = ( n26860 & n26865 ) | ( n26860 & ~n26870 ) | ( n26865 & ~n26870 ) ;
  assign n26872 = n25739 ^ n13172 ^ n3191 ;
  assign n26873 = n23090 ^ n12142 ^ n4117 ;
  assign n26874 = n26873 ^ n11479 ^ n5927 ;
  assign n26875 = n26874 ^ n22238 ^ n20104 ;
  assign n26876 = ( n5291 & ~n18842 ) | ( n5291 & n21651 ) | ( ~n18842 & n21651 ) ;
  assign n26877 = n5072 ^ n3254 ^ 1'b0 ;
  assign n26878 = n26876 | n26877 ;
  assign n26879 = n25897 ^ n934 ^ x56 ;
  assign n26880 = ( ~n7316 & n12257 ) | ( ~n7316 & n14185 ) | ( n12257 & n14185 ) ;
  assign n26881 = n26880 ^ n17119 ^ n6453 ;
  assign n26882 = ~n4832 & n16556 ;
  assign n26883 = n26882 ^ n24155 ^ n22085 ;
  assign n26884 = ( n10879 & n26881 ) | ( n10879 & ~n26883 ) | ( n26881 & ~n26883 ) ;
  assign n26885 = ~n23922 & n26884 ;
  assign n26886 = n26885 ^ n19491 ^ 1'b0 ;
  assign n26887 = n26886 ^ n13282 ^ n13068 ;
  assign n26891 = n18050 ^ n17221 ^ n17120 ;
  assign n26888 = n2618 & ~n8067 ;
  assign n26889 = n26888 ^ n7479 ^ 1'b0 ;
  assign n26890 = n26889 ^ n18815 ^ n13523 ;
  assign n26892 = n26891 ^ n26890 ^ 1'b0 ;
  assign n26893 = ~n298 & n2288 ;
  assign n26894 = n11812 ^ n5514 ^ n1663 ;
  assign n26895 = ( ~n16935 & n26893 ) | ( ~n16935 & n26894 ) | ( n26893 & n26894 ) ;
  assign n26896 = n5876 ^ n1763 ^ 1'b0 ;
  assign n26897 = n26896 ^ n25867 ^ n933 ;
  assign n26898 = n8642 & ~n26897 ;
  assign n26899 = ~n827 & n26898 ;
  assign n26900 = ( n4833 & n19394 ) | ( n4833 & n26899 ) | ( n19394 & n26899 ) ;
  assign n26901 = n5226 ^ n4086 ^ n2778 ;
  assign n26902 = n26901 ^ n16243 ^ n6972 ;
  assign n26903 = n26902 ^ n5884 ^ n1576 ;
  assign n26904 = n26903 ^ n22667 ^ 1'b0 ;
  assign n26907 = ( n502 & n11081 ) | ( n502 & n13016 ) | ( n11081 & n13016 ) ;
  assign n26905 = ( n1649 & ~n2785 ) | ( n1649 & n5257 ) | ( ~n2785 & n5257 ) ;
  assign n26906 = ~n5204 & n26905 ;
  assign n26908 = n26907 ^ n26906 ^ 1'b0 ;
  assign n26909 = n10671 ^ n8624 ^ n4376 ;
  assign n26910 = ( n18460 & n26908 ) | ( n18460 & ~n26909 ) | ( n26908 & ~n26909 ) ;
  assign n26911 = ( ~n11675 & n19142 ) | ( ~n11675 & n20570 ) | ( n19142 & n20570 ) ;
  assign n26912 = n26911 ^ n17468 ^ n1981 ;
  assign n26913 = ( n18919 & n21682 ) | ( n18919 & n26912 ) | ( n21682 & n26912 ) ;
  assign n26914 = n22430 ^ n18740 ^ n1690 ;
  assign n26915 = n18960 ^ x184 ^ 1'b0 ;
  assign n26916 = n26446 | n26915 ;
  assign n26917 = n10069 ^ n3958 ^ n2225 ;
  assign n26918 = ~n12551 & n26917 ;
  assign n26920 = n648 | n6609 ;
  assign n26919 = n24109 ^ n15892 ^ n2173 ;
  assign n26921 = n26920 ^ n26919 ^ n11817 ;
  assign n26922 = n16629 & ~n22797 ;
  assign n26923 = n26922 ^ n9112 ^ 1'b0 ;
  assign n26924 = n26923 ^ n7328 ^ 1'b0 ;
  assign n26925 = n26921 | n26924 ;
  assign n26926 = ( n26916 & n26918 ) | ( n26916 & ~n26925 ) | ( n26918 & ~n26925 ) ;
  assign n26927 = n26926 ^ n23559 ^ n6515 ;
  assign n26928 = ( ~n8268 & n26914 ) | ( ~n8268 & n26927 ) | ( n26914 & n26927 ) ;
  assign n26929 = n11347 & ~n16269 ;
  assign n26930 = n15387 & ~n26929 ;
  assign n26931 = n26930 ^ n10195 ^ 1'b0 ;
  assign n26941 = n14972 ^ n3607 ^ 1'b0 ;
  assign n26942 = ~n7184 & n26941 ;
  assign n26943 = ( n13284 & n14652 ) | ( n13284 & n26942 ) | ( n14652 & n26942 ) ;
  assign n26944 = ( n5178 & ~n19343 ) | ( n5178 & n26943 ) | ( ~n19343 & n26943 ) ;
  assign n26940 = n19491 ^ n15887 ^ 1'b0 ;
  assign n26945 = n26944 ^ n26940 ^ n19448 ;
  assign n26932 = n8812 ^ n3852 ^ 1'b0 ;
  assign n26933 = ~n14306 & n26932 ;
  assign n26934 = ( ~n2700 & n13067 ) | ( ~n2700 & n13553 ) | ( n13067 & n13553 ) ;
  assign n26935 = n10255 ^ n4864 ^ 1'b0 ;
  assign n26936 = n26935 ^ n10528 ^ n4709 ;
  assign n26937 = ( n10882 & n25280 ) | ( n10882 & n26936 ) | ( n25280 & n26936 ) ;
  assign n26938 = ( n4077 & n26934 ) | ( n4077 & ~n26937 ) | ( n26934 & ~n26937 ) ;
  assign n26939 = ( n26236 & ~n26933 ) | ( n26236 & n26938 ) | ( ~n26933 & n26938 ) ;
  assign n26946 = n26945 ^ n26939 ^ n17456 ;
  assign n26952 = n19231 ^ n13476 ^ n5931 ;
  assign n26947 = n8856 ^ n2822 ^ 1'b0 ;
  assign n26948 = n2023 | n26947 ;
  assign n26949 = n7518 & ~n26948 ;
  assign n26950 = n26949 ^ n18094 ^ n2254 ;
  assign n26951 = ( n6363 & ~n6394 ) | ( n6363 & n26950 ) | ( ~n6394 & n26950 ) ;
  assign n26953 = n26952 ^ n26951 ^ n6239 ;
  assign n26954 = ( n9333 & n12512 ) | ( n9333 & ~n13803 ) | ( n12512 & ~n13803 ) ;
  assign n26955 = n26954 ^ n20745 ^ n1439 ;
  assign n26956 = n10492 & n16700 ;
  assign n26957 = n3522 & n26956 ;
  assign n26966 = n9185 ^ n1807 ^ n1209 ;
  assign n26967 = ( ~n18057 & n26769 ) | ( ~n18057 & n26966 ) | ( n26769 & n26966 ) ;
  assign n26958 = n24165 ^ n9101 ^ 1'b0 ;
  assign n26959 = n12792 & n26958 ;
  assign n26960 = n12313 & n26959 ;
  assign n26961 = ( ~n1727 & n3281 ) | ( ~n1727 & n14997 ) | ( n3281 & n14997 ) ;
  assign n26962 = n26961 ^ n15727 ^ n7261 ;
  assign n26963 = n4540 & ~n6050 ;
  assign n26964 = ( ~n1707 & n26962 ) | ( ~n1707 & n26963 ) | ( n26962 & n26963 ) ;
  assign n26965 = ( n18188 & n26960 ) | ( n18188 & ~n26964 ) | ( n26960 & ~n26964 ) ;
  assign n26968 = n26967 ^ n26965 ^ n17421 ;
  assign n26969 = ( n3086 & n26957 ) | ( n3086 & n26968 ) | ( n26957 & n26968 ) ;
  assign n26970 = ( n1152 & n6133 ) | ( n1152 & ~n6639 ) | ( n6133 & ~n6639 ) ;
  assign n26971 = ( n748 & ~n13302 ) | ( n748 & n25119 ) | ( ~n13302 & n25119 ) ;
  assign n26972 = n26970 & n26971 ;
  assign n26973 = n26972 ^ n9441 ^ n1197 ;
  assign n26974 = ( n16544 & n21611 ) | ( n16544 & n26793 ) | ( n21611 & n26793 ) ;
  assign n26975 = n3959 | n5570 ;
  assign n26976 = n16239 & ~n26975 ;
  assign n26977 = n12418 ^ n8547 ^ n5032 ;
  assign n26978 = n26977 ^ n22796 ^ n414 ;
  assign n26979 = ( n6982 & n9077 ) | ( n6982 & ~n11597 ) | ( n9077 & ~n11597 ) ;
  assign n26980 = n26979 ^ n7375 ^ 1'b0 ;
  assign n26981 = n2488 | n26980 ;
  assign n26982 = n26981 ^ n22924 ^ n10452 ;
  assign n26985 = ( n9818 & n10042 ) | ( n9818 & ~n19219 ) | ( n10042 & ~n19219 ) ;
  assign n26983 = n1208 | n18278 ;
  assign n26984 = n23570 | n26983 ;
  assign n26986 = n26985 ^ n26984 ^ n15279 ;
  assign n26987 = ( n1011 & ~n1396 ) | ( n1011 & n2395 ) | ( ~n1396 & n2395 ) ;
  assign n26988 = n971 | n26987 ;
  assign n26989 = n26988 ^ n677 ^ 1'b0 ;
  assign n26990 = ( n13992 & n19674 ) | ( n13992 & n26989 ) | ( n19674 & n26989 ) ;
  assign n26991 = n9279 ^ n2965 ^ n1570 ;
  assign n26992 = ~n4235 & n26991 ;
  assign n26993 = ( n4144 & ~n7836 ) | ( n4144 & n24916 ) | ( ~n7836 & n24916 ) ;
  assign n26994 = ( ~n6299 & n24406 ) | ( ~n6299 & n26993 ) | ( n24406 & n26993 ) ;
  assign n26995 = n26994 ^ n3736 ^ n903 ;
  assign n26996 = ( n11590 & ~n15382 ) | ( n11590 & n17845 ) | ( ~n15382 & n17845 ) ;
  assign n27001 = n8617 ^ n840 ^ 1'b0 ;
  assign n27002 = n4402 & n27001 ;
  assign n27003 = n27002 ^ n21661 ^ n6064 ;
  assign n26997 = n10491 ^ n7365 ^ n1189 ;
  assign n26998 = ~n2788 & n6645 ;
  assign n26999 = n26997 & n26998 ;
  assign n27000 = n26999 ^ n23807 ^ n11419 ;
  assign n27004 = n27003 ^ n27000 ^ n6270 ;
  assign n27005 = n5725 & ~n8198 ;
  assign n27006 = ( n853 & n21540 ) | ( n853 & n24680 ) | ( n21540 & n24680 ) ;
  assign n27007 = ( n1052 & n6882 ) | ( n1052 & ~n10311 ) | ( n6882 & ~n10311 ) ;
  assign n27008 = n27007 ^ n23002 ^ n11183 ;
  assign n27009 = n27008 ^ n20545 ^ n7805 ;
  assign n27010 = ( ~n345 & n3014 ) | ( ~n345 & n11889 ) | ( n3014 & n11889 ) ;
  assign n27011 = ( ~n3816 & n25678 ) | ( ~n3816 & n27010 ) | ( n25678 & n27010 ) ;
  assign n27012 = x53 & n9277 ;
  assign n27013 = n18237 ^ n17345 ^ n17269 ;
  assign n27014 = ( ~n15148 & n27012 ) | ( ~n15148 & n27013 ) | ( n27012 & n27013 ) ;
  assign n27015 = n1049 & ~n11826 ;
  assign n27016 = ~n7774 & n27015 ;
  assign n27017 = n27016 ^ n24247 ^ n20350 ;
  assign n27018 = ( n27011 & ~n27014 ) | ( n27011 & n27017 ) | ( ~n27014 & n27017 ) ;
  assign n27019 = n13463 ^ n12967 ^ n6563 ;
  assign n27020 = ( n4075 & n11991 ) | ( n4075 & ~n27019 ) | ( n11991 & ~n27019 ) ;
  assign n27021 = n27020 ^ n20876 ^ n16969 ;
  assign n27022 = n7771 ^ n4462 ^ 1'b0 ;
  assign n27023 = n9203 ^ n8062 ^ n953 ;
  assign n27024 = ( ~n5752 & n10948 ) | ( ~n5752 & n20615 ) | ( n10948 & n20615 ) ;
  assign n27025 = ~n5573 & n14708 ;
  assign n27026 = n27024 & n27025 ;
  assign n27027 = n27023 & ~n27026 ;
  assign n27028 = n27027 ^ n4593 ^ 1'b0 ;
  assign n27029 = n8256 ^ n6517 ^ 1'b0 ;
  assign n27030 = n5419 & ~n27029 ;
  assign n27031 = n9346 ^ n2370 ^ 1'b0 ;
  assign n27032 = ( n11847 & n15104 ) | ( n11847 & n16023 ) | ( n15104 & n16023 ) ;
  assign n27033 = ~n27031 & n27032 ;
  assign n27034 = ~n27030 & n27033 ;
  assign n27035 = ( ~n7986 & n15905 ) | ( ~n7986 & n27034 ) | ( n15905 & n27034 ) ;
  assign n27036 = ( n2761 & n7377 ) | ( n2761 & n13206 ) | ( n7377 & n13206 ) ;
  assign n27037 = ~n3354 & n27036 ;
  assign n27038 = n26198 ^ n25358 ^ x36 ;
  assign n27039 = n20397 ^ n20326 ^ n3520 ;
  assign n27040 = n1281 | n10005 ;
  assign n27041 = n26725 | n27040 ;
  assign n27042 = n27041 ^ n22211 ^ n16653 ;
  assign n27043 = n258 & ~n15575 ;
  assign n27044 = n27042 & n27043 ;
  assign n27045 = n903 & n4025 ;
  assign n27046 = n27045 ^ n14705 ^ n5470 ;
  assign n27047 = n27046 ^ n21821 ^ n20567 ;
  assign n27048 = n26307 ^ n13867 ^ n8323 ;
  assign n27049 = n12855 ^ n8789 ^ n8690 ;
  assign n27054 = ( n3892 & n21309 ) | ( n3892 & n22671 ) | ( n21309 & n22671 ) ;
  assign n27050 = n10013 ^ n3120 ^ n2518 ;
  assign n27051 = n27050 ^ n21777 ^ n9048 ;
  assign n27052 = n22541 ^ n19971 ^ n18775 ;
  assign n27053 = ( n3477 & n27051 ) | ( n3477 & n27052 ) | ( n27051 & n27052 ) ;
  assign n27055 = n27054 ^ n27053 ^ n21731 ;
  assign n27056 = ( n11570 & ~n14497 ) | ( n11570 & n17986 ) | ( ~n14497 & n17986 ) ;
  assign n27057 = n27056 ^ n26754 ^ n16100 ;
  assign n27062 = n7177 ^ n2657 ^ n1546 ;
  assign n27060 = ( n830 & n1937 ) | ( n830 & n12108 ) | ( n1937 & n12108 ) ;
  assign n27058 = n18427 ^ n9052 ^ n6155 ;
  assign n27059 = n27058 ^ n18984 ^ n10410 ;
  assign n27061 = n27060 ^ n27059 ^ n5464 ;
  assign n27063 = n27062 ^ n27061 ^ n12218 ;
  assign n27064 = n12875 ^ n7873 ^ n300 ;
  assign n27065 = n23969 ^ n23556 ^ x83 ;
  assign n27066 = ~n14364 & n27065 ;
  assign n27067 = ~n27064 & n27066 ;
  assign n27068 = n10416 ^ n6207 ^ n3685 ;
  assign n27069 = ( ~n1445 & n8938 ) | ( ~n1445 & n27068 ) | ( n8938 & n27068 ) ;
  assign n27070 = n2022 & ~n16806 ;
  assign n27071 = ~n16467 & n27070 ;
  assign n27072 = ( n4342 & n9560 ) | ( n4342 & n27071 ) | ( n9560 & n27071 ) ;
  assign n27073 = ( n2862 & n7045 ) | ( n2862 & n17836 ) | ( n7045 & n17836 ) ;
  assign n27074 = ( n7448 & ~n19427 ) | ( n7448 & n27073 ) | ( ~n19427 & n27073 ) ;
  assign n27075 = n26188 ^ n14525 ^ n3005 ;
  assign n27076 = n16414 ^ n14760 ^ n9807 ;
  assign n27077 = ( n10257 & ~n27075 ) | ( n10257 & n27076 ) | ( ~n27075 & n27076 ) ;
  assign n27078 = n11910 & ~n21142 ;
  assign n27079 = ( ~n3427 & n4273 ) | ( ~n3427 & n6167 ) | ( n4273 & n6167 ) ;
  assign n27080 = ( n19778 & n26744 ) | ( n19778 & ~n27079 ) | ( n26744 & ~n27079 ) ;
  assign n27081 = n27080 ^ n4122 ^ 1'b0 ;
  assign n27082 = ~n3526 & n27081 ;
  assign n27083 = n18675 & ~n20910 ;
  assign n27084 = n15336 & n27083 ;
  assign n27085 = ( ~n1684 & n7940 ) | ( ~n1684 & n10624 ) | ( n7940 & n10624 ) ;
  assign n27086 = n27085 ^ n8460 ^ n7357 ;
  assign n27087 = n23449 & ~n24145 ;
  assign n27088 = ~n27086 & n27087 ;
  assign n27089 = ( n877 & ~n14804 ) | ( n877 & n27088 ) | ( ~n14804 & n27088 ) ;
  assign n27090 = n10082 & ~n17975 ;
  assign n27091 = n27090 ^ n26156 ^ n18230 ;
  assign n27092 = ( n3552 & n16436 ) | ( n3552 & n24254 ) | ( n16436 & n24254 ) ;
  assign n27093 = n16529 ^ n9523 ^ n4111 ;
  assign n27094 = ( ~n2776 & n8376 ) | ( ~n2776 & n13807 ) | ( n8376 & n13807 ) ;
  assign n27095 = n27094 ^ n13876 ^ n4197 ;
  assign n27096 = ( ~n3712 & n27093 ) | ( ~n3712 & n27095 ) | ( n27093 & n27095 ) ;
  assign n27097 = ( n6126 & n8301 ) | ( n6126 & ~n11552 ) | ( n8301 & ~n11552 ) ;
  assign n27098 = n27097 ^ x15 ^ 1'b0 ;
  assign n27099 = n10773 | n26151 ;
  assign n27100 = n27099 ^ n23846 ^ 1'b0 ;
  assign n27103 = n21682 ^ n14796 ^ n2155 ;
  assign n27102 = n10222 & ~n16547 ;
  assign n27104 = n27103 ^ n27102 ^ n18242 ;
  assign n27101 = ~n23116 & n24022 ;
  assign n27105 = n27104 ^ n27101 ^ 1'b0 ;
  assign n27106 = ( n585 & n19457 ) | ( n585 & n19803 ) | ( n19457 & n19803 ) ;
  assign n27107 = n27106 ^ n16105 ^ 1'b0 ;
  assign n27108 = n27107 ^ n12329 ^ 1'b0 ;
  assign n27109 = ( n3050 & ~n13058 ) | ( n3050 & n20620 ) | ( ~n13058 & n20620 ) ;
  assign n27110 = n27109 ^ n10804 ^ n2911 ;
  assign n27111 = n27110 ^ n26307 ^ n6408 ;
  assign n27112 = n27111 ^ n18880 ^ n8249 ;
  assign n27113 = ( n3819 & n10484 ) | ( n3819 & ~n25366 ) | ( n10484 & ~n25366 ) ;
  assign n27114 = ( ~n383 & n2029 ) | ( ~n383 & n27113 ) | ( n2029 & n27113 ) ;
  assign n27115 = n2042 & ~n4455 ;
  assign n27116 = n4424 & n27115 ;
  assign n27117 = n27116 ^ n2012 ^ n1420 ;
  assign n27118 = ( ~n8776 & n25206 ) | ( ~n8776 & n27117 ) | ( n25206 & n27117 ) ;
  assign n27119 = n27118 ^ n14127 ^ n11490 ;
  assign n27120 = n27119 ^ n14753 ^ n2891 ;
  assign n27122 = ( n17940 & n20644 ) | ( n17940 & n22394 ) | ( n20644 & n22394 ) ;
  assign n27121 = n10778 & ~n25653 ;
  assign n27123 = n27122 ^ n27121 ^ 1'b0 ;
  assign n27124 = ( ~n3375 & n4042 ) | ( ~n3375 & n9728 ) | ( n4042 & n9728 ) ;
  assign n27125 = n27124 ^ n3248 ^ 1'b0 ;
  assign n27126 = n15296 | n27125 ;
  assign n27127 = n10690 & ~n16240 ;
  assign n27128 = ~n11896 & n27127 ;
  assign n27129 = n25861 ^ n25415 ^ n8425 ;
  assign n27130 = ( x44 & ~n7737 ) | ( x44 & n11054 ) | ( ~n7737 & n11054 ) ;
  assign n27131 = n13005 | n19917 ;
  assign n27132 = n27131 ^ n8327 ^ 1'b0 ;
  assign n27133 = ( n15010 & n16237 ) | ( n15010 & n27132 ) | ( n16237 & n27132 ) ;
  assign n27134 = ( n12370 & ~n14337 ) | ( n12370 & n27133 ) | ( ~n14337 & n27133 ) ;
  assign n27135 = n27134 ^ n22777 ^ n13379 ;
  assign n27136 = ( n1548 & n27130 ) | ( n1548 & n27135 ) | ( n27130 & n27135 ) ;
  assign n27137 = n15160 ^ n1859 ^ n1814 ;
  assign n27138 = n27137 ^ n22014 ^ n9066 ;
  assign n27139 = n2867 & n22564 ;
  assign n27141 = n16606 ^ n3903 ^ n3091 ;
  assign n27140 = n1404 & ~n19894 ;
  assign n27142 = n27141 ^ n27140 ^ 1'b0 ;
  assign n27143 = n26984 ^ n2126 ^ 1'b0 ;
  assign n27144 = n27142 & n27143 ;
  assign n27145 = n26356 ^ x56 ^ 1'b0 ;
  assign n27146 = n3945 | n27145 ;
  assign n27147 = ( n8239 & n12558 ) | ( n8239 & n25579 ) | ( n12558 & n25579 ) ;
  assign n27148 = ( n341 & n5434 ) | ( n341 & ~n6858 ) | ( n5434 & ~n6858 ) ;
  assign n27149 = n7987 | n27148 ;
  assign n27150 = n17838 | n19675 ;
  assign n27151 = ( n1183 & ~n6758 ) | ( n1183 & n27150 ) | ( ~n6758 & n27150 ) ;
  assign n27152 = ( n7972 & n16853 ) | ( n7972 & ~n19156 ) | ( n16853 & ~n19156 ) ;
  assign n27153 = ( ~n2943 & n12613 ) | ( ~n2943 & n18902 ) | ( n12613 & n18902 ) ;
  assign n27154 = ( n9368 & n13548 ) | ( n9368 & n20102 ) | ( n13548 & n20102 ) ;
  assign n27155 = n27154 ^ n14364 ^ 1'b0 ;
  assign n27156 = n14274 | n27155 ;
  assign n27158 = n2406 & ~n11677 ;
  assign n27157 = ( ~n6073 & n18775 ) | ( ~n6073 & n19090 ) | ( n18775 & n19090 ) ;
  assign n27159 = n27158 ^ n27157 ^ n5269 ;
  assign n27160 = n15837 ^ n3820 ^ 1'b0 ;
  assign n27161 = ( n5991 & n6384 ) | ( n5991 & n18692 ) | ( n6384 & n18692 ) ;
  assign n27162 = n27161 ^ n17649 ^ n7911 ;
  assign n27163 = n17652 ^ n16021 ^ n13554 ;
  assign n27164 = n11687 ^ n5491 ^ n4074 ;
  assign n27166 = ( ~n5491 & n8737 ) | ( ~n5491 & n12594 ) | ( n8737 & n12594 ) ;
  assign n27165 = n19219 ^ n9759 ^ n5103 ;
  assign n27167 = n27166 ^ n27165 ^ n11930 ;
  assign n27168 = ( n7500 & n27164 ) | ( n7500 & ~n27167 ) | ( n27164 & ~n27167 ) ;
  assign n27169 = n22619 ^ n710 ^ 1'b0 ;
  assign n27170 = n374 & n27169 ;
  assign n27171 = n17561 & n27170 ;
  assign n27172 = ( n603 & n10209 ) | ( n603 & n17787 ) | ( n10209 & n17787 ) ;
  assign n27173 = n27172 ^ n20884 ^ n8079 ;
  assign n27174 = ( ~n3773 & n12164 ) | ( ~n3773 & n27173 ) | ( n12164 & n27173 ) ;
  assign n27176 = n23366 ^ n12605 ^ n2351 ;
  assign n27175 = n17443 ^ n15028 ^ n8925 ;
  assign n27177 = n27176 ^ n27175 ^ n23292 ;
  assign n27178 = n13788 ^ n13531 ^ n9588 ;
  assign n27179 = ( ~n5896 & n27177 ) | ( ~n5896 & n27178 ) | ( n27177 & n27178 ) ;
  assign n27180 = n21496 ^ n5244 ^ n2805 ;
  assign n27181 = n22591 ^ n18865 ^ n14611 ;
  assign n27182 = n27181 ^ n22165 ^ n14172 ;
  assign n27184 = ( n5079 & ~n7110 ) | ( n5079 & n15093 ) | ( ~n7110 & n15093 ) ;
  assign n27183 = n9157 ^ n8284 ^ n6982 ;
  assign n27185 = n27184 ^ n27183 ^ n19988 ;
  assign n27189 = ~n2996 & n8353 ;
  assign n27186 = n3859 ^ n3154 ^ n635 ;
  assign n27187 = ( n15134 & ~n20419 ) | ( n15134 & n27186 ) | ( ~n20419 & n27186 ) ;
  assign n27188 = n27187 ^ n27165 ^ n12762 ;
  assign n27190 = n27189 ^ n27188 ^ n26157 ;
  assign n27196 = ~n1762 & n11389 ;
  assign n27197 = n9505 & n27196 ;
  assign n27198 = n27197 ^ n20845 ^ 1'b0 ;
  assign n27199 = ( n6836 & ~n16358 ) | ( n6836 & n27198 ) | ( ~n16358 & n27198 ) ;
  assign n27194 = n7167 ^ n6074 ^ n3490 ;
  assign n27195 = n27194 ^ n23376 ^ n6384 ;
  assign n27191 = n22568 ^ n7049 ^ n2350 ;
  assign n27192 = n8775 & n27191 ;
  assign n27193 = n27192 ^ n4430 ^ n3654 ;
  assign n27200 = n27199 ^ n27195 ^ n27193 ;
  assign n27201 = n14002 ^ n7691 ^ n1658 ;
  assign n27202 = n27201 ^ n9425 ^ n8722 ;
  assign n27203 = n11694 ^ n4694 ^ n3767 ;
  assign n27204 = n27203 ^ n14415 ^ 1'b0 ;
  assign n27205 = n27202 & ~n27204 ;
  assign n27206 = n17178 ^ n15684 ^ n14857 ;
  assign n27207 = ( n3608 & n4220 ) | ( n3608 & n5649 ) | ( n4220 & n5649 ) ;
  assign n27208 = n2773 ^ n1469 ^ 1'b0 ;
  assign n27209 = ( ~n27206 & n27207 ) | ( ~n27206 & n27208 ) | ( n27207 & n27208 ) ;
  assign n27210 = ~n21789 & n27209 ;
  assign n27211 = n27210 ^ n10932 ^ 1'b0 ;
  assign n27212 = n26156 ^ n13140 ^ n13078 ;
  assign n27215 = n15006 ^ n13129 ^ 1'b0 ;
  assign n27213 = n17991 ^ n11564 ^ n9758 ;
  assign n27214 = n27213 ^ n22380 ^ n16762 ;
  assign n27216 = n27215 ^ n27214 ^ 1'b0 ;
  assign n27217 = n22413 ^ n19183 ^ n11925 ;
  assign n27218 = ( n970 & ~n3659 ) | ( n970 & n13728 ) | ( ~n3659 & n13728 ) ;
  assign n27219 = n20924 ^ n11046 ^ n9232 ;
  assign n27220 = ( n3958 & ~n11323 ) | ( n3958 & n27219 ) | ( ~n11323 & n27219 ) ;
  assign n27221 = n4077 ^ n2804 ^ n608 ;
  assign n27222 = ~n16868 & n27221 ;
  assign n27223 = n27222 ^ n6988 ^ 1'b0 ;
  assign n27224 = ( ~n11666 & n27220 ) | ( ~n11666 & n27223 ) | ( n27220 & n27223 ) ;
  assign n27225 = ( ~n26011 & n27218 ) | ( ~n26011 & n27224 ) | ( n27218 & n27224 ) ;
  assign n27226 = n27225 ^ n18254 ^ n3412 ;
  assign n27227 = ( n8071 & ~n16947 ) | ( n8071 & n20341 ) | ( ~n16947 & n20341 ) ;
  assign n27228 = n22300 | n27227 ;
  assign n27229 = n14979 ^ n6064 ^ n2711 ;
  assign n27230 = n9177 ^ n4166 ^ n2413 ;
  assign n27231 = ( n11452 & n16321 ) | ( n11452 & ~n27230 ) | ( n16321 & ~n27230 ) ;
  assign n27232 = ( n25140 & n25831 ) | ( n25140 & n27231 ) | ( n25831 & n27231 ) ;
  assign n27233 = ( n6907 & ~n11400 ) | ( n6907 & n13124 ) | ( ~n11400 & n13124 ) ;
  assign n27234 = ( n2856 & n19249 ) | ( n2856 & ~n27233 ) | ( n19249 & ~n27233 ) ;
  assign n27235 = ( n2540 & ~n13476 ) | ( n2540 & n27234 ) | ( ~n13476 & n27234 ) ;
  assign n27236 = n15162 ^ n13625 ^ n571 ;
  assign n27242 = ( ~n3263 & n5011 ) | ( ~n3263 & n17307 ) | ( n5011 & n17307 ) ;
  assign n27243 = n27242 ^ n6117 ^ n5368 ;
  assign n27237 = n14330 ^ n6347 ^ n4480 ;
  assign n27238 = n27237 ^ n12560 ^ n9538 ;
  assign n27239 = n27238 ^ n3291 ^ n1266 ;
  assign n27240 = ( ~n1762 & n3588 ) | ( ~n1762 & n27239 ) | ( n3588 & n27239 ) ;
  assign n27241 = n27240 ^ n17573 ^ n16758 ;
  assign n27244 = n27243 ^ n27241 ^ n10403 ;
  assign n27246 = n7290 ^ n6137 ^ n3107 ;
  assign n27245 = n12030 ^ n11426 ^ n2711 ;
  assign n27247 = n27246 ^ n27245 ^ n18832 ;
  assign n27248 = ( n937 & n2134 ) | ( n937 & ~n2612 ) | ( n2134 & ~n2612 ) ;
  assign n27249 = ( n4632 & ~n23684 ) | ( n4632 & n27248 ) | ( ~n23684 & n27248 ) ;
  assign n27250 = n27249 ^ n19466 ^ n11639 ;
  assign n27251 = n23219 ^ n20559 ^ n13064 ;
  assign n27253 = ( n3531 & n4782 ) | ( n3531 & ~n6377 ) | ( n4782 & ~n6377 ) ;
  assign n27252 = n11800 ^ n3384 ^ n3216 ;
  assign n27254 = n27253 ^ n27252 ^ n23884 ;
  assign n27255 = n10305 ^ n9655 ^ n3297 ;
  assign n27256 = ( n685 & n13679 ) | ( n685 & ~n27255 ) | ( n13679 & ~n27255 ) ;
  assign n27257 = n27254 | n27256 ;
  assign n27258 = ( n11142 & n27251 ) | ( n11142 & ~n27257 ) | ( n27251 & ~n27257 ) ;
  assign n27259 = n18667 ^ n8159 ^ n2263 ;
  assign n27262 = n9210 ^ n2575 ^ 1'b0 ;
  assign n27263 = n13764 & n27262 ;
  assign n27260 = n23553 ^ n13257 ^ 1'b0 ;
  assign n27261 = ( n8726 & n21817 ) | ( n8726 & ~n27260 ) | ( n21817 & ~n27260 ) ;
  assign n27264 = n27263 ^ n27261 ^ n6726 ;
  assign n27265 = n746 & ~n3815 ;
  assign n27266 = ( n18157 & ~n25602 ) | ( n18157 & n27265 ) | ( ~n25602 & n27265 ) ;
  assign n27268 = n9547 & ~n14222 ;
  assign n27269 = ~n5565 & n27268 ;
  assign n27267 = ( ~n9755 & n10746 ) | ( ~n9755 & n15515 ) | ( n10746 & n15515 ) ;
  assign n27270 = n27269 ^ n27267 ^ n469 ;
  assign n27271 = n27270 ^ n3169 ^ n1108 ;
  assign n27272 = ( n18046 & ~n21574 ) | ( n18046 & n27271 ) | ( ~n21574 & n27271 ) ;
  assign n27273 = ( n7655 & ~n27266 ) | ( n7655 & n27272 ) | ( ~n27266 & n27272 ) ;
  assign n27274 = n14101 ^ n9534 ^ n4789 ;
  assign n27275 = n18974 ^ n7064 ^ n6729 ;
  assign n27276 = n1944 & n4279 ;
  assign n27277 = n27275 & n27276 ;
  assign n27278 = ( n2158 & n6903 ) | ( n2158 & n26673 ) | ( n6903 & n26673 ) ;
  assign n27279 = n7941 ^ n3062 ^ n1849 ;
  assign n27280 = n27279 ^ n24289 ^ n7075 ;
  assign n27281 = n15179 ^ n7848 ^ 1'b0 ;
  assign n27288 = n14680 ^ n3763 ^ n2529 ;
  assign n27282 = n14018 | n22689 ;
  assign n27283 = ( n17092 & ~n21249 ) | ( n17092 & n22783 ) | ( ~n21249 & n22783 ) ;
  assign n27284 = ( n1662 & n6834 ) | ( n1662 & ~n27283 ) | ( n6834 & ~n27283 ) ;
  assign n27285 = ( n20417 & n27282 ) | ( n20417 & n27284 ) | ( n27282 & n27284 ) ;
  assign n27286 = n18770 ^ n16512 ^ 1'b0 ;
  assign n27287 = n27285 & n27286 ;
  assign n27289 = n27288 ^ n27287 ^ n6543 ;
  assign n27290 = n24911 ^ n23527 ^ 1'b0 ;
  assign n27291 = n17676 | n27290 ;
  assign n27292 = n11800 ^ n4374 ^ n4096 ;
  assign n27293 = n11619 ^ n4485 ^ n1489 ;
  assign n27294 = ( ~n18349 & n27292 ) | ( ~n18349 & n27293 ) | ( n27292 & n27293 ) ;
  assign n27295 = ( ~n10115 & n17795 ) | ( ~n10115 & n22002 ) | ( n17795 & n22002 ) ;
  assign n27296 = ( n8672 & n27294 ) | ( n8672 & ~n27295 ) | ( n27294 & ~n27295 ) ;
  assign n27300 = n10988 ^ n3926 ^ n3002 ;
  assign n27301 = n27300 ^ n15669 ^ n8707 ;
  assign n27297 = ( n5407 & n7737 ) | ( n5407 & n7933 ) | ( n7737 & n7933 ) ;
  assign n27298 = n8070 ^ n7930 ^ n1423 ;
  assign n27299 = ( ~n23174 & n27297 ) | ( ~n23174 & n27298 ) | ( n27297 & n27298 ) ;
  assign n27302 = n27301 ^ n27299 ^ n12517 ;
  assign n27303 = n27302 ^ n22340 ^ n1042 ;
  assign n27304 = ( n2557 & ~n22533 ) | ( n2557 & n23249 ) | ( ~n22533 & n23249 ) ;
  assign n27305 = ( n1849 & n3454 ) | ( n1849 & ~n12551 ) | ( n3454 & ~n12551 ) ;
  assign n27306 = n7842 ^ n7029 ^ 1'b0 ;
  assign n27307 = n14945 ^ n13631 ^ n2594 ;
  assign n27308 = ( n3503 & n27306 ) | ( n3503 & ~n27307 ) | ( n27306 & ~n27307 ) ;
  assign n27309 = n13043 | n27308 ;
  assign n27310 = n27309 ^ n14506 ^ 1'b0 ;
  assign n27311 = n26018 ^ n11168 ^ 1'b0 ;
  assign n27312 = n27311 ^ n25669 ^ n21675 ;
  assign n27313 = n18671 ^ n14545 ^ x152 ;
  assign n27314 = n568 & n27313 ;
  assign n27315 = ~n27312 & n27314 ;
  assign n27317 = ( n3589 & n10882 ) | ( n3589 & n17019 ) | ( n10882 & n17019 ) ;
  assign n27316 = n8193 ^ n7405 ^ 1'b0 ;
  assign n27318 = n27317 ^ n27316 ^ n17092 ;
  assign n27319 = n1662 & ~n21852 ;
  assign n27320 = n27319 ^ n3595 ^ 1'b0 ;
  assign n27321 = n27320 ^ n6185 ^ n2230 ;
  assign n27322 = n17553 ^ n12080 ^ n7599 ;
  assign n27323 = n8714 & n27322 ;
  assign n27324 = n27323 ^ n12698 ^ n10249 ;
  assign n27325 = ( n20095 & n20395 ) | ( n20095 & n24996 ) | ( n20395 & n24996 ) ;
  assign n27326 = ( n421 & n3133 ) | ( n421 & n9039 ) | ( n3133 & n9039 ) ;
  assign n27327 = ( ~n3132 & n14317 ) | ( ~n3132 & n22754 ) | ( n14317 & n22754 ) ;
  assign n27329 = n1317 | n8047 ;
  assign n27330 = n27329 ^ n9301 ^ 1'b0 ;
  assign n27328 = n7728 ^ n6895 ^ 1'b0 ;
  assign n27331 = n27330 ^ n27328 ^ n22713 ;
  assign n27332 = ( ~n23097 & n27327 ) | ( ~n23097 & n27331 ) | ( n27327 & n27331 ) ;
  assign n27333 = ( n8576 & ~n27326 ) | ( n8576 & n27332 ) | ( ~n27326 & n27332 ) ;
  assign n27334 = ( ~n266 & n5007 ) | ( ~n266 & n25359 ) | ( n5007 & n25359 ) ;
  assign n27335 = n27334 ^ n22472 ^ n9789 ;
  assign n27336 = ~n454 & n14673 ;
  assign n27337 = n4129 ^ n4074 ^ 1'b0 ;
  assign n27338 = n17290 & n27337 ;
  assign n27339 = ( ~n5111 & n23899 ) | ( ~n5111 & n27338 ) | ( n23899 & n27338 ) ;
  assign n27340 = ( n6192 & n14265 ) | ( n6192 & n27339 ) | ( n14265 & n27339 ) ;
  assign n27341 = n17954 ^ n8047 ^ n7010 ;
  assign n27343 = n14037 ^ n3893 ^ n1469 ;
  assign n27342 = n10663 ^ n2121 ^ n491 ;
  assign n27344 = n27343 ^ n27342 ^ n21465 ;
  assign n27345 = ~n1767 & n8614 ;
  assign n27347 = n21937 ^ n17061 ^ n3151 ;
  assign n27348 = n6239 & n16837 ;
  assign n27349 = n27347 & n27348 ;
  assign n27346 = n27177 ^ n27045 ^ n13108 ;
  assign n27350 = n27349 ^ n27346 ^ 1'b0 ;
  assign n27351 = ( x231 & n13961 ) | ( x231 & ~n17792 ) | ( n13961 & ~n17792 ) ;
  assign n27352 = ~n18229 & n27351 ;
  assign n27353 = n17119 & n27352 ;
  assign n27354 = n27353 ^ n20014 ^ 1'b0 ;
  assign n27355 = n27354 ^ n26705 ^ n26098 ;
  assign n27358 = ( n1677 & n3743 ) | ( n1677 & n3990 ) | ( n3743 & n3990 ) ;
  assign n27356 = ( n293 & ~n478 ) | ( n293 & n4103 ) | ( ~n478 & n4103 ) ;
  assign n27357 = ( n4153 & ~n10922 ) | ( n4153 & n27356 ) | ( ~n10922 & n27356 ) ;
  assign n27359 = n27358 ^ n27357 ^ 1'b0 ;
  assign n27360 = ~n10461 & n27359 ;
  assign n27361 = n27360 ^ n17365 ^ n3654 ;
  assign n27363 = ( n1519 & n6087 ) | ( n1519 & ~n8430 ) | ( n6087 & ~n8430 ) ;
  assign n27364 = n27363 ^ n23991 ^ n9017 ;
  assign n27362 = n17084 ^ n16768 ^ n10690 ;
  assign n27365 = n27364 ^ n27362 ^ n7712 ;
  assign n27366 = n14214 ^ n9108 ^ n2709 ;
  assign n27367 = ( n2735 & ~n12567 ) | ( n2735 & n27366 ) | ( ~n12567 & n27366 ) ;
  assign n27368 = n25910 ^ n24680 ^ n10055 ;
  assign n27373 = n12337 ^ n8260 ^ n7698 ;
  assign n27369 = ( n1074 & n2785 ) | ( n1074 & ~n17789 ) | ( n2785 & ~n17789 ) ;
  assign n27370 = n27369 ^ n19590 ^ n12513 ;
  assign n27371 = ( ~n4480 & n13229 ) | ( ~n4480 & n27370 ) | ( n13229 & n27370 ) ;
  assign n27372 = n27371 ^ n12050 ^ 1'b0 ;
  assign n27374 = n27373 ^ n27372 ^ n3616 ;
  assign n27375 = n27356 | n27374 ;
  assign n27376 = n27375 ^ n6659 ^ 1'b0 ;
  assign n27377 = ( n27367 & ~n27368 ) | ( n27367 & n27376 ) | ( ~n27368 & n27376 ) ;
  assign n27378 = ( ~n1448 & n27365 ) | ( ~n1448 & n27377 ) | ( n27365 & n27377 ) ;
  assign n27379 = n17276 ^ n6007 ^ n1460 ;
  assign n27380 = n17430 ^ n1063 ^ 1'b0 ;
  assign n27381 = n27380 ^ n12557 ^ n8338 ;
  assign n27382 = n21963 ^ n1512 ^ n1276 ;
  assign n27383 = n9375 & n22620 ;
  assign n27384 = ( n7646 & n27382 ) | ( n7646 & n27383 ) | ( n27382 & n27383 ) ;
  assign n27385 = n27384 ^ n12967 ^ n4085 ;
  assign n27386 = ( n27379 & n27381 ) | ( n27379 & n27385 ) | ( n27381 & n27385 ) ;
  assign n27392 = n6455 & n7931 ;
  assign n27393 = n27392 ^ x73 ^ 1'b0 ;
  assign n27390 = n8657 ^ n6708 ^ n5704 ;
  assign n27391 = n27390 ^ n11494 ^ n2487 ;
  assign n27388 = n25366 ^ n11208 ^ n9711 ;
  assign n27387 = n10211 ^ n2969 ^ n297 ;
  assign n27389 = n27388 ^ n27387 ^ n880 ;
  assign n27394 = n27393 ^ n27391 ^ n27389 ;
  assign n27395 = n21070 ^ n8357 ^ n8014 ;
  assign n27398 = ( ~n977 & n14972 ) | ( ~n977 & n16335 ) | ( n14972 & n16335 ) ;
  assign n27399 = ( ~n7027 & n15122 ) | ( ~n7027 & n27398 ) | ( n15122 & n27398 ) ;
  assign n27400 = ( n3621 & n17982 ) | ( n3621 & ~n27399 ) | ( n17982 & ~n27399 ) ;
  assign n27396 = n4118 ^ n3677 ^ n2277 ;
  assign n27397 = n27396 ^ n26307 ^ n17084 ;
  assign n27401 = n27400 ^ n27397 ^ n13932 ;
  assign n27402 = n27401 ^ n18735 ^ n2620 ;
  assign n27403 = ( n1929 & n2685 ) | ( n1929 & ~n8660 ) | ( n2685 & ~n8660 ) ;
  assign n27404 = n27403 ^ n6158 ^ 1'b0 ;
  assign n27405 = ~n18175 & n27404 ;
  assign n27406 = n27405 ^ n19039 ^ n17705 ;
  assign n27407 = n26850 ^ n23406 ^ n9983 ;
  assign n27408 = ( n11238 & n11816 ) | ( n11238 & ~n27407 ) | ( n11816 & ~n27407 ) ;
  assign n27409 = n27408 ^ n15784 ^ n5167 ;
  assign n27410 = n11588 ^ n6294 ^ n1194 ;
  assign n27411 = n27410 ^ n13209 ^ n4961 ;
  assign n27412 = ~n2964 & n9385 ;
  assign n27413 = n6851 & n27412 ;
  assign n27414 = x30 | n27413 ;
  assign n27415 = ( n4625 & ~n7095 ) | ( n4625 & n27414 ) | ( ~n7095 & n27414 ) ;
  assign n27416 = n27415 ^ n26881 ^ n21996 ;
  assign n27417 = n27416 ^ n25532 ^ n997 ;
  assign n27418 = ( n6605 & n11013 ) | ( n6605 & ~n12318 ) | ( n11013 & ~n12318 ) ;
  assign n27419 = ( ~n1127 & n4051 ) | ( ~n1127 & n22936 ) | ( n4051 & n22936 ) ;
  assign n27420 = n27419 ^ n7042 ^ n1164 ;
  assign n27421 = ( n5946 & ~n25059 ) | ( n5946 & n27420 ) | ( ~n25059 & n27420 ) ;
  assign n27422 = n12604 & n18053 ;
  assign n27423 = n27422 ^ n16863 ^ 1'b0 ;
  assign n27425 = ( n7786 & n10218 ) | ( n7786 & n16906 ) | ( n10218 & n16906 ) ;
  assign n27426 = ( n5169 & ~n17634 ) | ( n5169 & n21129 ) | ( ~n17634 & n21129 ) ;
  assign n27427 = ( n8666 & n27425 ) | ( n8666 & ~n27426 ) | ( n27425 & ~n27426 ) ;
  assign n27428 = ( n2817 & n16726 ) | ( n2817 & ~n27427 ) | ( n16726 & ~n27427 ) ;
  assign n27424 = n20619 ^ n12797 ^ n8985 ;
  assign n27429 = n27428 ^ n27424 ^ n8496 ;
  assign n27430 = n14540 ^ n992 ^ x212 ;
  assign n27431 = ( n13485 & n17735 ) | ( n13485 & ~n25823 ) | ( n17735 & ~n25823 ) ;
  assign n27432 = ( n22235 & ~n27198 ) | ( n22235 & n27431 ) | ( ~n27198 & n27431 ) ;
  assign n27433 = n5372 & n9322 ;
  assign n27434 = ( n6709 & n26954 ) | ( n6709 & n27433 ) | ( n26954 & n27433 ) ;
  assign n27435 = n27434 ^ n5660 ^ 1'b0 ;
  assign n27436 = ~n27432 & n27435 ;
  assign n27437 = ( n12912 & n27430 ) | ( n12912 & ~n27436 ) | ( n27430 & ~n27436 ) ;
  assign n27438 = n9401 & ~n27437 ;
  assign n27439 = n27438 ^ n22392 ^ 1'b0 ;
  assign n27440 = n1047 & n10030 ;
  assign n27441 = n27440 ^ n20107 ^ 1'b0 ;
  assign n27442 = n21595 ^ n1172 ^ 1'b0 ;
  assign n27443 = ( n21063 & n27224 ) | ( n21063 & n27442 ) | ( n27224 & n27442 ) ;
  assign n27444 = ( n5347 & n27441 ) | ( n5347 & ~n27443 ) | ( n27441 & ~n27443 ) ;
  assign n27445 = n25803 | n27243 ;
  assign n27446 = ( ~x203 & n20667 ) | ( ~x203 & n27445 ) | ( n20667 & n27445 ) ;
  assign n27454 = ( n498 & n1618 ) | ( n498 & n8601 ) | ( n1618 & n8601 ) ;
  assign n27448 = n24192 ^ n18563 ^ n16606 ;
  assign n27449 = n9909 | n27448 ;
  assign n27450 = n27449 ^ n10646 ^ 1'b0 ;
  assign n27451 = ( n11617 & n14625 ) | ( n11617 & n27450 ) | ( n14625 & n27450 ) ;
  assign n27447 = ( ~n8444 & n11941 ) | ( ~n8444 & n25673 ) | ( n11941 & n25673 ) ;
  assign n27452 = n27451 ^ n27447 ^ n21703 ;
  assign n27453 = n27452 ^ n21054 ^ 1'b0 ;
  assign n27455 = n27454 ^ n27453 ^ n12827 ;
  assign n27464 = n25729 ^ n1984 ^ n1629 ;
  assign n27465 = ( n7136 & n15274 ) | ( n7136 & ~n27464 ) | ( n15274 & ~n27464 ) ;
  assign n27461 = n848 & ~n11397 ;
  assign n27462 = n27461 ^ n5192 ^ 1'b0 ;
  assign n27463 = n27462 ^ n19500 ^ n5909 ;
  assign n27466 = n27465 ^ n27463 ^ 1'b0 ;
  assign n27456 = ( ~n1424 & n3922 ) | ( ~n1424 & n6379 ) | ( n3922 & n6379 ) ;
  assign n27457 = n23394 & ~n27456 ;
  assign n27458 = n27457 ^ n7666 ^ 1'b0 ;
  assign n27459 = n12612 | n27458 ;
  assign n27460 = ( n17130 & n21144 ) | ( n17130 & n27459 ) | ( n21144 & n27459 ) ;
  assign n27467 = n27466 ^ n27460 ^ n2938 ;
  assign n27468 = n7727 | n19475 ;
  assign n27469 = n27468 ^ n1825 ^ 1'b0 ;
  assign n27470 = ( n4980 & ~n8136 ) | ( n4980 & n27469 ) | ( ~n8136 & n27469 ) ;
  assign n27471 = ( n9869 & n12370 ) | ( n9869 & ~n27470 ) | ( n12370 & ~n27470 ) ;
  assign n27472 = ( n7442 & ~n13970 ) | ( n7442 & n20507 ) | ( ~n13970 & n20507 ) ;
  assign n27473 = n27472 ^ n9819 ^ n5833 ;
  assign n27474 = ( n9128 & n23206 ) | ( n9128 & ~n23922 ) | ( n23206 & ~n23922 ) ;
  assign n27475 = n18514 ^ n11965 ^ 1'b0 ;
  assign n27476 = n17711 ^ n3065 ^ n1668 ;
  assign n27477 = ( n4994 & ~n14663 ) | ( n4994 & n27476 ) | ( ~n14663 & n27476 ) ;
  assign n27478 = n19251 ^ n9807 ^ n5359 ;
  assign n27479 = n27183 & ~n27478 ;
  assign n27480 = ~n18039 & n27479 ;
  assign n27481 = n27480 ^ n22077 ^ n1048 ;
  assign n27482 = ( ~n13517 & n27477 ) | ( ~n13517 & n27481 ) | ( n27477 & n27481 ) ;
  assign n27484 = ( n2974 & n5857 ) | ( n2974 & ~n24082 ) | ( n5857 & ~n24082 ) ;
  assign n27483 = ( n2586 & n4157 ) | ( n2586 & ~n23835 ) | ( n4157 & ~n23835 ) ;
  assign n27485 = n27484 ^ n27483 ^ n9213 ;
  assign n27486 = ( n6620 & n7548 ) | ( n6620 & n27485 ) | ( n7548 & n27485 ) ;
  assign n27487 = n25710 ^ n10205 ^ n9708 ;
  assign n27494 = n20038 ^ n9855 ^ n9747 ;
  assign n27495 = n27494 ^ n13703 ^ n2538 ;
  assign n27496 = n3180 & n10447 ;
  assign n27497 = ~n27495 & n27496 ;
  assign n27492 = ( n923 & n2964 ) | ( n923 & ~n3494 ) | ( n2964 & ~n3494 ) ;
  assign n27493 = ( ~n8017 & n18088 ) | ( ~n8017 & n27492 ) | ( n18088 & n27492 ) ;
  assign n27488 = n21817 ^ n3206 ^ 1'b0 ;
  assign n27489 = ~n6409 & n27488 ;
  assign n27490 = n27489 ^ n19641 ^ n515 ;
  assign n27491 = n27490 ^ n25427 ^ n3170 ;
  assign n27498 = n27497 ^ n27493 ^ n27491 ;
  assign n27499 = n4029 ^ n2978 ^ 1'b0 ;
  assign n27500 = n4182 | n27499 ;
  assign n27501 = n5832 & n27500 ;
  assign n27502 = n27501 ^ n8931 ^ 1'b0 ;
  assign n27503 = ( n6336 & ~n19815 ) | ( n6336 & n27502 ) | ( ~n19815 & n27502 ) ;
  assign n27504 = n22352 ^ n19000 ^ n2513 ;
  assign n27505 = n27504 ^ n24331 ^ n10062 ;
  assign n27506 = n18079 ^ n13105 ^ n384 ;
  assign n27507 = ( n981 & ~n2261 ) | ( n981 & n27506 ) | ( ~n2261 & n27506 ) ;
  assign n27508 = n27507 ^ n24570 ^ n20559 ;
  assign n27509 = n18358 ^ n10948 ^ n1718 ;
  assign n27510 = ( n2072 & ~n12651 ) | ( n2072 & n27509 ) | ( ~n12651 & n27509 ) ;
  assign n27511 = n14612 & n19450 ;
  assign n27512 = n27511 ^ n12239 ^ 1'b0 ;
  assign n27513 = ( ~n26847 & n27510 ) | ( ~n26847 & n27512 ) | ( n27510 & n27512 ) ;
  assign n27514 = n27513 ^ n15234 ^ n13220 ;
  assign n27515 = n24066 ^ n16714 ^ n8754 ;
  assign n27516 = n27515 ^ n13135 ^ n6414 ;
  assign n27517 = n3815 ^ n2979 ^ 1'b0 ;
  assign n27518 = ~n2943 & n27517 ;
  assign n27519 = n27518 ^ n2007 ^ n1383 ;
  assign n27520 = n27519 ^ n13659 ^ n700 ;
  assign n27521 = n12766 ^ n1972 ^ 1'b0 ;
  assign n27522 = n27520 & n27521 ;
  assign n27523 = ~n8895 & n25471 ;
  assign n27524 = ~n27522 & n27523 ;
  assign n27525 = n19549 ^ n5607 ^ 1'b0 ;
  assign n27526 = n27524 | n27525 ;
  assign n27527 = n27526 ^ n21012 ^ n4965 ;
  assign n27528 = ( ~n4592 & n22554 ) | ( ~n4592 & n26701 ) | ( n22554 & n26701 ) ;
  assign n27529 = ( x185 & n2205 ) | ( x185 & n22282 ) | ( n2205 & n22282 ) ;
  assign n27530 = ( ~n9827 & n27528 ) | ( ~n9827 & n27529 ) | ( n27528 & n27529 ) ;
  assign n27534 = n12295 ^ n6934 ^ n2793 ;
  assign n27531 = n25728 ^ n19284 ^ n11140 ;
  assign n27532 = n27531 ^ n12433 ^ n8610 ;
  assign n27533 = ( n4500 & ~n7859 ) | ( n4500 & n27532 ) | ( ~n7859 & n27532 ) ;
  assign n27535 = n27534 ^ n27533 ^ n2221 ;
  assign n27536 = ( n13628 & n14259 ) | ( n13628 & ~n16459 ) | ( n14259 & ~n16459 ) ;
  assign n27537 = n27536 ^ n25206 ^ 1'b0 ;
  assign n27538 = n13004 ^ n3236 ^ n350 ;
  assign n27539 = n26035 ^ n21824 ^ 1'b0 ;
  assign n27540 = n582 | n9625 ;
  assign n27541 = n13067 | n27540 ;
  assign n27542 = n27541 ^ n19365 ^ 1'b0 ;
  assign n27543 = n26263 & n27542 ;
  assign n27544 = ( n1787 & n18152 ) | ( n1787 & n21795 ) | ( n18152 & n21795 ) ;
  assign n27545 = ( ~n3143 & n9873 ) | ( ~n3143 & n11672 ) | ( n9873 & n11672 ) ;
  assign n27546 = n27545 ^ n10849 ^ 1'b0 ;
  assign n27547 = ~n26971 & n27546 ;
  assign n27548 = ( n1861 & n27544 ) | ( n1861 & ~n27547 ) | ( n27544 & ~n27547 ) ;
  assign n27549 = n18043 ^ n5881 ^ n4169 ;
  assign n27550 = ( n14044 & n19484 ) | ( n14044 & ~n27549 ) | ( n19484 & ~n27549 ) ;
  assign n27551 = ( n9793 & n10793 ) | ( n9793 & ~n27550 ) | ( n10793 & ~n27550 ) ;
  assign n27552 = ( n1621 & n4968 ) | ( n1621 & ~n17990 ) | ( n4968 & ~n17990 ) ;
  assign n27553 = n27552 ^ n20733 ^ n2834 ;
  assign n27556 = ( n2454 & n11630 ) | ( n2454 & ~n25731 ) | ( n11630 & ~n25731 ) ;
  assign n27554 = n12172 ^ n1767 ^ 1'b0 ;
  assign n27555 = ~n9834 & n27554 ;
  assign n27557 = n27556 ^ n27555 ^ n1067 ;
  assign n27558 = ( n10335 & n16408 ) | ( n10335 & ~n22574 ) | ( n16408 & ~n22574 ) ;
  assign n27559 = n27558 ^ n12648 ^ n10377 ;
  assign n27560 = ( n7483 & n14954 ) | ( n7483 & n21712 ) | ( n14954 & n21712 ) ;
  assign n27561 = n27560 ^ n21073 ^ 1'b0 ;
  assign n27562 = n24178 | n27561 ;
  assign n27563 = ( n26316 & n27221 ) | ( n26316 & n27562 ) | ( n27221 & n27562 ) ;
  assign n27564 = n6302 ^ n2268 ^ n312 ;
  assign n27565 = n27564 ^ n7206 ^ n3123 ;
  assign n27566 = n8267 ^ n5061 ^ n1682 ;
  assign n27567 = n27566 ^ n9184 ^ n4594 ;
  assign n27568 = ( ~n836 & n3766 ) | ( ~n836 & n16428 ) | ( n3766 & n16428 ) ;
  assign n27569 = n5425 & n27568 ;
  assign n27570 = ( n27565 & ~n27567 ) | ( n27565 & n27569 ) | ( ~n27567 & n27569 ) ;
  assign n27571 = n27570 ^ n21422 ^ 1'b0 ;
  assign n27572 = n22485 ^ n22164 ^ n21033 ;
  assign n27573 = ( n6808 & ~n14212 ) | ( n6808 & n25123 ) | ( ~n14212 & n25123 ) ;
  assign n27574 = ( n1278 & ~n17264 ) | ( n1278 & n24174 ) | ( ~n17264 & n24174 ) ;
  assign n27575 = n27574 ^ n10203 ^ 1'b0 ;
  assign n27576 = n9659 ^ n498 ^ 1'b0 ;
  assign n27577 = n18273 & ~n27576 ;
  assign n27578 = ~n27575 & n27577 ;
  assign n27581 = n5086 ^ n1240 ^ 1'b0 ;
  assign n27582 = n27581 ^ n6362 ^ n5326 ;
  assign n27583 = n27582 ^ n27351 ^ n929 ;
  assign n27579 = n4602 & ~n26649 ;
  assign n27580 = n6397 & n27579 ;
  assign n27584 = n27583 ^ n27580 ^ n17535 ;
  assign n27585 = n15532 ^ n9092 ^ n6260 ;
  assign n27586 = ( n8050 & n20549 ) | ( n8050 & ~n27585 ) | ( n20549 & ~n27585 ) ;
  assign n27587 = ( ~n14658 & n17601 ) | ( ~n14658 & n25461 ) | ( n17601 & n25461 ) ;
  assign n27589 = ~n3726 & n23010 ;
  assign n27590 = ( ~n1464 & n5883 ) | ( ~n1464 & n8240 ) | ( n5883 & n8240 ) ;
  assign n27591 = ( n22293 & n27589 ) | ( n22293 & n27590 ) | ( n27589 & n27590 ) ;
  assign n27588 = n6539 | n18205 ;
  assign n27592 = n27591 ^ n27588 ^ 1'b0 ;
  assign n27593 = n27592 ^ n4900 ^ n4656 ;
  assign n27594 = ( n2347 & n6048 ) | ( n2347 & ~n6206 ) | ( n6048 & ~n6206 ) ;
  assign n27595 = n25205 ^ n5140 ^ n1169 ;
  assign n27596 = ( n20486 & n27594 ) | ( n20486 & n27595 ) | ( n27594 & n27595 ) ;
  assign n27597 = ( n21392 & ~n27593 ) | ( n21392 & n27596 ) | ( ~n27593 & n27596 ) ;
  assign n27598 = n26064 ^ n21554 ^ n4816 ;
  assign n27599 = n8912 | n27598 ;
  assign n27600 = ( n8790 & n18498 ) | ( n8790 & n27599 ) | ( n18498 & n27599 ) ;
  assign n27601 = n4873 | n18258 ;
  assign n27602 = n27601 ^ n16818 ^ 1'b0 ;
  assign n27603 = n27602 ^ n23790 ^ n14622 ;
  assign n27604 = ( n7206 & n17182 ) | ( n7206 & n25961 ) | ( n17182 & n25961 ) ;
  assign n27605 = n17770 ^ n10542 ^ n10054 ;
  assign n27606 = n6049 ^ n4867 ^ n521 ;
  assign n27607 = ( ~n702 & n5993 ) | ( ~n702 & n27606 ) | ( n5993 & n27606 ) ;
  assign n27608 = n12936 | n27607 ;
  assign n27609 = ( n288 & ~n9298 ) | ( n288 & n25510 ) | ( ~n9298 & n25510 ) ;
  assign n27610 = n19525 ^ n19081 ^ n2629 ;
  assign n27611 = n7476 | n26306 ;
  assign n27612 = n16097 ^ n8457 ^ n1975 ;
  assign n27613 = n22389 ^ n13147 ^ 1'b0 ;
  assign n27614 = ~n27612 & n27613 ;
  assign n27616 = n17707 ^ n11979 ^ 1'b0 ;
  assign n27615 = n12107 ^ n3011 ^ 1'b0 ;
  assign n27617 = n27616 ^ n27615 ^ 1'b0 ;
  assign n27618 = ~n11688 & n27617 ;
  assign n27619 = ( n2305 & n3686 ) | ( n2305 & ~n9447 ) | ( n3686 & ~n9447 ) ;
  assign n27620 = ( n7045 & n7837 ) | ( n7045 & ~n27619 ) | ( n7837 & ~n27619 ) ;
  assign n27621 = n27620 ^ n24771 ^ n24241 ;
  assign n27622 = n15723 ^ n15413 ^ n6921 ;
  assign n27623 = n9292 & n15435 ;
  assign n27624 = ~n9501 & n27623 ;
  assign n27625 = n27624 ^ n17864 ^ n17178 ;
  assign n27626 = n15081 ^ n2166 ^ 1'b0 ;
  assign n27627 = n2999 & ~n27626 ;
  assign n27628 = ~n27625 & n27627 ;
  assign n27630 = ( ~x213 & n6732 ) | ( ~x213 & n17307 ) | ( n6732 & n17307 ) ;
  assign n27629 = ( n809 & n3465 ) | ( n809 & n7849 ) | ( n3465 & n7849 ) ;
  assign n27631 = n27630 ^ n27629 ^ n2265 ;
  assign n27632 = ( ~n15315 & n21427 ) | ( ~n15315 & n24206 ) | ( n21427 & n24206 ) ;
  assign n27633 = ( n9254 & ~n9721 ) | ( n9254 & n27632 ) | ( ~n9721 & n27632 ) ;
  assign n27634 = n10820 ^ n2980 ^ n1157 ;
  assign n27635 = n27634 ^ n17680 ^ n5416 ;
  assign n27638 = ( n2788 & ~n8056 ) | ( n2788 & n8613 ) | ( ~n8056 & n8613 ) ;
  assign n27637 = ( n5117 & n7671 ) | ( n5117 & ~n11529 ) | ( n7671 & ~n11529 ) ;
  assign n27639 = n27638 ^ n27637 ^ n20536 ;
  assign n27636 = ( n3073 & n4356 ) | ( n3073 & n14489 ) | ( n4356 & n14489 ) ;
  assign n27640 = n27639 ^ n27636 ^ n22968 ;
  assign n27641 = n6137 & n27640 ;
  assign n27642 = n5515 & n6094 ;
  assign n27643 = ( ~n3120 & n21997 ) | ( ~n3120 & n27642 ) | ( n21997 & n27642 ) ;
  assign n27644 = n21950 ^ n14214 ^ n13078 ;
  assign n27645 = n27644 ^ n18296 ^ n7927 ;
  assign n27646 = n8913 ^ n7080 ^ n611 ;
  assign n27647 = n27646 ^ n8598 ^ n7943 ;
  assign n27648 = ( ~n4043 & n8399 ) | ( ~n4043 & n23862 ) | ( n8399 & n23862 ) ;
  assign n27649 = n27648 ^ n22324 ^ n2719 ;
  assign n27650 = n18048 ^ n6044 ^ n5703 ;
  assign n27651 = n27650 ^ n19733 ^ n10575 ;
  assign n27652 = n27651 ^ n21976 ^ 1'b0 ;
  assign n27653 = ~n19520 & n27652 ;
  assign n27654 = ( x98 & n453 ) | ( x98 & ~n10479 ) | ( n453 & ~n10479 ) ;
  assign n27655 = n27654 ^ n22214 ^ n16028 ;
  assign n27656 = ( ~n10428 & n20341 ) | ( ~n10428 & n27655 ) | ( n20341 & n27655 ) ;
  assign n27657 = ( ~n1485 & n10764 ) | ( ~n1485 & n12146 ) | ( n10764 & n12146 ) ;
  assign n27658 = n16875 & n20536 ;
  assign n27659 = n21364 & n27658 ;
  assign n27660 = ( n17857 & n19328 ) | ( n17857 & ~n24168 ) | ( n19328 & ~n24168 ) ;
  assign n27661 = ( ~n27657 & n27659 ) | ( ~n27657 & n27660 ) | ( n27659 & n27660 ) ;
  assign n27662 = n19544 ^ n4964 ^ n3385 ;
  assign n27663 = ( n6238 & n6276 ) | ( n6238 & n8171 ) | ( n6276 & n8171 ) ;
  assign n27664 = ( ~n2203 & n16927 ) | ( ~n2203 & n27663 ) | ( n16927 & n27663 ) ;
  assign n27665 = ( ~n21632 & n27662 ) | ( ~n21632 & n27664 ) | ( n27662 & n27664 ) ;
  assign n27666 = n19454 ^ n12783 ^ n9048 ;
  assign n27667 = n21393 ^ n10076 ^ n7236 ;
  assign n27668 = n10542 ^ n5184 ^ 1'b0 ;
  assign n27669 = ( ~n3182 & n27667 ) | ( ~n3182 & n27668 ) | ( n27667 & n27668 ) ;
  assign n27670 = n27669 ^ n21863 ^ n7704 ;
  assign n27671 = ( n4672 & ~n24815 ) | ( n4672 & n25738 ) | ( ~n24815 & n25738 ) ;
  assign n27672 = n27671 ^ n22281 ^ n1746 ;
  assign n27673 = ~n2886 & n27672 ;
  assign n27674 = ( n12859 & ~n13923 ) | ( n12859 & n24206 ) | ( ~n13923 & n24206 ) ;
  assign n27675 = ( ~n11150 & n12385 ) | ( ~n11150 & n27674 ) | ( n12385 & n27674 ) ;
  assign n27676 = n24503 | n27675 ;
  assign n27686 = n19314 ^ n6535 ^ n5594 ;
  assign n27687 = n27686 ^ n26439 ^ n9394 ;
  assign n27683 = n4275 & ~n15692 ;
  assign n27684 = n27683 ^ n14901 ^ 1'b0 ;
  assign n27679 = n5397 ^ n5042 ^ n1662 ;
  assign n27680 = n27679 ^ n9773 ^ 1'b0 ;
  assign n27681 = ~n9860 & n27680 ;
  assign n27682 = ( ~n1083 & n1250 ) | ( ~n1083 & n27681 ) | ( n1250 & n27681 ) ;
  assign n27677 = n10438 ^ n9461 ^ 1'b0 ;
  assign n27678 = n2311 & n27677 ;
  assign n27685 = n27684 ^ n27682 ^ n27678 ;
  assign n27688 = n27687 ^ n27685 ^ n27598 ;
  assign n27689 = n21780 ^ n13627 ^ n1035 ;
  assign n27690 = ( n2247 & ~n3412 ) | ( n2247 & n11770 ) | ( ~n3412 & n11770 ) ;
  assign n27691 = n27690 ^ n5759 ^ n4807 ;
  assign n27692 = n19769 ^ n17845 ^ 1'b0 ;
  assign n27693 = ( n27502 & n27691 ) | ( n27502 & ~n27692 ) | ( n27691 & ~n27692 ) ;
  assign n27696 = ( ~x143 & n716 ) | ( ~x143 & n17084 ) | ( n716 & n17084 ) ;
  assign n27697 = n27696 ^ n11706 ^ 1'b0 ;
  assign n27694 = ( n6510 & n12654 ) | ( n6510 & n19506 ) | ( n12654 & n19506 ) ;
  assign n27695 = n6361 & n27694 ;
  assign n27698 = n27697 ^ n27695 ^ 1'b0 ;
  assign n27699 = ( n5438 & ~n15321 ) | ( n5438 & n26462 ) | ( ~n15321 & n26462 ) ;
  assign n27700 = n25830 ^ n1374 ^ 1'b0 ;
  assign n27701 = n21691 & ~n27700 ;
  assign n27702 = n27699 & n27701 ;
  assign n27703 = n25138 ^ n22895 ^ 1'b0 ;
  assign n27704 = ( n1198 & ~n4630 ) | ( n1198 & n27703 ) | ( ~n4630 & n27703 ) ;
  assign n27705 = ( ~n2559 & n15196 ) | ( ~n2559 & n27704 ) | ( n15196 & n27704 ) ;
  assign n27706 = n7254 ^ n5540 ^ 1'b0 ;
  assign n27707 = ( n3807 & n26357 ) | ( n3807 & ~n27706 ) | ( n26357 & ~n27706 ) ;
  assign n27708 = n27707 ^ n16007 ^ n5567 ;
  assign n27709 = ( n4784 & n12080 ) | ( n4784 & n12399 ) | ( n12080 & n12399 ) ;
  assign n27710 = n14926 | n22096 ;
  assign n27711 = n20483 & ~n27710 ;
  assign n27712 = ( n10725 & n27709 ) | ( n10725 & ~n27711 ) | ( n27709 & ~n27711 ) ;
  assign n27713 = n27356 ^ n15861 ^ n3751 ;
  assign n27714 = n27713 ^ n15316 ^ n10348 ;
  assign n27715 = ( n3354 & n3446 ) | ( n3354 & n7941 ) | ( n3446 & n7941 ) ;
  assign n27716 = n27715 ^ n16252 ^ 1'b0 ;
  assign n27717 = n11513 & n27716 ;
  assign n27718 = n21513 ^ n8976 ^ n2628 ;
  assign n27719 = ( ~n1683 & n12646 ) | ( ~n1683 & n27718 ) | ( n12646 & n27718 ) ;
  assign n27720 = n10607 ^ n9191 ^ 1'b0 ;
  assign n27721 = n27720 ^ n22143 ^ n1349 ;
  assign n27722 = n27721 ^ n17509 ^ n8281 ;
  assign n27723 = n19704 ^ n12631 ^ 1'b0 ;
  assign n27724 = ( ~n389 & n9569 ) | ( ~n389 & n22666 ) | ( n9569 & n22666 ) ;
  assign n27725 = ( n5819 & n14466 ) | ( n5819 & n27724 ) | ( n14466 & n27724 ) ;
  assign n27726 = n8572 ^ n4065 ^ 1'b0 ;
  assign n27727 = ~n2625 & n27726 ;
  assign n27728 = ( ~n10538 & n13536 ) | ( ~n10538 & n27727 ) | ( n13536 & n27727 ) ;
  assign n27729 = n27728 ^ n8959 ^ 1'b0 ;
  assign n27730 = ~n21119 & n27729 ;
  assign n27733 = n24340 ^ n21559 ^ n17909 ;
  assign n27731 = n14420 ^ n7552 ^ n4218 ;
  assign n27732 = n12826 & n27731 ;
  assign n27734 = n27733 ^ n27732 ^ 1'b0 ;
  assign n27735 = ( n372 & ~n10258 ) | ( n372 & n22792 ) | ( ~n10258 & n22792 ) ;
  assign n27736 = ~n8815 & n27735 ;
  assign n27737 = n23756 ^ n20172 ^ n6435 ;
  assign n27738 = n27737 ^ n20809 ^ n4047 ;
  assign n27739 = n27738 ^ n14785 ^ n2231 ;
  assign n27740 = ( n8867 & n11183 ) | ( n8867 & ~n14136 ) | ( n11183 & ~n14136 ) ;
  assign n27741 = n27740 ^ n16167 ^ n11491 ;
  assign n27742 = n25482 ^ n18429 ^ n14816 ;
  assign n27743 = n27742 ^ n324 ^ x221 ;
  assign n27744 = n3150 | n8308 ;
  assign n27745 = ( n13212 & n16574 ) | ( n13212 & ~n27744 ) | ( n16574 & ~n27744 ) ;
  assign n27746 = n13577 ^ n12538 ^ n8636 ;
  assign n27747 = n4032 & ~n9277 ;
  assign n27748 = n27747 ^ n14652 ^ 1'b0 ;
  assign n27749 = ( n27745 & ~n27746 ) | ( n27745 & n27748 ) | ( ~n27746 & n27748 ) ;
  assign n27750 = n7415 & ~n19615 ;
  assign n27751 = n27750 ^ n2412 ^ 1'b0 ;
  assign n27752 = ( n5471 & ~n12200 ) | ( n5471 & n27751 ) | ( ~n12200 & n27751 ) ;
  assign n27753 = ( ~n15737 & n27749 ) | ( ~n15737 & n27752 ) | ( n27749 & n27752 ) ;
  assign n27754 = ( ~n1266 & n3550 ) | ( ~n1266 & n4381 ) | ( n3550 & n4381 ) ;
  assign n27755 = ( ~n2328 & n6494 ) | ( ~n2328 & n27754 ) | ( n6494 & n27754 ) ;
  assign n27756 = n2600 | n5095 ;
  assign n27757 = n27756 ^ n1710 ^ n1136 ;
  assign n27758 = n27757 ^ n15991 ^ n4443 ;
  assign n27761 = n4992 ^ n4236 ^ n3627 ;
  assign n27759 = ( n1210 & n3771 ) | ( n1210 & ~n4143 ) | ( n3771 & ~n4143 ) ;
  assign n27760 = n27759 ^ n10880 ^ n9462 ;
  assign n27762 = n27761 ^ n27760 ^ n5737 ;
  assign n27766 = ( n16358 & n18118 ) | ( n16358 & ~n18619 ) | ( n18118 & ~n18619 ) ;
  assign n27767 = ( n6251 & n16445 ) | ( n6251 & ~n27766 ) | ( n16445 & ~n27766 ) ;
  assign n27765 = n10096 ^ n7574 ^ n4148 ;
  assign n27763 = n17632 ^ n11015 ^ n5292 ;
  assign n27764 = n27763 ^ n2576 ^ n2342 ;
  assign n27768 = n27767 ^ n27765 ^ n27764 ;
  assign n27769 = n16872 ^ n9960 ^ n8848 ;
  assign n27770 = ( n4025 & n14779 ) | ( n4025 & n27769 ) | ( n14779 & n27769 ) ;
  assign n27771 = n20682 ^ n8668 ^ n5471 ;
  assign n27772 = ( n20419 & ~n27770 ) | ( n20419 & n27771 ) | ( ~n27770 & n27771 ) ;
  assign n27773 = n18448 ^ n6536 ^ n3962 ;
  assign n27774 = n27773 ^ n5452 ^ n4052 ;
  assign n27775 = n27774 ^ n4455 ^ 1'b0 ;
  assign n27776 = n27772 | n27775 ;
  assign n27777 = n13586 ^ n10861 ^ n7501 ;
  assign n27778 = n27777 ^ n10487 ^ 1'b0 ;
  assign n27779 = ( ~n869 & n18070 ) | ( ~n869 & n22523 ) | ( n18070 & n22523 ) ;
  assign n27780 = n24178 ^ n19794 ^ 1'b0 ;
  assign n27781 = ( n5833 & ~n18616 ) | ( n5833 & n20944 ) | ( ~n18616 & n20944 ) ;
  assign n27782 = n3610 | n12451 ;
  assign n27783 = n27782 ^ n4709 ^ 1'b0 ;
  assign n27786 = n23969 ^ n7528 ^ n772 ;
  assign n27784 = ( n3458 & ~n6529 ) | ( n3458 & n17650 ) | ( ~n6529 & n17650 ) ;
  assign n27785 = n27784 ^ n6915 ^ 1'b0 ;
  assign n27787 = n27786 ^ n27785 ^ n8641 ;
  assign n27788 = ( n7457 & n9974 ) | ( n7457 & ~n10170 ) | ( n9974 & ~n10170 ) ;
  assign n27789 = n27788 ^ n9495 ^ n2121 ;
  assign n27790 = n27789 ^ n27687 ^ n17620 ;
  assign n27791 = x176 & n718 ;
  assign n27792 = n16808 ^ n6337 ^ n4844 ;
  assign n27793 = n25666 ^ n22906 ^ x243 ;
  assign n27794 = n23865 ^ n12919 ^ n5755 ;
  assign n27795 = n3735 & ~n23795 ;
  assign n27796 = ( n27137 & n27794 ) | ( n27137 & ~n27795 ) | ( n27794 & ~n27795 ) ;
  assign n27802 = ( n7608 & ~n14960 ) | ( n7608 & n19781 ) | ( ~n14960 & n19781 ) ;
  assign n27803 = ( n1194 & n6912 ) | ( n1194 & n27802 ) | ( n6912 & n27802 ) ;
  assign n27797 = n4284 ^ n2543 ^ n1314 ;
  assign n27798 = n27797 ^ n19470 ^ n12980 ;
  assign n27799 = ( n8403 & n24155 ) | ( n8403 & n25481 ) | ( n24155 & n25481 ) ;
  assign n27800 = ~n7160 & n27799 ;
  assign n27801 = ( n4656 & n27798 ) | ( n4656 & n27800 ) | ( n27798 & n27800 ) ;
  assign n27804 = n27803 ^ n27801 ^ n11299 ;
  assign n27805 = n10323 ^ n8701 ^ n6685 ;
  assign n27809 = n11358 ^ n9661 ^ n2163 ;
  assign n27807 = n8196 ^ n7889 ^ n421 ;
  assign n27808 = n27807 ^ n7936 ^ n835 ;
  assign n27810 = n27809 ^ n27808 ^ n9501 ;
  assign n27806 = ( ~n9473 & n22117 ) | ( ~n9473 & n25733 ) | ( n22117 & n25733 ) ;
  assign n27811 = n27810 ^ n27806 ^ n878 ;
  assign n27812 = ( n2943 & n24047 ) | ( n2943 & ~n27811 ) | ( n24047 & ~n27811 ) ;
  assign n27813 = ( ~n13352 & n27805 ) | ( ~n13352 & n27812 ) | ( n27805 & n27812 ) ;
  assign n27814 = ( n1697 & n18473 ) | ( n1697 & ~n24649 ) | ( n18473 & ~n24649 ) ;
  assign n27817 = n14743 ^ n12418 ^ n2172 ;
  assign n27815 = ( n8162 & ~n16998 ) | ( n8162 & n23360 ) | ( ~n16998 & n23360 ) ;
  assign n27816 = n27815 ^ n27558 ^ n3522 ;
  assign n27818 = n27817 ^ n27816 ^ n2088 ;
  assign n27819 = n26339 ^ n19761 ^ n7367 ;
  assign n27820 = ( n27814 & ~n27818 ) | ( n27814 & n27819 ) | ( ~n27818 & n27819 ) ;
  assign n27821 = ( x20 & n8480 ) | ( x20 & ~n20778 ) | ( n8480 & ~n20778 ) ;
  assign n27824 = ( n3412 & ~n15791 ) | ( n3412 & n22090 ) | ( ~n15791 & n22090 ) ;
  assign n27825 = ( n4113 & ~n5321 ) | ( n4113 & n27824 ) | ( ~n5321 & n27824 ) ;
  assign n27822 = n8946 ^ n1312 ^ 1'b0 ;
  assign n27823 = n17072 & ~n27822 ;
  assign n27826 = n27825 ^ n27823 ^ n14594 ;
  assign n27829 = ~n2001 & n2586 ;
  assign n27830 = ~n4545 & n27829 ;
  assign n27827 = n3433 & n9053 ;
  assign n27828 = n27827 ^ n18460 ^ n14887 ;
  assign n27831 = n27830 ^ n27828 ^ n2502 ;
  assign n27832 = ~n3167 & n22125 ;
  assign n27833 = ( n1994 & n10484 ) | ( n1994 & ~n23250 ) | ( n10484 & ~n23250 ) ;
  assign n27834 = ( n2815 & ~n14053 ) | ( n2815 & n27833 ) | ( ~n14053 & n27833 ) ;
  assign n27835 = n11889 ^ n10237 ^ n6987 ;
  assign n27836 = ~n7921 & n27193 ;
  assign n27837 = ~n5541 & n27836 ;
  assign n27838 = n23713 ^ n21408 ^ n5265 ;
  assign n27839 = ( ~n9437 & n13316 ) | ( ~n9437 & n27838 ) | ( n13316 & n27838 ) ;
  assign n27840 = ( n8184 & ~n23388 ) | ( n8184 & n25415 ) | ( ~n23388 & n25415 ) ;
  assign n27841 = n8162 & n11180 ;
  assign n27842 = n27841 ^ n23286 ^ n3692 ;
  assign n27843 = n27842 ^ n6335 ^ n4625 ;
  assign n27844 = ( n5347 & n19702 ) | ( n5347 & ~n27843 ) | ( n19702 & ~n27843 ) ;
  assign n27850 = n9587 ^ n5669 ^ n661 ;
  assign n27845 = n17145 ^ n11988 ^ 1'b0 ;
  assign n27846 = n5087 & ~n27845 ;
  assign n27847 = ( ~n14440 & n17865 ) | ( ~n14440 & n27846 ) | ( n17865 & n27846 ) ;
  assign n27848 = ~n5262 & n27847 ;
  assign n27849 = n27848 ^ n12571 ^ n2822 ;
  assign n27851 = n27850 ^ n27849 ^ n20474 ;
  assign n27852 = ~n12238 & n20329 ;
  assign n27853 = n27852 ^ n13592 ^ n2255 ;
  assign n27854 = n27853 ^ n12348 ^ n3948 ;
  assign n27855 = n27854 ^ n13308 ^ n5301 ;
  assign n27856 = ( n3959 & n7358 ) | ( n3959 & n12138 ) | ( n7358 & n12138 ) ;
  assign n27862 = ( ~n1794 & n7574 ) | ( ~n1794 & n14976 ) | ( n7574 & n14976 ) ;
  assign n27863 = n27862 ^ n17030 ^ n6922 ;
  assign n27860 = ( n3320 & n12356 ) | ( n3320 & ~n18673 ) | ( n12356 & ~n18673 ) ;
  assign n27858 = n14449 ^ n11605 ^ n8421 ;
  assign n27857 = n15147 ^ n13738 ^ 1'b0 ;
  assign n27859 = n27858 ^ n27857 ^ n4500 ;
  assign n27861 = n27860 ^ n27859 ^ n648 ;
  assign n27864 = n27863 ^ n27861 ^ n27599 ;
  assign n27865 = ( n3423 & n6514 ) | ( n3423 & n7520 ) | ( n6514 & n7520 ) ;
  assign n27866 = n27865 ^ n24713 ^ 1'b0 ;
  assign n27867 = ( n2203 & n11089 ) | ( n2203 & ~n17611 ) | ( n11089 & ~n17611 ) ;
  assign n27868 = n27867 ^ n17551 ^ n8438 ;
  assign n27869 = ( ~n16574 & n23955 ) | ( ~n16574 & n27868 ) | ( n23955 & n27868 ) ;
  assign n27870 = n937 & n4844 ;
  assign n27871 = n27870 ^ n17415 ^ 1'b0 ;
  assign n27872 = n13882 & ~n27871 ;
  assign n27873 = n27872 ^ n12927 ^ 1'b0 ;
  assign n27874 = n27873 ^ n25947 ^ n9343 ;
  assign n27875 = n4213 & n7779 ;
  assign n27876 = ~n1489 & n27875 ;
  assign n27877 = n27876 ^ n23953 ^ 1'b0 ;
  assign n27878 = ( n3442 & n21404 ) | ( n3442 & ~n23458 ) | ( n21404 & ~n23458 ) ;
  assign n27879 = ( n10827 & ~n18535 ) | ( n10827 & n27878 ) | ( ~n18535 & n27878 ) ;
  assign n27882 = ( n14545 & n14586 ) | ( n14545 & n17727 ) | ( n14586 & n17727 ) ;
  assign n27880 = n19626 ^ n9357 ^ n3584 ;
  assign n27881 = n27880 ^ n21009 ^ n4973 ;
  assign n27883 = n27882 ^ n27881 ^ n8279 ;
  assign n27884 = ( n2521 & n11406 ) | ( n2521 & ~n13595 ) | ( n11406 & ~n13595 ) ;
  assign n27885 = ( n6114 & n8157 ) | ( n6114 & ~n25037 ) | ( n8157 & ~n25037 ) ;
  assign n27886 = n26966 | n27885 ;
  assign n27887 = n27886 ^ n6782 ^ 1'b0 ;
  assign n27888 = n19175 ^ n3254 ^ n1610 ;
  assign n27889 = n27888 ^ n21256 ^ n262 ;
  assign n27890 = n20026 ^ n3724 ^ n1432 ;
  assign n27891 = ( ~n10792 & n20031 ) | ( ~n10792 & n27890 ) | ( n20031 & n27890 ) ;
  assign n27892 = ( n11517 & ~n19689 ) | ( n11517 & n27891 ) | ( ~n19689 & n27891 ) ;
  assign n27893 = n27892 ^ n15103 ^ n1178 ;
  assign n27894 = ( n6654 & ~n18612 ) | ( n6654 & n26882 ) | ( ~n18612 & n26882 ) ;
  assign n27895 = n22463 ^ n9254 ^ n9116 ;
  assign n27896 = ( n4371 & n27894 ) | ( n4371 & n27895 ) | ( n27894 & n27895 ) ;
  assign n27897 = n6769 & n7453 ;
  assign n27898 = n27897 ^ n3983 ^ 1'b0 ;
  assign n27899 = n27896 | n27898 ;
  assign n27900 = n18960 ^ n18260 ^ 1'b0 ;
  assign n27901 = n27900 ^ n23604 ^ n8626 ;
  assign n27902 = n18253 ^ n16640 ^ n3538 ;
  assign n27903 = ( n4073 & ~n27901 ) | ( n4073 & n27902 ) | ( ~n27901 & n27902 ) ;
  assign n27904 = n13553 ^ n10345 ^ n784 ;
  assign n27905 = n27904 ^ n17280 ^ n3237 ;
  assign n27906 = n27905 ^ n25191 ^ n18518 ;
  assign n27907 = n22800 ^ n21243 ^ n12154 ;
  assign n27908 = n3278 ^ n2119 ^ 1'b0 ;
  assign n27909 = ~n27907 & n27908 ;
  assign n27910 = ( ~n4776 & n26677 ) | ( ~n4776 & n27909 ) | ( n26677 & n27909 ) ;
  assign n27911 = n12881 ^ n12115 ^ n11029 ;
  assign n27913 = ( n1230 & n3234 ) | ( n1230 & ~n9566 ) | ( n3234 & ~n9566 ) ;
  assign n27912 = ( n9081 & n20847 ) | ( n9081 & n27192 ) | ( n20847 & n27192 ) ;
  assign n27914 = n27913 ^ n27912 ^ n2809 ;
  assign n27915 = n23187 ^ n8663 ^ n5536 ;
  assign n27916 = ( n2011 & ~n7884 ) | ( n2011 & n8881 ) | ( ~n7884 & n8881 ) ;
  assign n27917 = ( n14695 & n23691 ) | ( n14695 & ~n27916 ) | ( n23691 & ~n27916 ) ;
  assign n27918 = ( n27914 & ~n27915 ) | ( n27914 & n27917 ) | ( ~n27915 & n27917 ) ;
  assign n27919 = ( ~n19005 & n27911 ) | ( ~n19005 & n27918 ) | ( n27911 & n27918 ) ;
  assign n27924 = ( n7692 & ~n14839 ) | ( n7692 & n18448 ) | ( ~n14839 & n18448 ) ;
  assign n27920 = n3057 & ~n6691 ;
  assign n27921 = ~n4554 & n27920 ;
  assign n27922 = n27921 ^ n20577 ^ n972 ;
  assign n27923 = ( n18375 & n21082 ) | ( n18375 & n27922 ) | ( n21082 & n27922 ) ;
  assign n27925 = n27924 ^ n27923 ^ n1892 ;
  assign n27926 = n14187 ^ n11239 ^ n10013 ;
  assign n27927 = ( n2782 & ~n8466 ) | ( n2782 & n11716 ) | ( ~n8466 & n11716 ) ;
  assign n27928 = n27927 ^ n19762 ^ 1'b0 ;
  assign n27929 = n27928 ^ n22867 ^ n21200 ;
  assign n27930 = n12584 ^ n5702 ^ n3833 ;
  assign n27932 = n3107 ^ n1595 ^ n556 ;
  assign n27931 = ( n14919 & n17002 ) | ( n14919 & ~n23807 ) | ( n17002 & ~n23807 ) ;
  assign n27933 = n27932 ^ n27931 ^ 1'b0 ;
  assign n27934 = n24211 | n27933 ;
  assign n27935 = n3842 & ~n27934 ;
  assign n27936 = n27930 & n27935 ;
  assign n27943 = n8157 ^ n726 ^ n600 ;
  assign n27942 = n27612 ^ n11349 ^ n8572 ;
  assign n27944 = n27943 ^ n27942 ^ n13638 ;
  assign n27940 = ( ~n4952 & n20935 ) | ( ~n4952 & n21267 ) | ( n20935 & n21267 ) ;
  assign n27938 = n22196 ^ n11871 ^ n1828 ;
  assign n27939 = ( n1917 & n8804 ) | ( n1917 & n27938 ) | ( n8804 & n27938 ) ;
  assign n27941 = n27940 ^ n27939 ^ n7147 ;
  assign n27945 = n27944 ^ n27941 ^ n11319 ;
  assign n27937 = n12582 ^ n7818 ^ n4593 ;
  assign n27946 = n27945 ^ n27937 ^ n5639 ;
  assign n27947 = n4623 & n9729 ;
  assign n27948 = n27947 ^ n5554 ^ 1'b0 ;
  assign n27949 = n27948 ^ n5433 ^ n3787 ;
  assign n27950 = n6218 | n14302 ;
  assign n27951 = n27949 | n27950 ;
  assign n27952 = ( n423 & ~n6511 ) | ( n423 & n27951 ) | ( ~n6511 & n27951 ) ;
  assign n27953 = ( ~n19251 & n21096 ) | ( ~n19251 & n27952 ) | ( n21096 & n27952 ) ;
  assign n27954 = n406 | n15518 ;
  assign n27959 = n5414 ^ n3256 ^ n2171 ;
  assign n27960 = n10956 ^ n10886 ^ n4862 ;
  assign n27961 = n27960 ^ n13010 ^ n4248 ;
  assign n27962 = ( n3770 & ~n14466 ) | ( n3770 & n27961 ) | ( ~n14466 & n27961 ) ;
  assign n27963 = ( n4774 & n27959 ) | ( n4774 & n27962 ) | ( n27959 & n27962 ) ;
  assign n27955 = n20628 ^ n17693 ^ n14853 ;
  assign n27956 = n15357 | n27955 ;
  assign n27957 = n27956 ^ n10711 ^ 1'b0 ;
  assign n27958 = ~n6020 & n27957 ;
  assign n27964 = n27963 ^ n27958 ^ 1'b0 ;
  assign n27965 = n6519 | n14738 ;
  assign n27966 = n1307 & ~n27965 ;
  assign n27967 = n17223 ^ n13337 ^ n1350 ;
  assign n27968 = ( n7609 & n22395 ) | ( n7609 & n27017 ) | ( n22395 & n27017 ) ;
  assign n27969 = ( ~n7408 & n11081 ) | ( ~n7408 & n13559 ) | ( n11081 & n13559 ) ;
  assign n27970 = n16312 ^ n10264 ^ 1'b0 ;
  assign n27971 = ~n27969 & n27970 ;
  assign n27972 = n27971 ^ n4963 ^ 1'b0 ;
  assign n27973 = n5321 & n27972 ;
  assign n27974 = n22151 ^ n10144 ^ n7912 ;
  assign n27975 = n27974 ^ n6354 ^ n1881 ;
  assign n27976 = ( ~n7816 & n9968 ) | ( ~n7816 & n17055 ) | ( n9968 & n17055 ) ;
  assign n27977 = n27976 ^ n20903 ^ n16447 ;
  assign n27978 = ( n656 & ~n27975 ) | ( n656 & n27977 ) | ( ~n27975 & n27977 ) ;
  assign n27979 = ( n21526 & n22268 ) | ( n21526 & ~n27370 ) | ( n22268 & ~n27370 ) ;
  assign n27980 = n14614 ^ n4757 ^ n3596 ;
  assign n27981 = n27907 ^ n15058 ^ n4791 ;
  assign n27982 = ~n5929 & n18261 ;
  assign n27983 = ( n3283 & n27981 ) | ( n3283 & ~n27982 ) | ( n27981 & ~n27982 ) ;
  assign n27984 = ( n14694 & n23251 ) | ( n14694 & n27983 ) | ( n23251 & n27983 ) ;
  assign n27985 = ( n26794 & n27980 ) | ( n26794 & ~n27984 ) | ( n27980 & ~n27984 ) ;
  assign n27986 = ( ~n1748 & n17145 ) | ( ~n1748 & n27985 ) | ( n17145 & n27985 ) ;
  assign n27987 = ( ~n1653 & n6975 ) | ( ~n1653 & n15184 ) | ( n6975 & n15184 ) ;
  assign n27988 = ( ~n14717 & n20627 ) | ( ~n14717 & n27987 ) | ( n20627 & n27987 ) ;
  assign n27989 = ( ~n4542 & n11637 ) | ( ~n4542 & n27988 ) | ( n11637 & n27988 ) ;
  assign n27990 = ( x48 & ~n2014 ) | ( x48 & n5154 ) | ( ~n2014 & n5154 ) ;
  assign n27991 = ( ~n3933 & n15019 ) | ( ~n3933 & n27990 ) | ( n15019 & n27990 ) ;
  assign n27992 = ( n5743 & n11234 ) | ( n5743 & ~n27991 ) | ( n11234 & ~n27991 ) ;
  assign n27993 = n27992 ^ n24685 ^ n3620 ;
  assign n27994 = n9024 ^ n8018 ^ n1905 ;
  assign n27995 = n27522 ^ n10242 ^ n974 ;
  assign n27996 = n7018 ^ n2152 ^ 1'b0 ;
  assign n27997 = n15383 & n27996 ;
  assign n27998 = ( ~n23942 & n27995 ) | ( ~n23942 & n27997 ) | ( n27995 & n27997 ) ;
  assign n27999 = n7199 ^ n3997 ^ n836 ;
  assign n28000 = ( n7240 & ~n27636 ) | ( n7240 & n27999 ) | ( ~n27636 & n27999 ) ;
  assign n28001 = n28000 ^ n12366 ^ n11368 ;
  assign n28002 = n14233 ^ n9898 ^ n8818 ;
  assign n28003 = ( ~n3737 & n7554 ) | ( ~n3737 & n28002 ) | ( n7554 & n28002 ) ;
  assign n28004 = n28003 ^ n27090 ^ n5947 ;
  assign n28005 = ( n3732 & n24976 ) | ( n3732 & ~n28004 ) | ( n24976 & ~n28004 ) ;
  assign n28006 = ( ~n5132 & n6017 ) | ( ~n5132 & n10411 ) | ( n6017 & n10411 ) ;
  assign n28007 = n11404 & n12766 ;
  assign n28008 = ( n6319 & n9291 ) | ( n6319 & n28007 ) | ( n9291 & n28007 ) ;
  assign n28009 = ( n15239 & n28006 ) | ( n15239 & ~n28008 ) | ( n28006 & ~n28008 ) ;
  assign n28010 = n2756 | n10340 ;
  assign n28011 = n28010 ^ n10635 ^ 1'b0 ;
  assign n28012 = ~n1864 & n24699 ;
  assign n28013 = n28012 ^ n15173 ^ 1'b0 ;
  assign n28014 = n28013 ^ n13061 ^ 1'b0 ;
  assign n28015 = ~n28011 & n28014 ;
  assign n28017 = n4807 ^ n2226 ^ 1'b0 ;
  assign n28016 = ( n4318 & n8311 ) | ( n4318 & ~n9219 ) | ( n8311 & ~n9219 ) ;
  assign n28018 = n28017 ^ n28016 ^ n19981 ;
  assign n28019 = n28018 ^ n24163 ^ n15170 ;
  assign n28020 = n16995 ^ n1546 ^ 1'b0 ;
  assign n28021 = n260 & ~n28020 ;
  assign n28022 = ( ~n2639 & n7113 ) | ( ~n2639 & n8946 ) | ( n7113 & n8946 ) ;
  assign n28023 = n28022 ^ n14561 ^ n7546 ;
  assign n28024 = ( ~n9066 & n22002 ) | ( ~n9066 & n28023 ) | ( n22002 & n28023 ) ;
  assign n28025 = ( ~n14685 & n28021 ) | ( ~n14685 & n28024 ) | ( n28021 & n28024 ) ;
  assign n28026 = ( n8293 & n10161 ) | ( n8293 & n28025 ) | ( n10161 & n28025 ) ;
  assign n28027 = n23051 ^ n12280 ^ 1'b0 ;
  assign n28028 = ~n28026 & n28027 ;
  assign n28029 = ( ~n931 & n1211 ) | ( ~n931 & n6370 ) | ( n1211 & n6370 ) ;
  assign n28030 = ( n7858 & ~n10475 ) | ( n7858 & n28029 ) | ( ~n10475 & n28029 ) ;
  assign n28031 = ( n507 & n4160 ) | ( n507 & n28030 ) | ( n4160 & n28030 ) ;
  assign n28032 = n9632 ^ n3168 ^ 1'b0 ;
  assign n28033 = ( n3726 & n10246 ) | ( n3726 & ~n28032 ) | ( n10246 & ~n28032 ) ;
  assign n28034 = ( n588 & n7154 ) | ( n588 & ~n28033 ) | ( n7154 & ~n28033 ) ;
  assign n28035 = ( ~n10085 & n28031 ) | ( ~n10085 & n28034 ) | ( n28031 & n28034 ) ;
  assign n28036 = ( n1907 & ~n9508 ) | ( n1907 & n11945 ) | ( ~n9508 & n11945 ) ;
  assign n28037 = ( n5200 & n5280 ) | ( n5200 & n28036 ) | ( n5280 & n28036 ) ;
  assign n28038 = n28037 ^ n2298 ^ n1249 ;
  assign n28041 = n3117 | n7103 ;
  assign n28042 = n28041 ^ n1833 ^ 1'b0 ;
  assign n28039 = ( ~n5762 & n18199 ) | ( ~n5762 & n19064 ) | ( n18199 & n19064 ) ;
  assign n28040 = n28039 ^ n25087 ^ n23482 ;
  assign n28043 = n28042 ^ n28040 ^ n9862 ;
  assign n28044 = ( n5095 & ~n18764 ) | ( n5095 & n22234 ) | ( ~n18764 & n22234 ) ;
  assign n28045 = ( ~n28038 & n28043 ) | ( ~n28038 & n28044 ) | ( n28043 & n28044 ) ;
  assign n28046 = n8976 ^ n6215 ^ n1806 ;
  assign n28047 = ( n4342 & n6489 ) | ( n4342 & n25097 ) | ( n6489 & n25097 ) ;
  assign n28048 = n3463 & ~n9492 ;
  assign n28049 = n21404 ^ n10660 ^ n2623 ;
  assign n28050 = ( ~n7867 & n28048 ) | ( ~n7867 & n28049 ) | ( n28048 & n28049 ) ;
  assign n28051 = n21411 ^ n8891 ^ 1'b0 ;
  assign n28052 = ( n3308 & n11822 ) | ( n3308 & n28051 ) | ( n11822 & n28051 ) ;
  assign n28053 = n16251 | n28052 ;
  assign n28054 = n28053 ^ n22095 ^ 1'b0 ;
  assign n28055 = ( n8254 & n17163 ) | ( n8254 & ~n18429 ) | ( n17163 & ~n18429 ) ;
  assign n28056 = n28055 ^ n785 ^ 1'b0 ;
  assign n28057 = ( n2036 & n5001 ) | ( n2036 & ~n14706 ) | ( n5001 & ~n14706 ) ;
  assign n28058 = ( ~n21096 & n21740 ) | ( ~n21096 & n28057 ) | ( n21740 & n28057 ) ;
  assign n28059 = ( ~n10293 & n10679 ) | ( ~n10293 & n14234 ) | ( n10679 & n14234 ) ;
  assign n28060 = n24958 ^ n22056 ^ n20888 ;
  assign n28061 = n26349 ^ n13937 ^ n9937 ;
  assign n28062 = ( n10629 & n10831 ) | ( n10629 & ~n26110 ) | ( n10831 & ~n26110 ) ;
  assign n28063 = n10919 | n28062 ;
  assign n28064 = n28061 & ~n28063 ;
  assign n28069 = ( ~n4173 & n24078 ) | ( ~n4173 & n25372 ) | ( n24078 & n25372 ) ;
  assign n28065 = ~n8145 & n10852 ;
  assign n28066 = ~n7784 & n28065 ;
  assign n28067 = n28066 ^ n16379 ^ n10167 ;
  assign n28068 = n13671 & n28067 ;
  assign n28070 = n28069 ^ n28068 ^ 1'b0 ;
  assign n28071 = n24666 ^ n14367 ^ n1393 ;
  assign n28074 = ( n4477 & n18586 ) | ( n4477 & n25101 ) | ( n18586 & n25101 ) ;
  assign n28072 = ( ~n2028 & n2720 ) | ( ~n2028 & n26185 ) | ( n2720 & n26185 ) ;
  assign n28073 = n1219 & ~n28072 ;
  assign n28075 = n28074 ^ n28073 ^ n7097 ;
  assign n28076 = ( n451 & n4199 ) | ( n451 & ~n23394 ) | ( n4199 & ~n23394 ) ;
  assign n28077 = ( n2168 & n7534 ) | ( n2168 & n28076 ) | ( n7534 & n28076 ) ;
  assign n28078 = ( n7673 & n14060 ) | ( n7673 & n28077 ) | ( n14060 & n28077 ) ;
  assign n28079 = n28078 ^ n15863 ^ n10608 ;
  assign n28080 = n13304 ^ n6344 ^ 1'b0 ;
  assign n28081 = n7737 ^ n2677 ^ 1'b0 ;
  assign n28082 = n28081 ^ n16714 ^ n6427 ;
  assign n28083 = ( n16110 & n24406 ) | ( n16110 & ~n28082 ) | ( n24406 & ~n28082 ) ;
  assign n28084 = n17930 ^ n17652 ^ n7861 ;
  assign n28085 = n28084 ^ n27175 ^ n9918 ;
  assign n28086 = n28085 ^ n13466 ^ n5689 ;
  assign n28087 = ( ~n1382 & n28083 ) | ( ~n1382 & n28086 ) | ( n28083 & n28086 ) ;
  assign n28088 = n28080 & ~n28087 ;
  assign n28089 = n28088 ^ n11038 ^ 1'b0 ;
  assign n28097 = n3202 ^ n1716 ^ 1'b0 ;
  assign n28098 = n28097 ^ n20070 ^ n10357 ;
  assign n28090 = n16288 ^ n2082 ^ n1458 ;
  assign n28091 = ( n9110 & ~n14901 ) | ( n9110 & n28090 ) | ( ~n14901 & n28090 ) ;
  assign n28092 = n28091 ^ n6076 ^ 1'b0 ;
  assign n28093 = ~n4094 & n28092 ;
  assign n28094 = ( n990 & n10021 ) | ( n990 & ~n28093 ) | ( n10021 & ~n28093 ) ;
  assign n28095 = ~n11574 & n28094 ;
  assign n28096 = n6639 & n28095 ;
  assign n28099 = n28098 ^ n28096 ^ n21839 ;
  assign n28100 = n19309 ^ n6216 ^ n2494 ;
  assign n28101 = n22511 ^ n21656 ^ n5414 ;
  assign n28103 = ( n1339 & n12738 ) | ( n1339 & n14285 ) | ( n12738 & n14285 ) ;
  assign n28102 = ( n1188 & n8235 ) | ( n1188 & n20707 ) | ( n8235 & n20707 ) ;
  assign n28104 = n28103 ^ n28102 ^ n19682 ;
  assign n28105 = n28104 ^ n19139 ^ n6706 ;
  assign n28106 = n8400 ^ n8369 ^ 1'b0 ;
  assign n28107 = ( n6317 & n15864 ) | ( n6317 & n28106 ) | ( n15864 & n28106 ) ;
  assign n28108 = n28107 ^ n18541 ^ 1'b0 ;
  assign n28109 = ( n7272 & n8914 ) | ( n7272 & n16084 ) | ( n8914 & n16084 ) ;
  assign n28110 = n24511 ^ n11228 ^ n6675 ;
  assign n28111 = n15490 ^ n6515 ^ n2160 ;
  assign n28112 = n28111 ^ n16308 ^ n14728 ;
  assign n28113 = n28112 ^ n24514 ^ n14849 ;
  assign n28114 = n20047 ^ n18224 ^ n10359 ;
  assign n28115 = n14180 ^ n13923 ^ n7203 ;
  assign n28116 = ( n9519 & n10650 ) | ( n9519 & n28115 ) | ( n10650 & n28115 ) ;
  assign n28117 = ( n5808 & n13469 ) | ( n5808 & n19946 ) | ( n13469 & n19946 ) ;
  assign n28118 = ( ~n3007 & n13785 ) | ( ~n3007 & n28117 ) | ( n13785 & n28117 ) ;
  assign n28119 = n19211 | n28118 ;
  assign n28120 = n28119 ^ n20605 ^ 1'b0 ;
  assign n28121 = ( n19858 & n28116 ) | ( n19858 & ~n28120 ) | ( n28116 & ~n28120 ) ;
  assign n28122 = n28121 ^ n4742 ^ x243 ;
  assign n28123 = n7583 & n10994 ;
  assign n28124 = ( n4471 & ~n9010 ) | ( n4471 & n15399 ) | ( ~n9010 & n15399 ) ;
  assign n28125 = n4123 & n22066 ;
  assign n28126 = n28125 ^ n1489 ^ 1'b0 ;
  assign n28127 = n28126 ^ n26525 ^ n25631 ;
  assign n28128 = ( ~n12546 & n28124 ) | ( ~n12546 & n28127 ) | ( n28124 & n28127 ) ;
  assign n28129 = n22981 ^ n12008 ^ n3023 ;
  assign n28130 = ( ~n1022 & n1167 ) | ( ~n1022 & n22104 ) | ( n1167 & n22104 ) ;
  assign n28131 = n10840 ^ n3870 ^ n3744 ;
  assign n28132 = ( n2986 & n4985 ) | ( n2986 & n28131 ) | ( n4985 & n28131 ) ;
  assign n28133 = n14566 | n24423 ;
  assign n28134 = n28133 ^ n23495 ^ n15551 ;
  assign n28135 = ( n1866 & n18410 ) | ( n1866 & n28134 ) | ( n18410 & n28134 ) ;
  assign n28147 = n9277 ^ n4286 ^ 1'b0 ;
  assign n28146 = n22797 ^ n12927 ^ n11332 ;
  assign n28148 = n28147 ^ n28146 ^ n13322 ;
  assign n28142 = n3507 & ~n18534 ;
  assign n28143 = n28142 ^ n13215 ^ 1'b0 ;
  assign n28144 = n28143 ^ n25243 ^ n1290 ;
  assign n28145 = n28144 ^ n3690 ^ n1350 ;
  assign n28136 = n8378 ^ n8259 ^ 1'b0 ;
  assign n28137 = n15549 ^ n14558 ^ n7969 ;
  assign n28138 = n28136 | n28137 ;
  assign n28139 = n28138 ^ n24270 ^ 1'b0 ;
  assign n28140 = ( n4717 & ~n8440 ) | ( n4717 & n15724 ) | ( ~n8440 & n15724 ) ;
  assign n28141 = ( n22741 & n28139 ) | ( n22741 & n28140 ) | ( n28139 & n28140 ) ;
  assign n28149 = n28148 ^ n28145 ^ n28141 ;
  assign n28150 = n20735 ^ n13556 ^ n728 ;
  assign n28151 = ( x18 & n6192 ) | ( x18 & n14513 ) | ( n6192 & n14513 ) ;
  assign n28152 = n6502 & ~n28151 ;
  assign n28153 = n28152 ^ n1499 ^ 1'b0 ;
  assign n28154 = n13702 ^ n12079 ^ n1246 ;
  assign n28155 = ( ~n6249 & n6901 ) | ( ~n6249 & n26284 ) | ( n6901 & n26284 ) ;
  assign n28156 = n28155 ^ n9488 ^ 1'b0 ;
  assign n28157 = n8160 ^ n6748 ^ n2047 ;
  assign n28158 = ( n10258 & n20960 ) | ( n10258 & n28157 ) | ( n20960 & n28157 ) ;
  assign n28159 = ( n11013 & ~n28156 ) | ( n11013 & n28158 ) | ( ~n28156 & n28158 ) ;
  assign n28160 = ( n3656 & ~n5426 ) | ( n3656 & n5463 ) | ( ~n5426 & n5463 ) ;
  assign n28161 = ( n1212 & ~n3168 ) | ( n1212 & n28160 ) | ( ~n3168 & n28160 ) ;
  assign n28162 = ( n16237 & n20095 ) | ( n16237 & n28161 ) | ( n20095 & n28161 ) ;
  assign n28163 = n28162 ^ n17862 ^ x237 ;
  assign n28164 = ( n1111 & ~n2007 ) | ( n1111 & n26072 ) | ( ~n2007 & n26072 ) ;
  assign n28165 = n16866 & ~n25748 ;
  assign n28166 = n28165 ^ n9754 ^ 1'b0 ;
  assign n28168 = ( ~x239 & n12421 ) | ( ~x239 & n23209 ) | ( n12421 & n23209 ) ;
  assign n28167 = ( n7357 & ~n11115 ) | ( n7357 & n16019 ) | ( ~n11115 & n16019 ) ;
  assign n28169 = n28168 ^ n28167 ^ n11232 ;
  assign n28170 = ( n16219 & n17708 ) | ( n16219 & ~n26375 ) | ( n17708 & ~n26375 ) ;
  assign n28171 = ( n16659 & n24248 ) | ( n16659 & ~n28170 ) | ( n24248 & ~n28170 ) ;
  assign n28172 = n21804 ^ n19646 ^ n17428 ;
  assign n28173 = n28172 ^ n13424 ^ n4900 ;
  assign n28174 = n6908 ^ n1162 ^ 1'b0 ;
  assign n28175 = n15100 ^ n12356 ^ n9171 ;
  assign n28176 = n28175 ^ n14280 ^ n9358 ;
  assign n28177 = n16890 & ~n28176 ;
  assign n28178 = n28177 ^ n6974 ^ n4419 ;
  assign n28179 = ( n514 & n1121 ) | ( n514 & ~n9412 ) | ( n1121 & ~n9412 ) ;
  assign n28180 = ( n4350 & n15905 ) | ( n4350 & n28179 ) | ( n15905 & n28179 ) ;
  assign n28181 = n28180 ^ n25670 ^ n22218 ;
  assign n28182 = n28181 ^ n9752 ^ n468 ;
  assign n28186 = n13162 ^ n7407 ^ n792 ;
  assign n28187 = ( n5444 & ~n5510 ) | ( n5444 & n28186 ) | ( ~n5510 & n28186 ) ;
  assign n28183 = n6231 ^ n5895 ^ n2408 ;
  assign n28184 = ( ~n8302 & n12264 ) | ( ~n8302 & n28183 ) | ( n12264 & n28183 ) ;
  assign n28185 = n9063 & ~n28184 ;
  assign n28188 = n28187 ^ n28185 ^ 1'b0 ;
  assign n28189 = x153 & n2077 ;
  assign n28190 = ~n13210 & n28189 ;
  assign n28191 = ( n533 & n1514 ) | ( n533 & ~n1863 ) | ( n1514 & ~n1863 ) ;
  assign n28192 = ( ~n8996 & n14100 ) | ( ~n8996 & n28191 ) | ( n14100 & n28191 ) ;
  assign n28193 = ( ~n4476 & n24845 ) | ( ~n4476 & n28192 ) | ( n24845 & n28192 ) ;
  assign n28194 = n28193 ^ n27897 ^ n14340 ;
  assign n28197 = n1213 ^ n885 ^ n784 ;
  assign n28198 = ( ~n6390 & n26292 ) | ( ~n6390 & n28197 ) | ( n26292 & n28197 ) ;
  assign n28195 = ( ~n4252 & n12824 ) | ( ~n4252 & n23212 ) | ( n12824 & n23212 ) ;
  assign n28196 = n19353 & n28195 ;
  assign n28199 = n28198 ^ n28196 ^ 1'b0 ;
  assign n28200 = ~n668 & n3445 ;
  assign n28201 = ( n944 & n22551 ) | ( n944 & n28200 ) | ( n22551 & n28200 ) ;
  assign n28202 = ( n3503 & ~n15072 ) | ( n3503 & n28201 ) | ( ~n15072 & n28201 ) ;
  assign n28203 = n14447 | n28202 ;
  assign n28204 = x207 | n28203 ;
  assign n28205 = n28204 ^ n14148 ^ 1'b0 ;
  assign n28206 = n4736 & n28205 ;
  assign n28207 = n28206 ^ n23231 ^ n3906 ;
  assign n28208 = n22683 ^ n6592 ^ n4056 ;
  assign n28209 = n24418 ^ n13842 ^ n10079 ;
  assign n28210 = ( n1670 & ~n28148 ) | ( n1670 & n28209 ) | ( ~n28148 & n28209 ) ;
  assign n28211 = ( n1024 & n3472 ) | ( n1024 & n5468 ) | ( n3472 & n5468 ) ;
  assign n28212 = ( n1118 & n10811 ) | ( n1118 & n28211 ) | ( n10811 & n28211 ) ;
  assign n28213 = ( n2105 & n24523 ) | ( n2105 & ~n28212 ) | ( n24523 & ~n28212 ) ;
  assign n28214 = n1337 ^ n1038 ^ 1'b0 ;
  assign n28215 = n28213 | n28214 ;
  assign n28216 = n28210 | n28215 ;
  assign n28217 = n28208 | n28216 ;
  assign n28218 = ( ~n623 & n2990 ) | ( ~n623 & n8050 ) | ( n2990 & n8050 ) ;
  assign n28219 = ( n6202 & n7234 ) | ( n6202 & n27075 ) | ( n7234 & n27075 ) ;
  assign n28220 = ( n3261 & n9455 ) | ( n3261 & n19937 ) | ( n9455 & n19937 ) ;
  assign n28221 = ( ~n28218 & n28219 ) | ( ~n28218 & n28220 ) | ( n28219 & n28220 ) ;
  assign n28224 = n2174 & ~n2422 ;
  assign n28225 = ~n1894 & n28224 ;
  assign n28226 = ( n8424 & n9044 ) | ( n8424 & n28225 ) | ( n9044 & n28225 ) ;
  assign n28223 = ( n8578 & ~n9383 ) | ( n8578 & n20745 ) | ( ~n9383 & n20745 ) ;
  assign n28222 = n23652 ^ n992 ^ 1'b0 ;
  assign n28227 = n28226 ^ n28223 ^ n28222 ;
  assign n28228 = n17728 ^ n6315 ^ n3959 ;
  assign n28229 = ( n4465 & n8496 ) | ( n4465 & ~n8687 ) | ( n8496 & ~n8687 ) ;
  assign n28230 = n28229 ^ n7408 ^ 1'b0 ;
  assign n28231 = ( n15754 & n28228 ) | ( n15754 & ~n28230 ) | ( n28228 & ~n28230 ) ;
  assign n28232 = n24498 ^ n16863 ^ n5401 ;
  assign n28233 = ( n18690 & n26843 ) | ( n18690 & n28232 ) | ( n26843 & n28232 ) ;
  assign n28234 = n15678 & ~n28233 ;
  assign n28235 = ( ~n2479 & n6928 ) | ( ~n2479 & n13229 ) | ( n6928 & n13229 ) ;
  assign n28236 = n28235 ^ n12120 ^ n1363 ;
  assign n28237 = n28236 ^ n12343 ^ n11473 ;
  assign n28238 = n17635 ^ n5291 ^ x168 ;
  assign n28239 = n28238 ^ n17586 ^ n11152 ;
  assign n28240 = ( ~n8817 & n11914 ) | ( ~n8817 & n28239 ) | ( n11914 & n28239 ) ;
  assign n28241 = n14030 & n28240 ;
  assign n28242 = ~n8246 & n28241 ;
  assign n28243 = n5456 & n11950 ;
  assign n28244 = n28242 & n28243 ;
  assign n28247 = n14652 ^ n13709 ^ n3682 ;
  assign n28245 = n17697 ^ n13208 ^ 1'b0 ;
  assign n28246 = n28245 ^ n24568 ^ n4387 ;
  assign n28248 = n28247 ^ n28246 ^ n7184 ;
  assign n28249 = n28212 ^ n17098 ^ n7968 ;
  assign n28250 = ( ~n7534 & n9968 ) | ( ~n7534 & n11181 ) | ( n9968 & n11181 ) ;
  assign n28251 = ( ~n9072 & n9148 ) | ( ~n9072 & n28250 ) | ( n9148 & n28250 ) ;
  assign n28252 = ( n3329 & ~n6250 ) | ( n3329 & n28251 ) | ( ~n6250 & n28251 ) ;
  assign n28253 = n22418 ^ n6608 ^ 1'b0 ;
  assign n28255 = n13897 ^ n4236 ^ 1'b0 ;
  assign n28254 = ( n8807 & ~n10309 ) | ( n8807 & n11991 ) | ( ~n10309 & n11991 ) ;
  assign n28256 = n28255 ^ n28254 ^ n9178 ;
  assign n28257 = ( n12781 & ~n26480 ) | ( n12781 & n28256 ) | ( ~n26480 & n28256 ) ;
  assign n28258 = n22263 ^ n11992 ^ n5072 ;
  assign n28259 = n2216 & n28258 ;
  assign n28260 = n28257 & n28259 ;
  assign n28261 = ( n7714 & ~n14350 ) | ( n7714 & n19000 ) | ( ~n14350 & n19000 ) ;
  assign n28262 = n10614 & n28261 ;
  assign n28263 = ~n27927 & n28262 ;
  assign n28264 = n28263 ^ n24517 ^ n17181 ;
  assign n28265 = n28264 ^ n17551 ^ n3347 ;
  assign n28266 = ( n3907 & n9066 ) | ( n3907 & n15937 ) | ( n9066 & n15937 ) ;
  assign n28267 = ( n5278 & n15984 ) | ( n5278 & n28266 ) | ( n15984 & n28266 ) ;
  assign n28268 = n18945 | n28267 ;
  assign n28269 = n23182 ^ n8402 ^ n2694 ;
  assign n28270 = ( n5099 & n23820 ) | ( n5099 & ~n25207 ) | ( n23820 & ~n25207 ) ;
  assign n28271 = ( n11035 & n28269 ) | ( n11035 & ~n28270 ) | ( n28269 & ~n28270 ) ;
  assign n28272 = ( n881 & n12150 ) | ( n881 & n15363 ) | ( n12150 & n15363 ) ;
  assign n28273 = n28272 ^ n4054 ^ n1454 ;
  assign n28274 = n11461 & ~n14733 ;
  assign n28275 = n28273 & n28274 ;
  assign n28276 = ( n1746 & n4033 ) | ( n1746 & ~n25591 ) | ( n4033 & ~n25591 ) ;
  assign n28277 = n14846 ^ n6270 ^ 1'b0 ;
  assign n28278 = n28277 ^ n10169 ^ n1622 ;
  assign n28279 = ( n9176 & ~n27300 ) | ( n9176 & n28278 ) | ( ~n27300 & n28278 ) ;
  assign n28280 = ( n11118 & n20043 ) | ( n11118 & ~n28279 ) | ( n20043 & ~n28279 ) ;
  assign n28281 = n28280 ^ n18745 ^ n13393 ;
  assign n28282 = ( n11431 & n28276 ) | ( n11431 & ~n28281 ) | ( n28276 & ~n28281 ) ;
  assign n28289 = ( n1275 & n1770 ) | ( n1275 & ~n13903 ) | ( n1770 & ~n13903 ) ;
  assign n28290 = ( ~n19246 & n19339 ) | ( ~n19246 & n28289 ) | ( n19339 & n28289 ) ;
  assign n28286 = n6200 & ~n18296 ;
  assign n28285 = n22429 ^ n15295 ^ n1223 ;
  assign n28287 = n28286 ^ n28285 ^ n3789 ;
  assign n28283 = n26446 ^ n22196 ^ n16811 ;
  assign n28284 = ~n21292 & n28283 ;
  assign n28288 = n28287 ^ n28284 ^ n6292 ;
  assign n28291 = n28290 ^ n28288 ^ n8641 ;
  assign n28292 = n12772 ^ n12437 ^ n7350 ;
  assign n28293 = n25502 ^ n17539 ^ n4849 ;
  assign n28294 = n28293 ^ n14647 ^ n12847 ;
  assign n28295 = ( ~n3522 & n11754 ) | ( ~n3522 & n26396 ) | ( n11754 & n26396 ) ;
  assign n28296 = ( n17421 & n22422 ) | ( n17421 & ~n28295 ) | ( n22422 & ~n28295 ) ;
  assign n28299 = ( n5609 & n6183 ) | ( n5609 & n15582 ) | ( n6183 & n15582 ) ;
  assign n28297 = n20206 ^ n7019 ^ n831 ;
  assign n28298 = n28297 ^ n9073 ^ n4321 ;
  assign n28300 = n28299 ^ n28298 ^ n5925 ;
  assign n28301 = n2606 & ~n7430 ;
  assign n28302 = ( n13218 & n14586 ) | ( n13218 & n22418 ) | ( n14586 & n22418 ) ;
  assign n28303 = ( n12527 & n28301 ) | ( n12527 & ~n28302 ) | ( n28301 & ~n28302 ) ;
  assign n28304 = ( ~n10222 & n13309 ) | ( ~n10222 & n17479 ) | ( n13309 & n17479 ) ;
  assign n28305 = ( n1306 & ~n15938 ) | ( n1306 & n28304 ) | ( ~n15938 & n28304 ) ;
  assign n28306 = n26027 ^ n7275 ^ 1'b0 ;
  assign n28307 = n4232 | n28306 ;
  assign n28308 = n746 & n16495 ;
  assign n28309 = n28308 ^ n19184 ^ n7202 ;
  assign n28310 = ~n5128 & n16447 ;
  assign n28311 = ( n1289 & n6898 ) | ( n1289 & ~n13700 ) | ( n6898 & ~n13700 ) ;
  assign n28313 = ~n1853 & n3458 ;
  assign n28314 = n25161 & n28313 ;
  assign n28315 = n28314 ^ n21610 ^ n13910 ;
  assign n28312 = n4674 & n27218 ;
  assign n28316 = n28315 ^ n28312 ^ 1'b0 ;
  assign n28317 = n13479 ^ n11688 ^ n3628 ;
  assign n28318 = n17307 ^ n13816 ^ n11672 ;
  assign n28319 = n26297 & ~n28318 ;
  assign n28320 = ( n3462 & n5715 ) | ( n3462 & ~n27346 ) | ( n5715 & ~n27346 ) ;
  assign n28321 = ( ~n9889 & n16116 ) | ( ~n9889 & n17150 ) | ( n16116 & n17150 ) ;
  assign n28322 = n27752 ^ n17037 ^ n6243 ;
  assign n28323 = ( n3618 & ~n18118 ) | ( n3618 & n22980 ) | ( ~n18118 & n22980 ) ;
  assign n28324 = n28323 ^ n1914 ^ 1'b0 ;
  assign n28325 = n23310 | n28324 ;
  assign n28326 = n16222 ^ n11538 ^ n5262 ;
  assign n28327 = ( ~n4560 & n18965 ) | ( ~n4560 & n28326 ) | ( n18965 & n28326 ) ;
  assign n28330 = n19640 ^ n11968 ^ 1'b0 ;
  assign n28331 = ~n3780 & n28330 ;
  assign n28328 = ( n2064 & n4794 ) | ( n2064 & n12859 ) | ( n4794 & n12859 ) ;
  assign n28329 = n28328 ^ n18326 ^ n6526 ;
  assign n28332 = n28331 ^ n28329 ^ n12285 ;
  assign n28333 = ( n4557 & n28327 ) | ( n4557 & n28332 ) | ( n28327 & n28332 ) ;
  assign n28334 = n28333 ^ n22973 ^ n2986 ;
  assign n28335 = ( n15048 & n18895 ) | ( n15048 & n19367 ) | ( n18895 & n19367 ) ;
  assign n28336 = ( n5370 & n24058 ) | ( n5370 & n28335 ) | ( n24058 & n28335 ) ;
  assign n28337 = ( ~n1742 & n18112 ) | ( ~n1742 & n24016 ) | ( n18112 & n24016 ) ;
  assign n28341 = ( n4384 & n10119 ) | ( n4384 & ~n26190 ) | ( n10119 & ~n26190 ) ;
  assign n28338 = n13802 ^ n8608 ^ n5621 ;
  assign n28339 = n28338 ^ n26415 ^ n13085 ;
  assign n28340 = n2893 & ~n28339 ;
  assign n28342 = n28341 ^ n28340 ^ 1'b0 ;
  assign n28343 = n8354 ^ n3592 ^ n2000 ;
  assign n28344 = n23016 & n28343 ;
  assign n28345 = n28344 ^ n3643 ^ 1'b0 ;
  assign n28346 = ( n4161 & n4863 ) | ( n4161 & ~n21906 ) | ( n4863 & ~n21906 ) ;
  assign n28347 = n14194 ^ n4148 ^ 1'b0 ;
  assign n28348 = n28347 ^ n22927 ^ n13059 ;
  assign n28349 = ( n4496 & n28346 ) | ( n4496 & n28348 ) | ( n28346 & n28348 ) ;
  assign n28350 = n16514 & ~n28349 ;
  assign n28351 = n28345 & n28350 ;
  assign n28352 = ( n4609 & n16187 ) | ( n4609 & ~n25269 ) | ( n16187 & ~n25269 ) ;
  assign n28353 = ( n2140 & n6548 ) | ( n2140 & ~n10618 ) | ( n6548 & ~n10618 ) ;
  assign n28355 = n21986 ^ n17413 ^ n10526 ;
  assign n28354 = ( n3373 & n5766 ) | ( n3373 & n19911 ) | ( n5766 & n19911 ) ;
  assign n28356 = n28355 ^ n28354 ^ n15321 ;
  assign n28357 = ( n4011 & n11259 ) | ( n4011 & n28356 ) | ( n11259 & n28356 ) ;
  assign n28358 = ( n1476 & ~n1884 ) | ( n1476 & n9877 ) | ( ~n1884 & n9877 ) ;
  assign n28359 = n28358 ^ n20973 ^ n2427 ;
  assign n28360 = ( n1384 & n24273 ) | ( n1384 & ~n27847 ) | ( n24273 & ~n27847 ) ;
  assign n28361 = n28360 ^ n22358 ^ n20473 ;
  assign n28362 = ( n21471 & ~n23479 ) | ( n21471 & n28361 ) | ( ~n23479 & n28361 ) ;
  assign n28363 = n28069 ^ n24698 ^ n10103 ;
  assign n28364 = n10990 ^ n9381 ^ 1'b0 ;
  assign n28365 = n4160 ^ n3560 ^ 1'b0 ;
  assign n28366 = ~n9329 & n28365 ;
  assign n28367 = ( n2156 & n2284 ) | ( n2156 & ~n4535 ) | ( n2284 & ~n4535 ) ;
  assign n28368 = ( n6610 & n8229 ) | ( n6610 & n28367 ) | ( n8229 & n28367 ) ;
  assign n28369 = n28368 ^ n23655 ^ 1'b0 ;
  assign n28370 = n28366 & n28369 ;
  assign n28371 = n28370 ^ n27399 ^ n11255 ;
  assign n28372 = ( n26302 & n28364 ) | ( n26302 & ~n28371 ) | ( n28364 & ~n28371 ) ;
  assign n28377 = n24610 ^ n14913 ^ n905 ;
  assign n28378 = ( n5141 & ~n10454 ) | ( n5141 & n28377 ) | ( ~n10454 & n28377 ) ;
  assign n28376 = ( n1674 & n21568 ) | ( n1674 & ~n23263 ) | ( n21568 & ~n23263 ) ;
  assign n28373 = ( ~n1725 & n4258 ) | ( ~n1725 & n11989 ) | ( n4258 & n11989 ) ;
  assign n28374 = n28373 ^ n6875 ^ n1188 ;
  assign n28375 = ( n6609 & n15871 ) | ( n6609 & ~n28374 ) | ( n15871 & ~n28374 ) ;
  assign n28379 = n28378 ^ n28376 ^ n28375 ;
  assign n28382 = ( n1484 & n2668 ) | ( n1484 & ~n12233 ) | ( n2668 & ~n12233 ) ;
  assign n28380 = ( n4191 & ~n10631 ) | ( n4191 & n12880 ) | ( ~n10631 & n12880 ) ;
  assign n28381 = n19724 & ~n28380 ;
  assign n28383 = n28382 ^ n28381 ^ 1'b0 ;
  assign n28386 = ( n14507 & n15828 ) | ( n14507 & n18376 ) | ( n15828 & n18376 ) ;
  assign n28384 = n11136 ^ n10330 ^ n5164 ;
  assign n28385 = ( n422 & n22146 ) | ( n422 & ~n28384 ) | ( n22146 & ~n28384 ) ;
  assign n28387 = n28386 ^ n28385 ^ n3593 ;
  assign n28388 = n19774 ^ n7541 ^ n3842 ;
  assign n28389 = n2591 & ~n16336 ;
  assign n28390 = ( n1443 & n13222 ) | ( n1443 & n28389 ) | ( n13222 & n28389 ) ;
  assign n28391 = ( n2514 & n4230 ) | ( n2514 & n7324 ) | ( n4230 & n7324 ) ;
  assign n28392 = ( n12858 & n21427 ) | ( n12858 & n28391 ) | ( n21427 & n28391 ) ;
  assign n28393 = n28392 ^ n25357 ^ n3725 ;
  assign n28394 = n23084 ^ n22643 ^ 1'b0 ;
  assign n28395 = ~n16915 & n28394 ;
  assign n28396 = n7962 | n24872 ;
  assign n28397 = n28396 ^ n14495 ^ 1'b0 ;
  assign n28398 = ~n2521 & n28397 ;
  assign n28399 = n28398 ^ n15762 ^ 1'b0 ;
  assign n28401 = n6490 ^ n4398 ^ n1963 ;
  assign n28402 = n28401 ^ n12540 ^ n6251 ;
  assign n28400 = n24454 ^ n10237 ^ n5768 ;
  assign n28403 = n28402 ^ n28400 ^ n24739 ;
  assign n28405 = ( n11114 & ~n15803 ) | ( n11114 & n17282 ) | ( ~n15803 & n17282 ) ;
  assign n28404 = ~n3363 & n16772 ;
  assign n28406 = n28405 ^ n28404 ^ n20522 ;
  assign n28407 = ( ~n6511 & n8172 ) | ( ~n6511 & n12247 ) | ( n8172 & n12247 ) ;
  assign n28408 = ( n3780 & n13844 ) | ( n3780 & ~n27663 ) | ( n13844 & ~n27663 ) ;
  assign n28409 = ( n3491 & n3997 ) | ( n3491 & n28408 ) | ( n3997 & n28408 ) ;
  assign n28410 = ( ~n23017 & n28407 ) | ( ~n23017 & n28409 ) | ( n28407 & n28409 ) ;
  assign n28411 = ( n5811 & n6844 ) | ( n5811 & ~n11577 ) | ( n6844 & ~n11577 ) ;
  assign n28412 = n28411 ^ n28175 ^ n16054 ;
  assign n28413 = n12398 ^ n2189 ^ n854 ;
  assign n28414 = ( ~n4725 & n28412 ) | ( ~n4725 & n28413 ) | ( n28412 & n28413 ) ;
  assign n28415 = n7650 ^ n5539 ^ n1117 ;
  assign n28416 = n2348 & ~n28415 ;
  assign n28417 = n28416 ^ n2698 ^ 1'b0 ;
  assign n28418 = n14675 ^ n7051 ^ n1895 ;
  assign n28419 = n28418 ^ n28037 ^ n13612 ;
  assign n28420 = ( n7674 & n16398 ) | ( n7674 & n23588 ) | ( n16398 & n23588 ) ;
  assign n28421 = ( n18295 & n27912 ) | ( n18295 & ~n28420 ) | ( n27912 & ~n28420 ) ;
  assign n28422 = ( ~n21659 & n28419 ) | ( ~n21659 & n28421 ) | ( n28419 & n28421 ) ;
  assign n28423 = ~n7409 & n8809 ;
  assign n28424 = n27696 ^ n13671 ^ n6628 ;
  assign n28425 = n5872 & ~n9961 ;
  assign n28426 = ( n4654 & ~n28424 ) | ( n4654 & n28425 ) | ( ~n28424 & n28425 ) ;
  assign n28427 = ( n12211 & ~n28423 ) | ( n12211 & n28426 ) | ( ~n28423 & n28426 ) ;
  assign n28428 = n20991 ^ n19618 ^ n4498 ;
  assign n28431 = n26949 ^ n8057 ^ n5729 ;
  assign n28430 = ~n3327 & n3412 ;
  assign n28432 = n28431 ^ n28430 ^ 1'b0 ;
  assign n28429 = n6354 & ~n9270 ;
  assign n28433 = n28432 ^ n28429 ^ 1'b0 ;
  assign n28434 = n28399 ^ n24864 ^ n7776 ;
  assign n28435 = n11146 ^ n1226 ^ n706 ;
  assign n28436 = n28435 ^ n21283 ^ 1'b0 ;
  assign n28437 = n21860 ^ n18492 ^ n8498 ;
  assign n28438 = ~n14796 & n28437 ;
  assign n28439 = ( ~n12616 & n22537 ) | ( ~n12616 & n28438 ) | ( n22537 & n28438 ) ;
  assign n28440 = n28439 ^ n27251 ^ n3734 ;
  assign n28443 = ( n3042 & ~n5261 ) | ( n3042 & n9463 ) | ( ~n5261 & n9463 ) ;
  assign n28444 = ( n8533 & ~n25652 ) | ( n8533 & n28443 ) | ( ~n25652 & n28443 ) ;
  assign n28445 = ( n4615 & ~n18382 ) | ( n4615 & n28444 ) | ( ~n18382 & n28444 ) ;
  assign n28441 = n9187 & ~n14838 ;
  assign n28442 = n28441 ^ n4617 ^ 1'b0 ;
  assign n28446 = n28445 ^ n28442 ^ n1686 ;
  assign n28447 = ( n3924 & ~n3986 ) | ( n3924 & n10227 ) | ( ~n3986 & n10227 ) ;
  assign n28448 = ( n9815 & ~n11267 ) | ( n9815 & n28447 ) | ( ~n11267 & n28447 ) ;
  assign n28449 = ~n1931 & n3608 ;
  assign n28450 = n15006 & n28449 ;
  assign n28451 = n28450 ^ n25199 ^ n10458 ;
  assign n28452 = ( n6085 & ~n28448 ) | ( n6085 & n28451 ) | ( ~n28448 & n28451 ) ;
  assign n28453 = n5402 | n15271 ;
  assign n28454 = ( ~n4214 & n18213 ) | ( ~n4214 & n28453 ) | ( n18213 & n28453 ) ;
  assign n28456 = n11005 ^ n9550 ^ n3047 ;
  assign n28455 = n9232 ^ n1833 ^ n1797 ;
  assign n28457 = n28456 ^ n28455 ^ 1'b0 ;
  assign n28458 = n9406 ^ n3825 ^ 1'b0 ;
  assign n28459 = n28458 ^ n27034 ^ n9420 ;
  assign n28460 = n2302 & ~n5605 ;
  assign n28461 = n28460 ^ n16124 ^ 1'b0 ;
  assign n28462 = ( n1987 & ~n6786 ) | ( n1987 & n28461 ) | ( ~n6786 & n28461 ) ;
  assign n28463 = ( n18575 & ~n27420 ) | ( n18575 & n28462 ) | ( ~n27420 & n28462 ) ;
  assign n28465 = ( n4176 & n5004 ) | ( n4176 & n11314 ) | ( n5004 & n11314 ) ;
  assign n28464 = n19812 ^ n2965 ^ 1'b0 ;
  assign n28466 = n28465 ^ n28464 ^ n18820 ;
  assign n28468 = ( n7423 & ~n9054 ) | ( n7423 & n15486 ) | ( ~n9054 & n15486 ) ;
  assign n28467 = n10144 & n14625 ;
  assign n28469 = n28468 ^ n28467 ^ n2624 ;
  assign n28470 = ( n5796 & ~n16799 ) | ( n5796 & n28469 ) | ( ~n16799 & n28469 ) ;
  assign n28471 = ( n19781 & n28466 ) | ( n19781 & n28470 ) | ( n28466 & n28470 ) ;
  assign n28472 = ( n6858 & ~n9863 ) | ( n6858 & n22535 ) | ( ~n9863 & n22535 ) ;
  assign n28473 = n7405 ^ n3156 ^ n1601 ;
  assign n28474 = ~n10979 & n27117 ;
  assign n28475 = n28473 & n28474 ;
  assign n28476 = ( ~n7577 & n28472 ) | ( ~n7577 & n28475 ) | ( n28472 & n28475 ) ;
  assign n28477 = n22082 ^ n14069 ^ n11221 ;
  assign n28478 = ( n6586 & n28476 ) | ( n6586 & n28477 ) | ( n28476 & n28477 ) ;
  assign n28483 = ( n953 & n3691 ) | ( n953 & ~n11938 ) | ( n3691 & ~n11938 ) ;
  assign n28484 = ( n3910 & n26413 ) | ( n3910 & ~n28483 ) | ( n26413 & ~n28483 ) ;
  assign n28480 = n22121 ^ n9197 ^ 1'b0 ;
  assign n28479 = n23081 ^ n21703 ^ n12830 ;
  assign n28481 = n28480 ^ n28479 ^ n820 ;
  assign n28482 = ( n9598 & n19869 ) | ( n9598 & ~n28481 ) | ( n19869 & ~n28481 ) ;
  assign n28485 = n28484 ^ n28482 ^ n26806 ;
  assign n28487 = n22591 ^ n11954 ^ n3182 ;
  assign n28486 = ( ~n7628 & n8317 ) | ( ~n7628 & n9165 ) | ( n8317 & n9165 ) ;
  assign n28488 = n28487 ^ n28486 ^ n12290 ;
  assign n28489 = n18552 ^ n12324 ^ n521 ;
  assign n28490 = ( n1524 & ~n27852 ) | ( n1524 & n28489 ) | ( ~n27852 & n28489 ) ;
  assign n28491 = n8142 ^ n3673 ^ 1'b0 ;
  assign n28492 = ( n2719 & n6205 ) | ( n2719 & ~n10192 ) | ( n6205 & ~n10192 ) ;
  assign n28493 = ( n28490 & n28491 ) | ( n28490 & n28492 ) | ( n28491 & n28492 ) ;
  assign n28494 = n10578 | n12042 ;
  assign n28495 = n28494 ^ n9966 ^ 1'b0 ;
  assign n28497 = n21906 ^ n7965 ^ n4968 ;
  assign n28496 = n9767 ^ n6655 ^ n4104 ;
  assign n28498 = n28497 ^ n28496 ^ n7182 ;
  assign n28499 = n28498 ^ n19994 ^ 1'b0 ;
  assign n28500 = n28495 & ~n28499 ;
  assign n28506 = ( ~n8686 & n10672 ) | ( ~n8686 & n25561 ) | ( n10672 & n25561 ) ;
  assign n28503 = n25425 ^ n15223 ^ 1'b0 ;
  assign n28504 = n4443 & n28503 ;
  assign n28505 = n28504 ^ n25918 ^ n3329 ;
  assign n28501 = n5682 & ~n23859 ;
  assign n28502 = n28501 ^ n26611 ^ 1'b0 ;
  assign n28507 = n28506 ^ n28505 ^ n28502 ;
  assign n28508 = n11774 | n28507 ;
  assign n28509 = n11869 & ~n28508 ;
  assign n28513 = ( n2642 & ~n5954 ) | ( n2642 & n12915 ) | ( ~n5954 & n12915 ) ;
  assign n28514 = n28513 ^ n25179 ^ n23816 ;
  assign n28510 = ( n12690 & ~n15437 ) | ( n12690 & n16230 ) | ( ~n15437 & n16230 ) ;
  assign n28511 = n28510 ^ n9971 ^ 1'b0 ;
  assign n28512 = ~n642 & n28511 ;
  assign n28515 = n28514 ^ n28512 ^ n416 ;
  assign n28516 = ( n5145 & n7663 ) | ( n5145 & ~n8103 ) | ( n7663 & ~n8103 ) ;
  assign n28517 = n28516 ^ n16748 ^ n12499 ;
  assign n28518 = ( ~n9186 & n28515 ) | ( ~n9186 & n28517 ) | ( n28515 & n28517 ) ;
  assign n28519 = n18112 ^ n15293 ^ n6974 ;
  assign n28520 = n22028 ^ n15293 ^ n14930 ;
  assign n28521 = n28520 ^ n17205 ^ 1'b0 ;
  assign n28522 = ( ~n1783 & n3366 ) | ( ~n1783 & n4384 ) | ( n3366 & n4384 ) ;
  assign n28523 = ( ~n3254 & n4528 ) | ( ~n3254 & n16709 ) | ( n4528 & n16709 ) ;
  assign n28524 = n6008 & n26684 ;
  assign n28525 = n28523 & n28524 ;
  assign n28526 = ( n11907 & n28522 ) | ( n11907 & ~n28525 ) | ( n28522 & ~n28525 ) ;
  assign n28527 = n7659 ^ n6663 ^ n3167 ;
  assign n28528 = ( n6158 & n21095 ) | ( n6158 & ~n28527 ) | ( n21095 & ~n28527 ) ;
  assign n28529 = n22799 ^ n21946 ^ n7196 ;
  assign n28530 = n1639 | n3984 ;
  assign n28531 = ( n17994 & n24658 ) | ( n17994 & ~n28530 ) | ( n24658 & ~n28530 ) ;
  assign n28532 = n28531 ^ n28239 ^ n15080 ;
  assign n28533 = ( n4355 & n7324 ) | ( n4355 & n28532 ) | ( n7324 & n28532 ) ;
  assign n28534 = n27201 ^ n16001 ^ 1'b0 ;
  assign n28535 = n28534 ^ n17582 ^ n11081 ;
  assign n28536 = n28535 ^ n19695 ^ n7680 ;
  assign n28537 = ( ~n2332 & n7378 ) | ( ~n2332 & n10620 ) | ( n7378 & n10620 ) ;
  assign n28538 = ( n2463 & ~n28283 ) | ( n2463 & n28537 ) | ( ~n28283 & n28537 ) ;
  assign n28539 = ~n24497 & n28538 ;
  assign n28540 = n28539 ^ n19516 ^ 1'b0 ;
  assign n28541 = n23605 ^ n11826 ^ n2708 ;
  assign n28542 = ( ~n9262 & n9269 ) | ( ~n9262 & n10770 ) | ( n9269 & n10770 ) ;
  assign n28543 = ( n2340 & n22306 ) | ( n2340 & n24224 ) | ( n22306 & n24224 ) ;
  assign n28544 = ( n7582 & n28542 ) | ( n7582 & n28543 ) | ( n28542 & n28543 ) ;
  assign n28545 = n25709 ^ n14883 ^ n4891 ;
  assign n28546 = ( ~n2790 & n15028 ) | ( ~n2790 & n17699 ) | ( n15028 & n17699 ) ;
  assign n28547 = ( ~n6895 & n9662 ) | ( ~n6895 & n28546 ) | ( n9662 & n28546 ) ;
  assign n28548 = n26674 ^ n11379 ^ n523 ;
  assign n28549 = n28548 ^ n10740 ^ n5713 ;
  assign n28558 = n9279 ^ x49 ^ 1'b0 ;
  assign n28556 = n17028 ^ n9580 ^ n1047 ;
  assign n28557 = ( n9370 & n16611 ) | ( n9370 & ~n28556 ) | ( n16611 & ~n28556 ) ;
  assign n28550 = ( n2336 & n2943 ) | ( n2336 & ~n11552 ) | ( n2943 & ~n11552 ) ;
  assign n28551 = n28550 ^ n8634 ^ n3828 ;
  assign n28552 = n6395 & ~n22971 ;
  assign n28553 = n18902 | n28552 ;
  assign n28554 = n2056 | n28553 ;
  assign n28555 = ( ~n13214 & n28551 ) | ( ~n13214 & n28554 ) | ( n28551 & n28554 ) ;
  assign n28559 = n28558 ^ n28557 ^ n28555 ;
  assign n28560 = n12067 & n21618 ;
  assign n28561 = n28560 ^ n19119 ^ n12947 ;
  assign n28562 = n28561 ^ n17540 ^ n14037 ;
  assign n28563 = n4645 ^ x154 ^ 1'b0 ;
  assign n28564 = ~n14457 & n28563 ;
  assign n28565 = ( n805 & ~n16436 ) | ( n805 & n18386 ) | ( ~n16436 & n18386 ) ;
  assign n28566 = ( n20728 & n26189 ) | ( n20728 & n28565 ) | ( n26189 & n28565 ) ;
  assign n28567 = n28566 ^ n20398 ^ n652 ;
  assign n28568 = n15647 & ~n20379 ;
  assign n28572 = n22869 ^ n12930 ^ n1589 ;
  assign n28569 = ( x17 & ~n6829 ) | ( x17 & n26966 ) | ( ~n6829 & n26966 ) ;
  assign n28570 = n18213 ^ n14439 ^ n7774 ;
  assign n28571 = ( ~n26431 & n28569 ) | ( ~n26431 & n28570 ) | ( n28569 & n28570 ) ;
  assign n28573 = n28572 ^ n28571 ^ n6207 ;
  assign n28574 = n9010 ^ n6898 ^ 1'b0 ;
  assign n28575 = n28574 ^ n17053 ^ n8403 ;
  assign n28576 = ( n17314 & ~n18467 ) | ( n17314 & n28575 ) | ( ~n18467 & n28575 ) ;
  assign n28577 = n28576 ^ n21257 ^ n10189 ;
  assign n28586 = ( ~n9963 & n11895 ) | ( ~n9963 & n23985 ) | ( n11895 & n23985 ) ;
  assign n28578 = n5298 ^ n2679 ^ 1'b0 ;
  assign n28579 = n9792 & n28578 ;
  assign n28580 = ( n14679 & n15302 ) | ( n14679 & ~n19585 ) | ( n15302 & ~n19585 ) ;
  assign n28581 = n28580 ^ n354 ^ 1'b0 ;
  assign n28582 = n21709 & n28581 ;
  assign n28583 = ( n14366 & n28579 ) | ( n14366 & ~n28582 ) | ( n28579 & ~n28582 ) ;
  assign n28584 = n28583 ^ n5218 ^ 1'b0 ;
  assign n28585 = ( n1039 & n1534 ) | ( n1039 & n28584 ) | ( n1534 & n28584 ) ;
  assign n28587 = n28586 ^ n28585 ^ 1'b0 ;
  assign n28588 = ( n3571 & ~n16834 ) | ( n3571 & n28197 ) | ( ~n16834 & n28197 ) ;
  assign n28589 = n28588 ^ n16306 ^ n14873 ;
  assign n28590 = n17819 ^ n15022 ^ 1'b0 ;
  assign n28591 = n13792 ^ n5386 ^ n1295 ;
  assign n28592 = ( n2127 & ~n16012 ) | ( n2127 & n28591 ) | ( ~n16012 & n28591 ) ;
  assign n28593 = ( ~n14104 & n19581 ) | ( ~n14104 & n28592 ) | ( n19581 & n28592 ) ;
  assign n28594 = ~n4013 & n9432 ;
  assign n28595 = ( ~n292 & n20900 ) | ( ~n292 & n28594 ) | ( n20900 & n28594 ) ;
  assign n28596 = ( n10340 & n10650 ) | ( n10340 & ~n28595 ) | ( n10650 & ~n28595 ) ;
  assign n28597 = n28596 ^ n14594 ^ n8919 ;
  assign n28598 = ~n14871 & n25689 ;
  assign n28599 = n28597 & n28598 ;
  assign n28600 = ( n13550 & n13728 ) | ( n13550 & n14874 ) | ( n13728 & n14874 ) ;
  assign n28601 = n28600 ^ n21821 ^ n19720 ;
  assign n28602 = ( n9668 & n16423 ) | ( n9668 & n28601 ) | ( n16423 & n28601 ) ;
  assign n28603 = n15668 ^ n5345 ^ n1036 ;
  assign n28606 = n26849 ^ n21156 ^ n5995 ;
  assign n28607 = n28606 ^ n17434 ^ n12140 ;
  assign n28604 = n20809 ^ n18502 ^ n9632 ;
  assign n28605 = n28604 ^ n25824 ^ n16233 ;
  assign n28608 = n28607 ^ n28605 ^ n25004 ;
  assign n28609 = n2989 | n10939 ;
  assign n28610 = n28609 ^ n10596 ^ 1'b0 ;
  assign n28611 = ( ~n17359 & n20095 ) | ( ~n17359 & n24388 ) | ( n20095 & n24388 ) ;
  assign n28612 = n22895 ^ n10171 ^ n2452 ;
  assign n28613 = n25399 ^ n23414 ^ n9132 ;
  assign n28614 = ( n28611 & n28612 ) | ( n28611 & ~n28613 ) | ( n28612 & ~n28613 ) ;
  assign n28615 = ( n13144 & n20545 ) | ( n13144 & ~n26819 ) | ( n20545 & ~n26819 ) ;
  assign n28616 = ( n1588 & ~n10103 ) | ( n1588 & n28615 ) | ( ~n10103 & n28615 ) ;
  assign n28617 = n28616 ^ n11091 ^ n1207 ;
  assign n28618 = ( n1627 & ~n23164 ) | ( n1627 & n28617 ) | ( ~n23164 & n28617 ) ;
  assign n28619 = n17470 ^ n6113 ^ n2796 ;
  assign n28620 = ~n301 & n28619 ;
  assign n28621 = ~n23053 & n28620 ;
  assign n28622 = ( n12640 & ~n17254 ) | ( n12640 & n27073 ) | ( ~n17254 & n27073 ) ;
  assign n28623 = n15881 ^ n14684 ^ n8970 ;
  assign n28624 = n28623 ^ n16165 ^ n14263 ;
  assign n28625 = ( n9245 & n10712 ) | ( n9245 & ~n15119 ) | ( n10712 & ~n15119 ) ;
  assign n28626 = n28625 ^ n27515 ^ n26598 ;
  assign n28630 = ( n9244 & n18795 ) | ( n9244 & n24706 ) | ( n18795 & n24706 ) ;
  assign n28631 = n28630 ^ n20377 ^ n16477 ;
  assign n28627 = n18662 ^ n3104 ^ 1'b0 ;
  assign n28628 = n2828 & n28627 ;
  assign n28629 = n18779 | n28628 ;
  assign n28632 = n28631 ^ n28629 ^ n10129 ;
  assign n28633 = n28632 ^ n18626 ^ n3954 ;
  assign n28634 = n28633 ^ n18239 ^ n577 ;
  assign n28635 = n24742 ^ n12687 ^ n11683 ;
  assign n28640 = n854 | n1428 ;
  assign n28641 = n8301 & ~n28640 ;
  assign n28636 = n14723 ^ n10618 ^ n9159 ;
  assign n28637 = n9915 | n12590 ;
  assign n28638 = n28637 ^ n7460 ^ n5575 ;
  assign n28639 = ( ~n14587 & n28636 ) | ( ~n14587 & n28638 ) | ( n28636 & n28638 ) ;
  assign n28642 = n28641 ^ n28639 ^ n20033 ;
  assign n28643 = n23560 & ~n28642 ;
  assign n28644 = n28643 ^ n5750 ^ x222 ;
  assign n28645 = n25451 ^ n13498 ^ n856 ;
  assign n28646 = ( n5606 & ~n6718 ) | ( n5606 & n14495 ) | ( ~n6718 & n14495 ) ;
  assign n28647 = n20397 ^ n6511 ^ 1'b0 ;
  assign n28648 = n11648 | n28647 ;
  assign n28649 = n7844 | n25362 ;
  assign n28650 = n25575 ^ n7840 ^ 1'b0 ;
  assign n28651 = n6510 | n28650 ;
  assign n28652 = n28651 ^ n19270 ^ n18946 ;
  assign n28653 = n16616 ^ n8815 ^ n3202 ;
  assign n28654 = n28653 ^ n6574 ^ 1'b0 ;
  assign n28655 = ( n22269 & n24460 ) | ( n22269 & ~n28654 ) | ( n24460 & ~n28654 ) ;
  assign n28656 = n12475 & ~n14722 ;
  assign n28657 = n8761 & n28656 ;
  assign n28658 = n28657 ^ n24288 ^ n5176 ;
  assign n28659 = n22047 ^ n21145 ^ n8582 ;
  assign n28660 = ( ~n1420 & n11716 ) | ( ~n1420 & n28659 ) | ( n11716 & n28659 ) ;
  assign n28661 = ( n16058 & n28658 ) | ( n16058 & ~n28660 ) | ( n28658 & ~n28660 ) ;
  assign n28662 = ( n17823 & n21097 ) | ( n17823 & n25900 ) | ( n21097 & n25900 ) ;
  assign n28663 = ( n17452 & ~n21815 ) | ( n17452 & n28662 ) | ( ~n21815 & n28662 ) ;
  assign n28664 = n1107 & n17612 ;
  assign n28665 = n28664 ^ n24665 ^ n8155 ;
  assign n28666 = n25635 ^ n6416 ^ 1'b0 ;
  assign n28667 = n8134 & n28666 ;
  assign n28668 = ~n4627 & n12333 ;
  assign n28672 = n364 | n1600 ;
  assign n28669 = ( ~x234 & n954 ) | ( ~x234 & n23475 ) | ( n954 & n23475 ) ;
  assign n28670 = ( n3977 & n19264 ) | ( n3977 & ~n28669 ) | ( n19264 & ~n28669 ) ;
  assign n28671 = n28670 ^ n21490 ^ n2756 ;
  assign n28673 = n28672 ^ n28671 ^ n11177 ;
  assign n28674 = ( ~n11543 & n16103 ) | ( ~n11543 & n16701 ) | ( n16103 & n16701 ) ;
  assign n28677 = ( ~n11776 & n12214 ) | ( ~n11776 & n16640 ) | ( n12214 & n16640 ) ;
  assign n28675 = ~n1586 & n4128 ;
  assign n28676 = n28675 ^ n19519 ^ n8697 ;
  assign n28678 = n28677 ^ n28676 ^ n20605 ;
  assign n28679 = n14156 & n28137 ;
  assign n28680 = ( n12919 & ~n20228 ) | ( n12919 & n28048 ) | ( ~n20228 & n28048 ) ;
  assign n28681 = ( ~n9877 & n22218 ) | ( ~n9877 & n28680 ) | ( n22218 & n28680 ) ;
  assign n28682 = ( n5836 & n28679 ) | ( n5836 & n28681 ) | ( n28679 & n28681 ) ;
  assign n28683 = ( ~n3753 & n10429 ) | ( ~n3753 & n22861 ) | ( n10429 & n22861 ) ;
  assign n28684 = n28683 ^ n15224 ^ n6129 ;
  assign n28685 = ( ~n13554 & n17394 ) | ( ~n13554 & n28684 ) | ( n17394 & n28684 ) ;
  assign n28692 = n15973 ^ n4373 ^ n493 ;
  assign n28686 = ( ~n10657 & n12342 ) | ( ~n10657 & n21415 ) | ( n12342 & n21415 ) ;
  assign n28687 = n28686 ^ n25604 ^ n1563 ;
  assign n28688 = ( ~n8307 & n10820 ) | ( ~n8307 & n22173 ) | ( n10820 & n22173 ) ;
  assign n28689 = ( n20928 & n28687 ) | ( n20928 & n28688 ) | ( n28687 & n28688 ) ;
  assign n28690 = n9607 ^ n7351 ^ n4816 ;
  assign n28691 = n28689 | n28690 ;
  assign n28693 = n28692 ^ n28691 ^ 1'b0 ;
  assign n28694 = ( n982 & n11663 ) | ( n982 & ~n16469 ) | ( n11663 & ~n16469 ) ;
  assign n28695 = n26384 ^ n18766 ^ n9042 ;
  assign n28696 = ( n13258 & n28694 ) | ( n13258 & n28695 ) | ( n28694 & n28695 ) ;
  assign n28697 = ( n3042 & n23083 ) | ( n3042 & n28696 ) | ( n23083 & n28696 ) ;
  assign n28698 = ( x195 & ~n19108 ) | ( x195 & n20800 ) | ( ~n19108 & n20800 ) ;
  assign n28699 = n9132 ^ n8914 ^ n6610 ;
  assign n28700 = ( n817 & n23140 ) | ( n817 & ~n28699 ) | ( n23140 & ~n28699 ) ;
  assign n28701 = ( ~n28405 & n28698 ) | ( ~n28405 & n28700 ) | ( n28698 & n28700 ) ;
  assign n28702 = n11669 & n17784 ;
  assign n28703 = n9865 & ~n21505 ;
  assign n28704 = ( n800 & n5649 ) | ( n800 & ~n19704 ) | ( n5649 & ~n19704 ) ;
  assign n28705 = n28704 ^ n5994 ^ n5087 ;
  assign n28706 = n12574 & n15496 ;
  assign n28707 = n1954 & n28706 ;
  assign n28708 = ( n12035 & ~n22293 ) | ( n12035 & n28707 ) | ( ~n22293 & n28707 ) ;
  assign n28709 = n6919 ^ x103 ^ 1'b0 ;
  assign n28710 = n16900 & n28709 ;
  assign n28711 = n28710 ^ n13354 ^ 1'b0 ;
  assign n28715 = n22484 ^ n16037 ^ n1929 ;
  assign n28716 = n28715 ^ n11092 ^ 1'b0 ;
  assign n28713 = n9939 | n17592 ;
  assign n28712 = ~n3628 & n21780 ;
  assign n28714 = n28713 ^ n28712 ^ n18653 ;
  assign n28717 = n28716 ^ n28714 ^ n17215 ;
  assign n28718 = ( n5298 & n17458 ) | ( n5298 & ~n22525 ) | ( n17458 & ~n22525 ) ;
  assign n28719 = n28718 ^ n12065 ^ 1'b0 ;
  assign n28720 = ( ~n3384 & n13073 ) | ( ~n3384 & n14130 ) | ( n13073 & n14130 ) ;
  assign n28721 = ( ~n7369 & n11692 ) | ( ~n7369 & n14321 ) | ( n11692 & n14321 ) ;
  assign n28722 = n28721 ^ n18953 ^ n3335 ;
  assign n28723 = ( n18078 & n28720 ) | ( n18078 & n28722 ) | ( n28720 & n28722 ) ;
  assign n28724 = ( n4519 & n12113 ) | ( n4519 & ~n24104 ) | ( n12113 & ~n24104 ) ;
  assign n28725 = n28724 ^ n23226 ^ n15637 ;
  assign n28726 = ( n4979 & ~n8228 ) | ( n4979 & n16028 ) | ( ~n8228 & n16028 ) ;
  assign n28727 = n28726 ^ n6479 ^ n1912 ;
  assign n28728 = n6974 & ~n13522 ;
  assign n28729 = n9960 & n28728 ;
  assign n28730 = n26305 ^ n22124 ^ n8645 ;
  assign n28731 = ( n1841 & ~n28729 ) | ( n1841 & n28730 ) | ( ~n28729 & n28730 ) ;
  assign n28732 = n16183 ^ n12676 ^ x148 ;
  assign n28733 = n28732 ^ n6300 ^ n6013 ;
  assign n28734 = ( n14587 & n18150 ) | ( n14587 & ~n28733 ) | ( n18150 & ~n28733 ) ;
  assign n28735 = n7651 ^ n3590 ^ 1'b0 ;
  assign n28736 = n15503 ^ n14349 ^ x53 ;
  assign n28737 = ( ~n3814 & n8953 ) | ( ~n3814 & n16732 ) | ( n8953 & n16732 ) ;
  assign n28738 = n4048 ^ n2176 ^ 1'b0 ;
  assign n28739 = n1382 & n28738 ;
  assign n28740 = n28739 ^ n9521 ^ n3868 ;
  assign n28741 = ( n4281 & n20268 ) | ( n4281 & ~n28740 ) | ( n20268 & ~n28740 ) ;
  assign n28742 = n28741 ^ n19621 ^ 1'b0 ;
  assign n28743 = ~n28737 & n28742 ;
  assign n28744 = n9724 ^ n4682 ^ n3998 ;
  assign n28745 = ( n9731 & ~n19684 ) | ( n9731 & n28744 ) | ( ~n19684 & n28744 ) ;
  assign n28746 = n28745 ^ n26725 ^ n3039 ;
  assign n28747 = n22145 ^ n2197 ^ 1'b0 ;
  assign n28748 = n13798 | n28747 ;
  assign n28749 = n4243 | n14539 ;
  assign n28750 = n28749 ^ n11765 ^ 1'b0 ;
  assign n28751 = n28748 & ~n28750 ;
  assign n28752 = n25561 ^ n16618 ^ n2395 ;
  assign n28753 = n28752 ^ n5678 ^ n2621 ;
  assign n28754 = ( n15878 & n16654 ) | ( n15878 & n28753 ) | ( n16654 & n28753 ) ;
  assign n28755 = n24969 ^ n23846 ^ 1'b0 ;
  assign n28756 = n13004 ^ n8036 ^ 1'b0 ;
  assign n28757 = n26038 ^ n16398 ^ 1'b0 ;
  assign n28758 = n28756 | n28757 ;
  assign n28759 = n26557 ^ n2053 ^ 1'b0 ;
  assign n28760 = n28759 ^ n22600 ^ n14690 ;
  assign n28764 = n23526 ^ n5201 ^ n340 ;
  assign n28763 = ( ~n3293 & n3742 ) | ( ~n3293 & n20913 ) | ( n3742 & n20913 ) ;
  assign n28761 = ( n3135 & n5953 ) | ( n3135 & ~n21098 ) | ( n5953 & ~n21098 ) ;
  assign n28762 = n28761 ^ n24972 ^ 1'b0 ;
  assign n28765 = n28764 ^ n28763 ^ n28762 ;
  assign n28766 = n8525 ^ n7295 ^ n5075 ;
  assign n28767 = ( n3691 & n11522 ) | ( n3691 & n28766 ) | ( n11522 & n28766 ) ;
  assign n28768 = ( x240 & n4368 ) | ( x240 & n18200 ) | ( n4368 & n18200 ) ;
  assign n28769 = ( n2394 & ~n4992 ) | ( n2394 & n12161 ) | ( ~n4992 & n12161 ) ;
  assign n28770 = ( ~n13763 & n25762 ) | ( ~n13763 & n28769 ) | ( n25762 & n28769 ) ;
  assign n28771 = ( n28767 & ~n28768 ) | ( n28767 & n28770 ) | ( ~n28768 & n28770 ) ;
  assign n28772 = n28771 ^ n11344 ^ n3730 ;
  assign n28773 = ( n4215 & n5574 ) | ( n4215 & ~n19009 ) | ( n5574 & ~n19009 ) ;
  assign n28774 = n27172 ^ n15718 ^ n8735 ;
  assign n28775 = n28774 ^ n25650 ^ n17784 ;
  assign n28776 = ( ~n4331 & n28773 ) | ( ~n4331 & n28775 ) | ( n28773 & n28775 ) ;
  assign n28777 = n18162 ^ n9601 ^ 1'b0 ;
  assign n28778 = n20505 & n28777 ;
  assign n28779 = n28778 ^ n28445 ^ n12362 ;
  assign n28780 = n2432 | n28779 ;
  assign n28781 = n11599 ^ n7828 ^ n806 ;
  assign n28782 = ( n1652 & n3319 ) | ( n1652 & n23185 ) | ( n3319 & n23185 ) ;
  assign n28783 = ( n4349 & n18315 ) | ( n4349 & ~n28782 ) | ( n18315 & ~n28782 ) ;
  assign n28784 = ( n28780 & ~n28781 ) | ( n28780 & n28783 ) | ( ~n28781 & n28783 ) ;
  assign n28785 = n1666 & n22889 ;
  assign n28786 = n3439 & n28785 ;
  assign n28787 = n7859 ^ n5251 ^ n3412 ;
  assign n28788 = n28575 ^ n13229 ^ 1'b0 ;
  assign n28789 = n28787 & n28788 ;
  assign n28790 = ( n4308 & n17381 ) | ( n4308 & ~n19702 ) | ( n17381 & ~n19702 ) ;
  assign n28791 = ( n17194 & ~n17553 ) | ( n17194 & n28790 ) | ( ~n17553 & n28790 ) ;
  assign n28792 = ( ~n7446 & n8794 ) | ( ~n7446 & n28791 ) | ( n8794 & n28791 ) ;
  assign n28794 = ( ~n292 & n15923 ) | ( ~n292 & n19287 ) | ( n15923 & n19287 ) ;
  assign n28793 = n11257 | n15444 ;
  assign n28795 = n28794 ^ n28793 ^ 1'b0 ;
  assign n28796 = ( n24460 & n28792 ) | ( n24460 & n28795 ) | ( n28792 & n28795 ) ;
  assign n28797 = n8500 | n21275 ;
  assign n28798 = n28797 ^ n26604 ^ 1'b0 ;
  assign n28799 = ( n3762 & n27332 ) | ( n3762 & n28798 ) | ( n27332 & n28798 ) ;
  assign n28800 = n25151 ^ n10073 ^ x169 ;
  assign n28801 = n6422 ^ n4597 ^ n1613 ;
  assign n28802 = n15980 & ~n28801 ;
  assign n28803 = n28802 ^ n19736 ^ n3028 ;
  assign n28804 = n5011 & n8485 ;
  assign n28805 = n28804 ^ n18261 ^ n13909 ;
  assign n28806 = n28754 | n28805 ;
  assign n28807 = n28806 ^ x216 ^ 1'b0 ;
  assign n28808 = n14858 ^ n14643 ^ n9647 ;
  assign n28809 = ~n3481 & n6148 ;
  assign n28810 = ( n1478 & ~n18003 ) | ( n1478 & n28809 ) | ( ~n18003 & n28809 ) ;
  assign n28811 = ( n22186 & n28808 ) | ( n22186 & ~n28810 ) | ( n28808 & ~n28810 ) ;
  assign n28812 = ( n6777 & ~n22556 ) | ( n6777 & n23549 ) | ( ~n22556 & n23549 ) ;
  assign n28813 = n27811 ^ n5401 ^ n3842 ;
  assign n28814 = n15430 ^ n14727 ^ n1005 ;
  assign n28815 = n13044 ^ n12848 ^ n6038 ;
  assign n28816 = ( n3448 & n28814 ) | ( n3448 & n28815 ) | ( n28814 & n28815 ) ;
  assign n28817 = n28816 ^ n13418 ^ n7383 ;
  assign n28818 = ( n574 & n4314 ) | ( n574 & ~n4443 ) | ( n4314 & ~n4443 ) ;
  assign n28821 = n2488 | n13985 ;
  assign n28822 = n25652 | n28821 ;
  assign n28819 = n11904 ^ n3387 ^ n2544 ;
  assign n28820 = n28819 ^ n26340 ^ n5366 ;
  assign n28823 = n28822 ^ n28820 ^ n3963 ;
  assign n28824 = n7922 & ~n18029 ;
  assign n28825 = n28824 ^ n24778 ^ 1'b0 ;
  assign n28826 = n24637 ^ n2641 ^ n1994 ;
  assign n28827 = n28825 | n28826 ;
  assign n28828 = n7486 & ~n28827 ;
  assign n28829 = n19708 ^ n11709 ^ n7447 ;
  assign n28831 = n11901 ^ n3100 ^ 1'b0 ;
  assign n28832 = n11047 & ~n28831 ;
  assign n28830 = ~n5761 & n9697 ;
  assign n28833 = n28832 ^ n28830 ^ n14708 ;
  assign n28834 = n15694 ^ n5798 ^ 1'b0 ;
  assign n28835 = n28834 ^ n2708 ^ 1'b0 ;
  assign n28836 = n6082 & n11566 ;
  assign n28837 = n26064 ^ n18334 ^ n17930 ;
  assign n28838 = ~n6850 & n28837 ;
  assign n28839 = n10277 | n18824 ;
  assign n28840 = n6974 | n28839 ;
  assign n28841 = ( n18892 & n28838 ) | ( n18892 & n28840 ) | ( n28838 & n28840 ) ;
  assign n28842 = ( n5115 & n6235 ) | ( n5115 & ~n8664 ) | ( n6235 & ~n8664 ) ;
  assign n28843 = ( n28836 & ~n28841 ) | ( n28836 & n28842 ) | ( ~n28841 & n28842 ) ;
  assign n28844 = ( n3314 & n4094 ) | ( n3314 & ~n25816 ) | ( n4094 & ~n25816 ) ;
  assign n28845 = ( x118 & ~n4247 ) | ( x118 & n12962 ) | ( ~n4247 & n12962 ) ;
  assign n28846 = ( n2278 & n20052 ) | ( n2278 & ~n28845 ) | ( n20052 & ~n28845 ) ;
  assign n28847 = n16547 ^ n12973 ^ n10919 ;
  assign n28848 = n28847 ^ n4342 ^ n2116 ;
  assign n28849 = n28848 ^ n23219 ^ n9112 ;
  assign n28850 = ( ~n9924 & n23929 ) | ( ~n9924 & n28849 ) | ( n23929 & n28849 ) ;
  assign n28851 = n21908 ^ n15870 ^ 1'b0 ;
  assign n28852 = n28851 ^ n24965 ^ n8490 ;
  assign n28853 = n28850 | n28852 ;
  assign n28854 = ( n28844 & ~n28846 ) | ( n28844 & n28853 ) | ( ~n28846 & n28853 ) ;
  assign n28855 = ( n7724 & n21200 ) | ( n7724 & n23776 ) | ( n21200 & n23776 ) ;
  assign n28856 = n25825 ^ n21116 ^ 1'b0 ;
  assign n28857 = n28855 & ~n28856 ;
  assign n28859 = ( ~n1670 & n2780 ) | ( ~n1670 & n23783 ) | ( n2780 & n23783 ) ;
  assign n28858 = n16514 ^ n15260 ^ n4675 ;
  assign n28860 = n28859 ^ n28858 ^ 1'b0 ;
  assign n28861 = n11386 & ~n28860 ;
  assign n28872 = n11214 ^ n11134 ^ n5568 ;
  assign n28870 = ( x148 & n10366 ) | ( x148 & ~n10977 ) | ( n10366 & ~n10977 ) ;
  assign n28866 = n6535 & ~n10719 ;
  assign n28867 = n28866 ^ n9107 ^ 1'b0 ;
  assign n28864 = ( n1590 & n2455 ) | ( n1590 & n22162 ) | ( n2455 & n22162 ) ;
  assign n28865 = ( n7837 & n13824 ) | ( n7837 & ~n28864 ) | ( n13824 & ~n28864 ) ;
  assign n28868 = n28867 ^ n28865 ^ n4564 ;
  assign n28869 = n3887 & ~n28868 ;
  assign n28871 = n28870 ^ n28869 ^ 1'b0 ;
  assign n28862 = ( n1095 & n4789 ) | ( n1095 & ~n11242 ) | ( n4789 & ~n11242 ) ;
  assign n28863 = ( n1176 & n20312 ) | ( n1176 & n28862 ) | ( n20312 & n28862 ) ;
  assign n28873 = n28872 ^ n28871 ^ n28863 ;
  assign n28874 = ( n5674 & n12893 ) | ( n5674 & ~n28348 ) | ( n12893 & ~n28348 ) ;
  assign n28875 = ( n4003 & ~n16180 ) | ( n4003 & n17407 ) | ( ~n16180 & n17407 ) ;
  assign n28876 = n580 & ~n18786 ;
  assign n28877 = n28876 ^ n1226 ^ 1'b0 ;
  assign n28878 = n6667 & ~n28877 ;
  assign n28879 = n28491 & n28878 ;
  assign n28880 = ( n14493 & ~n24016 ) | ( n14493 & n28879 ) | ( ~n24016 & n28879 ) ;
  assign n28881 = ( ~n12168 & n21426 ) | ( ~n12168 & n28880 ) | ( n21426 & n28880 ) ;
  assign n28882 = n14533 ^ n2725 ^ n669 ;
  assign n28883 = n18383 & n28882 ;
  assign n28894 = n21625 ^ n14256 ^ n12061 ;
  assign n28884 = n21839 ^ n10339 ^ n2807 ;
  assign n28885 = ( n4104 & n21018 ) | ( n4104 & n28884 ) | ( n21018 & n28884 ) ;
  assign n28886 = ~n3303 & n20020 ;
  assign n28887 = n14973 & ~n28886 ;
  assign n28888 = n25480 | n28887 ;
  assign n28889 = n15497 & ~n28888 ;
  assign n28890 = ( ~n12642 & n17789 ) | ( ~n12642 & n28889 ) | ( n17789 & n28889 ) ;
  assign n28891 = n20986 & ~n23579 ;
  assign n28892 = ( ~n18471 & n28890 ) | ( ~n18471 & n28891 ) | ( n28890 & n28891 ) ;
  assign n28893 = n28885 & ~n28892 ;
  assign n28895 = n28894 ^ n28893 ^ 1'b0 ;
  assign n28896 = n1085 & ~n12386 ;
  assign n28897 = n28896 ^ n8233 ^ 1'b0 ;
  assign n28898 = n28897 ^ n21503 ^ 1'b0 ;
  assign n28899 = ( n13933 & n18466 ) | ( n13933 & ~n21156 ) | ( n18466 & ~n21156 ) ;
  assign n28900 = ( n26340 & ~n28898 ) | ( n26340 & n28899 ) | ( ~n28898 & n28899 ) ;
  assign n28905 = n21791 ^ n8323 ^ n878 ;
  assign n28906 = n28905 ^ n16733 ^ n12360 ;
  assign n28901 = n25667 ^ n15500 ^ n1833 ;
  assign n28902 = n7247 & ~n28901 ;
  assign n28903 = ( n5801 & n24947 ) | ( n5801 & n28902 ) | ( n24947 & n28902 ) ;
  assign n28904 = n28903 ^ n24891 ^ n1580 ;
  assign n28907 = n28906 ^ n28904 ^ n26352 ;
  assign n28908 = n28094 ^ n4082 ^ n1379 ;
  assign n28909 = ( ~n8292 & n10091 ) | ( ~n8292 & n12570 ) | ( n10091 & n12570 ) ;
  assign n28910 = ( n5908 & n28908 ) | ( n5908 & ~n28909 ) | ( n28908 & ~n28909 ) ;
  assign n28911 = ( ~n19619 & n25234 ) | ( ~n19619 & n28910 ) | ( n25234 & n28910 ) ;
  assign n28912 = n6321 ^ n4758 ^ n1961 ;
  assign n28913 = n28912 ^ n7158 ^ 1'b0 ;
  assign n28914 = n17370 & n28913 ;
  assign n28915 = ( ~n1175 & n10670 ) | ( ~n1175 & n14480 ) | ( n10670 & n14480 ) ;
  assign n28916 = n17775 | n28915 ;
  assign n28917 = ( n13314 & n19598 ) | ( n13314 & ~n28916 ) | ( n19598 & ~n28916 ) ;
  assign n28927 = n6994 ^ n5546 ^ n1813 ;
  assign n28928 = n7610 & n28927 ;
  assign n28929 = ~n2143 & n28928 ;
  assign n28918 = n1662 & ~n18483 ;
  assign n28919 = n510 & n4942 ;
  assign n28920 = n6353 & n28919 ;
  assign n28921 = n835 & n16374 ;
  assign n28922 = ( n11159 & n28920 ) | ( n11159 & n28921 ) | ( n28920 & n28921 ) ;
  assign n28923 = n5563 & n15934 ;
  assign n28924 = n28923 ^ n2630 ^ 1'b0 ;
  assign n28925 = ( ~n23231 & n28922 ) | ( ~n23231 & n28924 ) | ( n28922 & n28924 ) ;
  assign n28926 = n28918 & n28925 ;
  assign n28930 = n28929 ^ n28926 ^ 1'b0 ;
  assign n28931 = ( n6802 & n9372 ) | ( n6802 & ~n11483 ) | ( n9372 & ~n11483 ) ;
  assign n28932 = n19260 ^ n15398 ^ n11893 ;
  assign n28933 = n4394 & ~n27260 ;
  assign n28934 = ( n1935 & n28932 ) | ( n1935 & n28933 ) | ( n28932 & n28933 ) ;
  assign n28935 = ( n28930 & ~n28931 ) | ( n28930 & n28934 ) | ( ~n28931 & n28934 ) ;
  assign n28936 = ( ~n380 & n2850 ) | ( ~n380 & n11659 ) | ( n2850 & n11659 ) ;
  assign n28937 = ~n19694 & n28936 ;
  assign n28938 = n28347 ^ n6593 ^ n5806 ;
  assign n28939 = ( n486 & n23616 ) | ( n486 & n28938 ) | ( n23616 & n28938 ) ;
  assign n28940 = ( ~n3716 & n20646 ) | ( ~n3716 & n28939 ) | ( n20646 & n28939 ) ;
  assign n28941 = ( n12228 & n24567 ) | ( n12228 & n28940 ) | ( n24567 & n28940 ) ;
  assign n28942 = n16990 ^ n10825 ^ n6299 ;
  assign n28943 = ( ~n7790 & n11411 ) | ( ~n7790 & n28942 ) | ( n11411 & n28942 ) ;
  assign n28944 = n28943 ^ n27654 ^ n2708 ;
  assign n28945 = ( n6747 & ~n15710 ) | ( n6747 & n21313 ) | ( ~n15710 & n21313 ) ;
  assign n28946 = n28945 ^ n24723 ^ n13169 ;
  assign n28947 = ( n16101 & ~n26690 ) | ( n16101 & n27326 ) | ( ~n26690 & n27326 ) ;
  assign n28948 = n21004 ^ n14842 ^ n3670 ;
  assign n28949 = ( n8746 & n16252 ) | ( n8746 & n28948 ) | ( n16252 & n28948 ) ;
  assign n28950 = n18001 ^ n11648 ^ n2017 ;
  assign n28951 = n28950 ^ n11996 ^ n2122 ;
  assign n28952 = ( x142 & n9607 ) | ( x142 & n11054 ) | ( n9607 & n11054 ) ;
  assign n28953 = ( ~n817 & n3003 ) | ( ~n817 & n13176 ) | ( n3003 & n13176 ) ;
  assign n28954 = n16939 ^ n12880 ^ n6543 ;
  assign n28955 = ( n9988 & ~n28953 ) | ( n9988 & n28954 ) | ( ~n28953 & n28954 ) ;
  assign n28956 = n28955 ^ n13364 ^ n11187 ;
  assign n28957 = ( n21325 & ~n28952 ) | ( n21325 & n28956 ) | ( ~n28952 & n28956 ) ;
  assign n28958 = n28957 ^ n2518 ^ 1'b0 ;
  assign n28959 = n28951 & ~n28958 ;
  assign n28960 = ( n1646 & ~n8903 ) | ( n1646 & n15707 ) | ( ~n8903 & n15707 ) ;
  assign n28961 = n11820 ^ n1934 ^ 1'b0 ;
  assign n28962 = n3320 & n28961 ;
  assign n28963 = n17815 & n28962 ;
  assign n28964 = n28963 ^ n15991 ^ 1'b0 ;
  assign n28965 = n8856 ^ n7524 ^ n6417 ;
  assign n28966 = ~n8761 & n28965 ;
  assign n28967 = ( n7010 & ~n28964 ) | ( n7010 & n28966 ) | ( ~n28964 & n28966 ) ;
  assign n28968 = n19367 & ~n23901 ;
  assign n28969 = ( n28960 & n28967 ) | ( n28960 & n28968 ) | ( n28967 & n28968 ) ;
  assign n28970 = n23180 ^ n15656 ^ n6170 ;
  assign n28971 = n28970 ^ n27873 ^ n26860 ;
  assign n28972 = ( ~n4651 & n6458 ) | ( ~n4651 & n16460 ) | ( n6458 & n16460 ) ;
  assign n28973 = ~n11034 & n28972 ;
  assign n28974 = n16263 & n28973 ;
  assign n28975 = n28974 ^ n22585 ^ n19291 ;
  assign n28976 = n581 | n28975 ;
  assign n28977 = n28976 ^ n17762 ^ n2602 ;
  assign n28982 = ( n3381 & n13387 ) | ( n3381 & ~n14190 ) | ( n13387 & ~n14190 ) ;
  assign n28983 = n28982 ^ n26002 ^ n6975 ;
  assign n28978 = ~n11590 & n20548 ;
  assign n28979 = n14697 | n16743 ;
  assign n28980 = ( n12763 & ~n16512 ) | ( n12763 & n28979 ) | ( ~n16512 & n28979 ) ;
  assign n28981 = n28978 | n28980 ;
  assign n28984 = n28983 ^ n28981 ^ n8935 ;
  assign n28985 = n28984 ^ n24083 ^ n9897 ;
  assign n28987 = n12039 ^ n8971 ^ n3169 ;
  assign n28988 = n28987 ^ n22509 ^ n14752 ;
  assign n28986 = n15660 ^ n2070 ^ n765 ;
  assign n28989 = n28988 ^ n28986 ^ n4775 ;
  assign n28990 = n18806 ^ n17103 ^ n8357 ;
  assign n28991 = n27849 ^ n9210 ^ n3158 ;
  assign n28992 = n28991 ^ n23597 ^ n7071 ;
  assign n28993 = ( n2131 & n14320 ) | ( n2131 & ~n14462 ) | ( n14320 & ~n14462 ) ;
  assign n28994 = ( n9003 & n20809 ) | ( n9003 & ~n28993 ) | ( n20809 & ~n28993 ) ;
  assign n28995 = n20833 ^ n10458 ^ n2883 ;
  assign n28996 = n17135 ^ n261 ^ x213 ;
  assign n28997 = ( n2015 & n16510 ) | ( n2015 & ~n28996 ) | ( n16510 & ~n28996 ) ;
  assign n28998 = n6646 & ~n28997 ;
  assign n28999 = ( n23102 & ~n28995 ) | ( n23102 & n28998 ) | ( ~n28995 & n28998 ) ;
  assign n29000 = n23635 ^ n8371 ^ n1552 ;
  assign n29001 = ( n4307 & n16770 ) | ( n4307 & ~n29000 ) | ( n16770 & ~n29000 ) ;
  assign n29002 = n14816 ^ n12013 ^ n9277 ;
  assign n29003 = n29002 ^ n10993 ^ 1'b0 ;
  assign n29004 = n7667 & n29003 ;
  assign n29005 = n29004 ^ n25134 ^ 1'b0 ;
  assign n29006 = n19749 | n20134 ;
  assign n29007 = n29006 ^ n3439 ^ 1'b0 ;
  assign n29009 = n24193 ^ n16969 ^ n7949 ;
  assign n29008 = ( n5341 & n11720 ) | ( n5341 & n25518 ) | ( n11720 & n25518 ) ;
  assign n29010 = n29009 ^ n29008 ^ 1'b0 ;
  assign n29013 = n24496 ^ n2551 ^ n1534 ;
  assign n29012 = n22268 ^ n18740 ^ n8506 ;
  assign n29014 = n29013 ^ n29012 ^ n7863 ;
  assign n29011 = ( n3511 & ~n5509 ) | ( n3511 & n25122 ) | ( ~n5509 & n25122 ) ;
  assign n29015 = n29014 ^ n29011 ^ n23275 ;
  assign n29016 = n13956 ^ n11499 ^ n964 ;
  assign n29017 = n29016 ^ n17302 ^ n12989 ;
  assign n29018 = ( n1788 & ~n16025 ) | ( n1788 & n29017 ) | ( ~n16025 & n29017 ) ;
  assign n29019 = n21474 ^ n8372 ^ n2603 ;
  assign n29020 = ( n9072 & n10083 ) | ( n9072 & n29019 ) | ( n10083 & n29019 ) ;
  assign n29021 = n29020 ^ n17859 ^ 1'b0 ;
  assign n29022 = n29021 ^ n9703 ^ n6960 ;
  assign n29023 = ( n3596 & n20883 ) | ( n3596 & n24697 ) | ( n20883 & n24697 ) ;
  assign n29024 = n22768 ^ n11450 ^ n1851 ;
  assign n29025 = n29024 ^ n15463 ^ n9587 ;
  assign n29026 = n23051 ^ n8539 ^ 1'b0 ;
  assign n29027 = ( n22685 & n29025 ) | ( n22685 & ~n29026 ) | ( n29025 & ~n29026 ) ;
  assign n29028 = n29027 ^ n22671 ^ n903 ;
  assign n29029 = ( n1459 & n10595 ) | ( n1459 & n29028 ) | ( n10595 & n29028 ) ;
  assign n29030 = x79 & ~n5897 ;
  assign n29031 = ~n13458 & n29030 ;
  assign n29032 = n10395 & ~n29031 ;
  assign n29033 = n14680 ^ n2786 ^ n2027 ;
  assign n29034 = n21013 ^ n4418 ^ n729 ;
  assign n29035 = n29034 ^ n13593 ^ 1'b0 ;
  assign n29036 = n25591 & n29035 ;
  assign n29037 = ( n15969 & n23356 ) | ( n15969 & ~n29036 ) | ( n23356 & ~n29036 ) ;
  assign n29038 = n17821 ^ n9752 ^ n5262 ;
  assign n29042 = ~n1627 & n5251 ;
  assign n29043 = ~n4080 & n29042 ;
  assign n29041 = n5459 & ~n9784 ;
  assign n29044 = n29043 ^ n29041 ^ 1'b0 ;
  assign n29040 = ~n18094 & n20744 ;
  assign n29045 = n29044 ^ n29040 ^ 1'b0 ;
  assign n29039 = ~n16721 & n19410 ;
  assign n29046 = n29045 ^ n29039 ^ n9440 ;
  assign n29047 = n22926 ^ n7447 ^ n1922 ;
  assign n29048 = ( n7282 & n9846 ) | ( n7282 & n21508 ) | ( n9846 & n21508 ) ;
  assign n29049 = n26558 ^ n14993 ^ 1'b0 ;
  assign n29050 = n7681 | n12015 ;
  assign n29051 = n2566 & ~n29050 ;
  assign n29052 = ( n3500 & n21864 ) | ( n3500 & ~n29051 ) | ( n21864 & ~n29051 ) ;
  assign n29053 = n7872 & ~n11124 ;
  assign n29054 = n20737 ^ n19711 ^ n15508 ;
  assign n29056 = ( n6955 & ~n9111 ) | ( n6955 & n9386 ) | ( ~n9111 & n9386 ) ;
  assign n29055 = ( n8240 & n19673 ) | ( n8240 & ~n24227 ) | ( n19673 & ~n24227 ) ;
  assign n29057 = n29056 ^ n29055 ^ n24015 ;
  assign n29059 = n18020 & n23872 ;
  assign n29058 = ( n6034 & n8415 ) | ( n6034 & ~n19716 ) | ( n8415 & ~n19716 ) ;
  assign n29060 = n29059 ^ n29058 ^ n11570 ;
  assign n29061 = n12129 ^ n8992 ^ n1748 ;
  assign n29062 = ( n18409 & ~n20845 ) | ( n18409 & n29061 ) | ( ~n20845 & n29061 ) ;
  assign n29063 = n20679 & ~n29062 ;
  assign n29064 = ~n5231 & n16311 ;
  assign n29065 = n6848 & n29064 ;
  assign n29066 = n9107 ^ n8058 ^ n6022 ;
  assign n29067 = n27017 ^ n23646 ^ n20572 ;
  assign n29068 = n10183 ^ n3808 ^ n3204 ;
  assign n29069 = n29068 ^ n7513 ^ n5443 ;
  assign n29070 = ( n1658 & n15212 ) | ( n1658 & ~n29069 ) | ( n15212 & ~n29069 ) ;
  assign n29071 = n25541 ^ n8314 ^ n511 ;
  assign n29072 = ( ~n7212 & n29070 ) | ( ~n7212 & n29071 ) | ( n29070 & n29071 ) ;
  assign n29073 = ( n14532 & n17233 ) | ( n14532 & ~n28489 ) | ( n17233 & ~n28489 ) ;
  assign n29074 = ( ~n16072 & n21231 ) | ( ~n16072 & n29073 ) | ( n21231 & n29073 ) ;
  assign n29075 = n29074 ^ n3590 ^ x1 ;
  assign n29076 = n23203 ^ n2780 ^ n2526 ;
  assign n29077 = ( n5721 & n5934 ) | ( n5721 & n6617 ) | ( n5934 & n6617 ) ;
  assign n29078 = n29077 ^ n4520 ^ n4145 ;
  assign n29079 = n14753 ^ n395 ^ 1'b0 ;
  assign n29080 = n29079 ^ n13236 ^ n10741 ;
  assign n29081 = n26632 ^ n21219 ^ n8725 ;
  assign n29085 = ( n2667 & ~n5397 ) | ( n2667 & n9355 ) | ( ~n5397 & n9355 ) ;
  assign n29086 = n3162 & n6416 ;
  assign n29087 = ( n5768 & ~n29085 ) | ( n5768 & n29086 ) | ( ~n29085 & n29086 ) ;
  assign n29082 = n25521 ^ n9419 ^ n3266 ;
  assign n29083 = ~n12601 & n29082 ;
  assign n29084 = n29083 ^ n5384 ^ 1'b0 ;
  assign n29088 = n29087 ^ n29084 ^ 1'b0 ;
  assign n29089 = n1008 | n25530 ;
  assign n29090 = n29089 ^ n13105 ^ 1'b0 ;
  assign n29091 = n29090 ^ n20788 ^ n3726 ;
  assign n29092 = ~n5267 & n23775 ;
  assign n29093 = n10188 | n15078 ;
  assign n29094 = n23201 & ~n29093 ;
  assign n29095 = n10904 ^ n1803 ^ 1'b0 ;
  assign n29096 = ( ~n16765 & n25876 ) | ( ~n16765 & n29095 ) | ( n25876 & n29095 ) ;
  assign n29097 = n29096 ^ n17061 ^ n3725 ;
  assign n29099 = n16291 ^ n3505 ^ n3048 ;
  assign n29100 = n29099 ^ n8957 ^ n3015 ;
  assign n29098 = n20226 ^ n19159 ^ n17269 ;
  assign n29101 = n29100 ^ n29098 ^ n10707 ;
  assign n29102 = n29101 ^ n11876 ^ n11866 ;
  assign n29103 = ( n6454 & n9946 ) | ( n6454 & ~n16058 ) | ( n9946 & ~n16058 ) ;
  assign n29104 = ( n14144 & ~n26497 ) | ( n14144 & n29103 ) | ( ~n26497 & n29103 ) ;
  assign n29105 = ( n1574 & n25695 ) | ( n1574 & n29104 ) | ( n25695 & n29104 ) ;
  assign n29106 = ( n21579 & n29102 ) | ( n21579 & ~n29105 ) | ( n29102 & ~n29105 ) ;
  assign n29107 = n18023 ^ n8738 ^ 1'b0 ;
  assign n29108 = n3750 ^ n2427 ^ x162 ;
  assign n29109 = n11643 ^ n2242 ^ 1'b0 ;
  assign n29110 = n29109 ^ n25123 ^ 1'b0 ;
  assign n29111 = n29110 ^ n23239 ^ n3916 ;
  assign n29112 = n12203 & n21097 ;
  assign n29113 = ( n17571 & n19293 ) | ( n17571 & n29112 ) | ( n19293 & n29112 ) ;
  assign n29114 = n24295 ^ n17871 ^ n8260 ;
  assign n29115 = n29114 ^ n13403 ^ n12780 ;
  assign n29116 = ( ~n1559 & n8859 ) | ( ~n1559 & n27489 ) | ( n8859 & n27489 ) ;
  assign n29117 = ( n9775 & ~n16567 ) | ( n9775 & n27142 ) | ( ~n16567 & n27142 ) ;
  assign n29118 = ( n22118 & ~n22678 ) | ( n22118 & n29117 ) | ( ~n22678 & n29117 ) ;
  assign n29121 = n2622 ^ n1921 ^ n677 ;
  assign n29122 = ( n1422 & n21187 ) | ( n1422 & n29121 ) | ( n21187 & n29121 ) ;
  assign n29123 = ( n3624 & n9361 ) | ( n3624 & n29122 ) | ( n9361 & n29122 ) ;
  assign n29124 = ( n11683 & ~n12927 ) | ( n11683 & n29123 ) | ( ~n12927 & n29123 ) ;
  assign n29119 = n18435 ^ n9229 ^ n3413 ;
  assign n29120 = ( n11734 & ~n15519 ) | ( n11734 & n29119 ) | ( ~n15519 & n29119 ) ;
  assign n29125 = n29124 ^ n29120 ^ n2062 ;
  assign n29126 = ( n7468 & ~n8563 ) | ( n7468 & n9151 ) | ( ~n8563 & n9151 ) ;
  assign n29127 = ( ~n2757 & n25377 ) | ( ~n2757 & n29126 ) | ( n25377 & n29126 ) ;
  assign n29128 = n29127 ^ n15155 ^ 1'b0 ;
  assign n29129 = n29125 & n29128 ;
  assign n29130 = ( n4964 & n5870 ) | ( n4964 & n13537 ) | ( n5870 & n13537 ) ;
  assign n29138 = n22296 ^ n5301 ^ n2775 ;
  assign n29139 = n29138 ^ n1802 ^ n587 ;
  assign n29136 = ( n7877 & ~n9943 ) | ( n7877 & n10671 ) | ( ~n9943 & n10671 ) ;
  assign n29137 = n29136 ^ n19831 ^ n5136 ;
  assign n29131 = ( n5206 & n10185 ) | ( n5206 & ~n12398 ) | ( n10185 & ~n12398 ) ;
  assign n29132 = n28137 ^ n16475 ^ 1'b0 ;
  assign n29133 = n29131 | n29132 ;
  assign n29134 = n29133 ^ n23682 ^ 1'b0 ;
  assign n29135 = ( ~n2713 & n16648 ) | ( ~n2713 & n29134 ) | ( n16648 & n29134 ) ;
  assign n29140 = n29139 ^ n29137 ^ n29135 ;
  assign n29142 = n21503 ^ n17853 ^ n11206 ;
  assign n29143 = ( ~n6917 & n27807 ) | ( ~n6917 & n29142 ) | ( n27807 & n29142 ) ;
  assign n29141 = ( ~n10040 & n20384 ) | ( ~n10040 & n22643 ) | ( n20384 & n22643 ) ;
  assign n29144 = n29143 ^ n29141 ^ n8369 ;
  assign n29145 = ( n7163 & ~n14905 ) | ( n7163 & n29043 ) | ( ~n14905 & n29043 ) ;
  assign n29151 = ( n3659 & ~n18608 ) | ( n3659 & n20407 ) | ( ~n18608 & n20407 ) ;
  assign n29148 = n14101 ^ n7606 ^ n2127 ;
  assign n29149 = n13651 ^ n11902 ^ n2781 ;
  assign n29150 = ( n8496 & ~n29148 ) | ( n8496 & n29149 ) | ( ~n29148 & n29149 ) ;
  assign n29146 = n23734 ^ n17631 ^ 1'b0 ;
  assign n29147 = n29146 ^ n14324 ^ n1922 ;
  assign n29152 = n29151 ^ n29150 ^ n29147 ;
  assign n29153 = n15702 ^ n4872 ^ n3117 ;
  assign n29154 = ( n5291 & n13574 ) | ( n5291 & ~n29153 ) | ( n13574 & ~n29153 ) ;
  assign n29155 = n29154 ^ n12357 ^ n11056 ;
  assign n29157 = n4748 ^ n3223 ^ n1093 ;
  assign n29156 = ( ~n15940 & n20939 ) | ( ~n15940 & n25381 ) | ( n20939 & n25381 ) ;
  assign n29158 = n29157 ^ n29156 ^ n2854 ;
  assign n29159 = n29158 ^ n16144 ^ n6014 ;
  assign n29160 = ( n13470 & n23403 ) | ( n13470 & n29159 ) | ( n23403 & n29159 ) ;
  assign n29161 = n7233 & ~n15836 ;
  assign n29162 = n29161 ^ n2101 ^ 1'b0 ;
  assign n29163 = ( n4587 & n9898 ) | ( n4587 & n29162 ) | ( n9898 & n29162 ) ;
  assign n29164 = n3155 & ~n4831 ;
  assign n29167 = ( n1631 & n6360 ) | ( n1631 & n16481 ) | ( n6360 & n16481 ) ;
  assign n29165 = ( x31 & n4900 ) | ( x31 & ~n9136 ) | ( n4900 & ~n9136 ) ;
  assign n29166 = n29165 ^ n27948 ^ x15 ;
  assign n29168 = n29167 ^ n29166 ^ n7583 ;
  assign n29169 = ( x31 & n641 ) | ( x31 & n8087 ) | ( n641 & n8087 ) ;
  assign n29170 = ( n17158 & ~n22098 ) | ( n17158 & n29169 ) | ( ~n22098 & n29169 ) ;
  assign n29171 = ( n8269 & n29168 ) | ( n8269 & ~n29170 ) | ( n29168 & ~n29170 ) ;
  assign n29172 = ( ~n23984 & n29164 ) | ( ~n23984 & n29171 ) | ( n29164 & n29171 ) ;
  assign n29173 = n26971 ^ n9395 ^ n8488 ;
  assign n29175 = n838 | n916 ;
  assign n29176 = n19974 | n29175 ;
  assign n29177 = ( ~n18796 & n19718 ) | ( ~n18796 & n29176 ) | ( n19718 & n29176 ) ;
  assign n29174 = ( ~n20802 & n20916 ) | ( ~n20802 & n21273 ) | ( n20916 & n21273 ) ;
  assign n29178 = n29177 ^ n29174 ^ n832 ;
  assign n29180 = ~n7368 & n7936 ;
  assign n29181 = ~n5826 & n29180 ;
  assign n29179 = n3436 & n7521 ;
  assign n29182 = n29181 ^ n29179 ^ n3652 ;
  assign n29183 = n7993 ^ n4041 ^ n3534 ;
  assign n29184 = n29183 ^ n13317 ^ n4531 ;
  assign n29185 = n15834 ^ n13788 ^ n8566 ;
  assign n29186 = n19938 ^ n13417 ^ n1880 ;
  assign n29187 = n29186 ^ n26214 ^ 1'b0 ;
  assign n29188 = ~n26277 & n29187 ;
  assign n29190 = n14204 ^ n7411 ^ n3385 ;
  assign n29191 = n29190 ^ n28996 ^ n14086 ;
  assign n29189 = n28120 ^ n5527 ^ 1'b0 ;
  assign n29192 = n29191 ^ n29189 ^ n17954 ;
  assign n29193 = ( n12912 & n14604 ) | ( n12912 & ~n24795 ) | ( n14604 & ~n24795 ) ;
  assign n29194 = ~n7084 & n22544 ;
  assign n29195 = n17218 ^ n9775 ^ n3250 ;
  assign n29196 = ( n4703 & n7855 ) | ( n4703 & n17982 ) | ( n7855 & n17982 ) ;
  assign n29197 = ( n2827 & ~n14924 ) | ( n2827 & n29196 ) | ( ~n14924 & n29196 ) ;
  assign n29198 = n19418 ^ n17662 ^ 1'b0 ;
  assign n29199 = n4413 & n29198 ;
  assign n29200 = ( ~n1575 & n8803 ) | ( ~n1575 & n29199 ) | ( n8803 & n29199 ) ;
  assign n29201 = ( n4708 & n12889 ) | ( n4708 & n25739 ) | ( n12889 & n25739 ) ;
  assign n29202 = ( n11904 & ~n13829 ) | ( n11904 & n20177 ) | ( ~n13829 & n20177 ) ;
  assign n29203 = n29202 ^ n26699 ^ n15563 ;
  assign n29204 = n22727 ^ n12302 ^ n2292 ;
  assign n29205 = n28427 ^ n27338 ^ 1'b0 ;
  assign n29206 = n29204 & ~n29205 ;
  assign n29208 = n5886 ^ n1336 ^ 1'b0 ;
  assign n29207 = ( n281 & n17057 ) | ( n281 & ~n28662 ) | ( n17057 & ~n28662 ) ;
  assign n29209 = n29208 ^ n29207 ^ n27218 ;
  assign n29213 = n14682 ^ n11666 ^ 1'b0 ;
  assign n29214 = ( n9428 & ~n10902 ) | ( n9428 & n29213 ) | ( ~n10902 & n29213 ) ;
  assign n29212 = n16847 ^ n14984 ^ n4115 ;
  assign n29215 = n29214 ^ n29212 ^ 1'b0 ;
  assign n29210 = n20570 ^ n16861 ^ n13466 ;
  assign n29211 = n29210 ^ n15156 ^ n14283 ;
  assign n29216 = n29215 ^ n29211 ^ 1'b0 ;
  assign n29218 = ( n2466 & n11871 ) | ( n2466 & n20088 ) | ( n11871 & n20088 ) ;
  assign n29217 = ( n1115 & n13760 ) | ( n1115 & n15515 ) | ( n13760 & n15515 ) ;
  assign n29219 = n29218 ^ n29217 ^ n13625 ;
  assign n29220 = n8676 ^ n4111 ^ 1'b0 ;
  assign n29221 = n2098 & ~n29220 ;
  assign n29222 = n15424 & n29221 ;
  assign n29223 = ~n12964 & n29222 ;
  assign n29224 = ( ~n608 & n24254 ) | ( ~n608 & n29054 ) | ( n24254 & n29054 ) ;
  assign n29225 = n23332 ^ n17867 ^ n9020 ;
  assign n29228 = n9480 ^ n7658 ^ 1'b0 ;
  assign n29229 = n22213 ^ n3548 ^ 1'b0 ;
  assign n29230 = ~n29228 & n29229 ;
  assign n29226 = ( n12491 & n13996 ) | ( n12491 & n27679 ) | ( n13996 & n27679 ) ;
  assign n29227 = n29226 ^ n25348 ^ n741 ;
  assign n29231 = n29230 ^ n29227 ^ n28461 ;
  assign n29233 = n10464 ^ n9626 ^ n5419 ;
  assign n29232 = ~n6388 & n22686 ;
  assign n29234 = n29233 ^ n29232 ^ 1'b0 ;
  assign n29235 = n12975 & ~n18973 ;
  assign n29236 = n29235 ^ n18053 ^ 1'b0 ;
  assign n29237 = ~n29234 & n29236 ;
  assign n29238 = n29237 ^ n15601 ^ n3366 ;
  assign n29239 = n22424 ^ n16480 ^ n3833 ;
  assign n29240 = n17562 ^ n9194 ^ n5089 ;
  assign n29241 = n29240 ^ n5450 ^ n306 ;
  assign n29242 = ( n2510 & n13581 ) | ( n2510 & ~n15552 ) | ( n13581 & ~n15552 ) ;
  assign n29243 = n29242 ^ n28431 ^ n20509 ;
  assign n29244 = n29243 ^ n19398 ^ n1471 ;
  assign n29245 = n26638 ^ n9446 ^ n5985 ;
  assign n29246 = n29245 ^ n6096 ^ n1121 ;
  assign n29247 = ( n27451 & n29244 ) | ( n27451 & ~n29246 ) | ( n29244 & ~n29246 ) ;
  assign n29252 = n4131 & n18033 ;
  assign n29253 = n29252 ^ n2400 ^ 1'b0 ;
  assign n29248 = ~n11812 & n25822 ;
  assign n29249 = n3304 & n29248 ;
  assign n29250 = n29249 ^ n5335 ^ n851 ;
  assign n29251 = ( n7408 & ~n10035 ) | ( n7408 & n29250 ) | ( ~n10035 & n29250 ) ;
  assign n29254 = n29253 ^ n29251 ^ n657 ;
  assign n29255 = n24635 ^ n4647 ^ 1'b0 ;
  assign n29256 = ( n2535 & n18797 ) | ( n2535 & ~n26184 ) | ( n18797 & ~n26184 ) ;
  assign n29257 = ( ~n14779 & n26044 ) | ( ~n14779 & n29256 ) | ( n26044 & n29256 ) ;
  assign n29258 = ( n7404 & ~n29255 ) | ( n7404 & n29257 ) | ( ~n29255 & n29257 ) ;
  assign n29259 = ( n1375 & ~n18539 ) | ( n1375 & n27591 ) | ( ~n18539 & n27591 ) ;
  assign n29260 = ( ~n12591 & n28988 ) | ( ~n12591 & n29259 ) | ( n28988 & n29259 ) ;
  assign n29263 = ( ~n5348 & n9000 ) | ( ~n5348 & n22145 ) | ( n9000 & n22145 ) ;
  assign n29261 = n23237 ^ n14126 ^ n5710 ;
  assign n29262 = n29261 ^ n22754 ^ x206 ;
  assign n29264 = n29263 ^ n29262 ^ n24067 ;
  assign n29265 = n17480 ^ n11513 ^ n4510 ;
  assign n29266 = ( ~n19190 & n20109 ) | ( ~n19190 & n27960 ) | ( n20109 & n27960 ) ;
  assign n29267 = n7034 & ~n29266 ;
  assign n29268 = n12247 & n29267 ;
  assign n29269 = ( ~n21965 & n28607 ) | ( ~n21965 & n29268 ) | ( n28607 & n29268 ) ;
  assign n29273 = n14368 ^ n6379 ^ n5239 ;
  assign n29270 = ( ~n5173 & n12262 ) | ( ~n5173 & n27478 ) | ( n12262 & n27478 ) ;
  assign n29271 = n14061 | n29270 ;
  assign n29272 = n2723 & n29271 ;
  assign n29274 = n29273 ^ n29272 ^ 1'b0 ;
  assign n29275 = n29274 ^ n26638 ^ n3862 ;
  assign n29276 = n26252 ^ n3121 ^ 1'b0 ;
  assign n29277 = n14876 ^ n9974 ^ 1'b0 ;
  assign n29278 = ( n14166 & n29276 ) | ( n14166 & ~n29277 ) | ( n29276 & ~n29277 ) ;
  assign n29279 = ( n7867 & ~n23275 ) | ( n7867 & n23956 ) | ( ~n23275 & n23956 ) ;
  assign n29280 = ( n2739 & n9289 ) | ( n2739 & n25879 ) | ( n9289 & n25879 ) ;
  assign n29281 = n1432 & ~n1440 ;
  assign n29282 = ( n9220 & n29280 ) | ( n9220 & ~n29281 ) | ( n29280 & ~n29281 ) ;
  assign n29283 = ( n21898 & n22095 ) | ( n21898 & n29282 ) | ( n22095 & n29282 ) ;
  assign n29285 = n19289 ^ n7506 ^ 1'b0 ;
  assign n29284 = ( ~n9789 & n10302 ) | ( ~n9789 & n19115 ) | ( n10302 & n19115 ) ;
  assign n29286 = n29285 ^ n29284 ^ n6690 ;
  assign n29287 = n9020 ^ n4002 ^ 1'b0 ;
  assign n29288 = n20424 ^ n15114 ^ n4171 ;
  assign n29289 = ( n13166 & ~n13936 ) | ( n13166 & n13958 ) | ( ~n13936 & n13958 ) ;
  assign n29290 = n29289 ^ n2870 ^ n2795 ;
  assign n29291 = ( n2947 & n13213 ) | ( n2947 & ~n29290 ) | ( n13213 & ~n29290 ) ;
  assign n29299 = ( ~n6859 & n10587 ) | ( ~n6859 & n27657 ) | ( n10587 & n27657 ) ;
  assign n29300 = n29299 ^ n12246 ^ n10299 ;
  assign n29294 = ~n2085 & n4087 ;
  assign n29295 = ~n11113 & n29294 ;
  assign n29296 = n3202 & ~n4639 ;
  assign n29297 = ( n10490 & ~n29295 ) | ( n10490 & n29296 ) | ( ~n29295 & n29296 ) ;
  assign n29292 = n1398 & n8938 ;
  assign n29293 = n29292 ^ n11368 ^ 1'b0 ;
  assign n29298 = n29297 ^ n29293 ^ n17069 ;
  assign n29301 = n29300 ^ n29298 ^ n7060 ;
  assign n29302 = ( ~n16031 & n29291 ) | ( ~n16031 & n29301 ) | ( n29291 & n29301 ) ;
  assign n29303 = ( ~n24098 & n29288 ) | ( ~n24098 & n29302 ) | ( n29288 & n29302 ) ;
  assign n29304 = ( n3642 & n9409 ) | ( n3642 & ~n10896 ) | ( n9409 & ~n10896 ) ;
  assign n29305 = n29304 ^ n17429 ^ n12466 ;
  assign n29306 = ( ~n6516 & n10002 ) | ( ~n6516 & n10976 ) | ( n10002 & n10976 ) ;
  assign n29307 = n14291 ^ n13272 ^ n12116 ;
  assign n29308 = n8632 ^ n927 ^ 1'b0 ;
  assign n29309 = n29308 ^ n14937 ^ n2207 ;
  assign n29310 = n14627 ^ n5874 ^ 1'b0 ;
  assign n29311 = n29309 & n29310 ;
  assign n29312 = ( n17662 & ~n29307 ) | ( n17662 & n29311 ) | ( ~n29307 & n29311 ) ;
  assign n29313 = ( n2427 & n29306 ) | ( n2427 & n29312 ) | ( n29306 & n29312 ) ;
  assign n29314 = n29305 & n29313 ;
  assign n29315 = n6366 ^ n3022 ^ 1'b0 ;
  assign n29316 = ( ~x90 & n2375 ) | ( ~x90 & n3570 ) | ( n2375 & n3570 ) ;
  assign n29317 = ( ~n2922 & n24869 ) | ( ~n2922 & n29316 ) | ( n24869 & n29316 ) ;
  assign n29318 = ( n4025 & n13030 ) | ( n4025 & n29317 ) | ( n13030 & n29317 ) ;
  assign n29319 = n28880 | n29318 ;
  assign n29320 = ( n6250 & n29315 ) | ( n6250 & ~n29319 ) | ( n29315 & ~n29319 ) ;
  assign n29321 = ( n4902 & n5177 ) | ( n4902 & n16210 ) | ( n5177 & n16210 ) ;
  assign n29322 = ( n810 & n2690 ) | ( n810 & n22493 ) | ( n2690 & n22493 ) ;
  assign n29323 = ~n4895 & n7156 ;
  assign n29324 = n11029 | n29323 ;
  assign n29325 = ( n2732 & n4734 ) | ( n2732 & ~n29324 ) | ( n4734 & ~n29324 ) ;
  assign n29326 = ( n3154 & ~n5065 ) | ( n3154 & n7554 ) | ( ~n5065 & n7554 ) ;
  assign n29327 = n29326 ^ n12047 ^ 1'b0 ;
  assign n29328 = n14337 | n29327 ;
  assign n29329 = ( n4772 & n13519 ) | ( n4772 & ~n16565 ) | ( n13519 & ~n16565 ) ;
  assign n29330 = n29329 ^ n24469 ^ n13007 ;
  assign n29331 = ( n13829 & n14633 ) | ( n13829 & ~n21983 ) | ( n14633 & ~n21983 ) ;
  assign n29332 = n9242 & ~n15898 ;
  assign n29333 = n29331 & n29332 ;
  assign n29334 = n29333 ^ n2319 ^ 1'b0 ;
  assign n29335 = n14868 ^ n6871 ^ n956 ;
  assign n29339 = ( n15030 & ~n20749 ) | ( n15030 & n23302 ) | ( ~n20749 & n23302 ) ;
  assign n29337 = x219 & ~n2245 ;
  assign n29338 = n19623 & n29337 ;
  assign n29340 = n29339 ^ n29338 ^ 1'b0 ;
  assign n29341 = ~n20792 & n29340 ;
  assign n29336 = ( n6962 & n9600 ) | ( n6962 & n18834 ) | ( n9600 & n18834 ) ;
  assign n29342 = n29341 ^ n29336 ^ n15757 ;
  assign n29343 = n29335 & ~n29342 ;
  assign n29344 = n11710 & n29343 ;
  assign n29345 = ( n16511 & n29334 ) | ( n16511 & ~n29344 ) | ( n29334 & ~n29344 ) ;
  assign n29346 = ( n9016 & n29330 ) | ( n9016 & ~n29345 ) | ( n29330 & ~n29345 ) ;
  assign n29347 = n26951 ^ n26351 ^ n8742 ;
  assign n29348 = n10009 & ~n19245 ;
  assign n29349 = n15079 ^ n2824 ^ n2617 ;
  assign n29350 = ( n4618 & n29348 ) | ( n4618 & ~n29349 ) | ( n29348 & ~n29349 ) ;
  assign n29351 = ( n8307 & n25851 ) | ( n8307 & n29350 ) | ( n25851 & n29350 ) ;
  assign n29352 = n5924 & ~n16765 ;
  assign n29353 = n29352 ^ n5130 ^ 1'b0 ;
  assign n29354 = n29353 ^ n22753 ^ n5304 ;
  assign n29355 = n27209 & ~n29354 ;
  assign n29356 = n29355 ^ n12207 ^ 1'b0 ;
  assign n29357 = n24373 ^ n17439 ^ n3561 ;
  assign n29358 = n29357 ^ n15664 ^ n6122 ;
  assign n29359 = n29358 ^ n13857 ^ n6233 ;
  assign n29360 = n28225 ^ n23774 ^ n19527 ;
  assign n29361 = n7812 ^ n3627 ^ 1'b0 ;
  assign n29362 = ~n8834 & n29361 ;
  assign n29363 = n29362 ^ n16988 ^ n10132 ;
  assign n29365 = ( x31 & n3237 ) | ( x31 & n8035 ) | ( n3237 & n8035 ) ;
  assign n29366 = ( n3742 & n5341 ) | ( n3742 & n29365 ) | ( n5341 & n29365 ) ;
  assign n29364 = n11877 ^ n10113 ^ n5528 ;
  assign n29367 = n29366 ^ n29364 ^ n10312 ;
  assign n29368 = n24197 ^ n13590 ^ n12335 ;
  assign n29369 = ( n7846 & ~n29367 ) | ( n7846 & n29368 ) | ( ~n29367 & n29368 ) ;
  assign n29370 = n13764 ^ n12973 ^ n12291 ;
  assign n29371 = n17281 ^ n6007 ^ n2917 ;
  assign n29372 = n29371 ^ n5956 ^ n4150 ;
  assign n29373 = ( ~n15503 & n29370 ) | ( ~n15503 & n29372 ) | ( n29370 & n29372 ) ;
  assign n29378 = ( n1030 & n4851 ) | ( n1030 & n25407 ) | ( n4851 & n25407 ) ;
  assign n29376 = n9504 ^ n2289 ^ 1'b0 ;
  assign n29377 = ( n7057 & n28639 ) | ( n7057 & ~n29376 ) | ( n28639 & ~n29376 ) ;
  assign n29374 = n13617 ^ n5730 ^ 1'b0 ;
  assign n29375 = ( n770 & ~n14560 ) | ( n770 & n29374 ) | ( ~n14560 & n29374 ) ;
  assign n29379 = n29378 ^ n29377 ^ n29375 ;
  assign n29380 = n24232 & n29379 ;
  assign n29381 = n18285 & n29380 ;
  assign n29382 = n29381 ^ n19749 ^ n10083 ;
  assign n29383 = ~n2249 & n11052 ;
  assign n29384 = n29383 ^ n12401 ^ 1'b0 ;
  assign n29385 = ( ~n18156 & n23617 ) | ( ~n18156 & n29384 ) | ( n23617 & n29384 ) ;
  assign n29386 = n29385 ^ n24821 ^ n12888 ;
  assign n29387 = ( ~n1382 & n3858 ) | ( ~n1382 & n11899 ) | ( n3858 & n11899 ) ;
  assign n29388 = n14611 ^ n14181 ^ n13530 ;
  assign n29389 = n29388 ^ n6137 ^ n2588 ;
  assign n29390 = n29389 ^ n8333 ^ 1'b0 ;
  assign n29391 = n29387 | n29390 ;
  assign n29395 = ( n22941 & ~n25238 ) | ( n22941 & n26534 ) | ( ~n25238 & n26534 ) ;
  assign n29393 = n26349 ^ n20365 ^ n7481 ;
  assign n29392 = n11170 ^ n5094 ^ n983 ;
  assign n29394 = n29393 ^ n29392 ^ n16329 ;
  assign n29396 = n29395 ^ n29394 ^ n2731 ;
  assign n29397 = ( x19 & n2775 ) | ( x19 & n19709 ) | ( n2775 & n19709 ) ;
  assign n29399 = ( n7408 & ~n25548 ) | ( n7408 & n26868 ) | ( ~n25548 & n26868 ) ;
  assign n29398 = ( n21829 & n25400 ) | ( n21829 & ~n25581 ) | ( n25400 & ~n25581 ) ;
  assign n29400 = n29399 ^ n29398 ^ n2943 ;
  assign n29401 = n20201 ^ n12244 ^ n11277 ;
  assign n29402 = ( ~n1651 & n3879 ) | ( ~n1651 & n7675 ) | ( n3879 & n7675 ) ;
  assign n29408 = n17278 ^ n16302 ^ n269 ;
  assign n29403 = n5768 ^ n331 ^ x59 ;
  assign n29404 = n29403 ^ n28038 ^ n487 ;
  assign n29405 = n11257 ^ n924 ^ 1'b0 ;
  assign n29406 = ~n29404 & n29405 ;
  assign n29407 = n29406 ^ n20251 ^ n5308 ;
  assign n29409 = n29408 ^ n29407 ^ n16104 ;
  assign n29410 = ( ~n5725 & n11466 ) | ( ~n5725 & n21906 ) | ( n11466 & n21906 ) ;
  assign n29411 = ( n3050 & ~n13484 ) | ( n3050 & n21585 ) | ( ~n13484 & n21585 ) ;
  assign n29412 = n11496 ^ n642 ^ 1'b0 ;
  assign n29413 = ~n13615 & n23174 ;
  assign n29414 = ( ~n12011 & n29412 ) | ( ~n12011 & n29413 ) | ( n29412 & n29413 ) ;
  assign n29415 = ( n5383 & n29411 ) | ( n5383 & n29414 ) | ( n29411 & n29414 ) ;
  assign n29416 = n9578 & ~n23268 ;
  assign n29417 = ~n2277 & n29416 ;
  assign n29418 = n10210 ^ n9124 ^ 1'b0 ;
  assign n29419 = n29418 ^ n21711 ^ n3826 ;
  assign n29420 = n29419 ^ n25565 ^ n2334 ;
  assign n29421 = ( n7584 & n15594 ) | ( n7584 & ~n29420 ) | ( n15594 & ~n29420 ) ;
  assign n29422 = ~n29417 & n29421 ;
  assign n29423 = n11352 ^ n6372 ^ n6102 ;
  assign n29424 = x222 & ~n25108 ;
  assign n29425 = n29424 ^ n11156 ^ n9160 ;
  assign n29426 = ( n13907 & n29329 ) | ( n13907 & n29425 ) | ( n29329 & n29425 ) ;
  assign n29427 = ( n4031 & n29423 ) | ( n4031 & n29426 ) | ( n29423 & n29426 ) ;
  assign n29428 = ~n3802 & n12407 ;
  assign n29429 = ~n15674 & n29428 ;
  assign n29430 = ( ~n17157 & n23893 ) | ( ~n17157 & n29429 ) | ( n23893 & n29429 ) ;
  assign n29431 = ( n20341 & ~n25674 ) | ( n20341 & n29430 ) | ( ~n25674 & n29430 ) ;
  assign n29432 = n7070 & n15588 ;
  assign n29433 = n18274 & n29432 ;
  assign n29434 = ( n14748 & n16821 ) | ( n14748 & ~n21287 ) | ( n16821 & ~n21287 ) ;
  assign n29438 = n2822 ^ n1709 ^ 1'b0 ;
  assign n29435 = n16606 ^ n12561 ^ n4234 ;
  assign n29436 = n29435 ^ n24214 ^ 1'b0 ;
  assign n29437 = ~n1912 & n29436 ;
  assign n29439 = n29438 ^ n29437 ^ 1'b0 ;
  assign n29440 = n29434 & n29439 ;
  assign n29441 = ( n14401 & n25607 ) | ( n14401 & ~n27799 ) | ( n25607 & ~n27799 ) ;
  assign n29445 = n6517 ^ n5701 ^ n2358 ;
  assign n29442 = n24657 ^ n7737 ^ n484 ;
  assign n29443 = n29442 ^ n6961 ^ 1'b0 ;
  assign n29444 = n23304 & ~n29443 ;
  assign n29446 = n29445 ^ n29444 ^ n16991 ;
  assign n29447 = n13970 ^ n10909 ^ n4965 ;
  assign n29454 = ( n13501 & n15155 ) | ( n13501 & n18222 ) | ( n15155 & n18222 ) ;
  assign n29451 = ( ~n6789 & n12927 ) | ( ~n6789 & n19375 ) | ( n12927 & n19375 ) ;
  assign n29452 = ( n2823 & n13760 ) | ( n2823 & n21645 ) | ( n13760 & n21645 ) ;
  assign n29453 = ( ~n11079 & n29451 ) | ( ~n11079 & n29452 ) | ( n29451 & n29452 ) ;
  assign n29448 = n24332 ^ n22863 ^ n8093 ;
  assign n29449 = ( ~n6164 & n20589 ) | ( ~n6164 & n29448 ) | ( n20589 & n29448 ) ;
  assign n29450 = n29449 ^ n11613 ^ n6487 ;
  assign n29455 = n29454 ^ n29453 ^ n29450 ;
  assign n29456 = n24327 ^ n15943 ^ n15812 ;
  assign n29457 = n29456 ^ n22466 ^ n3042 ;
  assign n29458 = n12461 ^ n6643 ^ n4927 ;
  assign n29459 = n29458 ^ n16935 ^ n11991 ;
  assign n29460 = ( ~n2620 & n21696 ) | ( ~n2620 & n29459 ) | ( n21696 & n29459 ) ;
  assign n29461 = n13744 ^ n5746 ^ n3222 ;
  assign n29462 = n7566 ^ n3724 ^ n2519 ;
  assign n29463 = n15230 ^ n3553 ^ 1'b0 ;
  assign n29464 = ( n6414 & n29462 ) | ( n6414 & n29463 ) | ( n29462 & n29463 ) ;
  assign n29465 = ( n3691 & n15705 ) | ( n3691 & n21213 ) | ( n15705 & n21213 ) ;
  assign n29466 = ( n7414 & n12707 ) | ( n7414 & n29465 ) | ( n12707 & n29465 ) ;
  assign n29467 = n29466 ^ n7505 ^ 1'b0 ;
  assign n29468 = n3261 | n28602 ;
  assign n29471 = ( n617 & n3512 ) | ( n617 & ~n7085 ) | ( n3512 & ~n7085 ) ;
  assign n29469 = ~n2470 & n3221 ;
  assign n29470 = ~n9603 & n29469 ;
  assign n29472 = n29471 ^ n29470 ^ n26160 ;
  assign n29473 = ( n21765 & n23126 ) | ( n21765 & n29472 ) | ( n23126 & n29472 ) ;
  assign n29475 = n23834 | n24586 ;
  assign n29474 = n29281 ^ n16995 ^ n4989 ;
  assign n29476 = n29475 ^ n29474 ^ n16063 ;
  assign n29477 = ( x237 & n11133 ) | ( x237 & ~n11389 ) | ( n11133 & ~n11389 ) ;
  assign n29478 = n11199 ^ n4560 ^ n3586 ;
  assign n29479 = n29478 ^ n5107 ^ n3956 ;
  assign n29483 = n26396 ^ n429 ^ 1'b0 ;
  assign n29480 = ( ~n6890 & n11327 ) | ( ~n6890 & n29103 ) | ( n11327 & n29103 ) ;
  assign n29481 = n29480 ^ n27261 ^ n22582 ;
  assign n29482 = n28422 & ~n29481 ;
  assign n29484 = n29483 ^ n29482 ^ 1'b0 ;
  assign n29485 = n1762 & n3715 ;
  assign n29486 = n29485 ^ n25853 ^ n21802 ;
  assign n29499 = n18501 ^ n8667 ^ 1'b0 ;
  assign n29500 = n23643 | n29499 ;
  assign n29501 = ( n10527 & ~n15454 ) | ( n10527 & n29500 ) | ( ~n15454 & n29500 ) ;
  assign n29494 = n9412 ^ n3733 ^ n2631 ;
  assign n29493 = ( n9059 & n15625 ) | ( n9059 & ~n21635 ) | ( n15625 & ~n21635 ) ;
  assign n29492 = n5064 ^ n2189 ^ 1'b0 ;
  assign n29495 = n29494 ^ n29493 ^ n29492 ;
  assign n29496 = n18603 ^ n6501 ^ 1'b0 ;
  assign n29497 = ( n7107 & n19417 ) | ( n7107 & ~n29496 ) | ( n19417 & ~n29496 ) ;
  assign n29498 = ( n854 & ~n29495 ) | ( n854 & n29497 ) | ( ~n29495 & n29497 ) ;
  assign n29487 = ~n5583 & n15179 ;
  assign n29488 = n24557 & n29487 ;
  assign n29489 = ~n8588 & n29488 ;
  assign n29490 = ( n14947 & ~n18787 ) | ( n14947 & n28076 ) | ( ~n18787 & n28076 ) ;
  assign n29491 = ( n15855 & n29489 ) | ( n15855 & ~n29490 ) | ( n29489 & ~n29490 ) ;
  assign n29502 = n29501 ^ n29498 ^ n29491 ;
  assign n29503 = n10977 ^ n10331 ^ n6565 ;
  assign n29504 = ( n16628 & n24671 ) | ( n16628 & ~n29503 ) | ( n24671 & ~n29503 ) ;
  assign n29505 = ( n6957 & ~n16474 ) | ( n6957 & n28239 ) | ( ~n16474 & n28239 ) ;
  assign n29506 = n17335 ^ n12754 ^ n5702 ;
  assign n29507 = n29506 ^ n29168 ^ n12448 ;
  assign n29508 = n12487 ^ n2441 ^ 1'b0 ;
  assign n29509 = n29508 ^ n2203 ^ n848 ;
  assign n29512 = ( n10111 & ~n11864 ) | ( n10111 & n18634 ) | ( ~n11864 & n18634 ) ;
  assign n29510 = n19864 & n24204 ;
  assign n29511 = n10731 & n29510 ;
  assign n29513 = n29512 ^ n29511 ^ n8833 ;
  assign n29522 = n8067 | n12524 ;
  assign n29523 = n29522 ^ n5042 ^ 1'b0 ;
  assign n29514 = n14276 ^ n7656 ^ n4439 ;
  assign n29515 = n20006 ^ n6182 ^ 1'b0 ;
  assign n29516 = n20503 & n29515 ;
  assign n29517 = ( n16047 & n29514 ) | ( n16047 & n29516 ) | ( n29514 & n29516 ) ;
  assign n29518 = n29517 ^ n319 ^ 1'b0 ;
  assign n29519 = n14752 | n29518 ;
  assign n29520 = n29519 ^ n1884 ^ 1'b0 ;
  assign n29521 = n29520 ^ n11900 ^ n7138 ;
  assign n29524 = n29523 ^ n29521 ^ n19643 ;
  assign n29525 = ( ~n2720 & n3851 ) | ( ~n2720 & n14649 ) | ( n3851 & n14649 ) ;
  assign n29526 = n3881 & ~n13232 ;
  assign n29527 = ( ~n1698 & n8891 ) | ( ~n1698 & n11679 ) | ( n8891 & n11679 ) ;
  assign n29528 = ( n18185 & n29526 ) | ( n18185 & ~n29527 ) | ( n29526 & ~n29527 ) ;
  assign n29529 = ~n29525 & n29528 ;
  assign n29530 = ( ~n7815 & n13687 ) | ( ~n7815 & n17111 ) | ( n13687 & n17111 ) ;
  assign n29531 = n13259 ^ n5572 ^ n2399 ;
  assign n29532 = ( n6061 & n29530 ) | ( n6061 & ~n29531 ) | ( n29530 & ~n29531 ) ;
  assign n29533 = n6812 & ~n27696 ;
  assign n29534 = n2523 & n29533 ;
  assign n29535 = n1082 | n21823 ;
  assign n29536 = ( ~n8204 & n11148 ) | ( ~n8204 & n26083 ) | ( n11148 & n26083 ) ;
  assign n29537 = n29536 ^ n29418 ^ n11887 ;
  assign n29538 = n29537 ^ n17822 ^ n11991 ;
  assign n29539 = n8031 ^ n1046 ^ x251 ;
  assign n29540 = n20933 & n29539 ;
  assign n29541 = ( n6462 & ~n19238 ) | ( n6462 & n29540 ) | ( ~n19238 & n29540 ) ;
  assign n29542 = ( n7011 & ~n15909 ) | ( n7011 & n29541 ) | ( ~n15909 & n29541 ) ;
  assign n29543 = ( ~n6068 & n6344 ) | ( ~n6068 & n9624 ) | ( n6344 & n9624 ) ;
  assign n29544 = ( ~n9823 & n17392 ) | ( ~n9823 & n29543 ) | ( n17392 & n29543 ) ;
  assign n29545 = n10886 & n29544 ;
  assign n29546 = n29542 & n29545 ;
  assign n29547 = ( n3864 & ~n12043 ) | ( n3864 & n18200 ) | ( ~n12043 & n18200 ) ;
  assign n29548 = n29547 ^ n4297 ^ n1446 ;
  assign n29549 = n28156 ^ n27167 ^ n6915 ;
  assign n29553 = n23176 & n24613 ;
  assign n29554 = ( ~n8604 & n13874 ) | ( ~n8604 & n29553 ) | ( n13874 & n29553 ) ;
  assign n29550 = ~n1006 & n8030 ;
  assign n29551 = n29550 ^ n17453 ^ n1581 ;
  assign n29552 = n29551 ^ n21695 ^ n8713 ;
  assign n29555 = n29554 ^ n29552 ^ n23611 ;
  assign n29561 = ( ~n8951 & n12247 ) | ( ~n8951 & n24705 ) | ( n12247 & n24705 ) ;
  assign n29556 = ( n7086 & n7605 ) | ( n7086 & ~n10034 ) | ( n7605 & ~n10034 ) ;
  assign n29557 = n29556 ^ n26063 ^ n7771 ;
  assign n29558 = ( n3670 & n15828 ) | ( n3670 & n29557 ) | ( n15828 & n29557 ) ;
  assign n29559 = n29558 ^ n9713 ^ n781 ;
  assign n29560 = n7179 | n29559 ;
  assign n29562 = n29561 ^ n29560 ^ n16075 ;
  assign n29563 = n15860 ^ n12257 ^ n10657 ;
  assign n29564 = ( x101 & ~n3972 ) | ( x101 & n23538 ) | ( ~n3972 & n23538 ) ;
  assign n29566 = n7224 ^ n6005 ^ n5379 ;
  assign n29565 = ~n6697 & n8085 ;
  assign n29567 = n29566 ^ n29565 ^ 1'b0 ;
  assign n29568 = n19190 ^ n10096 ^ 1'b0 ;
  assign n29569 = ( n3202 & ~n4718 ) | ( n3202 & n10644 ) | ( ~n4718 & n10644 ) ;
  assign n29570 = n29568 | n29569 ;
  assign n29571 = n20253 & n29570 ;
  assign n29572 = ~n29567 & n29571 ;
  assign n29573 = ( n1053 & ~n12583 ) | ( n1053 & n19079 ) | ( ~n12583 & n19079 ) ;
  assign n29574 = n29573 ^ n21043 ^ 1'b0 ;
  assign n29578 = n23553 ^ n19213 ^ n13535 ;
  assign n29579 = n14861 | n29578 ;
  assign n29580 = n29579 ^ n26368 ^ 1'b0 ;
  assign n29575 = ( n8959 & n13770 ) | ( n8959 & ~n18041 ) | ( n13770 & ~n18041 ) ;
  assign n29576 = ( ~n593 & n2186 ) | ( ~n593 & n28106 ) | ( n2186 & n28106 ) ;
  assign n29577 = ( n23225 & n29575 ) | ( n23225 & ~n29576 ) | ( n29575 & ~n29576 ) ;
  assign n29581 = n29580 ^ n29577 ^ n9793 ;
  assign n29582 = n7600 ^ n3903 ^ n1639 ;
  assign n29583 = n18180 & ~n29582 ;
  assign n29584 = n29583 ^ n9770 ^ 1'b0 ;
  assign n29587 = ( ~n1382 & n3130 ) | ( ~n1382 & n18301 ) | ( n3130 & n18301 ) ;
  assign n29585 = ( ~n685 & n3538 ) | ( ~n685 & n8171 ) | ( n3538 & n8171 ) ;
  assign n29586 = ( n13136 & n17627 ) | ( n13136 & n29585 ) | ( n17627 & n29585 ) ;
  assign n29588 = n29587 ^ n29586 ^ 1'b0 ;
  assign n29589 = ( n11792 & ~n27728 ) | ( n11792 & n29588 ) | ( ~n27728 & n29588 ) ;
  assign n29590 = ( n10649 & ~n16024 ) | ( n10649 & n20602 ) | ( ~n16024 & n20602 ) ;
  assign n29591 = n9370 | n25621 ;
  assign n29592 = n6332 | n10651 ;
  assign n29593 = n29591 | n29592 ;
  assign n29594 = n19945 ^ n3764 ^ 1'b0 ;
  assign n29595 = ( n7634 & n8641 ) | ( n7634 & n14847 ) | ( n8641 & n14847 ) ;
  assign n29596 = ( n878 & ~n4776 ) | ( n878 & n8268 ) | ( ~n4776 & n8268 ) ;
  assign n29597 = ( n19107 & n29536 ) | ( n19107 & ~n29596 ) | ( n29536 & ~n29596 ) ;
  assign n29598 = ( n9978 & n29595 ) | ( n9978 & n29597 ) | ( n29595 & n29597 ) ;
  assign n29599 = n3195 ^ n1258 ^ n1233 ;
  assign n29600 = n5740 | n28179 ;
  assign n29601 = n29600 ^ n26462 ^ 1'b0 ;
  assign n29602 = ( n5124 & ~n5865 ) | ( n5124 & n15136 ) | ( ~n5865 & n15136 ) ;
  assign n29603 = n29602 ^ n16465 ^ 1'b0 ;
  assign n29604 = n5439 & ~n29603 ;
  assign n29605 = x63 & n29604 ;
  assign n29606 = ( n945 & n15618 ) | ( n945 & ~n28437 ) | ( n15618 & ~n28437 ) ;
  assign n29607 = ( ~x244 & n1996 ) | ( ~x244 & n22796 ) | ( n1996 & n22796 ) ;
  assign n29608 = n23445 ^ n12944 ^ n7254 ;
  assign n29609 = ( n5262 & n29607 ) | ( n5262 & ~n29608 ) | ( n29607 & ~n29608 ) ;
  assign n29610 = n26889 ^ n24704 ^ n2969 ;
  assign n29612 = n26247 ^ n21859 ^ n12293 ;
  assign n29611 = n2841 & n23195 ;
  assign n29613 = n29612 ^ n29611 ^ 1'b0 ;
  assign n29614 = ( n19159 & n22285 ) | ( n19159 & ~n27598 ) | ( n22285 & ~n27598 ) ;
  assign n29615 = ( ~n16244 & n17797 ) | ( ~n16244 & n21919 ) | ( n17797 & n21919 ) ;
  assign n29616 = n29226 ^ n24663 ^ n1307 ;
  assign n29617 = ( n4135 & n7119 ) | ( n4135 & n8400 ) | ( n7119 & n8400 ) ;
  assign n29618 = n16236 ^ n4010 ^ n2341 ;
  assign n29619 = n29618 ^ n6508 ^ 1'b0 ;
  assign n29620 = ( n638 & ~n29617 ) | ( n638 & n29619 ) | ( ~n29617 & n29619 ) ;
  assign n29621 = ( n23644 & ~n29616 ) | ( n23644 & n29620 ) | ( ~n29616 & n29620 ) ;
  assign n29622 = n16150 ^ n8432 ^ n7296 ;
  assign n29623 = n12459 ^ n6437 ^ n1003 ;
  assign n29624 = ( n14008 & n29622 ) | ( n14008 & n29623 ) | ( n29622 & n29623 ) ;
  assign n29625 = ( n9197 & ~n28686 ) | ( n9197 & n29624 ) | ( ~n28686 & n29624 ) ;
  assign n29626 = ( ~n8915 & n18397 ) | ( ~n8915 & n29625 ) | ( n18397 & n29625 ) ;
  assign n29627 = ( ~n3630 & n5067 ) | ( ~n3630 & n23100 ) | ( n5067 & n23100 ) ;
  assign n29628 = n14868 ^ n11961 ^ 1'b0 ;
  assign n29629 = ~n25730 & n29628 ;
  assign n29630 = ( n13291 & ~n29627 ) | ( n13291 & n29629 ) | ( ~n29627 & n29629 ) ;
  assign n29631 = n13913 ^ n4917 ^ n3024 ;
  assign n29632 = n29631 ^ n22349 ^ n2214 ;
  assign n29633 = ( ~n1688 & n11073 ) | ( ~n1688 & n29632 ) | ( n11073 & n29632 ) ;
  assign n29634 = n9828 ^ n3266 ^ 1'b0 ;
  assign n29635 = ( n6284 & n20684 ) | ( n6284 & ~n21750 ) | ( n20684 & ~n21750 ) ;
  assign n29636 = ( n2258 & n10342 ) | ( n2258 & n19769 ) | ( n10342 & n19769 ) ;
  assign n29637 = n21537 ^ n18830 ^ n6454 ;
  assign n29638 = n29637 ^ n16179 ^ n15336 ;
  assign n29639 = n17111 ^ n5075 ^ 1'b0 ;
  assign n29640 = n14883 ^ n10044 ^ 1'b0 ;
  assign n29641 = n6540 & ~n29640 ;
  assign n29642 = ( n8233 & n18166 ) | ( n8233 & ~n29641 ) | ( n18166 & ~n29641 ) ;
  assign n29644 = ( n3773 & n4609 ) | ( n3773 & ~n7741 ) | ( n4609 & ~n7741 ) ;
  assign n29643 = n3661 & n26450 ;
  assign n29645 = n29644 ^ n29643 ^ 1'b0 ;
  assign n29646 = n29645 ^ n17362 ^ n10722 ;
  assign n29647 = n20272 ^ n14383 ^ n11831 ;
  assign n29648 = n20953 ^ n16091 ^ n6973 ;
  assign n29649 = ( ~n12940 & n18578 ) | ( ~n12940 & n22766 ) | ( n18578 & n22766 ) ;
  assign n29650 = n29649 ^ n12582 ^ n3160 ;
  assign n29652 = ( x152 & n1863 ) | ( x152 & ~n28864 ) | ( n1863 & ~n28864 ) ;
  assign n29651 = n26639 ^ n20351 ^ n17212 ;
  assign n29653 = n29652 ^ n29651 ^ n9650 ;
  assign n29654 = ( n13992 & n22467 ) | ( n13992 & n29653 ) | ( n22467 & n29653 ) ;
  assign n29655 = n29654 ^ n25859 ^ n705 ;
  assign n29656 = n22236 ^ x184 ^ 1'b0 ;
  assign n29657 = ( n18142 & n22622 ) | ( n18142 & n29656 ) | ( n22622 & n29656 ) ;
  assign n29658 = n17874 ^ n7031 ^ 1'b0 ;
  assign n29659 = n7818 ^ n505 ^ 1'b0 ;
  assign n29660 = n9048 | n29659 ;
  assign n29661 = ( n23176 & n29658 ) | ( n23176 & ~n29660 ) | ( n29658 & ~n29660 ) ;
  assign n29662 = n16668 ^ n5009 ^ n4986 ;
  assign n29663 = ( n17018 & ~n29661 ) | ( n17018 & n29662 ) | ( ~n29661 & n29662 ) ;
  assign n29664 = n18157 ^ n8390 ^ n4423 ;
  assign n29666 = n15157 ^ n11017 ^ n6885 ;
  assign n29665 = n428 ^ n297 ^ 1'b0 ;
  assign n29667 = n29666 ^ n29665 ^ n1388 ;
  assign n29668 = n19750 ^ n19532 ^ 1'b0 ;
  assign n29669 = n24017 | n29668 ;
  assign n29670 = n29669 ^ n23408 ^ n17994 ;
  assign n29674 = n19325 ^ n8835 ^ 1'b0 ;
  assign n29675 = n9218 & ~n29674 ;
  assign n29671 = ( n1149 & n10557 ) | ( n1149 & n16118 ) | ( n10557 & n16118 ) ;
  assign n29672 = ( n2532 & ~n5662 ) | ( n2532 & n29671 ) | ( ~n5662 & n29671 ) ;
  assign n29673 = n29672 ^ n26185 ^ 1'b0 ;
  assign n29676 = n29675 ^ n29673 ^ n6461 ;
  assign n29677 = ( n2258 & n9065 ) | ( n2258 & ~n18969 ) | ( n9065 & ~n18969 ) ;
  assign n29678 = n29677 ^ n11926 ^ n6309 ;
  assign n29679 = ( n5966 & n6468 ) | ( n5966 & n14242 ) | ( n6468 & n14242 ) ;
  assign n29683 = n9723 ^ n5695 ^ x125 ;
  assign n29684 = n29683 ^ n12643 ^ n9593 ;
  assign n29680 = ( n2555 & ~n14727 ) | ( n2555 & n17199 ) | ( ~n14727 & n17199 ) ;
  assign n29681 = n29680 ^ n21489 ^ n7279 ;
  assign n29682 = n29681 ^ n15118 ^ n13817 ;
  assign n29685 = n29684 ^ n29682 ^ n13622 ;
  assign n29686 = n978 & n5948 ;
  assign n29687 = ~n20537 & n29686 ;
  assign n29688 = n14648 ^ n4203 ^ 1'b0 ;
  assign n29689 = n10089 & n29688 ;
  assign n29690 = n27469 ^ n12896 ^ n3466 ;
  assign n29691 = n20917 ^ n12888 ^ n12551 ;
  assign n29692 = n9793 & ~n20931 ;
  assign n29693 = ( n15790 & n29691 ) | ( n15790 & n29692 ) | ( n29691 & n29692 ) ;
  assign n29694 = ( ~n7812 & n18183 ) | ( ~n7812 & n26894 ) | ( n18183 & n26894 ) ;
  assign n29697 = n16504 & n18333 ;
  assign n29698 = ~n12863 & n29697 ;
  assign n29695 = ( n902 & n3764 ) | ( n902 & n14274 ) | ( n3764 & n14274 ) ;
  assign n29696 = n7361 & ~n29695 ;
  assign n29699 = n29698 ^ n29696 ^ 1'b0 ;
  assign n29700 = ( n21266 & n29694 ) | ( n21266 & n29699 ) | ( n29694 & n29699 ) ;
  assign n29701 = n18101 ^ n13901 ^ n558 ;
  assign n29702 = ( n22236 & ~n29700 ) | ( n22236 & n29701 ) | ( ~n29700 & n29701 ) ;
  assign n29703 = ( ~n1475 & n17524 ) | ( ~n1475 & n23537 ) | ( n17524 & n23537 ) ;
  assign n29704 = n13841 ^ n5200 ^ n3694 ;
  assign n29705 = n1100 & ~n29704 ;
  assign n29706 = ~n20031 & n29705 ;
  assign n29707 = ( n8269 & n13319 ) | ( n8269 & n24182 ) | ( n13319 & n24182 ) ;
  assign n29708 = ( n24438 & n27252 ) | ( n24438 & ~n29707 ) | ( n27252 & ~n29707 ) ;
  assign n29709 = n29708 ^ n6676 ^ n3248 ;
  assign n29710 = n22303 ^ n18048 ^ n15488 ;
  assign n29711 = ( n2690 & n28766 ) | ( n2690 & n29710 ) | ( n28766 & n29710 ) ;
  assign n29712 = n10469 ^ n3952 ^ 1'b0 ;
  assign n29713 = x202 & ~n11482 ;
  assign n29714 = ~n18581 & n29713 ;
  assign n29718 = ( n4308 & ~n21681 ) | ( n4308 & n22323 ) | ( ~n21681 & n22323 ) ;
  assign n29716 = n29568 ^ n7921 ^ n6702 ;
  assign n29715 = ~n1963 & n7044 ;
  assign n29717 = n29716 ^ n29715 ^ 1'b0 ;
  assign n29719 = n29718 ^ n29717 ^ n24947 ;
  assign n29720 = n5659 ^ n2820 ^ 1'b0 ;
  assign n29721 = n29720 ^ n5545 ^ 1'b0 ;
  assign n29722 = ( n29714 & ~n29719 ) | ( n29714 & n29721 ) | ( ~n29719 & n29721 ) ;
  assign n29723 = n16262 ^ n7846 ^ n3084 ;
  assign n29724 = n21156 ^ n17463 ^ n3251 ;
  assign n29725 = n29724 ^ n16417 ^ 1'b0 ;
  assign n29726 = ( ~n733 & n10473 ) | ( ~n733 & n10546 ) | ( n10473 & n10546 ) ;
  assign n29727 = n13129 & ~n24634 ;
  assign n29728 = n23042 & n29727 ;
  assign n29729 = n21873 ^ n4986 ^ n3818 ;
  assign n29730 = n3773 ^ n1147 ^ 1'b0 ;
  assign n29731 = ( n11953 & n20379 ) | ( n11953 & n29730 ) | ( n20379 & n29730 ) ;
  assign n29732 = n28582 ^ n18695 ^ n2387 ;
  assign n29733 = ( n29729 & n29731 ) | ( n29729 & ~n29732 ) | ( n29731 & ~n29732 ) ;
  assign n29734 = n13579 ^ x214 ^ 1'b0 ;
  assign n29735 = ( n1935 & ~n1990 ) | ( n1935 & n7605 ) | ( ~n1990 & n7605 ) ;
  assign n29736 = n29735 ^ n5762 ^ n5351 ;
  assign n29737 = n29736 ^ n13915 ^ n13118 ;
  assign n29738 = ( x173 & n5442 ) | ( x173 & ~n29737 ) | ( n5442 & ~n29737 ) ;
  assign n29739 = ( ~n8842 & n29734 ) | ( ~n8842 & n29738 ) | ( n29734 & n29738 ) ;
  assign n29740 = n8299 ^ n5732 ^ 1'b0 ;
  assign n29741 = n28038 & n29740 ;
  assign n29742 = ( n11483 & n20113 ) | ( n11483 & n27766 ) | ( n20113 & n27766 ) ;
  assign n29743 = n29742 ^ n3544 ^ 1'b0 ;
  assign n29744 = ~n29741 & n29743 ;
  assign n29745 = ( n10302 & n17639 ) | ( n10302 & n19098 ) | ( n17639 & n19098 ) ;
  assign n29746 = n6694 ^ n719 ^ 1'b0 ;
  assign n29747 = n12323 | n29746 ;
  assign n29748 = n14991 ^ n13141 ^ n6479 ;
  assign n29749 = ( ~n27948 & n29747 ) | ( ~n27948 & n29748 ) | ( n29747 & n29748 ) ;
  assign n29750 = n20425 ^ n20017 ^ n16063 ;
  assign n29751 = ( n29745 & ~n29749 ) | ( n29745 & n29750 ) | ( ~n29749 & n29750 ) ;
  assign n29752 = n18602 ^ n5474 ^ n2768 ;
  assign n29753 = n29752 ^ n13536 ^ n11794 ;
  assign n29754 = n7231 ^ n4088 ^ n2564 ;
  assign n29755 = n10257 ^ n2432 ^ n1522 ;
  assign n29756 = ( n4986 & ~n29754 ) | ( n4986 & n29755 ) | ( ~n29754 & n29755 ) ;
  assign n29758 = n14724 ^ n12099 ^ n992 ;
  assign n29759 = n29758 ^ n12594 ^ n10398 ;
  assign n29757 = ( n13775 & n19134 ) | ( n13775 & n25410 ) | ( n19134 & n25410 ) ;
  assign n29760 = n29759 ^ n29757 ^ 1'b0 ;
  assign n29766 = n27885 ^ n21896 ^ n13567 ;
  assign n29761 = n2407 & n28988 ;
  assign n29762 = ~n3549 & n29761 ;
  assign n29763 = n6139 | n15074 ;
  assign n29764 = n29763 ^ n25290 ^ 1'b0 ;
  assign n29765 = ( n18125 & n29762 ) | ( n18125 & ~n29764 ) | ( n29762 & ~n29764 ) ;
  assign n29767 = n29766 ^ n29765 ^ n21180 ;
  assign n29768 = n11099 ^ n4437 ^ 1'b0 ;
  assign n29769 = n18929 & ~n29768 ;
  assign n29770 = n29769 ^ n19913 ^ n16587 ;
  assign n29771 = n29770 ^ n12407 ^ n3711 ;
  assign n29772 = ( ~n4369 & n4810 ) | ( ~n4369 & n6425 ) | ( n4810 & n6425 ) ;
  assign n29773 = n29772 ^ n25842 ^ n6351 ;
  assign n29774 = n29773 ^ n4910 ^ n1442 ;
  assign n29775 = n29774 ^ n17241 ^ n12623 ;
  assign n29776 = n29775 ^ n18780 ^ 1'b0 ;
  assign n29777 = n10357 & ~n29776 ;
  assign n29778 = ( n1355 & ~n2044 ) | ( n1355 & n23720 ) | ( ~n2044 & n23720 ) ;
  assign n29779 = ( ~n21106 & n26102 ) | ( ~n21106 & n29778 ) | ( n26102 & n29778 ) ;
  assign n29780 = ( n11821 & n24947 ) | ( n11821 & ~n29779 ) | ( n24947 & ~n29779 ) ;
  assign n29781 = n11128 ^ n1922 ^ 1'b0 ;
  assign n29782 = n7092 & n29781 ;
  assign n29783 = n29782 ^ n3567 ^ n1354 ;
  assign n29784 = ( n14822 & n21516 ) | ( n14822 & ~n29783 ) | ( n21516 & ~n29783 ) ;
  assign n29785 = n20343 ^ n18803 ^ n2106 ;
  assign n29786 = ( n2403 & n3490 ) | ( n2403 & n6398 ) | ( n3490 & n6398 ) ;
  assign n29787 = n18714 ^ n5339 ^ n3509 ;
  assign n29788 = n29787 ^ n11290 ^ n1741 ;
  assign n29789 = ( ~n16636 & n29786 ) | ( ~n16636 & n29788 ) | ( n29786 & n29788 ) ;
  assign n29790 = ( n3848 & n10194 ) | ( n3848 & ~n16796 ) | ( n10194 & ~n16796 ) ;
  assign n29791 = n29790 ^ n24108 ^ n5367 ;
  assign n29792 = ( n2292 & n29789 ) | ( n2292 & ~n29791 ) | ( n29789 & ~n29791 ) ;
  assign n29793 = ( n2809 & ~n4995 ) | ( n2809 & n29792 ) | ( ~n4995 & n29792 ) ;
  assign n29794 = ~n7655 & n7883 ;
  assign n29795 = ~n5649 & n29794 ;
  assign n29796 = n15343 | n29795 ;
  assign n29797 = n25594 & ~n29796 ;
  assign n29799 = ( n1180 & n1925 ) | ( n1180 & n25431 ) | ( n1925 & n25431 ) ;
  assign n29800 = ( n20511 & ~n25602 ) | ( n20511 & n29799 ) | ( ~n25602 & n29799 ) ;
  assign n29798 = n263 & n11113 ;
  assign n29801 = n29800 ^ n29798 ^ 1'b0 ;
  assign n29802 = n29801 ^ n11344 ^ n5688 ;
  assign n29803 = ( n7339 & n7363 ) | ( n7339 & ~n16569 ) | ( n7363 & ~n16569 ) ;
  assign n29804 = n6020 & ~n29803 ;
  assign n29805 = n29804 ^ n18270 ^ n3895 ;
  assign n29806 = n18428 ^ n8349 ^ n1963 ;
  assign n29807 = ( ~n22710 & n25372 ) | ( ~n22710 & n29806 ) | ( n25372 & n29806 ) ;
  assign n29808 = n22355 ^ n21794 ^ 1'b0 ;
  assign n29809 = n29808 ^ n15719 ^ n6763 ;
  assign n29810 = n29809 ^ n23611 ^ n3443 ;
  assign n29813 = ( n7002 & n16382 ) | ( n7002 & ~n25762 ) | ( n16382 & ~n25762 ) ;
  assign n29814 = n29813 ^ n25590 ^ n7584 ;
  assign n29811 = ( n273 & n4339 ) | ( n273 & n12285 ) | ( n4339 & n12285 ) ;
  assign n29812 = ~n7053 & n29811 ;
  assign n29815 = n29814 ^ n29812 ^ n19578 ;
  assign n29818 = ( n2714 & n16060 ) | ( n2714 & ~n17620 ) | ( n16060 & ~n17620 ) ;
  assign n29819 = n29818 ^ n18656 ^ 1'b0 ;
  assign n29817 = n4804 ^ n1687 ^ 1'b0 ;
  assign n29816 = ( ~n8555 & n12364 ) | ( ~n8555 & n16062 ) | ( n12364 & n16062 ) ;
  assign n29820 = n29819 ^ n29817 ^ n29816 ;
  assign n29821 = ~n8156 & n29820 ;
  assign n29822 = n29821 ^ n24916 ^ 1'b0 ;
  assign n29823 = n28425 ^ n15762 ^ n5804 ;
  assign n29824 = ( n3621 & n12401 ) | ( n3621 & n18156 ) | ( n12401 & n18156 ) ;
  assign n29826 = n11988 ^ n4322 ^ n874 ;
  assign n29825 = n14983 ^ n3989 ^ 1'b0 ;
  assign n29827 = n29826 ^ n29825 ^ n10746 ;
  assign n29828 = ( ~n11402 & n12952 ) | ( ~n11402 & n25562 ) | ( n12952 & n25562 ) ;
  assign n29829 = n29828 ^ n29215 ^ n5757 ;
  assign n29830 = ( n399 & ~n29827 ) | ( n399 & n29829 ) | ( ~n29827 & n29829 ) ;
  assign n29831 = n16095 & ~n23362 ;
  assign n29832 = ( ~n2803 & n9668 ) | ( ~n2803 & n12475 ) | ( n9668 & n12475 ) ;
  assign n29833 = n29832 ^ n12739 ^ 1'b0 ;
  assign n29834 = ( n1620 & n6580 ) | ( n1620 & n28755 ) | ( n6580 & n28755 ) ;
  assign n29843 = n18132 ^ n1304 ^ n1169 ;
  assign n29835 = ( n8920 & ~n13948 ) | ( n8920 & n28819 ) | ( ~n13948 & n28819 ) ;
  assign n29836 = n13509 ^ n7728 ^ n3410 ;
  assign n29837 = ( n2181 & n5075 ) | ( n2181 & n12103 ) | ( n5075 & n12103 ) ;
  assign n29838 = n29837 ^ n4060 ^ 1'b0 ;
  assign n29839 = ( n17264 & ~n29836 ) | ( n17264 & n29838 ) | ( ~n29836 & n29838 ) ;
  assign n29840 = n17057 & n29839 ;
  assign n29841 = ~n29835 & n29840 ;
  assign n29842 = n29841 ^ n22242 ^ n11634 ;
  assign n29844 = n29843 ^ n29842 ^ n14568 ;
  assign n29845 = n21082 ^ n15420 ^ n9622 ;
  assign n29846 = ~n604 & n12494 ;
  assign n29847 = n29846 ^ n3305 ^ 1'b0 ;
  assign n29848 = n29847 ^ n2675 ^ n1805 ;
  assign n29849 = ( n4400 & n5072 ) | ( n4400 & ~n29848 ) | ( n5072 & ~n29848 ) ;
  assign n29850 = n29845 & n29849 ;
  assign n29851 = ( n5076 & n6804 ) | ( n5076 & ~n20485 ) | ( n6804 & ~n20485 ) ;
  assign n29852 = ( ~n12130 & n13095 ) | ( ~n12130 & n29851 ) | ( n13095 & n29851 ) ;
  assign n29853 = n29852 ^ n2982 ^ n1726 ;
  assign n29854 = ( n29586 & n29850 ) | ( n29586 & n29853 ) | ( n29850 & n29853 ) ;
  assign n29855 = ( n3469 & ~n8390 ) | ( n3469 & n21568 ) | ( ~n8390 & n21568 ) ;
  assign n29856 = ( n8027 & n10793 ) | ( n8027 & ~n25459 ) | ( n10793 & ~n25459 ) ;
  assign n29857 = n18422 ^ n15151 ^ n5215 ;
  assign n29858 = ( ~n6079 & n29856 ) | ( ~n6079 & n29857 ) | ( n29856 & n29857 ) ;
  assign n29859 = n29858 ^ n17154 ^ n3024 ;
  assign n29860 = n28675 ^ n26972 ^ n5354 ;
  assign n29861 = n15591 & n28855 ;
  assign n29862 = ( n4133 & n29860 ) | ( n4133 & ~n29861 ) | ( n29860 & ~n29861 ) ;
  assign n29863 = ( n6340 & ~n6437 ) | ( n6340 & n14124 ) | ( ~n6437 & n14124 ) ;
  assign n29864 = ( ~n16239 & n23170 ) | ( ~n16239 & n29863 ) | ( n23170 & n29863 ) ;
  assign n29865 = ( ~n10135 & n15615 ) | ( ~n10135 & n20819 ) | ( n15615 & n20819 ) ;
  assign n29866 = n746 | n18462 ;
  assign n29867 = n773 & n29866 ;
  assign n29868 = n2129 & n3764 ;
  assign n29869 = n19173 & n29868 ;
  assign n29870 = ( ~n15255 & n23959 ) | ( ~n15255 & n26063 ) | ( n23959 & n26063 ) ;
  assign n29871 = n29870 ^ n21560 ^ n13962 ;
  assign n29872 = ( n4319 & n6045 ) | ( n4319 & n25907 ) | ( n6045 & n25907 ) ;
  assign n29873 = ( n9857 & n12375 ) | ( n9857 & n29872 ) | ( n12375 & n29872 ) ;
  assign n29874 = ( n1398 & n8834 ) | ( n1398 & n13304 ) | ( n8834 & n13304 ) ;
  assign n29875 = ( ~n15151 & n22598 ) | ( ~n15151 & n29874 ) | ( n22598 & n29874 ) ;
  assign n29876 = n3568 & n29875 ;
  assign n29877 = n29876 ^ n4954 ^ 1'b0 ;
  assign n29878 = n29877 ^ n23371 ^ n2802 ;
  assign n29879 = n707 & ~n19332 ;
  assign n29880 = n13725 & n29879 ;
  assign n29881 = n13696 ^ n11998 ^ 1'b0 ;
  assign n29882 = n4769 ^ n805 ^ 1'b0 ;
  assign n29883 = n29881 & n29882 ;
  assign n29884 = ( n3947 & n15762 ) | ( n3947 & n29883 ) | ( n15762 & n29883 ) ;
  assign n29885 = n12013 ^ n10452 ^ n7354 ;
  assign n29886 = ( n25122 & n29884 ) | ( n25122 & ~n29885 ) | ( n29884 & ~n29885 ) ;
  assign n29887 = n20025 ^ n17946 ^ n5502 ;
  assign n29888 = n28756 ^ n13219 ^ n308 ;
  assign n29889 = ( n4226 & n10707 ) | ( n4226 & ~n24723 ) | ( n10707 & ~n24723 ) ;
  assign n29890 = ( n7170 & ~n22215 ) | ( n7170 & n29889 ) | ( ~n22215 & n29889 ) ;
  assign n29893 = ( ~n626 & n12990 ) | ( ~n626 & n17045 ) | ( n12990 & n17045 ) ;
  assign n29891 = n15077 ^ n13489 ^ 1'b0 ;
  assign n29892 = n16764 & n29891 ;
  assign n29894 = n29893 ^ n29892 ^ x202 ;
  assign n29895 = n28592 ^ n20088 ^ n1192 ;
  assign n29896 = n12616 ^ n1730 ^ 1'b0 ;
  assign n29897 = ( n3467 & n4469 ) | ( n3467 & n9605 ) | ( n4469 & n9605 ) ;
  assign n29898 = n29897 ^ n8474 ^ n8305 ;
  assign n29899 = n13664 ^ n10115 ^ n1513 ;
  assign n29900 = n24053 & ~n29462 ;
  assign n29901 = n29900 ^ n25888 ^ 1'b0 ;
  assign n29902 = n27187 ^ n22449 ^ n2488 ;
  assign n29903 = n29714 ^ n18993 ^ n2827 ;
  assign n29904 = n27403 ^ n13507 ^ n3930 ;
  assign n29905 = n14320 & n29904 ;
  assign n29906 = n29905 ^ n7249 ^ 1'b0 ;
  assign n29907 = ( ~n10676 & n12413 ) | ( ~n10676 & n29906 ) | ( n12413 & n29906 ) ;
  assign n29910 = n7377 & n18842 ;
  assign n29911 = n29910 ^ n9840 ^ 1'b0 ;
  assign n29908 = ( n4304 & ~n14732 ) | ( n4304 & n29366 ) | ( ~n14732 & n29366 ) ;
  assign n29909 = n29908 ^ n18613 ^ n9866 ;
  assign n29912 = n29911 ^ n29909 ^ n4547 ;
  assign n29913 = ( ~n11552 & n26229 ) | ( ~n11552 & n29912 ) | ( n26229 & n29912 ) ;
  assign n29914 = ~n21310 & n22794 ;
  assign n29915 = ( ~n653 & n9608 ) | ( ~n653 & n12360 ) | ( n9608 & n12360 ) ;
  assign n29916 = n29915 ^ n15518 ^ n13659 ;
  assign n29917 = ( n2288 & n7302 ) | ( n2288 & n7649 ) | ( n7302 & n7649 ) ;
  assign n29918 = n26638 ^ n17150 ^ n14982 ;
  assign n29919 = ( n9565 & n23052 ) | ( n9565 & n29918 ) | ( n23052 & n29918 ) ;
  assign n29920 = n7325 & n8144 ;
  assign n29921 = ( ~n29917 & n29919 ) | ( ~n29917 & n29920 ) | ( n29919 & n29920 ) ;
  assign n29922 = n29921 ^ n26011 ^ n10424 ;
  assign n29923 = ( ~n1515 & n2036 ) | ( ~n1515 & n6315 ) | ( n2036 & n6315 ) ;
  assign n29924 = ( n9453 & ~n20297 ) | ( n9453 & n29923 ) | ( ~n20297 & n29923 ) ;
  assign n29925 = ( n12029 & n12842 ) | ( n12029 & n18906 ) | ( n12842 & n18906 ) ;
  assign n29926 = n25815 & ~n29925 ;
  assign n29927 = n29926 ^ n4594 ^ 1'b0 ;
  assign n29928 = n29296 ^ n21992 ^ n11785 ;
  assign n29929 = n29928 ^ n17992 ^ 1'b0 ;
  assign n29930 = n29927 & ~n29929 ;
  assign n29931 = ( n9502 & n18165 ) | ( n9502 & ~n19309 ) | ( n18165 & ~n19309 ) ;
  assign n29932 = n20847 ^ n12896 ^ n9047 ;
  assign n29933 = ( ~n15272 & n18492 ) | ( ~n15272 & n29932 ) | ( n18492 & n29932 ) ;
  assign n29934 = ~n4299 & n10148 ;
  assign n29935 = n4686 & n29934 ;
  assign n29936 = n19004 ^ n9662 ^ n6222 ;
  assign n29937 = ( ~n815 & n29935 ) | ( ~n815 & n29936 ) | ( n29935 & n29936 ) ;
  assign n29938 = n23839 ^ n20410 ^ n19965 ;
  assign n29939 = n11571 ^ n5203 ^ 1'b0 ;
  assign n29940 = n11344 | n29939 ;
  assign n29941 = n29940 ^ n27489 ^ n2020 ;
  assign n29942 = ( n6538 & n24329 ) | ( n6538 & ~n29941 ) | ( n24329 & ~n29941 ) ;
  assign n29943 = ( n7919 & n14991 ) | ( n7919 & n29942 ) | ( n14991 & n29942 ) ;
  assign n29945 = ( ~n5841 & n20485 ) | ( ~n5841 & n20688 ) | ( n20485 & n20688 ) ;
  assign n29946 = n5244 ^ n4389 ^ n4040 ;
  assign n29947 = ( n15984 & ~n29945 ) | ( n15984 & n29946 ) | ( ~n29945 & n29946 ) ;
  assign n29944 = n7907 & n23978 ;
  assign n29948 = n29947 ^ n29944 ^ 1'b0 ;
  assign n29950 = n19313 ^ n8988 ^ n4875 ;
  assign n29949 = n3059 | n5686 ;
  assign n29951 = n29950 ^ n29949 ^ 1'b0 ;
  assign n29952 = n21087 ^ n11816 ^ n8921 ;
  assign n29954 = n16786 ^ n2949 ^ x158 ;
  assign n29953 = ~n9010 & n18105 ;
  assign n29955 = n29954 ^ n29953 ^ n12882 ;
  assign n29956 = n21669 & ~n29955 ;
  assign n29957 = n29956 ^ n16483 ^ 1'b0 ;
  assign n29958 = ( n11034 & n29952 ) | ( n11034 & n29957 ) | ( n29952 & n29957 ) ;
  assign n29959 = n25296 ^ n17046 ^ n13948 ;
  assign n29960 = x245 & n899 ;
  assign n29961 = n10531 ^ n10391 ^ n8530 ;
  assign n29962 = n12852 ^ x234 ^ 1'b0 ;
  assign n29963 = n29961 | n29962 ;
  assign n29964 = n2978 ^ n2088 ^ x76 ;
  assign n29965 = ~n4031 & n4695 ;
  assign n29966 = ~n29964 & n29965 ;
  assign n29967 = ( n8777 & ~n18070 ) | ( n8777 & n29966 ) | ( ~n18070 & n29966 ) ;
  assign n29968 = ( ~n29960 & n29963 ) | ( ~n29960 & n29967 ) | ( n29963 & n29967 ) ;
  assign n29969 = ( n1627 & n28514 ) | ( n1627 & ~n29560 ) | ( n28514 & ~n29560 ) ;
  assign n29970 = ( n496 & ~n18142 ) | ( n496 & n27707 ) | ( ~n18142 & n27707 ) ;
  assign n29971 = ( n3864 & n10590 ) | ( n3864 & n18920 ) | ( n10590 & n18920 ) ;
  assign n29972 = n17228 ^ n5731 ^ 1'b0 ;
  assign n29973 = n19671 ^ n13399 ^ n11135 ;
  assign n29974 = n29973 ^ n16328 ^ 1'b0 ;
  assign n29975 = ~n29972 & n29974 ;
  assign n29976 = n2122 & n15846 ;
  assign n29977 = ~n1008 & n14518 ;
  assign n29978 = n5870 & n29977 ;
  assign n29979 = n29978 ^ n18259 ^ n14668 ;
  assign n29980 = n29587 ^ n27938 ^ n3182 ;
  assign n29981 = ( n29976 & n29979 ) | ( n29976 & n29980 ) | ( n29979 & n29980 ) ;
  assign n29982 = n17525 & ~n29841 ;
  assign n29983 = n4266 & n29982 ;
  assign n29984 = n23575 ^ n12948 ^ n9761 ;
  assign n29985 = n29984 ^ n17075 ^ x8 ;
  assign n29986 = n29786 ^ n6751 ^ 1'b0 ;
  assign n29987 = ~n585 & n28326 ;
  assign n29988 = ~n14903 & n29987 ;
  assign n29989 = ( ~n23202 & n29986 ) | ( ~n23202 & n29988 ) | ( n29986 & n29988 ) ;
  assign n29990 = ( n1919 & n5376 ) | ( n1919 & n8385 ) | ( n5376 & n8385 ) ;
  assign n29991 = ( n5573 & n11938 ) | ( n5573 & ~n17226 ) | ( n11938 & ~n17226 ) ;
  assign n29992 = ( ~n8186 & n12834 ) | ( ~n8186 & n29991 ) | ( n12834 & n29991 ) ;
  assign n29993 = x80 & ~n7371 ;
  assign n29994 = n29993 ^ n20533 ^ 1'b0 ;
  assign n29995 = ~n29992 & n29994 ;
  assign n29996 = n18868 ^ n13934 ^ n5695 ;
  assign n29997 = n7448 | n29996 ;
  assign n29998 = n29997 ^ n23271 ^ n16119 ;
  assign n29999 = ( n6145 & ~n26217 ) | ( n6145 & n29998 ) | ( ~n26217 & n29998 ) ;
  assign n30000 = n29999 ^ n26524 ^ n9036 ;
  assign n30001 = n24104 ^ n20148 ^ n9052 ;
  assign n30002 = ( n17924 & ~n18877 ) | ( n17924 & n30001 ) | ( ~n18877 & n30001 ) ;
  assign n30003 = n21579 ^ n19315 ^ n14394 ;
  assign n30005 = n28160 ^ n10198 ^ n302 ;
  assign n30006 = ( n5086 & ~n12540 ) | ( n5086 & n30005 ) | ( ~n12540 & n30005 ) ;
  assign n30004 = n18784 ^ n14104 ^ n2004 ;
  assign n30007 = n30006 ^ n30004 ^ n28191 ;
  assign n30009 = ( n3905 & n6321 ) | ( n3905 & n15803 ) | ( n6321 & n15803 ) ;
  assign n30008 = x179 & ~n18781 ;
  assign n30010 = n30009 ^ n30008 ^ 1'b0 ;
  assign n30014 = n5532 & ~n7967 ;
  assign n30012 = ( ~n5074 & n5778 ) | ( ~n5074 & n8937 ) | ( n5778 & n8937 ) ;
  assign n30013 = n30012 ^ n6319 ^ n3786 ;
  assign n30015 = n30014 ^ n30013 ^ n15007 ;
  assign n30011 = n14613 ^ n8329 ^ 1'b0 ;
  assign n30016 = n30015 ^ n30011 ^ n11965 ;
  assign n30017 = ( n9852 & ~n19344 ) | ( n9852 & n30016 ) | ( ~n19344 & n30016 ) ;
  assign n30018 = n27356 ^ n20094 ^ 1'b0 ;
  assign n30019 = n5514 & ~n30018 ;
  assign n30021 = n6211 ^ n650 ^ 1'b0 ;
  assign n30022 = n6812 & ~n30021 ;
  assign n30020 = n14290 | n15871 ;
  assign n30023 = n30022 ^ n30020 ^ 1'b0 ;
  assign n30024 = ( n2082 & n3950 ) | ( n2082 & ~n30023 ) | ( n3950 & ~n30023 ) ;
  assign n30025 = ( ~n25055 & n30019 ) | ( ~n25055 & n30024 ) | ( n30019 & n30024 ) ;
  assign n30026 = n30025 ^ n3356 ^ n1891 ;
  assign n30027 = n2410 | n10519 ;
  assign n30028 = ( n4852 & n7224 ) | ( n4852 & ~n17087 ) | ( n7224 & ~n17087 ) ;
  assign n30029 = ( n8611 & n30027 ) | ( n8611 & n30028 ) | ( n30027 & n30028 ) ;
  assign n30030 = ( n2042 & n2836 ) | ( n2042 & n15944 ) | ( n2836 & n15944 ) ;
  assign n30031 = ( n2152 & n23810 ) | ( n2152 & n30030 ) | ( n23810 & n30030 ) ;
  assign n30032 = n19960 ^ n16349 ^ n3995 ;
  assign n30033 = n4404 & n9105 ;
  assign n30034 = n30033 ^ n17788 ^ n11120 ;
  assign n30035 = n26354 ^ n13272 ^ n10772 ;
  assign n30036 = n20988 ^ n5268 ^ n301 ;
  assign n30037 = ( n8924 & n20913 ) | ( n8924 & ~n30036 ) | ( n20913 & ~n30036 ) ;
  assign n30038 = n25238 ^ n9626 ^ 1'b0 ;
  assign n30039 = n30038 ^ n11798 ^ n10689 ;
  assign n30040 = n30039 ^ n10389 ^ n2043 ;
  assign n30041 = n25367 ^ n8151 ^ 1'b0 ;
  assign n30042 = n30040 & n30041 ;
  assign n30043 = ( n8386 & n10405 ) | ( n8386 & ~n23931 ) | ( n10405 & ~n23931 ) ;
  assign n30047 = n29908 ^ n20070 ^ n7771 ;
  assign n30044 = n20104 ^ n19774 ^ n3224 ;
  assign n30045 = n30044 ^ n9849 ^ n2983 ;
  assign n30046 = ( n8474 & ~n24199 ) | ( n8474 & n30045 ) | ( ~n24199 & n30045 ) ;
  assign n30048 = n30047 ^ n30046 ^ 1'b0 ;
  assign n30049 = n25222 ^ n9441 ^ n8052 ;
  assign n30050 = n30049 ^ n28574 ^ n18386 ;
  assign n30051 = n30050 ^ n6664 ^ 1'b0 ;
  assign n30052 = ~n25101 & n30051 ;
  assign n30053 = ( n2477 & n4933 ) | ( n2477 & n14316 ) | ( n4933 & n14316 ) ;
  assign n30054 = ( n2962 & n13113 ) | ( n2962 & n30053 ) | ( n13113 & n30053 ) ;
  assign n30055 = ( ~n16976 & n22063 ) | ( ~n16976 & n30054 ) | ( n22063 & n30054 ) ;
  assign n30056 = ( n2479 & n30052 ) | ( n2479 & n30055 ) | ( n30052 & n30055 ) ;
  assign n30057 = n18931 & n30056 ;
  assign n30059 = n7607 ^ n7487 ^ n6303 ;
  assign n30058 = ~n1186 & n16666 ;
  assign n30060 = n30059 ^ n30058 ^ 1'b0 ;
  assign n30061 = ( n628 & n2163 ) | ( n628 & n25254 ) | ( n2163 & n25254 ) ;
  assign n30062 = n27012 ^ n7108 ^ n6674 ;
  assign n30065 = n4890 & ~n7772 ;
  assign n30063 = ( ~n5225 & n7138 ) | ( ~n5225 & n19974 ) | ( n7138 & n19974 ) ;
  assign n30064 = n30063 ^ n13983 ^ n6535 ;
  assign n30066 = n30065 ^ n30064 ^ n13812 ;
  assign n30067 = n8426 | n30066 ;
  assign n30068 = n16053 ^ n11992 ^ n8815 ;
  assign n30069 = ~n24178 & n26674 ;
  assign n30070 = n16374 & n30069 ;
  assign n30071 = n30070 ^ n19491 ^ n14324 ;
  assign n30072 = ( ~n17236 & n22430 ) | ( ~n17236 & n30071 ) | ( n22430 & n30071 ) ;
  assign n30073 = ( n11908 & n24060 ) | ( n11908 & ~n30072 ) | ( n24060 & ~n30072 ) ;
  assign n30075 = n2944 & ~n3409 ;
  assign n30074 = n20424 ^ n13039 ^ n2065 ;
  assign n30076 = n30075 ^ n30074 ^ n601 ;
  assign n30077 = n30076 ^ n8732 ^ n6126 ;
  assign n30080 = ( n6900 & n15036 ) | ( n6900 & n27031 ) | ( n15036 & n27031 ) ;
  assign n30081 = n30080 ^ n15002 ^ n6399 ;
  assign n30082 = ~n14876 & n19733 ;
  assign n30083 = ~n30081 & n30082 ;
  assign n30078 = ( n462 & ~n2298 ) | ( n462 & n5045 ) | ( ~n2298 & n5045 ) ;
  assign n30079 = ( n3045 & n10784 ) | ( n3045 & ~n30078 ) | ( n10784 & ~n30078 ) ;
  assign n30084 = n30083 ^ n30079 ^ n8260 ;
  assign n30085 = ( n9253 & n20251 ) | ( n9253 & ~n30084 ) | ( n20251 & ~n30084 ) ;
  assign n30086 = n25039 ^ n22416 ^ n13785 ;
  assign n30087 = n11619 ^ n8858 ^ n3720 ;
  assign n30088 = ( n4439 & ~n6446 ) | ( n4439 & n25207 ) | ( ~n6446 & n25207 ) ;
  assign n30089 = n16133 ^ n1762 ^ n1236 ;
  assign n30090 = n30089 ^ n8384 ^ n6132 ;
  assign n30091 = n12533 ^ n6711 ^ n2475 ;
  assign n30092 = ( n4170 & n8377 ) | ( n4170 & ~n22153 ) | ( n8377 & ~n22153 ) ;
  assign n30093 = ( n3580 & ~n5699 ) | ( n3580 & n30092 ) | ( ~n5699 & n30092 ) ;
  assign n30094 = ( n7799 & n30091 ) | ( n7799 & n30093 ) | ( n30091 & n30093 ) ;
  assign n30095 = ( n12079 & n15812 ) | ( n12079 & n30094 ) | ( n15812 & n30094 ) ;
  assign n30096 = ( n8886 & n13461 ) | ( n8886 & ~n30095 ) | ( n13461 & ~n30095 ) ;
  assign n30097 = n30090 & n30096 ;
  assign n30098 = n30097 ^ n20143 ^ 1'b0 ;
  assign n30099 = n18696 ^ n9823 ^ 1'b0 ;
  assign n30100 = ( n9182 & ~n11898 ) | ( n9182 & n30099 ) | ( ~n11898 & n30099 ) ;
  assign n30103 = n4525 | n22596 ;
  assign n30101 = n9336 & ~n24016 ;
  assign n30102 = ~n8586 & n30101 ;
  assign n30104 = n30103 ^ n30102 ^ n29695 ;
  assign n30105 = ( n938 & n14519 ) | ( n938 & ~n30104 ) | ( n14519 & ~n30104 ) ;
  assign n30106 = n30105 ^ n3100 ^ 1'b0 ;
  assign n30107 = n30106 ^ n16016 ^ n15654 ;
  assign n30108 = ~n10357 & n30107 ;
  assign n30109 = n15349 ^ n14848 ^ 1'b0 ;
  assign n30110 = ~n17023 & n30109 ;
  assign n30111 = n22615 ^ n20144 ^ n12090 ;
  assign n30112 = n30111 ^ n29419 ^ 1'b0 ;
  assign n30113 = n496 | n30112 ;
  assign n30114 = n30113 ^ n29208 ^ n8805 ;
  assign n30115 = n30110 & n30114 ;
  assign n30116 = n15492 ^ n11102 ^ n6928 ;
  assign n30117 = n7546 ^ n4503 ^ x103 ;
  assign n30118 = n30117 ^ n9578 ^ n7736 ;
  assign n30119 = n30118 ^ n12776 ^ 1'b0 ;
  assign n30120 = n30116 | n30119 ;
  assign n30121 = ( n12064 & n19740 ) | ( n12064 & n30120 ) | ( n19740 & n30120 ) ;
  assign n30122 = n16670 ^ n5346 ^ x205 ;
  assign n30123 = ( ~n11113 & n27218 ) | ( ~n11113 & n28467 ) | ( n27218 & n28467 ) ;
  assign n30124 = n30123 ^ n15487 ^ n781 ;
  assign n30125 = n30083 ^ n19627 ^ n2098 ;
  assign n30126 = ( n3968 & n17816 ) | ( n3968 & n18328 ) | ( n17816 & n18328 ) ;
  assign n30134 = ( ~n6121 & n9381 ) | ( ~n6121 & n23263 ) | ( n9381 & n23263 ) ;
  assign n30131 = n13669 ^ n8123 ^ n6069 ;
  assign n30132 = n30131 ^ n10034 ^ n5593 ;
  assign n30133 = n17923 & ~n30132 ;
  assign n30135 = n30134 ^ n30133 ^ n1984 ;
  assign n30127 = n11382 ^ n4261 ^ n1919 ;
  assign n30128 = n30127 ^ n19853 ^ 1'b0 ;
  assign n30129 = n27589 & ~n30128 ;
  assign n30130 = n30129 ^ n22999 ^ n9584 ;
  assign n30136 = n30135 ^ n30130 ^ n1056 ;
  assign n30139 = ( n1214 & ~n3058 ) | ( n1214 & n8231 ) | ( ~n3058 & n8231 ) ;
  assign n30140 = n3950 & ~n30139 ;
  assign n30141 = n12878 & n30140 ;
  assign n30137 = ( n21545 & n22181 ) | ( n21545 & n28579 ) | ( n22181 & n28579 ) ;
  assign n30138 = ( n11736 & n25678 ) | ( n11736 & n30137 ) | ( n25678 & n30137 ) ;
  assign n30142 = n30141 ^ n30138 ^ n17231 ;
  assign n30143 = ( n2875 & n12457 ) | ( n2875 & ~n15192 ) | ( n12457 & ~n15192 ) ;
  assign n30144 = n30143 ^ n1385 ^ n812 ;
  assign n30145 = n15224 ^ n11879 ^ 1'b0 ;
  assign n30146 = n24550 & ~n30145 ;
  assign n30147 = ( n5131 & n7460 ) | ( n5131 & n27568 ) | ( n7460 & n27568 ) ;
  assign n30148 = n30147 ^ n11422 ^ n8302 ;
  assign n30149 = ( n20485 & n25412 ) | ( n20485 & ~n30148 ) | ( n25412 & ~n30148 ) ;
  assign n30150 = n9985 ^ n8774 ^ 1'b0 ;
  assign n30151 = n1536 & n30150 ;
  assign n30152 = n30151 ^ n5656 ^ n2828 ;
  assign n30153 = ( ~n6496 & n25692 ) | ( ~n6496 & n30152 ) | ( n25692 & n30152 ) ;
  assign n30155 = n5204 ^ n3510 ^ n618 ;
  assign n30156 = n15439 ^ n15189 ^ 1'b0 ;
  assign n30157 = ( n22320 & ~n30155 ) | ( n22320 & n30156 ) | ( ~n30155 & n30156 ) ;
  assign n30154 = n15420 ^ n7628 ^ n1561 ;
  assign n30158 = n30157 ^ n30154 ^ n6062 ;
  assign n30159 = n30158 ^ n16899 ^ n13769 ;
  assign n30162 = n18023 ^ n5883 ^ n4226 ;
  assign n30160 = ( ~n2080 & n4953 ) | ( ~n2080 & n16855 ) | ( n4953 & n16855 ) ;
  assign n30161 = n30160 ^ n29954 ^ n13551 ;
  assign n30163 = n30162 ^ n30161 ^ n17057 ;
  assign n30164 = ( n13204 & ~n28840 ) | ( n13204 & n30163 ) | ( ~n28840 & n30163 ) ;
  assign n30165 = ( n17602 & ~n24358 ) | ( n17602 & n25738 ) | ( ~n24358 & n25738 ) ;
  assign n30166 = ( n1546 & ~n16092 ) | ( n1546 & n17949 ) | ( ~n16092 & n17949 ) ;
  assign n30168 = n7072 ^ n4071 ^ n1929 ;
  assign n30167 = n1645 ^ n1149 ^ n984 ;
  assign n30169 = n30168 ^ n30167 ^ n19065 ;
  assign n30170 = n30169 ^ n17882 ^ n3105 ;
  assign n30171 = n30170 ^ n11559 ^ n2751 ;
  assign n30172 = ( ~n25212 & n30166 ) | ( ~n25212 & n30171 ) | ( n30166 & n30171 ) ;
  assign n30173 = n9213 & n30172 ;
  assign n30174 = n3306 & n30173 ;
  assign n30175 = n8738 ^ n7989 ^ 1'b0 ;
  assign n30176 = n26989 ^ n10251 ^ n8095 ;
  assign n30177 = ( n784 & n7845 ) | ( n784 & n18990 ) | ( n7845 & n18990 ) ;
  assign n30178 = ( n905 & ~n15085 ) | ( n905 & n30177 ) | ( ~n15085 & n30177 ) ;
  assign n30179 = ( n2484 & ~n15767 ) | ( n2484 & n30178 ) | ( ~n15767 & n30178 ) ;
  assign n30180 = n17135 ^ n14324 ^ n7592 ;
  assign n30181 = ( ~n4444 & n10636 ) | ( ~n4444 & n30180 ) | ( n10636 & n30180 ) ;
  assign n30182 = n10689 & n24430 ;
  assign n30183 = n7847 & ~n26229 ;
  assign n30184 = n30183 ^ n27895 ^ 1'b0 ;
  assign n30185 = ~n14704 & n30184 ;
  assign n30186 = n30182 & n30185 ;
  assign n30187 = n18719 ^ n16272 ^ 1'b0 ;
  assign n30188 = n13129 & n30187 ;
  assign n30190 = n14887 ^ n9515 ^ x109 ;
  assign n30189 = n17631 ^ n8030 ^ n5455 ;
  assign n30191 = n30190 ^ n30189 ^ n19081 ;
  assign n30192 = ( n22365 & n28575 ) | ( n22365 & n30191 ) | ( n28575 & n30191 ) ;
  assign n30199 = n22510 ^ n22275 ^ n14868 ;
  assign n30193 = n8333 | n14240 ;
  assign n30194 = n30193 ^ n26208 ^ 1'b0 ;
  assign n30195 = n30194 ^ n1461 ^ 1'b0 ;
  assign n30196 = n3480 | n30195 ;
  assign n30197 = n30196 ^ n10886 ^ 1'b0 ;
  assign n30198 = ( ~n11431 & n16793 ) | ( ~n11431 & n30197 ) | ( n16793 & n30197 ) ;
  assign n30200 = n30199 ^ n30198 ^ n4196 ;
  assign n30201 = n30200 ^ n7720 ^ n5044 ;
  assign n30202 = ( n1343 & n1767 ) | ( n1343 & ~n17022 ) | ( n1767 & ~n17022 ) ;
  assign n30203 = n30016 ^ n9969 ^ n6128 ;
  assign n30204 = n28884 ^ n12247 ^ n5515 ;
  assign n30205 = n30204 ^ n23084 ^ n944 ;
  assign n30206 = ( ~n30202 & n30203 ) | ( ~n30202 & n30205 ) | ( n30203 & n30205 ) ;
  assign n30207 = ( n8281 & ~n12084 ) | ( n8281 & n12479 ) | ( ~n12084 & n12479 ) ;
  assign n30208 = n17043 ^ n4994 ^ 1'b0 ;
  assign n30209 = ~n30207 & n30208 ;
  assign n30210 = ( n5308 & n24995 ) | ( n5308 & n30209 ) | ( n24995 & n30209 ) ;
  assign n30211 = n30210 ^ n16528 ^ n12161 ;
  assign n30212 = n8835 & n26725 ;
  assign n30213 = n30212 ^ n27480 ^ n13492 ;
  assign n30214 = ( n3643 & ~n25206 ) | ( n3643 & n28613 ) | ( ~n25206 & n28613 ) ;
  assign n30216 = n2571 | n19527 ;
  assign n30215 = ( n5764 & n8748 ) | ( n5764 & n15177 ) | ( n8748 & n15177 ) ;
  assign n30217 = n30216 ^ n30215 ^ n27533 ;
  assign n30218 = ( n30213 & n30214 ) | ( n30213 & ~n30217 ) | ( n30214 & ~n30217 ) ;
  assign n30219 = ( n2139 & ~n3588 ) | ( n2139 & n28468 ) | ( ~n3588 & n28468 ) ;
  assign n30220 = n11473 ^ n11252 ^ n10230 ;
  assign n30221 = n18773 ^ n10407 ^ n810 ;
  assign n30222 = ( n2476 & n30220 ) | ( n2476 & n30221 ) | ( n30220 & n30221 ) ;
  assign n30223 = n30222 ^ n12266 ^ 1'b0 ;
  assign n30224 = n19506 & n30223 ;
  assign n30225 = n28424 ^ n1402 ^ 1'b0 ;
  assign n30226 = ( ~n3123 & n11538 ) | ( ~n3123 & n29825 ) | ( n11538 & n29825 ) ;
  assign n30227 = n30225 & n30226 ;
  assign n30228 = n30227 ^ n9445 ^ n4435 ;
  assign n30229 = n8843 & ~n16035 ;
  assign n30230 = n30229 ^ n3528 ^ 1'b0 ;
  assign n30231 = ( n266 & n9119 ) | ( n266 & n30230 ) | ( n9119 & n30230 ) ;
  assign n30232 = ( n5639 & n9362 ) | ( n5639 & ~n30231 ) | ( n9362 & ~n30231 ) ;
  assign n30233 = n30232 ^ n17313 ^ n17271 ;
  assign n30234 = n21898 ^ n18628 ^ n17627 ;
  assign n30235 = ( n14765 & n26053 ) | ( n14765 & ~n30234 ) | ( n26053 & ~n30234 ) ;
  assign n30236 = n19340 ^ n4427 ^ n2397 ;
  assign n30237 = ( ~n12558 & n14700 ) | ( ~n12558 & n20201 ) | ( n14700 & n20201 ) ;
  assign n30238 = ( n2875 & n3509 ) | ( n2875 & ~n6873 ) | ( n3509 & ~n6873 ) ;
  assign n30239 = ( n1472 & n22625 ) | ( n1472 & ~n24115 ) | ( n22625 & ~n24115 ) ;
  assign n30240 = n10019 ^ n6000 ^ n3731 ;
  assign n30241 = n30240 ^ n22615 ^ n13457 ;
  assign n30242 = ( n12070 & ~n18471 ) | ( n12070 & n30241 ) | ( ~n18471 & n30241 ) ;
  assign n30244 = n11436 ^ n9121 ^ 1'b0 ;
  assign n30245 = n1178 | n30244 ;
  assign n30243 = n7720 & n22795 ;
  assign n30246 = n30245 ^ n30243 ^ 1'b0 ;
  assign n30247 = n23856 ^ n18933 ^ n1214 ;
  assign n30248 = ~n14336 & n26014 ;
  assign n30249 = n30247 & n30248 ;
  assign n30250 = n18625 & ~n28085 ;
  assign n30254 = n3448 ^ n819 ^ 1'b0 ;
  assign n30253 = ~n1714 & n5165 ;
  assign n30255 = n30254 ^ n30253 ^ n20410 ;
  assign n30251 = ( ~n3074 & n3805 ) | ( ~n3074 & n16907 ) | ( n3805 & n16907 ) ;
  assign n30252 = n30251 ^ n17061 ^ n13519 ;
  assign n30256 = n30255 ^ n30252 ^ n6979 ;
  assign n30257 = ( n6029 & ~n13415 ) | ( n6029 & n15876 ) | ( ~n13415 & n15876 ) ;
  assign n30259 = n25366 ^ n5317 ^ n746 ;
  assign n30258 = ( n19623 & n24830 ) | ( n19623 & ~n26461 ) | ( n24830 & ~n26461 ) ;
  assign n30260 = n30259 ^ n30258 ^ n23274 ;
  assign n30261 = ( n14653 & n27878 ) | ( n14653 & n30260 ) | ( n27878 & n30260 ) ;
  assign n30262 = n30261 ^ n27433 ^ n17442 ;
  assign n30263 = n6049 ^ n5165 ^ 1'b0 ;
  assign n30264 = ~n5369 & n30263 ;
  assign n30265 = n30264 ^ n13772 ^ 1'b0 ;
  assign n30266 = n20796 | n23505 ;
  assign n30267 = n30265 | n30266 ;
  assign n30268 = ( ~n1155 & n19036 ) | ( ~n1155 & n30267 ) | ( n19036 & n30267 ) ;
  assign n30269 = n16899 & n30268 ;
  assign n30270 = n22413 & n30269 ;
  assign n30271 = n20346 ^ n4787 ^ 1'b0 ;
  assign n30272 = n28391 & n30271 ;
  assign n30273 = ( n2165 & n17394 ) | ( n2165 & ~n19198 ) | ( n17394 & ~n19198 ) ;
  assign n30275 = n23521 ^ n22160 ^ n12913 ;
  assign n30276 = n30275 ^ n28238 ^ n21076 ;
  assign n30274 = n10991 ^ n7303 ^ n2390 ;
  assign n30277 = n30276 ^ n30274 ^ n15862 ;
  assign n30278 = n25692 ^ n18617 ^ 1'b0 ;
  assign n30279 = n26822 ^ n26450 ^ n1377 ;
  assign n30280 = n5093 ^ x26 ^ 1'b0 ;
  assign n30281 = n16799 ^ n7049 ^ n3157 ;
  assign n30282 = ( n13554 & ~n30280 ) | ( n13554 & n30281 ) | ( ~n30280 & n30281 ) ;
  assign n30283 = n12782 ^ n1282 ^ n744 ;
  assign n30284 = n10993 & n20538 ;
  assign n30285 = n30284 ^ n11257 ^ 1'b0 ;
  assign n30286 = ( ~n23102 & n30283 ) | ( ~n23102 & n30285 ) | ( n30283 & n30285 ) ;
  assign n30287 = ( n11030 & n25282 ) | ( n11030 & ~n30286 ) | ( n25282 & ~n30286 ) ;
  assign n30288 = ( n7264 & ~n30282 ) | ( n7264 & n30287 ) | ( ~n30282 & n30287 ) ;
  assign n30289 = n18670 ^ n12171 ^ n9497 ;
  assign n30290 = n30289 ^ n28405 ^ 1'b0 ;
  assign n30291 = n25713 ^ n22098 ^ 1'b0 ;
  assign n30292 = ( n11327 & n30290 ) | ( n11327 & ~n30291 ) | ( n30290 & ~n30291 ) ;
  assign n30293 = ( ~n10150 & n13252 ) | ( ~n10150 & n30292 ) | ( n13252 & n30292 ) ;
  assign n30294 = n1235 & ~n11688 ;
  assign n30295 = n16608 & n30294 ;
  assign n30296 = n4174 ^ n3664 ^ n1023 ;
  assign n30297 = n30296 ^ n10702 ^ n3070 ;
  assign n30298 = ( n11475 & n15564 ) | ( n11475 & n30297 ) | ( n15564 & n30297 ) ;
  assign n30299 = n23707 ^ n16565 ^ 1'b0 ;
  assign n30300 = ( n10372 & n13984 ) | ( n10372 & n30299 ) | ( n13984 & n30299 ) ;
  assign n30301 = n30298 | n30300 ;
  assign n30302 = ( n14707 & n19212 ) | ( n14707 & ~n30301 ) | ( n19212 & ~n30301 ) ;
  assign n30303 = n26836 ^ n9865 ^ n4498 ;
  assign n30304 = ( n3712 & ~n10376 ) | ( n3712 & n26669 ) | ( ~n10376 & n26669 ) ;
  assign n30305 = ( n4551 & n24563 ) | ( n4551 & n30304 ) | ( n24563 & n30304 ) ;
  assign n30306 = ( n3284 & n4236 ) | ( n3284 & n30305 ) | ( n4236 & n30305 ) ;
  assign n30307 = n30306 ^ n24177 ^ n3870 ;
  assign n30308 = n23873 ^ n10083 ^ n4927 ;
  assign n30309 = ( ~n3968 & n20815 ) | ( ~n3968 & n30308 ) | ( n20815 & n30308 ) ;
  assign n30310 = n30309 ^ n28281 ^ n19721 ;
  assign n30311 = n17110 ^ n8609 ^ 1'b0 ;
  assign n30312 = n15647 & n30311 ;
  assign n30313 = ( n5578 & n15141 ) | ( n5578 & ~n30312 ) | ( n15141 & ~n30312 ) ;
  assign n30314 = n26763 ^ n25145 ^ n1175 ;
  assign n30319 = n14731 ^ n12843 ^ n11580 ;
  assign n30315 = n8500 ^ n3092 ^ 1'b0 ;
  assign n30316 = ( n855 & n16771 ) | ( n855 & n20210 ) | ( n16771 & n20210 ) ;
  assign n30317 = ( n8369 & ~n30315 ) | ( n8369 & n30316 ) | ( ~n30315 & n30316 ) ;
  assign n30318 = x170 & n30317 ;
  assign n30320 = n30319 ^ n30318 ^ 1'b0 ;
  assign n30321 = n22365 ^ n11374 ^ n6717 ;
  assign n30322 = ( ~n5201 & n6810 ) | ( ~n5201 & n30321 ) | ( n6810 & n30321 ) ;
  assign n30323 = n21922 ^ n11809 ^ n8891 ;
  assign n30324 = ( n10060 & n13705 ) | ( n10060 & n14896 ) | ( n13705 & n14896 ) ;
  assign n30325 = ( ~n8029 & n16624 ) | ( ~n8029 & n30324 ) | ( n16624 & n30324 ) ;
  assign n30326 = ( n4549 & n13190 ) | ( n4549 & ~n19312 ) | ( n13190 & ~n19312 ) ;
  assign n30328 = n4460 & ~n14808 ;
  assign n30329 = n30328 ^ n15676 ^ 1'b0 ;
  assign n30327 = ( n3487 & ~n3964 ) | ( n3487 & n6567 ) | ( ~n3964 & n6567 ) ;
  assign n30330 = n30329 ^ n30327 ^ n27157 ;
  assign n30331 = n24251 & n25639 ;
  assign n30332 = ( n22024 & n25112 ) | ( n22024 & ~n28339 ) | ( n25112 & ~n28339 ) ;
  assign n30333 = n21547 ^ n20163 ^ 1'b0 ;
  assign n30334 = ( n4097 & n18292 ) | ( n4097 & n30333 ) | ( n18292 & n30333 ) ;
  assign n30335 = n24872 ^ n5996 ^ n3072 ;
  assign n30336 = n24733 & n30335 ;
  assign n30337 = ( n851 & n1650 ) | ( n851 & ~n13147 ) | ( n1650 & ~n13147 ) ;
  assign n30338 = n24442 ^ n4817 ^ n1901 ;
  assign n30339 = ( n601 & n8090 ) | ( n601 & ~n30338 ) | ( n8090 & ~n30338 ) ;
  assign n30340 = n30339 ^ n20293 ^ n5598 ;
  assign n30341 = n8895 | n30340 ;
  assign n30342 = n30337 & ~n30341 ;
  assign n30343 = n1628 | n16623 ;
  assign n30344 = n30343 ^ n12989 ^ n10168 ;
  assign n30346 = ( n9054 & n13162 ) | ( n9054 & ~n18820 ) | ( n13162 & ~n18820 ) ;
  assign n30347 = n30346 ^ n23487 ^ n12183 ;
  assign n30345 = n22974 ^ n11721 ^ n987 ;
  assign n30348 = n30347 ^ n30345 ^ n29772 ;
  assign n30351 = ( n6743 & ~n6763 ) | ( n6743 & n23991 ) | ( ~n6763 & n23991 ) ;
  assign n30352 = n3855 | n7938 ;
  assign n30353 = n30351 & ~n30352 ;
  assign n30354 = n30353 ^ n17808 ^ n8897 ;
  assign n30350 = ( n3636 & n5286 ) | ( n3636 & n14042 ) | ( n5286 & n14042 ) ;
  assign n30349 = n16329 ^ n16169 ^ n13592 ;
  assign n30355 = n30354 ^ n30350 ^ n30349 ;
  assign n30356 = n15895 ^ n991 ^ 1'b0 ;
  assign n30359 = n17309 ^ n11834 ^ n5944 ;
  assign n30357 = n20503 ^ n10447 ^ n5209 ;
  assign n30358 = ( n4584 & ~n19490 ) | ( n4584 & n30357 ) | ( ~n19490 & n30357 ) ;
  assign n30360 = n30359 ^ n30358 ^ n13740 ;
  assign n30361 = n16114 ^ n2846 ^ 1'b0 ;
  assign n30362 = ~n8646 & n30361 ;
  assign n30363 = n13665 ^ n8655 ^ 1'b0 ;
  assign n30364 = n30362 & n30363 ;
  assign n30365 = n30364 ^ n19530 ^ n13430 ;
  assign n30366 = ( n14159 & n17735 ) | ( n14159 & n30365 ) | ( n17735 & n30365 ) ;
  assign n30367 = n13837 | n18172 ;
  assign n30368 = n30367 ^ n29745 ^ n3002 ;
  assign n30369 = ( n15474 & n22406 ) | ( n15474 & ~n30368 ) | ( n22406 & ~n30368 ) ;
  assign n30370 = ( ~n5403 & n7085 ) | ( ~n5403 & n8564 ) | ( n7085 & n8564 ) ;
  assign n30371 = n18402 ^ n10565 ^ 1'b0 ;
  assign n30372 = n30371 ^ n25823 ^ 1'b0 ;
  assign n30373 = n30370 | n30372 ;
  assign n30374 = ( n2422 & n10263 ) | ( n2422 & ~n30353 ) | ( n10263 & ~n30353 ) ;
  assign n30375 = n30374 ^ n14871 ^ n10763 ;
  assign n30376 = ( n12884 & ~n20762 ) | ( n12884 & n30375 ) | ( ~n20762 & n30375 ) ;
  assign n30377 = n30376 ^ n14085 ^ 1'b0 ;
  assign n30378 = ( x178 & n7685 ) | ( x178 & ~n7847 ) | ( n7685 & ~n7847 ) ;
  assign n30379 = ( ~n4604 & n5769 ) | ( ~n4604 & n30378 ) | ( n5769 & n30378 ) ;
  assign n30380 = ~n8451 & n23181 ;
  assign n30381 = ( ~n5041 & n14821 ) | ( ~n5041 & n15593 ) | ( n14821 & n15593 ) ;
  assign n30384 = n18051 ^ n13557 ^ n3808 ;
  assign n30382 = n21468 ^ n5235 ^ n1517 ;
  assign n30383 = ( n8914 & n15113 ) | ( n8914 & ~n30382 ) | ( n15113 & ~n30382 ) ;
  assign n30385 = n30384 ^ n30383 ^ n25216 ;
  assign n30386 = ( n4631 & n5294 ) | ( n4631 & ~n30385 ) | ( n5294 & ~n30385 ) ;
  assign n30387 = ( n14067 & ~n14322 ) | ( n14067 & n22263 ) | ( ~n14322 & n22263 ) ;
  assign n30388 = n27842 ^ n20470 ^ n9954 ;
  assign n30389 = ( n3673 & n4862 ) | ( n3673 & ~n16535 ) | ( n4862 & ~n16535 ) ;
  assign n30390 = ( n9598 & n17497 ) | ( n9598 & n28368 ) | ( n17497 & n28368 ) ;
  assign n30391 = ( n19874 & n20700 ) | ( n19874 & ~n30390 ) | ( n20700 & ~n30390 ) ;
  assign n30392 = ( n7998 & ~n13775 ) | ( n7998 & n20364 ) | ( ~n13775 & n20364 ) ;
  assign n30393 = ( n4778 & n11167 ) | ( n4778 & ~n30392 ) | ( n11167 & ~n30392 ) ;
  assign n30394 = ~n2478 & n30393 ;
  assign n30395 = n10687 & n30394 ;
  assign n30398 = ( n1594 & n2233 ) | ( n1594 & ~n2684 ) | ( n2233 & ~n2684 ) ;
  assign n30396 = ( x49 & ~n6086 ) | ( x49 & n20859 ) | ( ~n6086 & n20859 ) ;
  assign n30397 = n30396 ^ n7882 ^ n6127 ;
  assign n30399 = n30398 ^ n30397 ^ n7083 ;
  assign n30400 = n25114 ^ n20641 ^ n3174 ;
  assign n30401 = ( n4675 & ~n30399 ) | ( n4675 & n30400 ) | ( ~n30399 & n30400 ) ;
  assign n30402 = n30401 ^ n6061 ^ 1'b0 ;
  assign n30403 = ( ~n6160 & n10139 ) | ( ~n6160 & n26453 ) | ( n10139 & n26453 ) ;
  assign n30404 = n13903 | n30403 ;
  assign n30405 = n4930 | n30404 ;
  assign n30410 = n26950 ^ n11740 ^ x136 ;
  assign n30411 = n30410 ^ n14484 ^ n10865 ;
  assign n30409 = n30297 ^ n30127 ^ n3405 ;
  assign n30406 = n21809 ^ n13831 ^ n2640 ;
  assign n30407 = ( n6942 & n15947 ) | ( n6942 & n30406 ) | ( n15947 & n30406 ) ;
  assign n30408 = n30407 ^ n6373 ^ n3813 ;
  assign n30412 = n30411 ^ n30409 ^ n30408 ;
  assign n30413 = ( ~n6392 & n7691 ) | ( ~n6392 & n12819 ) | ( n7691 & n12819 ) ;
  assign n30414 = ( n2449 & n4090 ) | ( n2449 & n26579 ) | ( n4090 & n26579 ) ;
  assign n30415 = ( n23896 & n27566 ) | ( n23896 & ~n30414 ) | ( n27566 & ~n30414 ) ;
  assign n30416 = n25201 ^ n24608 ^ n15279 ;
  assign n30417 = ( n1594 & ~n13169 ) | ( n1594 & n22491 ) | ( ~n13169 & n22491 ) ;
  assign n30418 = ( n11854 & ~n12269 ) | ( n11854 & n25360 ) | ( ~n12269 & n25360 ) ;
  assign n30419 = n30418 ^ n22586 ^ n19639 ;
  assign n30420 = ( n18000 & n28778 ) | ( n18000 & ~n28993 ) | ( n28778 & ~n28993 ) ;
  assign n30421 = ( n1549 & n3036 ) | ( n1549 & n20497 ) | ( n3036 & n20497 ) ;
  assign n30422 = n30421 ^ n3737 ^ 1'b0 ;
  assign n30423 = n27328 | n30422 ;
  assign n30424 = n30423 ^ n11071 ^ 1'b0 ;
  assign n30425 = n21888 ^ n7732 ^ 1'b0 ;
  assign n30426 = n7557 & ~n30425 ;
  assign n30427 = ( ~n10131 & n28007 ) | ( ~n10131 & n30426 ) | ( n28007 & n30426 ) ;
  assign n30428 = n25292 ^ n6016 ^ n5473 ;
  assign n30429 = n30428 ^ n24168 ^ n17401 ;
  assign n30430 = ( n5989 & ~n26278 ) | ( n5989 & n29852 ) | ( ~n26278 & n29852 ) ;
  assign n30431 = ( ~n12689 & n25319 ) | ( ~n12689 & n30430 ) | ( n25319 & n30430 ) ;
  assign n30432 = n28951 ^ n5611 ^ n1469 ;
  assign n30433 = ( n2948 & n3194 ) | ( n2948 & n9546 ) | ( n3194 & n9546 ) ;
  assign n30434 = n13940 ^ n12937 ^ n7162 ;
  assign n30435 = ( n11803 & ~n16851 ) | ( n11803 & n30434 ) | ( ~n16851 & n30434 ) ;
  assign n30436 = n22020 & n30162 ;
  assign n30437 = n30436 ^ n21402 ^ n2443 ;
  assign n30438 = ( n21984 & n30435 ) | ( n21984 & ~n30437 ) | ( n30435 & ~n30437 ) ;
  assign n30439 = ( ~x7 & n2573 ) | ( ~x7 & n8766 ) | ( n2573 & n8766 ) ;
  assign n30440 = n10318 ^ n3349 ^ 1'b0 ;
  assign n30441 = n30439 | n30440 ;
  assign n30442 = n895 & ~n5383 ;
  assign n30443 = n387 & n30442 ;
  assign n30444 = ( n10515 & ~n30441 ) | ( n10515 & n30443 ) | ( ~n30441 & n30443 ) ;
  assign n30445 = ~n6080 & n26034 ;
  assign n30446 = ( n26246 & ~n30364 ) | ( n26246 & n30445 ) | ( ~n30364 & n30445 ) ;
  assign n30447 = n30446 ^ n25597 ^ n22765 ;
  assign n30448 = ( n18745 & n27728 ) | ( n18745 & n30447 ) | ( n27728 & n30447 ) ;
  assign n30449 = n16693 ^ n483 ^ x126 ;
  assign n30450 = ( n3453 & n19586 ) | ( n3453 & ~n30449 ) | ( n19586 & ~n30449 ) ;
  assign n30451 = n10772 ^ n9701 ^ 1'b0 ;
  assign n30452 = n30451 ^ n22471 ^ n7316 ;
  assign n30453 = n30452 ^ n22082 ^ n5234 ;
  assign n30454 = n23567 & n27529 ;
  assign n30455 = ( n6355 & n13259 ) | ( n6355 & ~n14243 ) | ( n13259 & ~n14243 ) ;
  assign n30456 = n30455 ^ n5856 ^ n1600 ;
  assign n30457 = n5799 | n16131 ;
  assign n30458 = ( n9873 & n25316 ) | ( n9873 & ~n30457 ) | ( n25316 & ~n30457 ) ;
  assign n30459 = n30458 ^ n18826 ^ n3199 ;
  assign n30460 = ( ~n22137 & n30456 ) | ( ~n22137 & n30459 ) | ( n30456 & n30459 ) ;
  assign n30461 = ( n2596 & ~n22904 ) | ( n2596 & n24388 ) | ( ~n22904 & n24388 ) ;
  assign n30462 = ( n4364 & ~n10583 ) | ( n4364 & n29308 ) | ( ~n10583 & n29308 ) ;
  assign n30463 = n9817 ^ n3757 ^ x140 ;
  assign n30464 = ( n4377 & ~n8227 ) | ( n4377 & n13354 ) | ( ~n8227 & n13354 ) ;
  assign n30465 = ( n10653 & n30463 ) | ( n10653 & n30464 ) | ( n30463 & n30464 ) ;
  assign n30466 = ( ~n6316 & n7147 ) | ( ~n6316 & n30465 ) | ( n7147 & n30465 ) ;
  assign n30467 = ( n2661 & n30462 ) | ( n2661 & ~n30466 ) | ( n30462 & ~n30466 ) ;
  assign n30468 = n11840 ^ n5652 ^ 1'b0 ;
  assign n30470 = ( n772 & ~n3138 ) | ( n772 & n6326 ) | ( ~n3138 & n6326 ) ;
  assign n30469 = n30285 ^ n23016 ^ n9542 ;
  assign n30471 = n30470 ^ n30469 ^ n14876 ;
  assign n30472 = ( n1255 & n7556 ) | ( n1255 & ~n8209 ) | ( n7556 & ~n8209 ) ;
  assign n30473 = n30472 ^ n8506 ^ 1'b0 ;
  assign n30474 = n23984 & ~n30473 ;
  assign n30475 = n10776 ^ n6309 ^ n849 ;
  assign n30476 = n30475 ^ n20955 ^ n14728 ;
  assign n30477 = n30476 ^ n17553 ^ n10580 ;
  assign n30478 = n22246 ^ n15271 ^ n2342 ;
  assign n30479 = ( n1240 & ~n28714 ) | ( n1240 & n30478 ) | ( ~n28714 & n30478 ) ;
  assign n30480 = ( n1136 & n16909 ) | ( n1136 & ~n30479 ) | ( n16909 & ~n30479 ) ;
  assign n30481 = ( n5121 & ~n17832 ) | ( n5121 & n30480 ) | ( ~n17832 & n30480 ) ;
  assign n30483 = n14379 ^ n10637 ^ n9035 ;
  assign n30482 = n25689 ^ n17211 ^ n14302 ;
  assign n30484 = n30483 ^ n30482 ^ 1'b0 ;
  assign n30485 = n19009 ^ n18509 ^ n18101 ;
  assign n30486 = n17331 ^ n8122 ^ n479 ;
  assign n30487 = ( n1394 & n1586 ) | ( n1394 & ~n6824 ) | ( n1586 & ~n6824 ) ;
  assign n30488 = ( n18143 & n30486 ) | ( n18143 & n30487 ) | ( n30486 & n30487 ) ;
  assign n30490 = ( ~n11206 & n14900 ) | ( ~n11206 & n18469 ) | ( n14900 & n18469 ) ;
  assign n30489 = ( n671 & n19312 ) | ( n671 & ~n19898 ) | ( n19312 & ~n19898 ) ;
  assign n30491 = n30490 ^ n30489 ^ n11922 ;
  assign n30492 = n1986 & n13311 ;
  assign n30493 = ~n16270 & n30492 ;
  assign n30494 = n23051 ^ n16466 ^ n1817 ;
  assign n30495 = ~n2566 & n30494 ;
  assign n30496 = n30495 ^ n4024 ^ 1'b0 ;
  assign n30497 = ( n13839 & ~n30493 ) | ( n13839 & n30496 ) | ( ~n30493 & n30496 ) ;
  assign n30498 = n7368 ^ n4646 ^ n855 ;
  assign n30499 = ~n4021 & n4722 ;
  assign n30500 = ~n2398 & n30499 ;
  assign n30501 = ( n23647 & ~n30498 ) | ( n23647 & n30500 ) | ( ~n30498 & n30500 ) ;
  assign n30503 = n14269 ^ n2486 ^ n1078 ;
  assign n30502 = n8802 ^ n7783 ^ n3054 ;
  assign n30504 = n30503 ^ n30502 ^ n1622 ;
  assign n30505 = ( n5377 & n27090 ) | ( n5377 & n30504 ) | ( n27090 & n30504 ) ;
  assign n30508 = n20270 ^ n16522 ^ n2098 ;
  assign n30509 = ( ~n6162 & n7122 ) | ( ~n6162 & n30508 ) | ( n7122 & n30508 ) ;
  assign n30506 = ( n6391 & ~n7531 ) | ( n6391 & n9602 ) | ( ~n7531 & n9602 ) ;
  assign n30507 = n30506 ^ n9729 ^ 1'b0 ;
  assign n30510 = n30509 ^ n30507 ^ n11342 ;
  assign n30511 = ( n7872 & ~n18015 ) | ( n7872 & n20671 ) | ( ~n18015 & n20671 ) ;
  assign n30512 = ( n13264 & n16779 ) | ( n13264 & n30511 ) | ( n16779 & n30511 ) ;
  assign n30513 = n8371 ^ n4221 ^ n2205 ;
  assign n30514 = ( n21731 & n24473 ) | ( n21731 & ~n30513 ) | ( n24473 & ~n30513 ) ;
  assign n30515 = n7522 ^ x47 ^ 1'b0 ;
  assign n30516 = n30515 ^ n11687 ^ n9464 ;
  assign n30517 = n30516 ^ n24524 ^ n4358 ;
  assign n30518 = ( n15299 & ~n18197 ) | ( n15299 & n28815 ) | ( ~n18197 & n28815 ) ;
  assign n30519 = n10579 | n30518 ;
  assign n30520 = n2807 & ~n14429 ;
  assign n30523 = n18412 ^ n5827 ^ n837 ;
  assign n30521 = ~n8612 & n11202 ;
  assign n30522 = n3705 & n30521 ;
  assign n30524 = n30523 ^ n30522 ^ n17327 ;
  assign n30525 = n27363 ^ n18619 ^ n5164 ;
  assign n30526 = ( n9773 & ~n19123 ) | ( n9773 & n19194 ) | ( ~n19123 & n19194 ) ;
  assign n30527 = n8113 ^ n665 ^ x99 ;
  assign n30529 = n8358 ^ n3070 ^ n1200 ;
  assign n30528 = ( ~n1688 & n6626 ) | ( ~n1688 & n16991 ) | ( n6626 & n16991 ) ;
  assign n30530 = n30529 ^ n30528 ^ n3489 ;
  assign n30531 = ( n4307 & n30527 ) | ( n4307 & ~n30530 ) | ( n30527 & ~n30530 ) ;
  assign n30532 = n20305 & ~n30531 ;
  assign n30533 = n30532 ^ n8837 ^ 1'b0 ;
  assign n30534 = n16240 | n22838 ;
  assign n30535 = n1612 | n30534 ;
  assign n30536 = n15138 ^ n7853 ^ n3816 ;
  assign n30537 = n20302 ^ n10746 ^ 1'b0 ;
  assign n30538 = n13311 & ~n30537 ;
  assign n30539 = n30538 ^ n12041 ^ 1'b0 ;
  assign n30540 = n30536 & n30539 ;
  assign n30541 = ( n11664 & n15848 ) | ( n11664 & n19203 ) | ( n15848 & n19203 ) ;
  assign n30542 = ~n14268 & n15770 ;
  assign n30543 = n30542 ^ n18967 ^ n16619 ;
  assign n30544 = n30541 | n30543 ;
  assign n30545 = n30359 | n30544 ;
  assign n30546 = ( n30535 & ~n30540 ) | ( n30535 & n30545 ) | ( ~n30540 & n30545 ) ;
  assign n30547 = n15986 ^ n9846 ^ n5654 ;
  assign n30548 = ( n4767 & n10553 ) | ( n4767 & n25129 ) | ( n10553 & n25129 ) ;
  assign n30549 = n30548 ^ n26882 ^ n13933 ;
  assign n30550 = ( n20192 & ~n30547 ) | ( n20192 & n30549 ) | ( ~n30547 & n30549 ) ;
  assign n30551 = n6727 & n10261 ;
  assign n30552 = n14180 & n30551 ;
  assign n30553 = ( n11315 & n26073 ) | ( n11315 & ~n30552 ) | ( n26073 & ~n30552 ) ;
  assign n30554 = ( ~n5269 & n6959 ) | ( ~n5269 & n14392 ) | ( n6959 & n14392 ) ;
  assign n30555 = ( n7526 & n23198 ) | ( n7526 & ~n30554 ) | ( n23198 & ~n30554 ) ;
  assign n30556 = n10683 & ~n16801 ;
  assign n30557 = ( ~n8160 & n30555 ) | ( ~n8160 & n30556 ) | ( n30555 & n30556 ) ;
  assign n30558 = n20977 & ~n22914 ;
  assign n30559 = ( n24115 & n24701 ) | ( n24115 & ~n30558 ) | ( n24701 & ~n30558 ) ;
  assign n30560 = ( ~n10218 & n18009 ) | ( ~n10218 & n30559 ) | ( n18009 & n30559 ) ;
  assign n30561 = n4910 | n15846 ;
  assign n30562 = n30561 ^ n7107 ^ 1'b0 ;
  assign n30563 = ( n4223 & ~n16636 ) | ( n4223 & n30562 ) | ( ~n16636 & n30562 ) ;
  assign n30564 = ( n2986 & n10742 ) | ( n2986 & n30563 ) | ( n10742 & n30563 ) ;
  assign n30565 = ( n376 & n14009 ) | ( n376 & ~n30564 ) | ( n14009 & ~n30564 ) ;
  assign n30566 = n30565 ^ n17923 ^ n11474 ;
  assign n30567 = n11725 ^ n1158 ^ 1'b0 ;
  assign n30568 = n21821 & ~n30567 ;
  assign n30569 = ( n19692 & n24589 ) | ( n19692 & n26051 ) | ( n24589 & n26051 ) ;
  assign n30570 = n22636 ^ n6294 ^ n3676 ;
  assign n30571 = ( n6279 & ~n12456 ) | ( n6279 & n30570 ) | ( ~n12456 & n30570 ) ;
  assign n30572 = ( n8350 & n19300 ) | ( n8350 & ~n30571 ) | ( n19300 & ~n30571 ) ;
  assign n30573 = ( n272 & ~n6972 ) | ( n272 & n15302 ) | ( ~n6972 & n15302 ) ;
  assign n30574 = n18121 ^ n11655 ^ n7484 ;
  assign n30575 = ( n5587 & ~n11292 ) | ( n5587 & n30574 ) | ( ~n11292 & n30574 ) ;
  assign n30576 = ( ~n10635 & n30573 ) | ( ~n10635 & n30575 ) | ( n30573 & n30575 ) ;
  assign n30577 = n23216 ^ n7947 ^ 1'b0 ;
  assign n30578 = n17115 & n30577 ;
  assign n30579 = ( n1583 & n5167 ) | ( n1583 & n17334 ) | ( n5167 & n17334 ) ;
  assign n30580 = ( n9018 & ~n20298 ) | ( n9018 & n20524 ) | ( ~n20298 & n20524 ) ;
  assign n30581 = ( ~n9609 & n30579 ) | ( ~n9609 & n30580 ) | ( n30579 & n30580 ) ;
  assign n30582 = ( n12791 & ~n27248 ) | ( n12791 & n29904 ) | ( ~n27248 & n29904 ) ;
  assign n30583 = n30582 ^ n20845 ^ n11157 ;
  assign n30584 = n19480 ^ n1974 ^ 1'b0 ;
  assign n30585 = ( n23654 & n30583 ) | ( n23654 & n30584 ) | ( n30583 & n30584 ) ;
  assign n30586 = ( ~n8634 & n10163 ) | ( ~n8634 & n30585 ) | ( n10163 & n30585 ) ;
  assign n30587 = ( ~n2545 & n30581 ) | ( ~n2545 & n30586 ) | ( n30581 & n30586 ) ;
  assign n30588 = n29478 ^ n12943 ^ n4239 ;
  assign n30589 = n30588 ^ n18270 ^ n16710 ;
  assign n30590 = n28820 ^ n18898 ^ n18418 ;
  assign n30591 = ( n1274 & n18691 ) | ( n1274 & n30590 ) | ( n18691 & n30590 ) ;
  assign n30592 = n14330 ^ n9386 ^ n7322 ;
  assign n30593 = n23406 ^ n13916 ^ n799 ;
  assign n30594 = ( n4482 & ~n20987 ) | ( n4482 & n30593 ) | ( ~n20987 & n30593 ) ;
  assign n30595 = ( n3515 & n10224 ) | ( n3515 & n30594 ) | ( n10224 & n30594 ) ;
  assign n30596 = n30592 & n30595 ;
  assign n30597 = ~n11498 & n30596 ;
  assign n30598 = n30597 ^ n18809 ^ n2224 ;
  assign n30599 = n9969 ^ n7237 ^ 1'b0 ;
  assign n30600 = ~n5586 & n30599 ;
  assign n30601 = n30600 ^ n11073 ^ n2160 ;
  assign n30602 = n10295 ^ n929 ^ 1'b0 ;
  assign n30603 = n18519 & ~n30602 ;
  assign n30604 = ( n9438 & n14748 ) | ( n9438 & ~n30603 ) | ( n14748 & ~n30603 ) ;
  assign n30605 = n16939 ^ n8567 ^ x178 ;
  assign n30606 = n30605 ^ n5910 ^ n5084 ;
  assign n30607 = n11590 | n15448 ;
  assign n30608 = n30606 & ~n30607 ;
  assign n30609 = ( n30601 & n30604 ) | ( n30601 & n30608 ) | ( n30604 & n30608 ) ;
  assign n30610 = n24575 ^ n4631 ^ 1'b0 ;
  assign n30611 = n21818 & ~n30610 ;
  assign n30612 = ( n11587 & n30609 ) | ( n11587 & ~n30611 ) | ( n30609 & ~n30611 ) ;
  assign n30613 = n30612 ^ n4614 ^ 1'b0 ;
  assign n30614 = ( ~n5719 & n15732 ) | ( ~n5719 & n25864 ) | ( n15732 & n25864 ) ;
  assign n30615 = ( n3514 & n8126 ) | ( n3514 & n10096 ) | ( n8126 & n10096 ) ;
  assign n30616 = n19403 ^ n14455 ^ n14178 ;
  assign n30617 = ~n30615 & n30616 ;
  assign n30618 = n19196 ^ n13824 ^ n2238 ;
  assign n30619 = n30618 ^ n25726 ^ n25409 ;
  assign n30620 = n4521 | n6252 ;
  assign n30621 = n30620 ^ n19238 ^ n6895 ;
  assign n30622 = n8846 & ~n30621 ;
  assign n30623 = ( n17187 & n21293 ) | ( n17187 & ~n23221 ) | ( n21293 & ~n23221 ) ;
  assign n30624 = ~n6336 & n11199 ;
  assign n30625 = n30624 ^ n13306 ^ n8681 ;
  assign n30626 = n20768 ^ n19070 ^ n10038 ;
  assign n30627 = n4396 & ~n5192 ;
  assign n30628 = ( n16004 & ~n23514 ) | ( n16004 & n30627 ) | ( ~n23514 & n30627 ) ;
  assign n30629 = n13298 ^ n10558 ^ n471 ;
  assign n30630 = n12857 ^ n12286 ^ n10799 ;
  assign n30631 = n30630 ^ n23121 ^ n9477 ;
  assign n30632 = ( n30628 & n30629 ) | ( n30628 & n30631 ) | ( n30629 & n30631 ) ;
  assign n30636 = n18939 ^ n9025 ^ n1278 ;
  assign n30633 = ( ~n5262 & n10935 ) | ( ~n5262 & n14087 ) | ( n10935 & n14087 ) ;
  assign n30634 = ( n10697 & n18732 ) | ( n10697 & n30633 ) | ( n18732 & n30633 ) ;
  assign n30635 = n30634 ^ n22828 ^ n7955 ;
  assign n30637 = n30636 ^ n30635 ^ n16767 ;
  assign n30638 = n21697 ^ n1712 ^ n289 ;
  assign n30639 = n19313 | n30638 ;
  assign n30640 = n15447 | n30639 ;
  assign n30641 = ( ~n343 & n11249 ) | ( ~n343 & n30640 ) | ( n11249 & n30640 ) ;
  assign n30642 = ( ~n9287 & n10692 ) | ( ~n9287 & n30005 ) | ( n10692 & n30005 ) ;
  assign n30643 = n30642 ^ n28527 ^ n27034 ;
  assign n30644 = n20548 ^ n18626 ^ 1'b0 ;
  assign n30645 = n30643 & ~n30644 ;
  assign n30646 = ( n2250 & n5140 ) | ( n2250 & ~n14623 ) | ( n5140 & ~n14623 ) ;
  assign n30647 = n21595 ^ n17524 ^ n14331 ;
  assign n30648 = ( n6880 & ~n30646 ) | ( n6880 & n30647 ) | ( ~n30646 & n30647 ) ;
  assign n30649 = ( n8837 & n29026 ) | ( n8837 & ~n30648 ) | ( n29026 & ~n30648 ) ;
  assign n30650 = ( n1989 & n10095 ) | ( n1989 & n11392 ) | ( n10095 & n11392 ) ;
  assign n30651 = n30650 ^ n20103 ^ n17443 ;
  assign n30652 = ( n9040 & ~n14104 ) | ( n9040 & n30651 ) | ( ~n14104 & n30651 ) ;
  assign n30653 = n6802 ^ n4887 ^ 1'b0 ;
  assign n30654 = n14699 ^ n6995 ^ n4553 ;
  assign n30655 = ( x244 & ~n11923 ) | ( x244 & n12482 ) | ( ~n11923 & n12482 ) ;
  assign n30656 = ( ~n17899 & n23301 ) | ( ~n17899 & n30655 ) | ( n23301 & n30655 ) ;
  assign n30657 = ( ~n569 & n30654 ) | ( ~n569 & n30656 ) | ( n30654 & n30656 ) ;
  assign n30658 = ( x167 & ~n13067 ) | ( x167 & n20888 ) | ( ~n13067 & n20888 ) ;
  assign n30659 = ( n7772 & ~n12364 ) | ( n7772 & n30658 ) | ( ~n12364 & n30658 ) ;
  assign n30660 = ( n1427 & ~n5215 ) | ( n1427 & n8944 ) | ( ~n5215 & n8944 ) ;
  assign n30661 = ( n6250 & n30319 ) | ( n6250 & n30660 ) | ( n30319 & n30660 ) ;
  assign n30662 = ( ~n11032 & n17608 ) | ( ~n11032 & n30661 ) | ( n17608 & n30661 ) ;
  assign n30663 = n16201 | n21780 ;
  assign n30664 = ( n577 & n22689 ) | ( n577 & n30663 ) | ( n22689 & n30663 ) ;
  assign n30665 = n30664 ^ n21992 ^ n11630 ;
  assign n30666 = n11722 & ~n21053 ;
  assign n30667 = n30665 & n30666 ;
  assign n30673 = n24929 ^ n20464 ^ n17398 ;
  assign n30668 = n16169 ^ n14191 ^ n7919 ;
  assign n30669 = n30668 ^ n13258 ^ 1'b0 ;
  assign n30670 = n13686 & ~n30669 ;
  assign n30671 = n9729 ^ x25 ^ 1'b0 ;
  assign n30672 = n30670 & n30671 ;
  assign n30674 = n30673 ^ n30672 ^ n17902 ;
  assign n30675 = ( n6546 & n8106 ) | ( n6546 & n13541 ) | ( n8106 & n13541 ) ;
  assign n30676 = n30675 ^ n24461 ^ n675 ;
  assign n30677 = n15513 ^ n8214 ^ n449 ;
  assign n30678 = n23090 ^ n14168 ^ n10039 ;
  assign n30679 = ( x159 & n1296 ) | ( x159 & ~n30678 ) | ( n1296 & ~n30678 ) ;
  assign n30680 = ~n10620 & n23680 ;
  assign n30681 = ~n18912 & n30680 ;
  assign n30682 = ( n1276 & ~n4344 ) | ( n1276 & n11667 ) | ( ~n4344 & n11667 ) ;
  assign n30683 = n30682 ^ n27443 ^ 1'b0 ;
  assign n30684 = ~n30681 & n30683 ;
  assign n30685 = ( ~n5198 & n7365 ) | ( ~n5198 & n13047 ) | ( n7365 & n13047 ) ;
  assign n30686 = ( n3082 & ~n4323 ) | ( n3082 & n12396 ) | ( ~n4323 & n12396 ) ;
  assign n30687 = ( ~n9083 & n24582 ) | ( ~n9083 & n30686 ) | ( n24582 & n30686 ) ;
  assign n30688 = n25860 ^ n10839 ^ n9010 ;
  assign n30689 = ( ~n22732 & n30687 ) | ( ~n22732 & n30688 ) | ( n30687 & n30688 ) ;
  assign n30690 = n28891 ^ n18464 ^ n10776 ;
  assign n30691 = n30690 ^ n24839 ^ n1117 ;
  assign n30692 = ( ~n4576 & n9573 ) | ( ~n4576 & n18526 ) | ( n9573 & n18526 ) ;
  assign n30693 = n30692 ^ n5923 ^ n4734 ;
  assign n30694 = ( n2118 & ~n30691 ) | ( n2118 & n30693 ) | ( ~n30691 & n30693 ) ;
  assign n30695 = n30694 ^ n26439 ^ n18107 ;
  assign n30696 = ( n8943 & n25063 ) | ( n8943 & n30695 ) | ( n25063 & n30695 ) ;
  assign n30697 = n9280 ^ n3189 ^ 1'b0 ;
  assign n30699 = n19213 ^ n9849 ^ 1'b0 ;
  assign n30700 = n30699 ^ n21496 ^ n6957 ;
  assign n30701 = n30700 ^ n26270 ^ n4728 ;
  assign n30698 = ( ~n8887 & n19945 ) | ( ~n8887 & n23553 ) | ( n19945 & n23553 ) ;
  assign n30702 = n30701 ^ n30698 ^ n26950 ;
  assign n30703 = ( n3763 & n18836 ) | ( n3763 & ~n25488 ) | ( n18836 & ~n25488 ) ;
  assign n30704 = ( n30697 & n30702 ) | ( n30697 & ~n30703 ) | ( n30702 & ~n30703 ) ;
  assign n30705 = ( n12050 & n25188 ) | ( n12050 & ~n30463 ) | ( n25188 & ~n30463 ) ;
  assign n30706 = n19844 ^ n9359 ^ n912 ;
  assign n30707 = ( n1511 & ~n5699 ) | ( n1511 & n26106 ) | ( ~n5699 & n26106 ) ;
  assign n30708 = ~n23486 & n30707 ;
  assign n30709 = n30708 ^ n18591 ^ 1'b0 ;
  assign n30710 = ( n813 & n1928 ) | ( n813 & n9495 ) | ( n1928 & n9495 ) ;
  assign n30711 = n30710 ^ n25960 ^ n5567 ;
  assign n30712 = n30709 & ~n30711 ;
  assign n30713 = ~n30706 & n30712 ;
  assign n30714 = n29695 ^ n16842 ^ n15921 ;
  assign n30715 = ( ~n539 & n25083 ) | ( ~n539 & n30714 ) | ( n25083 & n30714 ) ;
  assign n30716 = ( n2752 & ~n6463 ) | ( n2752 & n6819 ) | ( ~n6463 & n6819 ) ;
  assign n30717 = n20962 & n30716 ;
  assign n30718 = n30715 & n30717 ;
  assign n30719 = n14968 ^ n11231 ^ n6882 ;
  assign n30720 = n30719 ^ n22669 ^ n16815 ;
  assign n30721 = ( n13532 & n15984 ) | ( n13532 & n28538 ) | ( n15984 & n28538 ) ;
  assign n30722 = n14942 & n16535 ;
  assign n30723 = ( n612 & n10094 ) | ( n612 & ~n13994 ) | ( n10094 & ~n13994 ) ;
  assign n30724 = n7130 & ~n28908 ;
  assign n30725 = ~n30723 & n30724 ;
  assign n30726 = n6362 | n30725 ;
  assign n30727 = n24986 | n30726 ;
  assign n30728 = n4713 & n30727 ;
  assign n30729 = n30722 & n30728 ;
  assign n30730 = ( n819 & n20142 ) | ( n819 & n30729 ) | ( n20142 & n30729 ) ;
  assign n30731 = ( ~n14455 & n24282 ) | ( ~n14455 & n30730 ) | ( n24282 & n30730 ) ;
  assign n30733 = x73 & ~n8371 ;
  assign n30732 = n12517 ^ n5321 ^ n5105 ;
  assign n30734 = n30733 ^ n30732 ^ n858 ;
  assign n30735 = ( x47 & n8097 ) | ( x47 & n22974 ) | ( n8097 & n22974 ) ;
  assign n30736 = ( n9259 & n28975 ) | ( n9259 & n30735 ) | ( n28975 & n30735 ) ;
  assign n30737 = n21542 ^ n1276 ^ 1'b0 ;
  assign n30738 = ( n6545 & n21873 ) | ( n6545 & n30737 ) | ( n21873 & n30737 ) ;
  assign n30747 = ( n3051 & n7077 ) | ( n3051 & ~n15505 ) | ( n7077 & ~n15505 ) ;
  assign n30745 = n29724 ^ n21117 ^ n9262 ;
  assign n30739 = n13099 & ~n14883 ;
  assign n30740 = ~n26708 & n30739 ;
  assign n30741 = n18923 ^ n11338 ^ n7118 ;
  assign n30742 = n7463 | n13717 ;
  assign n30743 = n30741 & ~n30742 ;
  assign n30744 = ( n2292 & n30740 ) | ( n2292 & ~n30743 ) | ( n30740 & ~n30743 ) ;
  assign n30746 = n30745 ^ n30744 ^ n6853 ;
  assign n30748 = n30747 ^ n30746 ^ n17430 ;
  assign n30750 = n18888 ^ n6823 ^ 1'b0 ;
  assign n30749 = n13722 ^ n9679 ^ n6252 ;
  assign n30751 = n30750 ^ n30749 ^ 1'b0 ;
  assign n30752 = n20054 ^ n12367 ^ 1'b0 ;
  assign n30756 = ( n6261 & ~n6596 ) | ( n6261 & n7822 ) | ( ~n6596 & n7822 ) ;
  assign n30755 = ( ~n5753 & n5769 ) | ( ~n5753 & n6105 ) | ( n5769 & n6105 ) ;
  assign n30753 = n9964 & n13674 ;
  assign n30754 = ~n8341 & n30753 ;
  assign n30757 = n30756 ^ n30755 ^ n30754 ;
  assign n30758 = ( ~n2720 & n9184 ) | ( ~n2720 & n23325 ) | ( n9184 & n23325 ) ;
  assign n30759 = n24988 ^ n8260 ^ n7000 ;
  assign n30760 = ( n9422 & ~n30758 ) | ( n9422 & n30759 ) | ( ~n30758 & n30759 ) ;
  assign n30761 = ( n7168 & ~n18454 ) | ( n7168 & n21208 ) | ( ~n18454 & n21208 ) ;
  assign n30762 = n30761 ^ n20777 ^ 1'b0 ;
  assign n30763 = ( n1018 & n7030 ) | ( n1018 & ~n14177 ) | ( n7030 & ~n14177 ) ;
  assign n30764 = n4117 & ~n10655 ;
  assign n30765 = n30763 & n30764 ;
  assign n30766 = n2334 & ~n30765 ;
  assign n30767 = n30766 ^ n16359 ^ 1'b0 ;
  assign n30768 = n30767 ^ n24502 ^ n18280 ;
  assign n30769 = n19689 ^ n13848 ^ 1'b0 ;
  assign n30770 = ( n5910 & n12439 ) | ( n5910 & ~n30769 ) | ( n12439 & ~n30769 ) ;
  assign n30772 = n23268 ^ n6697 ^ n4502 ;
  assign n30771 = ( n7611 & ~n19787 ) | ( n7611 & n24818 ) | ( ~n19787 & n24818 ) ;
  assign n30773 = n30772 ^ n30771 ^ n25230 ;
  assign n30774 = n11668 & ~n29770 ;
  assign n30775 = n30774 ^ n15658 ^ 1'b0 ;
  assign n30776 = n13158 ^ n12744 ^ n4141 ;
  assign n30777 = n30776 ^ n20883 ^ 1'b0 ;
  assign n30778 = n5498 & n30777 ;
  assign n30780 = n3352 ^ n2166 ^ n835 ;
  assign n30779 = ( n8617 & n9857 ) | ( n8617 & ~n16514 ) | ( n9857 & ~n16514 ) ;
  assign n30781 = n30780 ^ n30779 ^ n27797 ;
  assign n30782 = n21339 ^ n7643 ^ x108 ;
  assign n30783 = ( n3271 & ~n8030 ) | ( n3271 & n26006 ) | ( ~n8030 & n26006 ) ;
  assign n30784 = ( n8444 & n13256 ) | ( n8444 & ~n20186 ) | ( n13256 & ~n20186 ) ;
  assign n30785 = ( ~n6093 & n30783 ) | ( ~n6093 & n30784 ) | ( n30783 & n30784 ) ;
  assign n30787 = n9447 ^ n6924 ^ n6180 ;
  assign n30786 = n4534 | n23258 ;
  assign n30788 = n30787 ^ n30786 ^ 1'b0 ;
  assign n30789 = ( n5160 & n16764 ) | ( n5160 & ~n19329 ) | ( n16764 & ~n19329 ) ;
  assign n30790 = n4662 & n15757 ;
  assign n30791 = n4484 & n30790 ;
  assign n30792 = n30791 ^ n28116 ^ 1'b0 ;
  assign n30793 = n30792 ^ n19435 ^ n18984 ;
  assign n30794 = ( ~n4863 & n17788 ) | ( ~n4863 & n21036 ) | ( n17788 & n21036 ) ;
  assign n30795 = n13128 ^ n7742 ^ n769 ;
  assign n30796 = n16855 ^ n6254 ^ 1'b0 ;
  assign n30797 = n2072 & n30796 ;
  assign n30798 = ( n4442 & n10642 ) | ( n4442 & ~n30797 ) | ( n10642 & ~n30797 ) ;
  assign n30799 = n30798 ^ n7571 ^ 1'b0 ;
  assign n30800 = n30795 & ~n30799 ;
  assign n30801 = n17051 ^ n16814 ^ n13606 ;
  assign n30802 = n30801 ^ n19997 ^ n6155 ;
  assign n30803 = ( ~n4518 & n11015 ) | ( ~n4518 & n19988 ) | ( n11015 & n19988 ) ;
  assign n30804 = n24569 ^ n8109 ^ n4544 ;
  assign n30805 = n10021 & n11411 ;
  assign n30806 = ( ~n5509 & n12146 ) | ( ~n5509 & n19212 ) | ( n12146 & n19212 ) ;
  assign n30807 = n30806 ^ n26929 ^ n6939 ;
  assign n30808 = ( n23358 & n30805 ) | ( n23358 & ~n30807 ) | ( n30805 & ~n30807 ) ;
  assign n30809 = ( ~n23668 & n30804 ) | ( ~n23668 & n30808 ) | ( n30804 & n30808 ) ;
  assign n30817 = n21355 ^ n7977 ^ n6479 ;
  assign n30811 = n18715 ^ n6572 ^ n5972 ;
  assign n30812 = n17481 ^ n6201 ^ 1'b0 ;
  assign n30813 = n30811 & ~n30812 ;
  assign n30814 = ~n5434 & n30813 ;
  assign n30815 = n30814 ^ n17620 ^ 1'b0 ;
  assign n30810 = ( ~n4844 & n9003 ) | ( ~n4844 & n27073 ) | ( n9003 & n27073 ) ;
  assign n30816 = n30815 ^ n30810 ^ n2777 ;
  assign n30818 = n30817 ^ n30816 ^ n1007 ;
  assign n30819 = n28051 ^ n16588 ^ 1'b0 ;
  assign n30820 = n3943 & ~n30819 ;
  assign n30821 = ( ~n11901 & n11940 ) | ( ~n11901 & n30820 ) | ( n11940 & n30820 ) ;
  assign n30822 = n1472 & n3014 ;
  assign n30823 = n3270 & ~n18775 ;
  assign n30824 = n4111 ^ n2937 ^ n448 ;
  assign n30826 = ( ~n1509 & n1666 ) | ( ~n1509 & n10935 ) | ( n1666 & n10935 ) ;
  assign n30825 = n17345 & ~n24177 ;
  assign n30827 = n30826 ^ n30825 ^ 1'b0 ;
  assign n30828 = n30827 ^ n27520 ^ n19147 ;
  assign n30829 = ( n14783 & n30824 ) | ( n14783 & ~n30828 ) | ( n30824 & ~n30828 ) ;
  assign n30830 = ~n1874 & n30829 ;
  assign n30831 = ( n30822 & ~n30823 ) | ( n30822 & n30830 ) | ( ~n30823 & n30830 ) ;
  assign n30832 = n17022 ^ n12724 ^ n7283 ;
  assign n30833 = ( n451 & n3329 ) | ( n451 & n30832 ) | ( n3329 & n30832 ) ;
  assign n30834 = ( n24448 & ~n28534 ) | ( n24448 & n30833 ) | ( ~n28534 & n30833 ) ;
  assign n30835 = ( ~n24640 & n27678 ) | ( ~n24640 & n30834 ) | ( n27678 & n30834 ) ;
  assign n30836 = n27103 ^ n16051 ^ n7766 ;
  assign n30837 = ( n8924 & ~n12347 ) | ( n8924 & n30836 ) | ( ~n12347 & n30836 ) ;
  assign n30838 = n30837 ^ n28778 ^ n597 ;
  assign n30839 = n9000 ^ n6131 ^ n4783 ;
  assign n30840 = n30839 ^ n14100 ^ n12698 ;
  assign n30841 = n30840 ^ n9792 ^ n1502 ;
  assign n30842 = n30841 ^ n12631 ^ 1'b0 ;
  assign n30848 = n11104 ^ n9868 ^ n4282 ;
  assign n30849 = n30848 ^ n13862 ^ n4199 ;
  assign n30844 = ( ~n10386 & n18153 ) | ( ~n10386 & n26959 ) | ( n18153 & n26959 ) ;
  assign n30845 = n12262 ^ n4460 ^ 1'b0 ;
  assign n30846 = n3063 & ~n30845 ;
  assign n30847 = ( n5854 & n30844 ) | ( n5854 & n30846 ) | ( n30844 & n30846 ) ;
  assign n30843 = n20003 ^ n9797 ^ n1779 ;
  assign n30850 = n30849 ^ n30847 ^ n30843 ;
  assign n30851 = n6166 & n11216 ;
  assign n30852 = ~n3589 & n30851 ;
  assign n30853 = ( n8632 & n13445 ) | ( n8632 & n30852 ) | ( n13445 & n30852 ) ;
  assign n30854 = n24334 | n30853 ;
  assign n30855 = n7734 & ~n30854 ;
  assign n30856 = ( n273 & n3495 ) | ( n273 & n30855 ) | ( n3495 & n30855 ) ;
  assign n30857 = ( ~n819 & n4782 ) | ( ~n819 & n11315 ) | ( n4782 & n11315 ) ;
  assign n30858 = n30857 ^ n2678 ^ n1846 ;
  assign n30859 = ( n8523 & n9535 ) | ( n8523 & n16097 ) | ( n9535 & n16097 ) ;
  assign n30860 = n30859 ^ n13871 ^ n11406 ;
  assign n30861 = n30860 ^ n20018 ^ n14141 ;
  assign n30862 = ( n6374 & ~n19373 ) | ( n6374 & n30861 ) | ( ~n19373 & n30861 ) ;
  assign n30863 = ( n1272 & ~n1381 ) | ( n1272 & n7857 ) | ( ~n1381 & n7857 ) ;
  assign n30864 = ( n3439 & n5408 ) | ( n3439 & ~n6845 ) | ( n5408 & ~n6845 ) ;
  assign n30865 = ( ~n3801 & n30863 ) | ( ~n3801 & n30864 ) | ( n30863 & n30864 ) ;
  assign n30866 = ( ~n1879 & n2599 ) | ( ~n1879 & n30865 ) | ( n2599 & n30865 ) ;
  assign n30867 = ( n11365 & n23190 ) | ( n11365 & ~n30866 ) | ( n23190 & ~n30866 ) ;
  assign n30868 = ~n4142 & n8241 ;
  assign n30869 = n399 & n30868 ;
  assign n30870 = n3403 | n30869 ;
  assign n30871 = n11182 | n30870 ;
  assign n30872 = ( ~n2212 & n18152 ) | ( ~n2212 & n20740 ) | ( n18152 & n20740 ) ;
  assign n30873 = ( ~n8233 & n23341 ) | ( ~n8233 & n30872 ) | ( n23341 & n30872 ) ;
  assign n30874 = ( n4738 & ~n7358 ) | ( n4738 & n9326 ) | ( ~n7358 & n9326 ) ;
  assign n30875 = n3763 & ~n8732 ;
  assign n30876 = n6835 & ~n30875 ;
  assign n30877 = n30876 ^ n15940 ^ n11470 ;
  assign n30878 = ( n10339 & n10941 ) | ( n10339 & ~n30877 ) | ( n10941 & ~n30877 ) ;
  assign n30879 = ( n680 & ~n10043 ) | ( n680 & n30878 ) | ( ~n10043 & n30878 ) ;
  assign n30880 = ( n1555 & n9946 ) | ( n1555 & n30843 ) | ( n9946 & n30843 ) ;
  assign n30881 = n29339 ^ n19361 ^ n15378 ;
  assign n30882 = n30881 ^ n27650 ^ n27253 ;
  assign n30887 = n27358 ^ n17585 ^ n7712 ;
  assign n30883 = n22372 ^ n2325 ^ 1'b0 ;
  assign n30884 = n12567 & n30883 ;
  assign n30885 = n30884 ^ n16796 ^ 1'b0 ;
  assign n30886 = n21353 & ~n30885 ;
  assign n30888 = n30887 ^ n30886 ^ 1'b0 ;
  assign n30889 = ~n8897 & n30888 ;
  assign n30890 = n1282 & n4699 ;
  assign n30891 = n30890 ^ n6477 ^ 1'b0 ;
  assign n30892 = ( x237 & ~n8405 ) | ( x237 & n30891 ) | ( ~n8405 & n30891 ) ;
  assign n30893 = ( n7302 & n27420 ) | ( n7302 & n30892 ) | ( n27420 & n30892 ) ;
  assign n30894 = n29889 ^ n21932 ^ n8974 ;
  assign n30897 = n18406 ^ n17696 ^ n11373 ;
  assign n30895 = ( n9870 & ~n14478 ) | ( n9870 & n30315 ) | ( ~n14478 & n30315 ) ;
  assign n30896 = ( n9599 & n17155 ) | ( n9599 & ~n30895 ) | ( n17155 & ~n30895 ) ;
  assign n30898 = n30897 ^ n30896 ^ n8081 ;
  assign n30899 = ~n8595 & n20576 ;
  assign n30900 = n30899 ^ n15905 ^ n1911 ;
  assign n30901 = ( ~n1270 & n3392 ) | ( ~n1270 & n6462 ) | ( n3392 & n6462 ) ;
  assign n30902 = n30901 ^ n6626 ^ n3692 ;
  assign n30903 = ( n17629 & n26774 ) | ( n17629 & ~n26849 ) | ( n26774 & ~n26849 ) ;
  assign n30904 = ( n8027 & n17464 ) | ( n8027 & ~n29716 ) | ( n17464 & ~n29716 ) ;
  assign n30905 = ( n30902 & n30903 ) | ( n30902 & n30904 ) | ( n30903 & n30904 ) ;
  assign n30906 = n13601 ^ n5447 ^ 1'b0 ;
  assign n30907 = n30906 ^ n23592 ^ n20364 ;
  assign n30908 = n30907 ^ n23635 ^ n14001 ;
  assign n30909 = n19591 ^ n8216 ^ n4341 ;
  assign n30910 = n18226 | n23553 ;
  assign n30911 = n8407 | n30910 ;
  assign n30912 = n30911 ^ n26857 ^ n24590 ;
  assign n30913 = n30912 ^ n19544 ^ n13769 ;
  assign n30914 = ( n30009 & n30909 ) | ( n30009 & n30913 ) | ( n30909 & n30913 ) ;
  assign n30915 = ( ~n2960 & n7334 ) | ( ~n2960 & n23302 ) | ( n7334 & n23302 ) ;
  assign n30916 = n30915 ^ n21224 ^ n16338 ;
  assign n30917 = n15989 ^ n2677 ^ n266 ;
  assign n30918 = ( n5442 & ~n9647 ) | ( n5442 & n30917 ) | ( ~n9647 & n30917 ) ;
  assign n30919 = ( n6678 & n30916 ) | ( n6678 & ~n30918 ) | ( n30916 & ~n30918 ) ;
  assign n30920 = ( ~n10216 & n11502 ) | ( ~n10216 & n11554 ) | ( n11502 & n11554 ) ;
  assign n30921 = n18196 ^ n11797 ^ n650 ;
  assign n30922 = n30921 ^ n26340 ^ n18667 ;
  assign n30923 = ( n22175 & n30920 ) | ( n22175 & n30922 ) | ( n30920 & n30922 ) ;
  assign n30924 = ( ~n24114 & n26608 ) | ( ~n24114 & n28951 ) | ( n26608 & n28951 ) ;
  assign n30925 = n28432 ^ n16958 ^ n15504 ;
  assign n30926 = ( ~n15088 & n20928 ) | ( ~n15088 & n30275 ) | ( n20928 & n30275 ) ;
  assign n30927 = ( n2629 & n8856 ) | ( n2629 & ~n16400 ) | ( n8856 & ~n16400 ) ;
  assign n30928 = ( n1315 & ~n22550 ) | ( n1315 & n30927 ) | ( ~n22550 & n30927 ) ;
  assign n30931 = ( n5025 & n5379 ) | ( n5025 & n10431 ) | ( n5379 & n10431 ) ;
  assign n30929 = n26229 ^ n24410 ^ 1'b0 ;
  assign n30930 = n10814 & n30929 ;
  assign n30932 = n30931 ^ n30930 ^ n14603 ;
  assign n30933 = n26542 ^ n9588 ^ 1'b0 ;
  assign n30934 = n8017 | n30933 ;
  assign n30936 = ( ~n2963 & n5042 ) | ( ~n2963 & n15084 ) | ( n5042 & n15084 ) ;
  assign n30935 = n17020 ^ n1282 ^ n423 ;
  assign n30937 = n30936 ^ n30935 ^ n3835 ;
  assign n30938 = ( n8338 & ~n11840 ) | ( n8338 & n15836 ) | ( ~n11840 & n15836 ) ;
  assign n30939 = n30938 ^ n23337 ^ 1'b0 ;
  assign n30940 = n23442 & n30939 ;
  assign n30941 = ( n10765 & n25790 ) | ( n10765 & n30940 ) | ( n25790 & n30940 ) ;
  assign n30942 = ( n9374 & ~n30937 ) | ( n9374 & n30941 ) | ( ~n30937 & n30941 ) ;
  assign n30943 = n30942 ^ n15952 ^ x211 ;
  assign n30944 = n11150 & n19212 ;
  assign n30945 = ( n6259 & ~n8487 ) | ( n6259 & n23615 ) | ( ~n8487 & n23615 ) ;
  assign n30946 = ( ~n21281 & n30944 ) | ( ~n21281 & n30945 ) | ( n30944 & n30945 ) ;
  assign n30947 = ( n832 & n6463 ) | ( n832 & n29806 ) | ( n6463 & n29806 ) ;
  assign n30951 = n26961 ^ n13092 ^ n9994 ;
  assign n30948 = n25928 ^ n2195 ^ n826 ;
  assign n30949 = n30948 ^ n14032 ^ 1'b0 ;
  assign n30950 = n29952 & n30949 ;
  assign n30952 = n30951 ^ n30950 ^ n21411 ;
  assign n30953 = n12430 & n17420 ;
  assign n30954 = n5811 & n30953 ;
  assign n30955 = ( n3293 & ~n14736 ) | ( n3293 & n30954 ) | ( ~n14736 & n30954 ) ;
  assign n30956 = ( n1326 & ~n25745 ) | ( n1326 & n30364 ) | ( ~n25745 & n30364 ) ;
  assign n30957 = ( n8029 & ~n30955 ) | ( n8029 & n30956 ) | ( ~n30955 & n30956 ) ;
  assign n30958 = ( n18185 & ~n24762 ) | ( n18185 & n30957 ) | ( ~n24762 & n30957 ) ;
  assign n30959 = ( n12616 & n13998 ) | ( n12616 & ~n27368 ) | ( n13998 & ~n27368 ) ;
  assign n30960 = n28600 ^ n19891 ^ n2592 ;
  assign n30961 = n11168 ^ n11038 ^ n7638 ;
  assign n30962 = n30961 ^ n24435 ^ 1'b0 ;
  assign n30963 = n22547 ^ n4536 ^ n2154 ;
  assign n30964 = n3384 | n11805 ;
  assign n30965 = n30964 ^ n30719 ^ 1'b0 ;
  assign n30966 = n30965 ^ n29242 ^ n9129 ;
  assign n30967 = ( ~n14136 & n30963 ) | ( ~n14136 & n30966 ) | ( n30963 & n30966 ) ;
  assign n30968 = ( n30960 & n30962 ) | ( n30960 & ~n30967 ) | ( n30962 & ~n30967 ) ;
  assign n30969 = n7734 ^ n569 ^ 1'b0 ;
  assign n30970 = ( n15867 & ~n15917 ) | ( n15867 & n26028 ) | ( ~n15917 & n26028 ) ;
  assign n30971 = n30642 ^ n18440 ^ n14708 ;
  assign n30972 = ( ~n14586 & n21412 ) | ( ~n14586 & n23231 ) | ( n21412 & n23231 ) ;
  assign n30973 = n22741 ^ n14353 ^ n11926 ;
  assign n30974 = ( n19334 & n21009 ) | ( n19334 & ~n30973 ) | ( n21009 & ~n30973 ) ;
  assign n30975 = n30974 ^ n25157 ^ n16591 ;
  assign n30977 = n14466 ^ n8548 ^ n5044 ;
  assign n30978 = n30977 ^ n23506 ^ n12733 ;
  assign n30979 = ( n18001 & ~n22954 ) | ( n18001 & n30978 ) | ( ~n22954 & n30978 ) ;
  assign n30976 = n13055 & ~n24478 ;
  assign n30980 = n30979 ^ n30976 ^ 1'b0 ;
  assign n30981 = n21752 ^ n20985 ^ n19970 ;
  assign n30983 = ( x80 & n1260 ) | ( x80 & n6683 ) | ( n1260 & n6683 ) ;
  assign n30982 = ( n1893 & n7537 ) | ( n1893 & ~n29074 ) | ( n7537 & ~n29074 ) ;
  assign n30984 = n30983 ^ n30982 ^ n12714 ;
  assign n30988 = n16192 ^ n12016 ^ n3266 ;
  assign n30989 = n30988 ^ n9124 ^ n8301 ;
  assign n30985 = n6014 ^ n5625 ^ n4642 ;
  assign n30986 = ( ~n12766 & n13181 ) | ( ~n12766 & n30985 ) | ( n13181 & n30985 ) ;
  assign n30987 = n30986 ^ n18576 ^ n7146 ;
  assign n30990 = n30989 ^ n30987 ^ n10745 ;
  assign n30991 = ( n1435 & n2651 ) | ( n1435 & n19511 ) | ( n2651 & n19511 ) ;
  assign n30992 = ( n6277 & n22974 ) | ( n6277 & ~n30991 ) | ( n22974 & ~n30991 ) ;
  assign n30993 = ( ~n5009 & n13824 ) | ( ~n5009 & n24424 ) | ( n13824 & n24424 ) ;
  assign n30994 = n21650 ^ n2920 ^ 1'b0 ;
  assign n30995 = ~n9781 & n30994 ;
  assign n30996 = ( n8183 & ~n17736 ) | ( n8183 & n30995 ) | ( ~n17736 & n30995 ) ;
  assign n30997 = ( ~n17833 & n30993 ) | ( ~n17833 & n30996 ) | ( n30993 & n30996 ) ;
  assign n31001 = n14848 ^ n10688 ^ n6697 ;
  assign n31002 = n6277 | n18393 ;
  assign n31003 = n6027 | n31002 ;
  assign n31004 = ( n15663 & n31001 ) | ( n15663 & n31003 ) | ( n31001 & n31003 ) ;
  assign n30998 = ( n905 & n914 ) | ( n905 & n9138 ) | ( n914 & n9138 ) ;
  assign n30999 = n30998 ^ n28022 ^ n22666 ;
  assign n31000 = n30999 ^ n6136 ^ n6007 ;
  assign n31005 = n31004 ^ n31000 ^ n15295 ;
  assign n31006 = ( x105 & n4205 ) | ( x105 & ~n30723 ) | ( n4205 & ~n30723 ) ;
  assign n31007 = n31006 ^ n28586 ^ 1'b0 ;
  assign n31008 = n31005 & n31007 ;
  assign n31009 = x133 & ~n16190 ;
  assign n31010 = n20835 ^ n7320 ^ 1'b0 ;
  assign n31011 = n16969 & n31010 ;
  assign n31012 = ( ~n16876 & n22977 ) | ( ~n16876 & n31011 ) | ( n22977 & n31011 ) ;
  assign n31013 = n31012 ^ n16571 ^ n8101 ;
  assign n31016 = ( n4573 & ~n9076 ) | ( n4573 & n10476 ) | ( ~n9076 & n10476 ) ;
  assign n31017 = ( n7187 & n8186 ) | ( n7187 & n31016 ) | ( n8186 & n31016 ) ;
  assign n31014 = n6330 ^ n3744 ^ n349 ;
  assign n31015 = n31014 ^ n14919 ^ x97 ;
  assign n31018 = n31017 ^ n31015 ^ n17758 ;
  assign n31019 = n12749 ^ n7820 ^ 1'b0 ;
  assign n31025 = n8815 ^ n2823 ^ n351 ;
  assign n31026 = ( n257 & n3675 ) | ( n257 & n31025 ) | ( n3675 & n31025 ) ;
  assign n31024 = n8468 | n12989 ;
  assign n31027 = n31026 ^ n31024 ^ n14352 ;
  assign n31023 = n14139 & ~n18276 ;
  assign n31028 = n31027 ^ n31023 ^ 1'b0 ;
  assign n31020 = n27591 ^ n8125 ^ n7844 ;
  assign n31021 = ( ~n9176 & n23366 ) | ( ~n9176 & n31020 ) | ( n23366 & n31020 ) ;
  assign n31022 = n31021 ^ n13865 ^ n8904 ;
  assign n31029 = n31028 ^ n31022 ^ 1'b0 ;
  assign n31030 = ~n6864 & n31029 ;
  assign n31031 = ( n13559 & n19468 ) | ( n13559 & ~n31030 ) | ( n19468 & ~n31030 ) ;
  assign n31032 = ~n13865 & n17030 ;
  assign n31035 = n15848 ^ n2694 ^ n1458 ;
  assign n31036 = n31035 ^ n28542 ^ n17214 ;
  assign n31037 = n996 & ~n31036 ;
  assign n31038 = n14094 ^ n3616 ^ 1'b0 ;
  assign n31039 = n31038 ^ n11290 ^ n1090 ;
  assign n31040 = n31039 ^ n19995 ^ n17125 ;
  assign n31041 = ( n7659 & n31037 ) | ( n7659 & n31040 ) | ( n31037 & n31040 ) ;
  assign n31033 = ( ~n7225 & n8849 ) | ( ~n7225 & n20546 ) | ( n8849 & n20546 ) ;
  assign n31034 = n31033 ^ n7294 ^ n7101 ;
  assign n31042 = n31041 ^ n31034 ^ n29578 ;
  assign n31043 = n19510 ^ n8103 ^ n2809 ;
  assign n31044 = ( n12212 & n21275 ) | ( n12212 & n31043 ) | ( n21275 & n31043 ) ;
  assign n31045 = ( ~n15818 & n22495 ) | ( ~n15818 & n23899 ) | ( n22495 & n23899 ) ;
  assign n31053 = n19091 ^ n16808 ^ n4826 ;
  assign n31048 = ~n574 & n9337 ;
  assign n31046 = ( n12966 & ~n13469 ) | ( n12966 & n23043 ) | ( ~n13469 & n23043 ) ;
  assign n31047 = n31046 ^ n16583 ^ n7666 ;
  assign n31049 = n31048 ^ n31047 ^ n4440 ;
  assign n31050 = n3335 & ~n31049 ;
  assign n31051 = n31050 ^ n11182 ^ 1'b0 ;
  assign n31052 = n31051 ^ n26143 ^ n12415 ;
  assign n31054 = n31053 ^ n31052 ^ x205 ;
  assign n31055 = n11967 & ~n11976 ;
  assign n31056 = ~n12171 & n31055 ;
  assign n31057 = n12847 ^ n11500 ^ n727 ;
  assign n31058 = n4137 & ~n18821 ;
  assign n31059 = n21193 & n31058 ;
  assign n31060 = ( ~n12030 & n31057 ) | ( ~n12030 & n31059 ) | ( n31057 & n31059 ) ;
  assign n31061 = ( n8739 & n15938 ) | ( n8739 & n31060 ) | ( n15938 & n31060 ) ;
  assign n31062 = n9566 ^ n7926 ^ n2968 ;
  assign n31063 = n31062 ^ n16034 ^ n7958 ;
  assign n31064 = ( n4215 & n11576 ) | ( n4215 & ~n19814 ) | ( n11576 & ~n19814 ) ;
  assign n31065 = ( ~n24663 & n27937 ) | ( ~n24663 & n28891 ) | ( n27937 & n28891 ) ;
  assign n31066 = ( ~n904 & n10171 ) | ( ~n904 & n31065 ) | ( n10171 & n31065 ) ;
  assign n31067 = n26857 ^ n21887 ^ n20619 ;
  assign n31068 = n13146 ^ n4385 ^ n3862 ;
  assign n31069 = ~n26371 & n31068 ;
  assign n31070 = ~n31067 & n31069 ;
  assign n31071 = ( ~n5492 & n29874 ) | ( ~n5492 & n31070 ) | ( n29874 & n31070 ) ;
  assign n31072 = n20415 ^ n13567 ^ n3947 ;
  assign n31073 = n31072 ^ n25125 ^ n10642 ;
  assign n31074 = n20508 ^ n7433 ^ 1'b0 ;
  assign n31075 = n12617 ^ n3908 ^ 1'b0 ;
  assign n31076 = n31075 ^ n30695 ^ n24152 ;
  assign n31077 = n29852 ^ n26587 ^ n3103 ;
  assign n31086 = ( n11135 & n12385 ) | ( n11135 & n14530 ) | ( n12385 & n14530 ) ;
  assign n31087 = ( n4581 & n5027 ) | ( n4581 & ~n31086 ) | ( n5027 & ~n31086 ) ;
  assign n31088 = ( n15558 & n19209 ) | ( n15558 & ~n31087 ) | ( n19209 & ~n31087 ) ;
  assign n31081 = ( n794 & ~n1120 ) | ( n794 & n7578 ) | ( ~n1120 & n7578 ) ;
  assign n31082 = n27051 ^ n21695 ^ 1'b0 ;
  assign n31083 = n7661 & n31082 ;
  assign n31084 = n15961 & n31083 ;
  assign n31085 = ( n23753 & n31081 ) | ( n23753 & n31084 ) | ( n31081 & n31084 ) ;
  assign n31079 = n2754 | n4771 ;
  assign n31078 = ( n6423 & n7537 ) | ( n6423 & n22219 ) | ( n7537 & n22219 ) ;
  assign n31080 = n31079 ^ n31078 ^ n4483 ;
  assign n31089 = n31088 ^ n31085 ^ n31080 ;
  assign n31090 = ( n4602 & n5768 ) | ( n4602 & n28200 ) | ( n5768 & n28200 ) ;
  assign n31091 = n2682 & ~n31090 ;
  assign n31092 = ~n31089 & n31091 ;
  assign n31093 = n31092 ^ n12235 ^ n527 ;
  assign n31094 = n28486 ^ n24857 ^ 1'b0 ;
  assign n31095 = n29211 ^ n21725 ^ n12460 ;
  assign n31096 = n11508 ^ n10524 ^ n3984 ;
  assign n31097 = n16641 ^ n15927 ^ n12482 ;
  assign n31098 = ( n4322 & n31096 ) | ( n4322 & n31097 ) | ( n31096 & n31097 ) ;
  assign n31099 = n28067 ^ n19976 ^ n14124 ;
  assign n31100 = n18430 ^ n4569 ^ 1'b0 ;
  assign n31101 = ~n4923 & n31100 ;
  assign n31102 = n18978 ^ n10878 ^ 1'b0 ;
  assign n31103 = ( ~n15088 & n31101 ) | ( ~n15088 & n31102 ) | ( n31101 & n31102 ) ;
  assign n31104 = n31103 ^ n10188 ^ n496 ;
  assign n31105 = ( n2783 & n13898 ) | ( n2783 & n22029 ) | ( n13898 & n22029 ) ;
  assign n31106 = n16805 ^ n3338 ^ n2655 ;
  assign n31107 = ( ~n14010 & n25238 ) | ( ~n14010 & n26461 ) | ( n25238 & n26461 ) ;
  assign n31108 = ( n2492 & n24134 ) | ( n2492 & n31107 ) | ( n24134 & n31107 ) ;
  assign n31109 = n15453 & ~n31108 ;
  assign n31110 = ( ~n3383 & n9263 ) | ( ~n3383 & n24984 ) | ( n9263 & n24984 ) ;
  assign n31111 = ( n19209 & n21471 ) | ( n19209 & ~n31110 ) | ( n21471 & ~n31110 ) ;
  assign n31116 = ( n4570 & n6680 ) | ( n4570 & ~n7066 ) | ( n6680 & ~n7066 ) ;
  assign n31115 = n28779 ^ n17918 ^ n12474 ;
  assign n31112 = n3869 & n22861 ;
  assign n31113 = n31112 ^ n27454 ^ 1'b0 ;
  assign n31114 = ( n1658 & ~n23522 ) | ( n1658 & n31113 ) | ( ~n23522 & n31113 ) ;
  assign n31117 = n31116 ^ n31115 ^ n31114 ;
  assign n31118 = n17588 ^ n11631 ^ 1'b0 ;
  assign n31119 = n19343 & ~n31118 ;
  assign n31120 = ( n371 & n4616 ) | ( n371 & ~n10251 ) | ( n4616 & ~n10251 ) ;
  assign n31121 = ( n1944 & ~n30396 ) | ( n1944 & n31120 ) | ( ~n30396 & n31120 ) ;
  assign n31122 = n6243 & ~n16158 ;
  assign n31123 = n25113 & n31122 ;
  assign n31124 = ~n31121 & n31123 ;
  assign n31127 = n20987 ^ n10449 ^ n6490 ;
  assign n31126 = ( n1402 & ~n5741 ) | ( n1402 & n22174 ) | ( ~n5741 & n22174 ) ;
  assign n31128 = n31127 ^ n31126 ^ n16091 ;
  assign n31125 = ( n4246 & n17481 ) | ( n4246 & n19843 ) | ( n17481 & n19843 ) ;
  assign n31129 = n31128 ^ n31125 ^ n20635 ;
  assign n31130 = n11900 ^ n4376 ^ 1'b0 ;
  assign n31131 = ( n6879 & ~n7259 ) | ( n6879 & n11362 ) | ( ~n7259 & n11362 ) ;
  assign n31132 = n13498 ^ n10445 ^ n9091 ;
  assign n31133 = n31132 ^ n26733 ^ n7960 ;
  assign n31134 = ( ~n11200 & n19003 ) | ( ~n11200 & n31133 ) | ( n19003 & n31133 ) ;
  assign n31135 = n31134 ^ n14142 ^ n12166 ;
  assign n31136 = n31135 ^ n28934 ^ n16350 ;
  assign n31137 = n31136 ^ n23552 ^ n13717 ;
  assign n31138 = n30337 ^ n8200 ^ 1'b0 ;
  assign n31139 = ( n5826 & n22727 ) | ( n5826 & ~n31138 ) | ( n22727 & ~n31138 ) ;
  assign n31140 = n25022 ^ n14281 ^ n3891 ;
  assign n31147 = ( n10826 & ~n12171 ) | ( n10826 & n26342 ) | ( ~n12171 & n26342 ) ;
  assign n31144 = n10818 ^ n9341 ^ n5679 ;
  assign n31145 = n31144 ^ n8151 ^ n8073 ;
  assign n31146 = n3056 & ~n31145 ;
  assign n31142 = ( ~n693 & n12437 ) | ( ~n693 & n24969 ) | ( n12437 & n24969 ) ;
  assign n31141 = n27254 ^ n26536 ^ n14839 ;
  assign n31143 = n31142 ^ n31141 ^ n24555 ;
  assign n31148 = n31147 ^ n31146 ^ n31143 ;
  assign n31153 = ( x21 & n8666 ) | ( x21 & ~n12783 ) | ( n8666 & ~n12783 ) ;
  assign n31149 = n8681 ^ n4289 ^ 1'b0 ;
  assign n31150 = n31149 ^ n15960 ^ n7813 ;
  assign n31151 = ( n6060 & n26493 ) | ( n6060 & ~n31150 ) | ( n26493 & ~n31150 ) ;
  assign n31152 = n31151 ^ n30841 ^ n13175 ;
  assign n31154 = n31153 ^ n31152 ^ n2890 ;
  assign n31155 = n26970 ^ n18434 ^ n10629 ;
  assign n31156 = n21426 ^ n14611 ^ n5737 ;
  assign n31161 = n9114 ^ n3919 ^ n2230 ;
  assign n31162 = ( n9949 & n22171 ) | ( n9949 & ~n31161 ) | ( n22171 & ~n31161 ) ;
  assign n31163 = n31162 ^ n22600 ^ n9796 ;
  assign n31157 = n27948 ^ n18129 ^ n4307 ;
  assign n31158 = ( n16950 & n20901 ) | ( n16950 & n30437 ) | ( n20901 & n30437 ) ;
  assign n31159 = ( ~n30091 & n31157 ) | ( ~n30091 & n31158 ) | ( n31157 & n31158 ) ;
  assign n31160 = ( n10504 & ~n20030 ) | ( n10504 & n31159 ) | ( ~n20030 & n31159 ) ;
  assign n31164 = n31163 ^ n31160 ^ n14747 ;
  assign n31168 = n6859 ^ n6752 ^ n2555 ;
  assign n31165 = n12244 ^ n6583 ^ n5339 ;
  assign n31166 = n25094 & n31165 ;
  assign n31167 = n31166 ^ n12324 ^ 1'b0 ;
  assign n31169 = n31168 ^ n31167 ^ 1'b0 ;
  assign n31170 = ( n11431 & ~n18222 ) | ( n11431 & n25203 ) | ( ~n18222 & n25203 ) ;
  assign n31171 = n31170 ^ n812 ^ 1'b0 ;
  assign n31172 = n28324 | n31171 ;
  assign n31173 = ( n7274 & ~n10424 ) | ( n7274 & n24878 ) | ( ~n10424 & n24878 ) ;
  assign n31174 = n2947 & n31173 ;
  assign n31175 = n31174 ^ x224 ^ 1'b0 ;
  assign n31178 = ( ~n762 & n2201 ) | ( ~n762 & n7923 ) | ( n2201 & n7923 ) ;
  assign n31176 = ( ~n9566 & n23213 ) | ( ~n9566 & n29103 ) | ( n23213 & n29103 ) ;
  assign n31177 = n31176 ^ n17277 ^ n5498 ;
  assign n31179 = n31178 ^ n31177 ^ n18651 ;
  assign n31180 = ( x223 & n4424 ) | ( x223 & n9819 ) | ( n4424 & n9819 ) ;
  assign n31181 = n31180 ^ n26925 ^ n2948 ;
  assign n31182 = n8198 ^ n5233 ^ n3863 ;
  assign n31183 = n12455 ^ n1141 ^ 1'b0 ;
  assign n31184 = n31183 ^ n19980 ^ n14431 ;
  assign n31185 = n26847 & n31184 ;
  assign n31186 = n31185 ^ n17296 ^ 1'b0 ;
  assign n31187 = n18814 ^ n18151 ^ n4294 ;
  assign n31188 = ( n2220 & n19232 ) | ( n2220 & ~n31187 ) | ( n19232 & ~n31187 ) ;
  assign n31189 = n31188 ^ n10352 ^ n4981 ;
  assign n31190 = ( ~n309 & n6286 ) | ( ~n309 & n14065 ) | ( n6286 & n14065 ) ;
  assign n31191 = ( n6525 & ~n15641 ) | ( n6525 & n31190 ) | ( ~n15641 & n31190 ) ;
  assign n31192 = n31191 ^ n6135 ^ n4637 ;
  assign n31193 = n23642 ^ n20811 ^ n7464 ;
  assign n31197 = n21540 ^ n16245 ^ n14715 ;
  assign n31194 = n3954 & ~n24672 ;
  assign n31195 = n31194 ^ n2587 ^ 1'b0 ;
  assign n31196 = n31195 ^ n10631 ^ n6806 ;
  assign n31198 = n31197 ^ n31196 ^ n18520 ;
  assign n31199 = ( ~n26544 & n27678 ) | ( ~n26544 & n31198 ) | ( n27678 & n31198 ) ;
  assign n31200 = n27638 ^ n15519 ^ n5915 ;
  assign n31201 = ( n14499 & ~n15180 ) | ( n14499 & n31200 ) | ( ~n15180 & n31200 ) ;
  assign n31202 = n9179 ^ n6911 ^ n4921 ;
  assign n31203 = n14261 & ~n28036 ;
  assign n31204 = ( n9337 & n9543 ) | ( n9337 & n31203 ) | ( n9543 & n31203 ) ;
  assign n31205 = n31202 | n31204 ;
  assign n31206 = n31205 ^ n10159 ^ n7895 ;
  assign n31207 = n23324 ^ n8489 ^ 1'b0 ;
  assign n31208 = n8178 & ~n31207 ;
  assign n31209 = ( n7600 & ~n18637 ) | ( n7600 & n31208 ) | ( ~n18637 & n31208 ) ;
  assign n31210 = ( ~n4837 & n5857 ) | ( ~n4837 & n31209 ) | ( n5857 & n31209 ) ;
  assign n31212 = n26773 ^ n8639 ^ n5780 ;
  assign n31211 = ( n7129 & ~n10775 ) | ( n7129 & n16786 ) | ( ~n10775 & n16786 ) ;
  assign n31213 = n31212 ^ n31211 ^ n21826 ;
  assign n31214 = ( ~n14063 & n31210 ) | ( ~n14063 & n31213 ) | ( n31210 & n31213 ) ;
  assign n31215 = ( n18964 & n28768 ) | ( n18964 & ~n31214 ) | ( n28768 & ~n31214 ) ;
  assign n31216 = n4274 & n28638 ;
  assign n31217 = n31216 ^ n14769 ^ 1'b0 ;
  assign n31218 = x95 & ~n7380 ;
  assign n31219 = ~n8279 & n31218 ;
  assign n31220 = ( ~n11311 & n17284 ) | ( ~n11311 & n31219 ) | ( n17284 & n31219 ) ;
  assign n31221 = n22424 & ~n31220 ;
  assign n31222 = n31221 ^ n7945 ^ 1'b0 ;
  assign n31223 = n31222 ^ n15965 ^ n11279 ;
  assign n31224 = ( n3698 & n6722 ) | ( n3698 & n8816 ) | ( n6722 & n8816 ) ;
  assign n31225 = n13472 & ~n31224 ;
  assign n31226 = ~n31223 & n31225 ;
  assign n31227 = n27246 ^ n14639 ^ n4257 ;
  assign n31228 = n31227 ^ n8004 ^ n3595 ;
  assign n31229 = n17821 ^ n10504 ^ n5874 ;
  assign n31230 = n31229 ^ n23845 ^ n20786 ;
  assign n31232 = ( ~n13600 & n17712 ) | ( ~n13600 & n24749 ) | ( n17712 & n24749 ) ;
  assign n31231 = n25669 ^ n25484 ^ n17784 ;
  assign n31233 = n31232 ^ n31231 ^ n8588 ;
  assign n31234 = ( n2930 & n22188 ) | ( n2930 & ~n22971 ) | ( n22188 & ~n22971 ) ;
  assign n31235 = ( n5339 & n9576 ) | ( n5339 & n31234 ) | ( n9576 & n31234 ) ;
  assign n31236 = n31235 ^ n26630 ^ n25530 ;
  assign n31237 = ( n1335 & n12070 ) | ( n1335 & n31236 ) | ( n12070 & n31236 ) ;
  assign n31238 = n3639 & n6435 ;
  assign n31239 = n31238 ^ n6208 ^ 1'b0 ;
  assign n31240 = ( ~n18511 & n20253 ) | ( ~n18511 & n31239 ) | ( n20253 & n31239 ) ;
  assign n31241 = ( n3317 & n19976 ) | ( n3317 & n31240 ) | ( n19976 & n31240 ) ;
  assign n31242 = ( n4341 & n6896 ) | ( n4341 & n7182 ) | ( n6896 & n7182 ) ;
  assign n31243 = n31242 ^ n19674 ^ n5976 ;
  assign n31244 = ( n1409 & n7431 ) | ( n1409 & n31243 ) | ( n7431 & n31243 ) ;
  assign n31245 = n25930 ^ n23544 ^ n11283 ;
  assign n31246 = n23279 ^ n21086 ^ n9659 ;
  assign n31247 = n31246 ^ n10226 ^ n9581 ;
  assign n31251 = ( ~n9189 & n16441 ) | ( ~n9189 & n17275 ) | ( n16441 & n17275 ) ;
  assign n31248 = ( ~n1449 & n3147 ) | ( ~n1449 & n16445 ) | ( n3147 & n16445 ) ;
  assign n31249 = n31248 ^ n11038 ^ 1'b0 ;
  assign n31250 = n8178 & n31249 ;
  assign n31252 = n31251 ^ n31250 ^ 1'b0 ;
  assign n31253 = n24223 | n31252 ;
  assign n31254 = ( ~n993 & n1345 ) | ( ~n993 & n5850 ) | ( n1345 & n5850 ) ;
  assign n31255 = ( n10767 & ~n27243 ) | ( n10767 & n31254 ) | ( ~n27243 & n31254 ) ;
  assign n31256 = ( n2791 & n6544 ) | ( n2791 & ~n7072 ) | ( n6544 & ~n7072 ) ;
  assign n31257 = ( ~n12213 & n17976 ) | ( ~n12213 & n31256 ) | ( n17976 & n31256 ) ;
  assign n31261 = ( n910 & ~n4273 ) | ( n910 & n17492 ) | ( ~n4273 & n17492 ) ;
  assign n31258 = ( n2433 & n15550 ) | ( n2433 & ~n18675 ) | ( n15550 & ~n18675 ) ;
  assign n31259 = n16356 | n19261 ;
  assign n31260 = n31258 & ~n31259 ;
  assign n31262 = n31261 ^ n31260 ^ n16056 ;
  assign n31263 = n27256 ^ n10808 ^ n717 ;
  assign n31264 = n22027 ^ n4352 ^ 1'b0 ;
  assign n31265 = n6805 & ~n11970 ;
  assign n31266 = ~n31264 & n31265 ;
  assign n31267 = n31266 ^ n28867 ^ n13649 ;
  assign n31268 = n9806 & ~n12215 ;
  assign n31269 = n26774 ^ n25721 ^ n8260 ;
  assign n31270 = n23741 ^ n4630 ^ n4438 ;
  assign n31271 = n31270 ^ n11802 ^ n6966 ;
  assign n31272 = ( n1452 & n12921 ) | ( n1452 & n15550 ) | ( n12921 & n15550 ) ;
  assign n31273 = n17504 ^ n12002 ^ n9108 ;
  assign n31274 = n31272 & ~n31273 ;
  assign n31275 = n31274 ^ n18187 ^ 1'b0 ;
  assign n31276 = ( ~n8029 & n31271 ) | ( ~n8029 & n31275 ) | ( n31271 & n31275 ) ;
  assign n31277 = n25666 ^ n6377 ^ n2839 ;
  assign n31278 = ( ~n1172 & n8474 ) | ( ~n1172 & n15057 ) | ( n8474 & n15057 ) ;
  assign n31279 = n31278 ^ n12336 ^ 1'b0 ;
  assign n31280 = ( n2733 & n15857 ) | ( n2733 & n18448 ) | ( n15857 & n18448 ) ;
  assign n31281 = n31280 ^ n12184 ^ n7948 ;
  assign n31282 = n29374 ^ n19420 ^ n6454 ;
  assign n31283 = n31282 ^ n12927 ^ n11839 ;
  assign n31284 = ( n17006 & ~n19353 ) | ( n17006 & n31283 ) | ( ~n19353 & n31283 ) ;
  assign n31285 = n6970 & n21778 ;
  assign n31286 = n31284 & n31285 ;
  assign n31287 = n31286 ^ x33 ^ 1'b0 ;
  assign n31288 = ( n7669 & ~n21223 ) | ( n7669 & n29935 ) | ( ~n21223 & n29935 ) ;
  assign n31289 = n3576 & ~n16576 ;
  assign n31290 = n31289 ^ n18275 ^ n7304 ;
  assign n31291 = n19500 ^ n18304 ^ n1847 ;
  assign n31292 = ( n17207 & ~n26989 ) | ( n17207 & n31291 ) | ( ~n26989 & n31291 ) ;
  assign n31293 = n10915 ^ n6672 ^ n4202 ;
  assign n31294 = n31293 ^ n22271 ^ n11569 ;
  assign n31295 = n31294 ^ n17840 ^ 1'b0 ;
  assign n31297 = ( n1488 & n3436 ) | ( n1488 & ~n8670 ) | ( n3436 & ~n8670 ) ;
  assign n31296 = ( n12240 & n26858 ) | ( n12240 & n29379 ) | ( n26858 & n29379 ) ;
  assign n31298 = n31297 ^ n31296 ^ n8887 ;
  assign n31299 = ( n3167 & n9122 ) | ( n3167 & ~n29856 ) | ( n9122 & ~n29856 ) ;
  assign n31300 = n21871 & ~n31299 ;
  assign n31301 = n9183 & n16297 ;
  assign n31302 = ( n17873 & n31300 ) | ( n17873 & ~n31301 ) | ( n31300 & ~n31301 ) ;
  assign n31303 = ( n5800 & ~n9252 ) | ( n5800 & n19013 ) | ( ~n9252 & n19013 ) ;
  assign n31304 = n31303 ^ n18333 ^ n3994 ;
  assign n31305 = n3937 ^ n1691 ^ 1'b0 ;
  assign n31306 = n31304 | n31305 ;
  assign n31307 = ( n4078 & ~n15500 ) | ( n4078 & n21250 ) | ( ~n15500 & n21250 ) ;
  assign n31308 = ( n663 & n10973 ) | ( n663 & ~n31307 ) | ( n10973 & ~n31307 ) ;
  assign n31309 = n6332 ^ n2542 ^ 1'b0 ;
  assign n31310 = n20597 ^ n512 ^ 1'b0 ;
  assign n31311 = ( n5295 & n10791 ) | ( n5295 & ~n24388 ) | ( n10791 & ~n24388 ) ;
  assign n31312 = n31311 ^ n23458 ^ n1236 ;
  assign n31313 = n13227 ^ n1056 ^ 1'b0 ;
  assign n31316 = n11896 ^ n11710 ^ 1'b0 ;
  assign n31314 = n12274 ^ n3742 ^ n2704 ;
  assign n31315 = ~n14007 & n31314 ;
  assign n31317 = n31316 ^ n31315 ^ 1'b0 ;
  assign n31318 = n13806 ^ n13300 ^ n4693 ;
  assign n31319 = n21526 & ~n31318 ;
  assign n31320 = ~n31317 & n31319 ;
  assign n31321 = ( n3294 & n17916 ) | ( n3294 & ~n21440 ) | ( n17916 & ~n21440 ) ;
  assign n31322 = ( n1476 & n21029 ) | ( n1476 & ~n26957 ) | ( n21029 & ~n26957 ) ;
  assign n31323 = ( n16016 & n17481 ) | ( n16016 & n31322 ) | ( n17481 & n31322 ) ;
  assign n31324 = n15307 ^ n10130 ^ n8088 ;
  assign n31325 = ( n12481 & ~n19847 ) | ( n12481 & n31324 ) | ( ~n19847 & n31324 ) ;
  assign n31326 = ( n6492 & n9394 ) | ( n6492 & ~n24373 ) | ( n9394 & ~n24373 ) ;
  assign n31327 = ( n11966 & n18768 ) | ( n11966 & ~n31326 ) | ( n18768 & ~n31326 ) ;
  assign n31328 = n26064 ^ n13166 ^ n11098 ;
  assign n31329 = n31328 ^ n17446 ^ 1'b0 ;
  assign n31330 = ( n31325 & ~n31327 ) | ( n31325 & n31329 ) | ( ~n31327 & n31329 ) ;
  assign n31331 = ( n4029 & n11680 ) | ( n4029 & n29966 ) | ( n11680 & n29966 ) ;
  assign n31332 = n31331 ^ n31120 ^ n21337 ;
  assign n31335 = n11069 ^ n11068 ^ n3507 ;
  assign n31334 = n18429 ^ n14452 ^ n849 ;
  assign n31333 = ( n3244 & n8226 ) | ( n3244 & n23615 ) | ( n8226 & n23615 ) ;
  assign n31336 = n31335 ^ n31334 ^ n31333 ;
  assign n31337 = n31336 ^ n25043 ^ n9863 ;
  assign n31338 = n18665 ^ n8943 ^ 1'b0 ;
  assign n31339 = ( ~n7991 & n17611 ) | ( ~n7991 & n31338 ) | ( n17611 & n31338 ) ;
  assign n31340 = n31339 ^ n28263 ^ n18711 ;
  assign n31341 = ( ~n1586 & n6921 ) | ( ~n1586 & n13258 ) | ( n6921 & n13258 ) ;
  assign n31342 = n31341 ^ n15314 ^ n658 ;
  assign n31343 = n10264 & n18967 ;
  assign n31344 = n31343 ^ n13385 ^ 1'b0 ;
  assign n31345 = n24543 ^ n17865 ^ n1900 ;
  assign n31346 = n31345 ^ n25474 ^ n25352 ;
  assign n31347 = ( n1341 & n3492 ) | ( n1341 & n4191 ) | ( n3492 & n4191 ) ;
  assign n31348 = n6273 ^ n1370 ^ 1'b0 ;
  assign n31349 = n27371 | n31348 ;
  assign n31350 = n31349 ^ n16114 ^ n6492 ;
  assign n31351 = ( n30365 & n31347 ) | ( n30365 & ~n31350 ) | ( n31347 & ~n31350 ) ;
  assign n31352 = n31351 ^ n25804 ^ 1'b0 ;
  assign n31353 = n4051 & ~n31352 ;
  assign n31354 = n25205 ^ n8101 ^ 1'b0 ;
  assign n31355 = n31354 ^ n27414 ^ n22957 ;
  assign n31356 = n23505 ^ n9364 ^ n482 ;
  assign n31357 = ( n3325 & n5283 ) | ( n3325 & ~n26638 ) | ( n5283 & ~n26638 ) ;
  assign n31358 = ( n2221 & n19671 ) | ( n2221 & ~n31357 ) | ( n19671 & ~n31357 ) ;
  assign n31359 = ( n2781 & ~n5291 ) | ( n2781 & n7552 ) | ( ~n5291 & n7552 ) ;
  assign n31360 = n4950 | n31359 ;
  assign n31361 = ( n505 & ~n950 ) | ( n505 & n8587 ) | ( ~n950 & n8587 ) ;
  assign n31362 = ( n5895 & n17179 ) | ( n5895 & n31361 ) | ( n17179 & n31361 ) ;
  assign n31367 = ( n10114 & ~n16520 ) | ( n10114 & n28495 ) | ( ~n16520 & n28495 ) ;
  assign n31368 = n31367 ^ n7814 ^ 1'b0 ;
  assign n31363 = n1282 & n7750 ;
  assign n31364 = n31363 ^ n7283 ^ 1'b0 ;
  assign n31365 = ~n20819 & n31364 ;
  assign n31366 = n27897 & n31365 ;
  assign n31369 = n31368 ^ n31366 ^ n21594 ;
  assign n31370 = ~n31362 & n31369 ;
  assign n31371 = n26172 ^ n12538 ^ 1'b0 ;
  assign n31372 = n24174 & ~n31371 ;
  assign n31373 = n21771 ^ n21471 ^ n9347 ;
  assign n31374 = n31373 ^ n13710 ^ n4387 ;
  assign n31375 = ( n1025 & ~n29110 ) | ( n1025 & n31374 ) | ( ~n29110 & n31374 ) ;
  assign n31376 = ( n434 & n906 ) | ( n434 & n3974 ) | ( n906 & n3974 ) ;
  assign n31377 = n14041 ^ n1945 ^ n1819 ;
  assign n31378 = n31377 ^ n30089 ^ n10484 ;
  assign n31379 = ( n7732 & ~n26907 ) | ( n7732 & n31378 ) | ( ~n26907 & n31378 ) ;
  assign n31380 = ( ~n28247 & n31376 ) | ( ~n28247 & n31379 ) | ( n31376 & n31379 ) ;
  assign n31382 = n17364 & n18526 ;
  assign n31381 = n24722 ^ n2807 ^ n569 ;
  assign n31383 = n31382 ^ n31381 ^ n13052 ;
  assign n31384 = n31383 ^ n29261 ^ n8617 ;
  assign n31385 = n27045 ^ n12566 ^ n2454 ;
  assign n31386 = ( n13179 & n25824 ) | ( n13179 & ~n31385 ) | ( n25824 & ~n31385 ) ;
  assign n31389 = n7184 ^ n4286 ^ n1108 ;
  assign n31388 = n7788 | n18309 ;
  assign n31390 = n31389 ^ n31388 ^ n10672 ;
  assign n31387 = ( n5787 & n12879 ) | ( n5787 & n30030 ) | ( n12879 & n30030 ) ;
  assign n31391 = n31390 ^ n31387 ^ n20784 ;
  assign n31392 = ( n6891 & ~n21445 ) | ( n6891 & n22218 ) | ( ~n21445 & n22218 ) ;
  assign n31393 = n24023 ^ n17164 ^ 1'b0 ;
  assign n31394 = x98 & n31393 ;
  assign n31395 = ( n8735 & ~n10611 ) | ( n8735 & n12311 ) | ( ~n10611 & n12311 ) ;
  assign n31396 = ( ~n14953 & n17246 ) | ( ~n14953 & n31395 ) | ( n17246 & n31395 ) ;
  assign n31397 = ( ~n1578 & n6133 ) | ( ~n1578 & n18734 ) | ( n6133 & n18734 ) ;
  assign n31398 = n31397 ^ n11768 ^ n2233 ;
  assign n31399 = n31398 ^ n20725 ^ n16091 ;
  assign n31400 = n12892 ^ n5997 ^ n1614 ;
  assign n31401 = n11506 ^ n5979 ^ n3755 ;
  assign n31402 = n31401 ^ n15433 ^ x247 ;
  assign n31403 = ( n3257 & n12848 ) | ( n3257 & ~n30202 ) | ( n12848 & ~n30202 ) ;
  assign n31404 = n28885 ^ n11224 ^ n5819 ;
  assign n31405 = ( ~n24688 & n31403 ) | ( ~n24688 & n31404 ) | ( n31403 & n31404 ) ;
  assign n31408 = n25309 ^ n9915 ^ n3068 ;
  assign n31406 = ( ~n2287 & n6656 ) | ( ~n2287 & n20517 ) | ( n6656 & n20517 ) ;
  assign n31407 = n31406 ^ n20490 ^ n19556 ;
  assign n31409 = n31408 ^ n31407 ^ n31210 ;
  assign n31410 = n31409 ^ n22735 ^ 1'b0 ;
  assign n31411 = n31405 | n31410 ;
  assign n31412 = ( x236 & n16050 ) | ( x236 & ~n23960 ) | ( n16050 & ~n23960 ) ;
  assign n31413 = n31412 ^ n26601 ^ n8240 ;
  assign n31414 = n26034 ^ n19445 ^ 1'b0 ;
  assign n31415 = ( ~n8670 & n20097 ) | ( ~n8670 & n31414 ) | ( n20097 & n31414 ) ;
  assign n31416 = ( n7066 & ~n20996 ) | ( n7066 & n31415 ) | ( ~n20996 & n31415 ) ;
  assign n31418 = ( n1700 & n13542 ) | ( n1700 & ~n28465 ) | ( n13542 & ~n28465 ) ;
  assign n31419 = n31418 ^ n16413 ^ n2122 ;
  assign n31420 = n31419 ^ n18544 ^ n13413 ;
  assign n31417 = ( n6455 & ~n15431 ) | ( n6455 & n20777 ) | ( ~n15431 & n20777 ) ;
  assign n31421 = n31420 ^ n31417 ^ n27485 ;
  assign n31422 = ( ~n2082 & n19729 ) | ( ~n2082 & n20679 ) | ( n19729 & n20679 ) ;
  assign n31423 = n12292 & ~n26302 ;
  assign n31424 = n31423 ^ n704 ^ 1'b0 ;
  assign n31425 = n31422 & ~n31424 ;
  assign n31426 = ~n14253 & n31425 ;
  assign n31428 = n20188 ^ n14692 ^ n9041 ;
  assign n31427 = n20326 ^ n16117 ^ n4858 ;
  assign n31429 = n31428 ^ n31427 ^ n21210 ;
  assign n31430 = n7855 ^ n3641 ^ n2612 ;
  assign n31431 = ( ~n15445 & n21013 ) | ( ~n15445 & n31430 ) | ( n21013 & n31430 ) ;
  assign n31432 = ( ~n983 & n14917 ) | ( ~n983 & n31431 ) | ( n14917 & n31431 ) ;
  assign n31433 = ( n21760 & ~n31429 ) | ( n21760 & n31432 ) | ( ~n31429 & n31432 ) ;
  assign n31435 = ( n8289 & n14805 ) | ( n8289 & n17942 ) | ( n14805 & n17942 ) ;
  assign n31434 = ( n10452 & ~n19451 ) | ( n10452 & n23885 ) | ( ~n19451 & n23885 ) ;
  assign n31436 = n31435 ^ n31434 ^ n10419 ;
  assign n31439 = ( n513 & n15282 ) | ( n513 & ~n17895 ) | ( n15282 & ~n17895 ) ;
  assign n31437 = ( n780 & n2447 ) | ( n780 & ~n10516 ) | ( n2447 & ~n10516 ) ;
  assign n31438 = n31437 ^ n25647 ^ n14440 ;
  assign n31440 = n31439 ^ n31438 ^ n11335 ;
  assign n31441 = ( ~n13317 & n23560 ) | ( ~n13317 & n31440 ) | ( n23560 & n31440 ) ;
  assign n31442 = n31441 ^ n25704 ^ n6631 ;
  assign n31443 = n21804 ^ n14423 ^ n939 ;
  assign n31444 = ( n932 & n6527 ) | ( n932 & ~n9673 ) | ( n6527 & ~n9673 ) ;
  assign n31445 = ( n9328 & n23138 ) | ( n9328 & ~n31444 ) | ( n23138 & ~n31444 ) ;
  assign n31446 = n31445 ^ n30163 ^ n28657 ;
  assign n31447 = n31446 ^ n9704 ^ n2074 ;
  assign n31448 = ( ~n10562 & n14661 ) | ( ~n10562 & n30911 ) | ( n14661 & n30911 ) ;
  assign n31449 = n31448 ^ n2532 ^ 1'b0 ;
  assign n31450 = n31449 ^ n28938 ^ n5261 ;
  assign n31451 = n11247 ^ n7418 ^ 1'b0 ;
  assign n31452 = n31451 ^ n31092 ^ n12103 ;
  assign n31453 = n27640 ^ n25852 ^ n20037 ;
  assign n31454 = ( ~n1169 & n21364 ) | ( ~n1169 & n30828 ) | ( n21364 & n30828 ) ;
  assign n31455 = n31454 ^ n27828 ^ n268 ;
  assign n31456 = ( n2773 & n11139 ) | ( n2773 & n30426 ) | ( n11139 & n30426 ) ;
  assign n31457 = n12125 | n20896 ;
  assign n31458 = ( n7077 & n11282 ) | ( n7077 & n26669 ) | ( n11282 & n26669 ) ;
  assign n31459 = n13017 ^ n6586 ^ 1'b0 ;
  assign n31460 = n31458 & n31459 ;
  assign n31461 = ~n31457 & n31460 ;
  assign n31462 = ( n10039 & ~n31456 ) | ( n10039 & n31461 ) | ( ~n31456 & n31461 ) ;
  assign n31463 = n27308 ^ n23592 ^ n5378 ;
  assign n31464 = ( n1280 & n5629 ) | ( n1280 & n15524 ) | ( n5629 & n15524 ) ;
  assign n31467 = ( n1763 & n22582 ) | ( n1763 & ~n23368 ) | ( n22582 & ~n23368 ) ;
  assign n31465 = n22612 ^ n14074 ^ 1'b0 ;
  assign n31466 = n31465 ^ n29085 ^ n16845 ;
  assign n31468 = n31467 ^ n31466 ^ n16299 ;
  assign n31469 = n13792 ^ n10192 ^ n1808 ;
  assign n31470 = n31469 ^ n22244 ^ n527 ;
  assign n31471 = n1205 & n6580 ;
  assign n31472 = n31471 ^ n6631 ^ 1'b0 ;
  assign n31473 = n8713 & ~n21252 ;
  assign n31474 = n31473 ^ n5801 ^ 1'b0 ;
  assign n31475 = n31472 & ~n31474 ;
  assign n31476 = n22299 ^ n11357 ^ n5654 ;
  assign n31477 = n31476 ^ n25048 ^ n2131 ;
  assign n31478 = n31477 ^ n28741 ^ 1'b0 ;
  assign n31479 = ~n31475 & n31478 ;
  assign n31480 = n11715 & ~n17533 ;
  assign n31481 = n18084 & n31480 ;
  assign n31482 = n24436 & ~n31481 ;
  assign n31483 = n31482 ^ n4924 ^ 1'b0 ;
  assign n31484 = n2523 ^ n824 ^ 1'b0 ;
  assign n31485 = ( ~n10114 & n24798 ) | ( ~n10114 & n31484 ) | ( n24798 & n31484 ) ;
  assign n31490 = n14975 | n22638 ;
  assign n31491 = n30013 & ~n31490 ;
  assign n31492 = ( n18306 & n27544 ) | ( n18306 & ~n31491 ) | ( n27544 & ~n31491 ) ;
  assign n31486 = n4871 & ~n9833 ;
  assign n31487 = ~n20818 & n31486 ;
  assign n31488 = n21166 ^ n12827 ^ n8055 ;
  assign n31489 = ( n1491 & n31487 ) | ( n1491 & ~n31488 ) | ( n31487 & ~n31488 ) ;
  assign n31493 = n31492 ^ n31489 ^ n3137 ;
  assign n31494 = ( n4212 & n9894 ) | ( n4212 & n14368 ) | ( n9894 & n14368 ) ;
  assign n31495 = n28747 ^ n26985 ^ 1'b0 ;
  assign n31496 = ( n15520 & n30050 ) | ( n15520 & n31495 ) | ( n30050 & n31495 ) ;
  assign n31497 = n31496 ^ n15719 ^ n2016 ;
  assign n31498 = n9968 | n15353 ;
  assign n31499 = n31498 ^ n7979 ^ 1'b0 ;
  assign n31500 = ( ~n10758 & n14008 ) | ( ~n10758 & n31499 ) | ( n14008 & n31499 ) ;
  assign n31501 = ( n6034 & n11552 ) | ( n6034 & ~n31500 ) | ( n11552 & ~n31500 ) ;
  assign n31502 = ( ~n2623 & n4882 ) | ( ~n2623 & n18252 ) | ( n4882 & n18252 ) ;
  assign n31503 = n31502 ^ n22174 ^ n21514 ;
  assign n31504 = n19953 & ~n24071 ;
  assign n31505 = ~n2512 & n31504 ;
  assign n31506 = n6238 | n19186 ;
  assign n31507 = ~n3117 & n6581 ;
  assign n31508 = ( n6369 & n7335 ) | ( n6369 & n20162 ) | ( n7335 & n20162 ) ;
  assign n31509 = n1159 & ~n31508 ;
  assign n31510 = n31509 ^ n2515 ^ n562 ;
  assign n31511 = x27 & ~n31510 ;
  assign n31512 = n31511 ^ n9352 ^ 1'b0 ;
  assign n31513 = ( n1263 & n27413 ) | ( n1263 & ~n31512 ) | ( n27413 & ~n31512 ) ;
  assign n31514 = n31513 ^ n6245 ^ n1041 ;
  assign n31517 = ( n3843 & n8065 ) | ( n3843 & ~n22985 ) | ( n8065 & ~n22985 ) ;
  assign n31518 = ( n3800 & n7234 ) | ( n3800 & ~n9718 ) | ( n7234 & ~n9718 ) ;
  assign n31519 = ( ~n24779 & n31517 ) | ( ~n24779 & n31518 ) | ( n31517 & n31518 ) ;
  assign n31515 = n27650 ^ n21055 ^ n5869 ;
  assign n31516 = n31515 ^ n30304 ^ n15530 ;
  assign n31520 = n31519 ^ n31516 ^ n4340 ;
  assign n31521 = ( ~n31507 & n31514 ) | ( ~n31507 & n31520 ) | ( n31514 & n31520 ) ;
  assign n31522 = ( n972 & n8447 ) | ( n972 & ~n28636 ) | ( n8447 & ~n28636 ) ;
  assign n31523 = n5975 & ~n31522 ;
  assign n31524 = n9472 & ~n31523 ;
  assign n31525 = n31524 ^ n20141 ^ 1'b0 ;
  assign n31526 = ~n1757 & n5364 ;
  assign n31527 = n3472 & n31526 ;
  assign n31528 = n5040 & n31527 ;
  assign n31529 = n31528 ^ n26343 ^ n9362 ;
  assign n31530 = n31529 ^ n21700 ^ x34 ;
  assign n31531 = ( ~n27287 & n28680 ) | ( ~n27287 & n31530 ) | ( n28680 & n31530 ) ;
  assign n31534 = n8235 ^ n7031 ^ n4018 ;
  assign n31532 = n17758 ^ n15969 ^ 1'b0 ;
  assign n31533 = n12757 & n31532 ;
  assign n31535 = n31534 ^ n31533 ^ n9781 ;
  assign n31536 = n16978 ^ n4931 ^ n2046 ;
  assign n31537 = n31334 ^ n13291 ^ n1417 ;
  assign n31538 = ( n12132 & n31536 ) | ( n12132 & n31537 ) | ( n31536 & n31537 ) ;
  assign n31539 = n18570 ^ n4551 ^ 1'b0 ;
  assign n31540 = ~n28002 & n31539 ;
  assign n31541 = n19037 ^ n16219 ^ n16202 ;
  assign n31542 = n16927 ^ n11769 ^ n10352 ;
  assign n31543 = n21954 ^ n11678 ^ 1'b0 ;
  assign n31545 = n22974 ^ n11160 ^ n6076 ;
  assign n31546 = n31545 ^ n914 ^ n502 ;
  assign n31544 = ( n1243 & n21769 ) | ( n1243 & n30852 ) | ( n21769 & n30852 ) ;
  assign n31547 = n31546 ^ n31544 ^ n7253 ;
  assign n31548 = n31547 ^ n1749 ^ 1'b0 ;
  assign n31549 = n26199 ^ n9870 ^ n8858 ;
  assign n31550 = n8722 & n10785 ;
  assign n31551 = n31550 ^ n23771 ^ n11618 ;
  assign n31552 = n31551 ^ n30633 ^ 1'b0 ;
  assign n31553 = n30385 & ~n31552 ;
  assign n31554 = ~n9907 & n25148 ;
  assign n31555 = n31554 ^ n1680 ^ 1'b0 ;
  assign n31556 = ( n5994 & ~n12407 ) | ( n5994 & n31555 ) | ( ~n12407 & n31555 ) ;
  assign n31560 = n24699 ^ n1591 ^ n857 ;
  assign n31557 = ( n2899 & n14358 ) | ( n2899 & n17395 ) | ( n14358 & n17395 ) ;
  assign n31558 = n12731 & ~n31557 ;
  assign n31559 = n31558 ^ n13829 ^ 1'b0 ;
  assign n31561 = n31560 ^ n31559 ^ n24005 ;
  assign n31562 = n7350 ^ n6205 ^ x120 ;
  assign n31563 = ( n10972 & n16255 ) | ( n10972 & ~n31562 ) | ( n16255 & ~n31562 ) ;
  assign n31564 = ( n3425 & n12765 ) | ( n3425 & ~n31563 ) | ( n12765 & ~n31563 ) ;
  assign n31565 = n16054 ^ x253 ^ 1'b0 ;
  assign n31566 = n25887 ^ n11815 ^ n3791 ;
  assign n31567 = ( n7696 & n17305 ) | ( n7696 & ~n24657 ) | ( n17305 & ~n24657 ) ;
  assign n31569 = n18272 ^ n17500 ^ n7473 ;
  assign n31568 = ( n11823 & n16321 ) | ( n11823 & n18657 ) | ( n16321 & n18657 ) ;
  assign n31570 = n31569 ^ n31568 ^ n13108 ;
  assign n31571 = ( n14355 & n31567 ) | ( n14355 & n31570 ) | ( n31567 & n31570 ) ;
  assign n31572 = n8558 & n31397 ;
  assign n31573 = ( n9412 & n14675 ) | ( n9412 & ~n31572 ) | ( n14675 & ~n31572 ) ;
  assign n31574 = n31573 ^ n16900 ^ n7066 ;
  assign n31575 = n31574 ^ n12482 ^ 1'b0 ;
  assign n31576 = x244 & ~n9955 ;
  assign n31577 = n2340 ^ n1775 ^ 1'b0 ;
  assign n31578 = n3735 | n31577 ;
  assign n31579 = ( n4864 & ~n31576 ) | ( n4864 & n31578 ) | ( ~n31576 & n31578 ) ;
  assign n31580 = n24176 ^ n11851 ^ 1'b0 ;
  assign n31582 = n13492 ^ n9987 ^ n9711 ;
  assign n31581 = ( n9846 & ~n10337 ) | ( n9846 & n11425 ) | ( ~n10337 & n11425 ) ;
  assign n31583 = n31582 ^ n31581 ^ n20894 ;
  assign n31584 = n31583 ^ n4846 ^ n4627 ;
  assign n31585 = ( ~n1583 & n5181 ) | ( ~n1583 & n25558 ) | ( n5181 & n25558 ) ;
  assign n31586 = n31585 ^ n24123 ^ n7895 ;
  assign n31588 = n2930 | n8230 ;
  assign n31589 = n4308 | n31588 ;
  assign n31587 = n26673 ^ n14835 ^ n10464 ;
  assign n31590 = n31589 ^ n31587 ^ 1'b0 ;
  assign n31591 = ( n17777 & n31586 ) | ( n17777 & ~n31590 ) | ( n31586 & ~n31590 ) ;
  assign n31592 = ( n2771 & n5406 ) | ( n2771 & ~n11393 ) | ( n5406 & ~n11393 ) ;
  assign n31593 = ( n1732 & n18891 ) | ( n1732 & n31592 ) | ( n18891 & n31592 ) ;
  assign n31595 = n20425 ^ n7783 ^ n2972 ;
  assign n31596 = n31595 ^ n29243 ^ n16302 ;
  assign n31597 = ( n2273 & n6686 ) | ( n2273 & ~n31596 ) | ( n6686 & ~n31596 ) ;
  assign n31594 = n6535 & ~n14135 ;
  assign n31598 = n31597 ^ n31594 ^ 1'b0 ;
  assign n31603 = ( n13856 & n14198 ) | ( n13856 & ~n31529 ) | ( n14198 & ~n31529 ) ;
  assign n31600 = ( n1222 & ~n2546 ) | ( n1222 & n5624 ) | ( ~n2546 & n5624 ) ;
  assign n31601 = n31600 ^ n7828 ^ n2086 ;
  assign n31599 = ( ~n774 & n10429 ) | ( ~n774 & n26792 ) | ( n10429 & n26792 ) ;
  assign n31602 = n31601 ^ n31599 ^ n29715 ;
  assign n31604 = n31603 ^ n31602 ^ n25629 ;
  assign n31605 = ( n2922 & n24550 ) | ( n2922 & n31604 ) | ( n24550 & n31604 ) ;
  assign n31607 = ( ~n3674 & n7347 ) | ( ~n3674 & n16130 ) | ( n7347 & n16130 ) ;
  assign n31608 = n31607 ^ n10404 ^ 1'b0 ;
  assign n31609 = n7170 & n31608 ;
  assign n31606 = n28131 ^ n9665 ^ n1343 ;
  assign n31610 = n31609 ^ n31606 ^ n22397 ;
  assign n31611 = n24726 ^ n13441 ^ n4463 ;
  assign n31612 = n8546 | n19659 ;
  assign n31613 = n31612 ^ n742 ^ 1'b0 ;
  assign n31614 = n31613 ^ n9328 ^ n5023 ;
  assign n31619 = n898 ^ x213 ^ x174 ;
  assign n31615 = n11854 ^ n8226 ^ n6482 ;
  assign n31616 = ( n11620 & n12068 ) | ( n11620 & ~n31615 ) | ( n12068 & ~n31615 ) ;
  assign n31617 = n9730 & ~n31616 ;
  assign n31618 = ( ~n27187 & n31126 ) | ( ~n27187 & n31617 ) | ( n31126 & n31617 ) ;
  assign n31620 = n31619 ^ n31618 ^ n5109 ;
  assign n31621 = ( ~n595 & n13383 ) | ( ~n595 & n19984 ) | ( n13383 & n19984 ) ;
  assign n31622 = ( n4285 & n10527 ) | ( n4285 & n31621 ) | ( n10527 & n31621 ) ;
  assign n31623 = ( n11522 & n12612 ) | ( n11522 & n31622 ) | ( n12612 & n31622 ) ;
  assign n31624 = n31623 ^ n29651 ^ n9971 ;
  assign n31625 = ( ~n5078 & n11672 ) | ( ~n5078 & n13664 ) | ( n11672 & n13664 ) ;
  assign n31626 = ( n2559 & n5821 ) | ( n2559 & n8146 ) | ( n5821 & n8146 ) ;
  assign n31627 = ~n13388 & n31626 ;
  assign n31628 = ( n16134 & n31625 ) | ( n16134 & n31627 ) | ( n31625 & n31627 ) ;
  assign n31629 = n5842 & ~n8148 ;
  assign n31630 = n31629 ^ n20973 ^ 1'b0 ;
  assign n31631 = n31630 ^ n29585 ^ n13771 ;
  assign n31632 = n16991 | n31631 ;
  assign n31633 = ( n3947 & ~n5027 ) | ( n3947 & n5601 ) | ( ~n5027 & n5601 ) ;
  assign n31634 = n31633 ^ n20293 ^ n13081 ;
  assign n31635 = n9030 ^ n2804 ^ n2466 ;
  assign n31636 = ( ~n12854 & n20090 ) | ( ~n12854 & n31635 ) | ( n20090 & n31635 ) ;
  assign n31637 = ( n7145 & n7333 ) | ( n7145 & ~n9410 ) | ( n7333 & ~n9410 ) ;
  assign n31638 = n10141 ^ n9755 ^ n6235 ;
  assign n31639 = ( n5804 & ~n31637 ) | ( n5804 & n31638 ) | ( ~n31637 & n31638 ) ;
  assign n31640 = n31639 ^ n24830 ^ n14662 ;
  assign n31641 = n31640 ^ n22133 ^ n1355 ;
  assign n31642 = n24090 ^ n23926 ^ n12876 ;
  assign n31643 = ( n12418 & ~n27442 ) | ( n12418 & n31642 ) | ( ~n27442 & n31642 ) ;
  assign n31644 = n26589 ^ n20997 ^ n9788 ;
  assign n31645 = n2018 & ~n31644 ;
  assign n31646 = ~n9892 & n31645 ;
  assign n31648 = ( n9347 & n17309 ) | ( n9347 & ~n29883 ) | ( n17309 & ~n29883 ) ;
  assign n31649 = n31648 ^ n25457 ^ n304 ;
  assign n31647 = n16567 ^ n6649 ^ 1'b0 ;
  assign n31650 = n31649 ^ n31647 ^ n21625 ;
  assign n31651 = n31650 ^ n5027 ^ 1'b0 ;
  assign n31652 = n27497 ^ n22545 ^ n17931 ;
  assign n31653 = n26580 ^ n6151 ^ n4091 ;
  assign n31654 = n31653 ^ n25863 ^ n25243 ;
  assign n31655 = n2559 | n12121 ;
  assign n31656 = ( n16614 & ~n31654 ) | ( n16614 & n31655 ) | ( ~n31654 & n31655 ) ;
  assign n31657 = n24311 ^ n23481 ^ n5099 ;
  assign n31658 = n31657 ^ n29456 ^ n17251 ;
  assign n31659 = ( ~n4893 & n12150 ) | ( ~n4893 & n31658 ) | ( n12150 & n31658 ) ;
  assign n31660 = n4849 ^ n1821 ^ 1'b0 ;
  assign n31661 = n31660 ^ n14435 ^ n3130 ;
  assign n31662 = n557 & ~n31661 ;
  assign n31663 = ( n7836 & n22694 ) | ( n7836 & ~n31662 ) | ( n22694 & ~n31662 ) ;
  assign n31666 = ( ~n758 & n11337 ) | ( ~n758 & n16129 ) | ( n11337 & n16129 ) ;
  assign n31664 = ( n1804 & n9966 ) | ( n1804 & n15304 ) | ( n9966 & n15304 ) ;
  assign n31665 = n31664 ^ n19163 ^ n7980 ;
  assign n31667 = n31666 ^ n31665 ^ n23721 ;
  assign n31668 = ( ~n6145 & n24760 ) | ( ~n6145 & n31667 ) | ( n24760 & n31667 ) ;
  assign n31669 = n24275 ^ n17946 ^ n16836 ;
  assign n31670 = ( ~n13655 & n23681 ) | ( ~n13655 & n31669 ) | ( n23681 & n31669 ) ;
  assign n31671 = n31668 | n31670 ;
  assign n31672 = n10087 | n10734 ;
  assign n31673 = n10793 & ~n31672 ;
  assign n31674 = ~n6706 & n31673 ;
  assign n31675 = ( n3140 & n10492 ) | ( n3140 & ~n10874 ) | ( n10492 & ~n10874 ) ;
  assign n31676 = n31675 ^ n20665 ^ n2526 ;
  assign n31677 = n31676 ^ n3370 ^ 1'b0 ;
  assign n31678 = ( n6145 & ~n15140 ) | ( n6145 & n25025 ) | ( ~n15140 & n25025 ) ;
  assign n31679 = n9924 ^ n639 ^ 1'b0 ;
  assign n31680 = ~n18779 & n31679 ;
  assign n31681 = ( ~n12660 & n22966 ) | ( ~n12660 & n31680 ) | ( n22966 & n31680 ) ;
  assign n31682 = ( ~n5255 & n23683 ) | ( ~n5255 & n31681 ) | ( n23683 & n31681 ) ;
  assign n31683 = n18721 ^ n5696 ^ n3801 ;
  assign n31684 = n6593 & n31683 ;
  assign n31685 = n31684 ^ n1928 ^ 1'b0 ;
  assign n31686 = ( n9934 & ~n14446 ) | ( n9934 & n31685 ) | ( ~n14446 & n31685 ) ;
  assign n31687 = n25842 ^ n19030 ^ 1'b0 ;
  assign n31688 = n31687 ^ n31381 ^ 1'b0 ;
  assign n31689 = n19501 ^ n3972 ^ 1'b0 ;
  assign n31693 = n6462 ^ n3614 ^ n1583 ;
  assign n31692 = ( n3256 & n7451 ) | ( n3256 & ~n29365 ) | ( n7451 & ~n29365 ) ;
  assign n31690 = ( n1855 & ~n11184 ) | ( n1855 & n17731 ) | ( ~n11184 & n17731 ) ;
  assign n31691 = n31690 ^ n5051 ^ n4819 ;
  assign n31694 = n31693 ^ n31692 ^ n31691 ;
  assign n31695 = ( n14203 & ~n31689 ) | ( n14203 & n31694 ) | ( ~n31689 & n31694 ) ;
  assign n31696 = n29087 ^ n2244 ^ 1'b0 ;
  assign n31697 = n17122 & n31696 ;
  assign n31698 = n31697 ^ n25095 ^ n12550 ;
  assign n31699 = ( ~n17328 & n17767 ) | ( ~n17328 & n23070 ) | ( n17767 & n23070 ) ;
  assign n31700 = n31699 ^ n25554 ^ n22837 ;
  assign n31701 = x160 & n14026 ;
  assign n31702 = n31701 ^ n29165 ^ 1'b0 ;
  assign n31703 = n7316 ^ n6667 ^ n3495 ;
  assign n31704 = n31703 ^ n18814 ^ 1'b0 ;
  assign n31705 = ~n31702 & n31704 ;
  assign n31707 = n16337 ^ n7497 ^ 1'b0 ;
  assign n31708 = n6610 | n31707 ;
  assign n31706 = n31586 ^ n24438 ^ n6517 ;
  assign n31709 = n31708 ^ n31706 ^ n23023 ;
  assign n31710 = n31709 ^ n23468 ^ n10418 ;
  assign n31711 = n16651 ^ n10705 ^ n6251 ;
  assign n31713 = n27558 ^ n19682 ^ n14009 ;
  assign n31712 = n16805 | n23178 ;
  assign n31714 = n31713 ^ n31712 ^ n31661 ;
  assign n31715 = n21002 ^ n12546 ^ 1'b0 ;
  assign n31716 = n16382 | n16765 ;
  assign n31717 = n18877 ^ n3050 ^ 1'b0 ;
  assign n31718 = n3409 | n31717 ;
  assign n31719 = ( n6816 & ~n8232 ) | ( n6816 & n18723 ) | ( ~n8232 & n18723 ) ;
  assign n31720 = ( n10451 & ~n31718 ) | ( n10451 & n31719 ) | ( ~n31718 & n31719 ) ;
  assign n31721 = ( n3297 & n12321 ) | ( n3297 & n31720 ) | ( n12321 & n31720 ) ;
  assign n31722 = ( n7627 & n18958 ) | ( n7627 & ~n31721 ) | ( n18958 & ~n31721 ) ;
  assign n31723 = n31716 | n31722 ;
  assign n31724 = n22819 ^ n14303 ^ n11511 ;
  assign n31725 = n31724 ^ n20299 ^ n7016 ;
  assign n31726 = n29904 ^ n984 ^ 1'b0 ;
  assign n31727 = n1806 & ~n31726 ;
  assign n31728 = n23282 ^ n8378 ^ 1'b0 ;
  assign n31729 = n17640 | n31728 ;
  assign n31730 = n814 & ~n31729 ;
  assign n31731 = ( n16626 & ~n31727 ) | ( n16626 & n31730 ) | ( ~n31727 & n31730 ) ;
  assign n31732 = n17016 & n19668 ;
  assign n31733 = n31732 ^ n30974 ^ 1'b0 ;
  assign n31737 = n3405 & n12868 ;
  assign n31738 = ~n31079 & n31737 ;
  assign n31734 = ( n1276 & n4698 ) | ( n1276 & n6468 ) | ( n4698 & n6468 ) ;
  assign n31735 = n31734 ^ n17110 ^ n9429 ;
  assign n31736 = n31735 ^ n20745 ^ n6213 ;
  assign n31739 = n31738 ^ n31736 ^ n2327 ;
  assign n31740 = ( ~n727 & n29345 ) | ( ~n727 & n31739 ) | ( n29345 & n31739 ) ;
  assign n31741 = ( ~n2833 & n13398 ) | ( ~n2833 & n23711 ) | ( n13398 & n23711 ) ;
  assign n31742 = n31741 ^ n21071 ^ n8405 ;
  assign n31743 = n31742 ^ n25006 ^ n15421 ;
  assign n31744 = n17291 ^ n3596 ^ n786 ;
  assign n31745 = n23528 ^ n16025 ^ n1975 ;
  assign n31746 = ( n10826 & ~n12348 ) | ( n10826 & n14175 ) | ( ~n12348 & n14175 ) ;
  assign n31747 = ( n31744 & n31745 ) | ( n31744 & n31746 ) | ( n31745 & n31746 ) ;
  assign n31748 = ( n3742 & ~n5374 ) | ( n3742 & n31747 ) | ( ~n5374 & n31747 ) ;
  assign n31749 = ( n7981 & ~n10636 ) | ( n7981 & n31748 ) | ( ~n10636 & n31748 ) ;
  assign n31750 = n3509 & n3564 ;
  assign n31751 = ( ~n4514 & n11405 ) | ( ~n4514 & n31750 ) | ( n11405 & n31750 ) ;
  assign n31752 = n31751 ^ n17481 ^ n6580 ;
  assign n31753 = n31752 ^ n27713 ^ n3255 ;
  assign n31754 = ( n1941 & n24527 ) | ( n1941 & ~n31753 ) | ( n24527 & ~n31753 ) ;
  assign n31755 = n31754 ^ n20293 ^ n13375 ;
  assign n31756 = ( n12460 & n12654 ) | ( n12460 & n25239 ) | ( n12654 & n25239 ) ;
  assign n31759 = n19025 ^ n18610 ^ 1'b0 ;
  assign n31760 = n9905 & n31759 ;
  assign n31761 = n31760 ^ n8998 ^ 1'b0 ;
  assign n31757 = n4346 & n12297 ;
  assign n31758 = n31757 ^ n18651 ^ n14719 ;
  assign n31762 = n31761 ^ n31758 ^ n8533 ;
  assign n31763 = ( n5391 & n10893 ) | ( n5391 & n30074 ) | ( n10893 & n30074 ) ;
  assign n31764 = n28778 ^ n26698 ^ 1'b0 ;
  assign n31765 = n31764 ^ n13141 ^ n5612 ;
  assign n31766 = ( n17652 & n18304 ) | ( n17652 & ~n26963 ) | ( n18304 & ~n26963 ) ;
  assign n31771 = n26349 ^ n13353 ^ n9471 ;
  assign n31768 = ( n2255 & ~n3059 ) | ( n2255 & n3458 ) | ( ~n3059 & n3458 ) ;
  assign n31769 = n8553 & n31768 ;
  assign n31770 = n31769 ^ n3151 ^ 1'b0 ;
  assign n31767 = n25822 ^ n18868 ^ n15349 ;
  assign n31772 = n31771 ^ n31770 ^ n31767 ;
  assign n31776 = n18373 ^ n13561 ^ n8208 ;
  assign n31773 = ( n2190 & n10181 ) | ( n2190 & n15508 ) | ( n10181 & n15508 ) ;
  assign n31774 = n29425 ^ n2237 ^ 1'b0 ;
  assign n31775 = ( ~n5204 & n31773 ) | ( ~n5204 & n31774 ) | ( n31773 & n31774 ) ;
  assign n31777 = n31776 ^ n31775 ^ n14859 ;
  assign n31779 = n28137 ^ n8257 ^ n7905 ;
  assign n31780 = ~n8765 & n31779 ;
  assign n31778 = ( n8097 & n22992 ) | ( n8097 & n23576 ) | ( n22992 & n23576 ) ;
  assign n31781 = n31780 ^ n31778 ^ n19288 ;
  assign n31782 = n18224 ^ n5024 ^ n2036 ;
  assign n31783 = ( x82 & ~n4583 ) | ( x82 & n10711 ) | ( ~n4583 & n10711 ) ;
  assign n31784 = n31783 ^ n20977 ^ n2107 ;
  assign n31785 = ( n1408 & n31782 ) | ( n1408 & n31784 ) | ( n31782 & n31784 ) ;
  assign n31786 = n9968 ^ n8721 ^ n2698 ;
  assign n31787 = n24732 ^ n17122 ^ n3835 ;
  assign n31788 = n8189 ^ n6400 ^ n2945 ;
  assign n31789 = n31788 ^ n12143 ^ 1'b0 ;
  assign n31790 = ( ~n31786 & n31787 ) | ( ~n31786 & n31789 ) | ( n31787 & n31789 ) ;
  assign n31791 = ( ~n9772 & n11089 ) | ( ~n9772 & n17705 ) | ( n11089 & n17705 ) ;
  assign n31792 = n30579 ^ n27544 ^ 1'b0 ;
  assign n31793 = n31791 & ~n31792 ;
  assign n31794 = n31793 ^ n24206 ^ n10161 ;
  assign n31795 = ( x158 & n8576 ) | ( x158 & ~n31794 ) | ( n8576 & ~n31794 ) ;
  assign n31796 = n16103 ^ n12341 ^ n9167 ;
  assign n31797 = n31796 ^ n17255 ^ n9796 ;
  assign n31798 = n4414 ^ n2796 ^ 1'b0 ;
  assign n31799 = n9950 & ~n31798 ;
  assign n31800 = n26731 ^ n21712 ^ n18005 ;
  assign n31801 = ( n29556 & n31799 ) | ( n29556 & ~n31800 ) | ( n31799 & ~n31800 ) ;
  assign n31804 = ~n679 & n14082 ;
  assign n31805 = ~n9796 & n31804 ;
  assign n31802 = n12783 ^ n9364 ^ n993 ;
  assign n31803 = n31802 ^ n22411 ^ n6955 ;
  assign n31806 = n31805 ^ n31803 ^ n3539 ;
  assign n31807 = ( n1737 & ~n3182 ) | ( n1737 & n13272 ) | ( ~n3182 & n13272 ) ;
  assign n31808 = ( n3303 & ~n24775 ) | ( n3303 & n31807 ) | ( ~n24775 & n31807 ) ;
  assign n31809 = ( n5253 & ~n20694 ) | ( n5253 & n31808 ) | ( ~n20694 & n31808 ) ;
  assign n31810 = ( n2114 & n3237 ) | ( n2114 & n9081 ) | ( n3237 & n9081 ) ;
  assign n31812 = ( n2850 & ~n3036 ) | ( n2850 & n11006 ) | ( ~n3036 & n11006 ) ;
  assign n31811 = n1258 ^ x199 ^ 1'b0 ;
  assign n31813 = n31812 ^ n31811 ^ n22750 ;
  assign n31814 = ( n14859 & ~n31810 ) | ( n14859 & n31813 ) | ( ~n31810 & n31813 ) ;
  assign n31815 = n18033 ^ n4096 ^ n1359 ;
  assign n31816 = n25752 ^ n12153 ^ 1'b0 ;
  assign n31817 = n31815 | n31816 ;
  assign n31818 = ( n6231 & ~n16882 ) | ( n6231 & n27292 ) | ( ~n16882 & n27292 ) ;
  assign n31819 = x141 & ~n24145 ;
  assign n31820 = ~n3245 & n31819 ;
  assign n31821 = n11648 | n31820 ;
  assign n31822 = n31821 ^ n14214 ^ 1'b0 ;
  assign n31823 = n2113 | n31822 ;
  assign n31824 = n10320 | n11962 ;
  assign n31825 = n27737 & n31824 ;
  assign n31826 = ( ~n29435 & n31823 ) | ( ~n29435 & n31825 ) | ( n31823 & n31825 ) ;
  assign n31827 = n29503 ^ n23512 ^ n22073 ;
  assign n31828 = n12359 ^ n6552 ^ 1'b0 ;
  assign n31829 = n10556 & n30118 ;
  assign n31830 = ( n8922 & n22330 ) | ( n8922 & ~n27914 ) | ( n22330 & ~n27914 ) ;
  assign n31831 = ( ~n1634 & n24606 ) | ( ~n1634 & n31830 ) | ( n24606 & n31830 ) ;
  assign n31832 = ~n6066 & n24845 ;
  assign n31833 = ~n24193 & n31832 ;
  assign n31834 = ( ~n5231 & n9750 ) | ( ~n5231 & n12224 ) | ( n9750 & n12224 ) ;
  assign n31835 = n31834 ^ n28541 ^ n24420 ;
  assign n31839 = n7626 ^ x221 ^ 1'b0 ;
  assign n31840 = ( n13160 & ~n28872 ) | ( n13160 & n31839 ) | ( ~n28872 & n31839 ) ;
  assign n31837 = n4794 ^ n1949 ^ x121 ;
  assign n31838 = n31837 ^ n24815 ^ n8892 ;
  assign n31836 = n7740 & n28962 ;
  assign n31841 = n31840 ^ n31838 ^ n31836 ;
  assign n31842 = ( ~n18586 & n21661 ) | ( ~n18586 & n21920 ) | ( n21661 & n21920 ) ;
  assign n31843 = ( n6191 & ~n19749 ) | ( n6191 & n25061 ) | ( ~n19749 & n25061 ) ;
  assign n31844 = ( n355 & n16428 ) | ( n355 & n23223 ) | ( n16428 & n23223 ) ;
  assign n31845 = n31844 ^ n24893 ^ n17412 ;
  assign n31846 = n12420 ^ n3675 ^ n2216 ;
  assign n31847 = ( ~n13387 & n14793 ) | ( ~n13387 & n31846 ) | ( n14793 & n31846 ) ;
  assign n31848 = n25590 ^ n11937 ^ 1'b0 ;
  assign n31849 = n10264 & n31848 ;
  assign n31850 = n31849 ^ n25691 ^ n11460 ;
  assign n31851 = n20537 ^ n2233 ^ 1'b0 ;
  assign n31852 = n21127 ^ n5208 ^ 1'b0 ;
  assign n31853 = n18260 & ~n31852 ;
  assign n31854 = ( ~n865 & n31851 ) | ( ~n865 & n31853 ) | ( n31851 & n31853 ) ;
  assign n31855 = ( n13192 & n14442 ) | ( n13192 & ~n17563 ) | ( n14442 & ~n17563 ) ;
  assign n31856 = ( n14871 & ~n20088 ) | ( n14871 & n31855 ) | ( ~n20088 & n31855 ) ;
  assign n31857 = ~n12996 & n31856 ;
  assign n31858 = n7829 ^ n547 ^ n532 ;
  assign n31859 = ( ~n12484 & n31857 ) | ( ~n12484 & n31858 ) | ( n31857 & n31858 ) ;
  assign n31860 = ( ~n2192 & n14091 ) | ( ~n2192 & n20953 ) | ( n14091 & n20953 ) ;
  assign n31861 = ( n9280 & ~n23124 ) | ( n9280 & n31655 ) | ( ~n23124 & n31655 ) ;
  assign n31862 = ( n23659 & n31860 ) | ( n23659 & ~n31861 ) | ( n31860 & ~n31861 ) ;
  assign n31863 = n10663 ^ n3534 ^ n1902 ;
  assign n31864 = n21178 ^ n8179 ^ n3042 ;
  assign n31865 = ( n544 & n16072 ) | ( n544 & n31864 ) | ( n16072 & n31864 ) ;
  assign n31866 = ( n15768 & n18133 ) | ( n15768 & ~n31865 ) | ( n18133 & ~n31865 ) ;
  assign n31867 = ( n18719 & n31863 ) | ( n18719 & ~n31866 ) | ( n31863 & ~n31866 ) ;
  assign n31868 = n22621 ^ n10039 ^ n5307 ;
  assign n31869 = n31868 ^ n29344 ^ n9530 ;
  assign n31870 = n4019 | n31869 ;
  assign n31871 = n13285 ^ n11567 ^ n1423 ;
  assign n31872 = ( n2506 & ~n27478 ) | ( n2506 & n31871 ) | ( ~n27478 & n31871 ) ;
  assign n31873 = n31872 ^ n20830 ^ n3932 ;
  assign n31874 = ( n909 & n990 ) | ( n909 & n28450 ) | ( n990 & n28450 ) ;
  assign n31875 = n25153 ^ n13388 ^ n1132 ;
  assign n31876 = n30455 ^ n14805 ^ n4638 ;
  assign n31877 = ( n29259 & n31875 ) | ( n29259 & n31876 ) | ( n31875 & n31876 ) ;
  assign n31879 = ( n5419 & ~n10457 ) | ( n5419 & n10564 ) | ( ~n10457 & n10564 ) ;
  assign n31878 = n4104 & ~n26413 ;
  assign n31880 = n31879 ^ n31878 ^ n27861 ;
  assign n31883 = n9425 | n27283 ;
  assign n31884 = n31883 ^ n20054 ^ 1'b0 ;
  assign n31881 = ( n22980 & n23480 ) | ( n22980 & n23929 ) | ( n23480 & n23929 ) ;
  assign n31882 = ( n4420 & n20789 ) | ( n4420 & ~n31881 ) | ( n20789 & ~n31881 ) ;
  assign n31885 = n31884 ^ n31882 ^ n4693 ;
  assign n31886 = ( ~n3571 & n5253 ) | ( ~n3571 & n13258 ) | ( n5253 & n13258 ) ;
  assign n31887 = n31886 ^ n10136 ^ n9869 ;
  assign n31888 = n4374 & n13270 ;
  assign n31889 = n31887 & n31888 ;
  assign n31890 = ( n3052 & n8027 ) | ( n3052 & n8056 ) | ( n8027 & n8056 ) ;
  assign n31891 = ( ~n2127 & n8668 ) | ( ~n2127 & n31890 ) | ( n8668 & n31890 ) ;
  assign n31892 = n13063 ^ n8819 ^ n6509 ;
  assign n31893 = ( ~n427 & n20126 ) | ( ~n427 & n31892 ) | ( n20126 & n31892 ) ;
  assign n31894 = n30682 ^ n10502 ^ n1401 ;
  assign n31897 = ( n5611 & ~n8505 ) | ( n5611 & n11871 ) | ( ~n8505 & n11871 ) ;
  assign n31895 = ~n6769 & n11159 ;
  assign n31896 = n24557 & n31895 ;
  assign n31898 = n31897 ^ n31896 ^ n10948 ;
  assign n31899 = n20252 ^ n19453 ^ n341 ;
  assign n31900 = n31899 ^ n13928 ^ n3428 ;
  assign n31901 = ( n3065 & n12855 ) | ( n3065 & ~n19178 ) | ( n12855 & ~n19178 ) ;
  assign n31902 = ( ~n1662 & n6323 ) | ( ~n1662 & n31901 ) | ( n6323 & n31901 ) ;
  assign n31903 = n9339 & ~n31902 ;
  assign n31904 = ~n30134 & n31903 ;
  assign n31905 = n25343 ^ n22937 ^ x49 ;
  assign n31906 = ( ~n5619 & n6589 ) | ( ~n5619 & n31905 ) | ( n6589 & n31905 ) ;
  assign n31907 = ( n3278 & n21253 ) | ( n3278 & n21563 ) | ( n21253 & n21563 ) ;
  assign n31908 = ( n1409 & n11130 ) | ( n1409 & n31907 ) | ( n11130 & n31907 ) ;
  assign n31909 = n1571 & n2449 ;
  assign n31910 = ( n4961 & n22029 ) | ( n4961 & n31909 ) | ( n22029 & n31909 ) ;
  assign n31911 = ( n1401 & n6321 ) | ( n1401 & n10175 ) | ( n6321 & n10175 ) ;
  assign n31912 = n25678 ^ n2516 ^ 1'b0 ;
  assign n31913 = ~n5809 & n31912 ;
  assign n31917 = n2753 | n7098 ;
  assign n31918 = n4844 & ~n31917 ;
  assign n31914 = ( n863 & ~n2256 ) | ( n863 & n3158 ) | ( ~n2256 & n3158 ) ;
  assign n31915 = ( n6825 & n14818 ) | ( n6825 & ~n31914 ) | ( n14818 & ~n31914 ) ;
  assign n31916 = n31915 ^ n28619 ^ n28531 ;
  assign n31919 = n31918 ^ n31916 ^ n19848 ;
  assign n31925 = n21675 ^ n9988 ^ n2685 ;
  assign n31920 = n18785 ^ n11180 ^ n5779 ;
  assign n31921 = ~n7265 & n26396 ;
  assign n31922 = n31921 ^ n3915 ^ 1'b0 ;
  assign n31923 = n10650 | n17103 ;
  assign n31924 = ( n31920 & ~n31922 ) | ( n31920 & n31923 ) | ( ~n31922 & n31923 ) ;
  assign n31926 = n31925 ^ n31924 ^ x0 ;
  assign n31927 = n21633 ^ n10305 ^ n5125 ;
  assign n31928 = ~n4246 & n15712 ;
  assign n31929 = n31928 ^ n21954 ^ n20373 ;
  assign n31930 = ( ~n28950 & n31927 ) | ( ~n28950 & n31929 ) | ( n31927 & n31929 ) ;
  assign n31931 = n18247 ^ n5164 ^ n258 ;
  assign n31932 = n11367 ^ n9707 ^ n3491 ;
  assign n31933 = ( n4494 & ~n11614 ) | ( n4494 & n20551 ) | ( ~n11614 & n20551 ) ;
  assign n31934 = n26917 & n31933 ;
  assign n31935 = n31934 ^ n7359 ^ 1'b0 ;
  assign n31936 = ( n11155 & ~n17259 ) | ( n11155 & n31935 ) | ( ~n17259 & n31935 ) ;
  assign n31937 = n26061 ^ n16668 ^ n12876 ;
  assign n31938 = n24827 & n31937 ;
  assign n31939 = n31936 | n31938 ;
  assign n31940 = n951 & n7833 ;
  assign n31941 = n30530 ^ n13843 ^ 1'b0 ;
  assign n31942 = ( ~n9900 & n31940 ) | ( ~n9900 & n31941 ) | ( n31940 & n31941 ) ;
  assign n31943 = n31815 ^ n24409 ^ n8945 ;
  assign n31944 = ( ~n4948 & n12497 ) | ( ~n4948 & n18125 ) | ( n12497 & n18125 ) ;
  assign n31945 = ( n5516 & ~n11869 ) | ( n5516 & n14460 ) | ( ~n11869 & n14460 ) ;
  assign n31946 = ( ~n11276 & n11280 ) | ( ~n11276 & n12545 ) | ( n11280 & n12545 ) ;
  assign n31947 = n31946 ^ n19847 ^ n12306 ;
  assign n31948 = n31947 ^ n7137 ^ n4349 ;
  assign n31951 = ( n13233 & n14540 ) | ( n13233 & n16975 ) | ( n14540 & n16975 ) ;
  assign n31949 = n6118 ^ n4387 ^ n874 ;
  assign n31950 = n31949 ^ n3395 ^ 1'b0 ;
  assign n31952 = n31951 ^ n31950 ^ 1'b0 ;
  assign n31953 = ( n2369 & ~n16081 ) | ( n2369 & n17201 ) | ( ~n16081 & n17201 ) ;
  assign n31954 = ( n17240 & n29837 ) | ( n17240 & n31953 ) | ( n29837 & n31953 ) ;
  assign n31955 = ( n27283 & n30578 ) | ( n27283 & ~n31954 ) | ( n30578 & ~n31954 ) ;
  assign n31956 = ( n1080 & n5970 ) | ( n1080 & n31955 ) | ( n5970 & n31955 ) ;
  assign n31958 = ( n6222 & n13175 ) | ( n6222 & ~n16602 ) | ( n13175 & ~n16602 ) ;
  assign n31957 = n24568 | n25015 ;
  assign n31959 = n31958 ^ n31957 ^ 1'b0 ;
  assign n31960 = n31959 ^ n19232 ^ x238 ;
  assign n31963 = n7818 & n17718 ;
  assign n31964 = n31963 ^ n23707 ^ 1'b0 ;
  assign n31965 = ( n14844 & n15078 ) | ( n14844 & ~n31964 ) | ( n15078 & ~n31964 ) ;
  assign n31961 = ( n10555 & ~n17758 ) | ( n10555 & n29256 ) | ( ~n17758 & n29256 ) ;
  assign n31962 = n31961 ^ n26065 ^ n895 ;
  assign n31966 = n31965 ^ n31962 ^ n17668 ;
  assign n31967 = ( n22906 & n31960 ) | ( n22906 & n31966 ) | ( n31960 & n31966 ) ;
  assign n31968 = ~n7323 & n26329 ;
  assign n31969 = n31968 ^ n9895 ^ 1'b0 ;
  assign n31970 = n31969 ^ n5935 ^ n3618 ;
  assign n31971 = n21254 ^ n7010 ^ 1'b0 ;
  assign n31972 = ( n8060 & n9368 ) | ( n8060 & ~n21327 ) | ( n9368 & ~n21327 ) ;
  assign n31973 = ( n16606 & n20684 ) | ( n16606 & n31972 ) | ( n20684 & n31972 ) ;
  assign n31974 = ( n4427 & n31971 ) | ( n4427 & ~n31973 ) | ( n31971 & ~n31973 ) ;
  assign n31975 = n28576 ^ n18525 ^ n6976 ;
  assign n31979 = n12550 ^ n10760 ^ n1409 ;
  assign n31980 = n31979 ^ n22550 ^ n18473 ;
  assign n31976 = ( n320 & n3172 ) | ( n320 & n8070 ) | ( n3172 & n8070 ) ;
  assign n31977 = ( n2506 & ~n28692 ) | ( n2506 & n31976 ) | ( ~n28692 & n31976 ) ;
  assign n31978 = ( n11485 & n13640 ) | ( n11485 & n31977 ) | ( n13640 & n31977 ) ;
  assign n31981 = n31980 ^ n31978 ^ n5247 ;
  assign n31983 = ( n2144 & n2641 ) | ( n2144 & ~n22567 ) | ( n2641 & ~n22567 ) ;
  assign n31982 = n26356 ^ n12901 ^ n9232 ;
  assign n31984 = n31983 ^ n31982 ^ n11619 ;
  assign n31985 = n27255 ^ n10633 ^ 1'b0 ;
  assign n31986 = ( n555 & n23232 ) | ( n555 & n31985 ) | ( n23232 & n31985 ) ;
  assign n31987 = n31986 ^ n13504 ^ n12048 ;
  assign n31988 = n1741 ^ n1712 ^ 1'b0 ;
  assign n31989 = ( n10822 & n31987 ) | ( n10822 & n31988 ) | ( n31987 & n31988 ) ;
  assign n31990 = n12294 & n31989 ;
  assign n31991 = ( n13894 & ~n15208 ) | ( n13894 & n24384 ) | ( ~n15208 & n24384 ) ;
  assign n31992 = ( n3840 & n14001 ) | ( n3840 & n20985 ) | ( n14001 & n20985 ) ;
  assign n31993 = ( n31799 & n31991 ) | ( n31799 & ~n31992 ) | ( n31991 & ~n31992 ) ;
  assign n31994 = n27385 ^ n5053 ^ n4013 ;
  assign n31995 = n31994 ^ n23328 ^ n2925 ;
  assign n31996 = n1640 | n11005 ;
  assign n31997 = n5297 | n31996 ;
  assign n31998 = n23122 ^ n21346 ^ 1'b0 ;
  assign n31999 = ( n1041 & ~n3222 ) | ( n1041 & n13261 ) | ( ~n3222 & n13261 ) ;
  assign n32000 = n31999 ^ n6381 ^ n1056 ;
  assign n32001 = ( n31997 & n31998 ) | ( n31997 & ~n32000 ) | ( n31998 & ~n32000 ) ;
  assign n32004 = n6004 ^ n5959 ^ 1'b0 ;
  assign n32005 = ~n23042 & n32004 ;
  assign n32006 = n29250 & n32005 ;
  assign n32002 = n2304 | n9828 ;
  assign n32003 = n11041 | n32002 ;
  assign n32007 = n32006 ^ n32003 ^ n30295 ;
  assign n32008 = n29827 ^ n25471 ^ n2117 ;
  assign n32009 = n4337 ^ n3962 ^ n1752 ;
  assign n32010 = n32009 ^ n11135 ^ n6885 ;
  assign n32011 = n15922 ^ n4067 ^ n3168 ;
  assign n32012 = ( n485 & n10549 ) | ( n485 & ~n11083 ) | ( n10549 & ~n11083 ) ;
  assign n32013 = n32012 ^ n1103 ^ 1'b0 ;
  assign n32014 = ( ~n2271 & n4941 ) | ( ~n2271 & n5768 ) | ( n4941 & n5768 ) ;
  assign n32017 = ( n3826 & n15001 ) | ( n3826 & n29462 ) | ( n15001 & n29462 ) ;
  assign n32015 = ( n1805 & n1928 ) | ( n1805 & n6908 ) | ( n1928 & n6908 ) ;
  assign n32016 = n6081 & n32015 ;
  assign n32018 = n32017 ^ n32016 ^ 1'b0 ;
  assign n32019 = n5115 | n24212 ;
  assign n32020 = n32019 ^ n28147 ^ n19511 ;
  assign n32021 = n6234 | n32020 ;
  assign n32022 = n32021 ^ n30747 ^ 1'b0 ;
  assign n32024 = n20401 ^ n6674 ^ 1'b0 ;
  assign n32025 = n19695 & ~n32024 ;
  assign n32026 = ( n7477 & n12387 ) | ( n7477 & ~n32025 ) | ( n12387 & ~n32025 ) ;
  assign n32023 = n10320 | n14743 ;
  assign n32027 = n32026 ^ n32023 ^ 1'b0 ;
  assign n32028 = ( n7971 & ~n27080 ) | ( n7971 & n32027 ) | ( ~n27080 & n32027 ) ;
  assign n32029 = ( ~n32018 & n32022 ) | ( ~n32018 & n32028 ) | ( n32022 & n32028 ) ;
  assign n32030 = n32014 & ~n32029 ;
  assign n32031 = n7110 & n9527 ;
  assign n32032 = ~n6975 & n32031 ;
  assign n32033 = ( n6625 & n15559 ) | ( n6625 & ~n18349 ) | ( n15559 & ~n18349 ) ;
  assign n32034 = ( ~n300 & n7102 ) | ( ~n300 & n10786 ) | ( n7102 & n10786 ) ;
  assign n32035 = n5672 ^ n1232 ^ 1'b0 ;
  assign n32036 = n265 & n31653 ;
  assign n32037 = ~n21650 & n32036 ;
  assign n32038 = n28405 ^ n18253 ^ n16359 ;
  assign n32039 = n32038 ^ n20141 ^ n9813 ;
  assign n32040 = n9786 ^ n4462 ^ 1'b0 ;
  assign n32041 = n10079 ^ n4288 ^ 1'b0 ;
  assign n32042 = n19121 & ~n32041 ;
  assign n32043 = n32042 ^ n18107 ^ 1'b0 ;
  assign n32044 = ( n1811 & n32040 ) | ( n1811 & ~n32043 ) | ( n32040 & ~n32043 ) ;
  assign n32045 = ( n28906 & n32039 ) | ( n28906 & n32044 ) | ( n32039 & n32044 ) ;
  assign n32046 = n20417 ^ n15526 ^ n8232 ;
  assign n32047 = n32046 ^ n11048 ^ n4331 ;
  assign n32048 = n32047 ^ n24386 ^ n10272 ;
  assign n32049 = n1350 & ~n4832 ;
  assign n32050 = ( n424 & n7724 ) | ( n424 & ~n12247 ) | ( n7724 & ~n12247 ) ;
  assign n32051 = n2089 | n16607 ;
  assign n32052 = n32051 ^ n1226 ^ 1'b0 ;
  assign n32053 = n32052 ^ n31637 ^ n13971 ;
  assign n32054 = ( n4127 & n4156 ) | ( n4127 & ~n4863 ) | ( n4156 & ~n4863 ) ;
  assign n32055 = n10062 ^ n7029 ^ 1'b0 ;
  assign n32056 = ( ~n32053 & n32054 ) | ( ~n32053 & n32055 ) | ( n32054 & n32055 ) ;
  assign n32057 = n32056 ^ n29845 ^ n11237 ;
  assign n32058 = ( n25416 & ~n32050 ) | ( n25416 & n32057 ) | ( ~n32050 & n32057 ) ;
  assign n32059 = ( n569 & n10305 ) | ( n569 & n11063 ) | ( n10305 & n11063 ) ;
  assign n32060 = n32059 ^ n14604 ^ n14219 ;
  assign n32061 = n30291 ^ n25803 ^ n14271 ;
  assign n32062 = n29442 ^ n20547 ^ 1'b0 ;
  assign n32063 = n11958 | n32062 ;
  assign n32064 = n32063 ^ n7288 ^ n4428 ;
  assign n32065 = n32064 ^ n30317 ^ 1'b0 ;
  assign n32066 = n24083 ^ n15990 ^ n6782 ;
  assign n32067 = n32066 ^ n31458 ^ n27583 ;
  assign n32068 = n22252 ^ n1797 ^ n663 ;
  assign n32069 = ( n756 & n17000 ) | ( n756 & ~n21061 ) | ( n17000 & ~n21061 ) ;
  assign n32070 = ( ~n9106 & n16970 ) | ( ~n9106 & n32069 ) | ( n16970 & n32069 ) ;
  assign n32071 = ( n22313 & n23708 ) | ( n22313 & ~n32070 ) | ( n23708 & ~n32070 ) ;
  assign n32072 = ( n24961 & n25687 ) | ( n24961 & n31209 ) | ( n25687 & n31209 ) ;
  assign n32073 = n32072 ^ n18750 ^ n8776 ;
  assign n32074 = ( ~n22402 & n27056 ) | ( ~n22402 & n32073 ) | ( n27056 & n32073 ) ;
  assign n32077 = n15413 ^ n916 ^ n702 ;
  assign n32075 = n30483 ^ n20035 ^ n19272 ;
  assign n32076 = n32075 ^ n8331 ^ n1003 ;
  assign n32078 = n32077 ^ n32076 ^ 1'b0 ;
  assign n32079 = ( n6033 & ~n8522 ) | ( n6033 & n14344 ) | ( ~n8522 & n14344 ) ;
  assign n32080 = n32079 ^ n29556 ^ 1'b0 ;
  assign n32081 = n19140 & n32080 ;
  assign n32082 = ( n11493 & n30374 ) | ( n11493 & n32081 ) | ( n30374 & n32081 ) ;
  assign n32083 = n14411 | n32082 ;
  assign n32084 = n32083 ^ n13903 ^ 1'b0 ;
  assign n32085 = n32084 ^ n13720 ^ n4860 ;
  assign n32086 = n25696 ^ n13094 ^ 1'b0 ;
  assign n32087 = ~n25335 & n32086 ;
  assign n32088 = n32087 ^ n27931 ^ n19452 ;
  assign n32093 = ( n11304 & ~n20988 ) | ( n11304 & n26654 ) | ( ~n20988 & n26654 ) ;
  assign n32094 = n20459 ^ n12619 ^ 1'b0 ;
  assign n32095 = ~n22204 & n32094 ;
  assign n32096 = ( n9224 & n32093 ) | ( n9224 & ~n32095 ) | ( n32093 & ~n32095 ) ;
  assign n32089 = ( n5536 & ~n11939 ) | ( n5536 & n22300 ) | ( ~n11939 & n22300 ) ;
  assign n32090 = n1933 | n16568 ;
  assign n32091 = n32089 | n32090 ;
  assign n32092 = ( n5943 & n14205 ) | ( n5943 & ~n32091 ) | ( n14205 & ~n32091 ) ;
  assign n32097 = n32096 ^ n32092 ^ n4076 ;
  assign n32098 = ( n4632 & ~n6537 ) | ( n4632 & n9071 ) | ( ~n6537 & n9071 ) ;
  assign n32099 = n6462 ^ n4979 ^ n966 ;
  assign n32100 = ( n341 & ~n1544 ) | ( n341 & n32099 ) | ( ~n1544 & n32099 ) ;
  assign n32101 = n1977 & ~n32100 ;
  assign n32102 = ~n32098 & n32101 ;
  assign n32103 = n32102 ^ n21379 ^ n14914 ;
  assign n32105 = ( n768 & n1102 ) | ( n768 & n2550 ) | ( n1102 & n2550 ) ;
  assign n32104 = ~n3710 & n14459 ;
  assign n32106 = n32105 ^ n32104 ^ 1'b0 ;
  assign n32107 = n16148 ^ n7642 ^ n3575 ;
  assign n32108 = n32107 ^ n29002 ^ n2781 ;
  assign n32109 = n32108 ^ n27818 ^ n5636 ;
  assign n32110 = n11865 ^ n9713 ^ 1'b0 ;
  assign n32111 = n29358 & n32110 ;
  assign n32112 = n32111 ^ n3391 ^ n2975 ;
  assign n32113 = ( n3966 & n12456 ) | ( n3966 & ~n14050 ) | ( n12456 & ~n14050 ) ;
  assign n32114 = n19306 ^ n13663 ^ n6285 ;
  assign n32115 = n29683 ^ n10808 ^ n4663 ;
  assign n32116 = ( ~n32113 & n32114 ) | ( ~n32113 & n32115 ) | ( n32114 & n32115 ) ;
  assign n32117 = ( n6237 & n10426 ) | ( n6237 & ~n32116 ) | ( n10426 & ~n32116 ) ;
  assign n32118 = n5001 & ~n28858 ;
  assign n32119 = n8495 & n32118 ;
  assign n32120 = n15126 ^ n12231 ^ n1548 ;
  assign n32121 = n32120 ^ n24969 ^ n14663 ;
  assign n32122 = n18604 ^ n11242 ^ n2804 ;
  assign n32125 = n30605 ^ n26035 ^ n21008 ;
  assign n32123 = n4379 ^ n4015 ^ 1'b0 ;
  assign n32124 = n22496 & ~n32123 ;
  assign n32126 = n32125 ^ n32124 ^ n7348 ;
  assign n32127 = n21449 ^ n15286 ^ 1'b0 ;
  assign n32128 = n11464 & n32127 ;
  assign n32129 = ( n732 & n18929 ) | ( n732 & n32128 ) | ( n18929 & n32128 ) ;
  assign n32130 = n14030 ^ n9341 ^ n7001 ;
  assign n32131 = ( ~n3426 & n17818 ) | ( ~n3426 & n32130 ) | ( n17818 & n32130 ) ;
  assign n32132 = ( ~n4174 & n21482 ) | ( ~n4174 & n32131 ) | ( n21482 & n32131 ) ;
  assign n32133 = ( n17884 & n24350 ) | ( n17884 & n26944 ) | ( n24350 & n26944 ) ;
  assign n32134 = n11876 ^ n10808 ^ n2685 ;
  assign n32135 = n32134 ^ n29872 ^ n14451 ;
  assign n32136 = n26039 ^ n23200 ^ n22306 ;
  assign n32137 = n32136 ^ n29903 ^ 1'b0 ;
  assign n32138 = n11487 | n32137 ;
  assign n32139 = ( n6120 & n9702 ) | ( n6120 & ~n18973 ) | ( n9702 & ~n18973 ) ;
  assign n32140 = ( n18276 & n23443 ) | ( n18276 & ~n32139 ) | ( n23443 & ~n32139 ) ;
  assign n32141 = ( n26250 & n32061 ) | ( n26250 & n32140 ) | ( n32061 & n32140 ) ;
  assign n32142 = n26619 ^ n25309 ^ n8556 ;
  assign n32143 = n32142 ^ n20403 ^ n5596 ;
  assign n32144 = ( n6155 & n15673 ) | ( n6155 & ~n32143 ) | ( n15673 & ~n32143 ) ;
  assign n32145 = ~n1581 & n9155 ;
  assign n32146 = n32145 ^ n22835 ^ 1'b0 ;
  assign n32147 = n27356 ^ n3510 ^ n2183 ;
  assign n32148 = n12686 | n32147 ;
  assign n32149 = n32148 ^ n3548 ^ 1'b0 ;
  assign n32154 = n19265 ^ n5932 ^ 1'b0 ;
  assign n32150 = n2891 & ~n20028 ;
  assign n32151 = n2795 & n32150 ;
  assign n32152 = ( ~n7591 & n10509 ) | ( ~n7591 & n32151 ) | ( n10509 & n32151 ) ;
  assign n32153 = n32152 ^ n17888 ^ 1'b0 ;
  assign n32155 = n32154 ^ n32153 ^ n15281 ;
  assign n32156 = ( x51 & n8766 ) | ( x51 & n9978 ) | ( n8766 & n9978 ) ;
  assign n32157 = n26214 ^ n11112 ^ n8265 ;
  assign n32158 = n2588 & n7661 ;
  assign n32159 = n32158 ^ n29277 ^ 1'b0 ;
  assign n32160 = ( n1718 & ~n11959 ) | ( n1718 & n25988 ) | ( ~n11959 & n25988 ) ;
  assign n32161 = ( n1443 & n6837 ) | ( n1443 & n13614 ) | ( n6837 & n13614 ) ;
  assign n32162 = ( ~n15212 & n30106 ) | ( ~n15212 & n32161 ) | ( n30106 & n32161 ) ;
  assign n32163 = ( ~n611 & n10044 ) | ( ~n611 & n32162 ) | ( n10044 & n32162 ) ;
  assign n32164 = ( n22389 & n32160 ) | ( n22389 & ~n32163 ) | ( n32160 & ~n32163 ) ;
  assign n32165 = n9289 ^ n5796 ^ n3219 ;
  assign n32166 = n22678 ^ n20241 ^ n2646 ;
  assign n32167 = ( n16034 & n32165 ) | ( n16034 & n32166 ) | ( n32165 & n32166 ) ;
  assign n32168 = n26418 ^ n22294 ^ n6245 ;
  assign n32169 = n2224 & ~n3182 ;
  assign n32170 = n32168 & n32169 ;
  assign n32171 = n32170 ^ n3836 ^ n3715 ;
  assign n32172 = ( ~n955 & n15288 ) | ( ~n955 & n19324 ) | ( n15288 & n19324 ) ;
  assign n32173 = n14292 ^ n13360 ^ n10269 ;
  assign n32174 = n8835 ^ n4515 ^ 1'b0 ;
  assign n32175 = n32174 ^ n22483 ^ n13427 ;
  assign n32176 = ( n8854 & n20365 ) | ( n8854 & n32066 ) | ( n20365 & n32066 ) ;
  assign n32183 = n1677 | n7851 ;
  assign n32179 = n23682 ^ n6391 ^ 1'b0 ;
  assign n32180 = n4041 & n32179 ;
  assign n32178 = ( n1143 & n2659 ) | ( n1143 & ~n6999 ) | ( n2659 & ~n6999 ) ;
  assign n32181 = n32180 ^ n32178 ^ n4099 ;
  assign n32177 = ( n402 & n9033 ) | ( n402 & n22219 ) | ( n9033 & n22219 ) ;
  assign n32182 = n32181 ^ n32177 ^ n11902 ;
  assign n32184 = n32183 ^ n32182 ^ n10293 ;
  assign n32185 = n32184 ^ n14310 ^ n6656 ;
  assign n32186 = n20166 ^ n16090 ^ x241 ;
  assign n32187 = ( n16239 & n19767 ) | ( n16239 & n32186 ) | ( n19767 & n32186 ) ;
  assign n32188 = n8363 ^ n5435 ^ 1'b0 ;
  assign n32189 = ( n2796 & n3451 ) | ( n2796 & n15132 ) | ( n3451 & n15132 ) ;
  assign n32190 = n29077 ^ n16719 ^ n10622 ;
  assign n32191 = ( n32188 & n32189 ) | ( n32188 & n32190 ) | ( n32189 & n32190 ) ;
  assign n32192 = ( n4860 & ~n25207 ) | ( n4860 & n32191 ) | ( ~n25207 & n32191 ) ;
  assign n32193 = n16730 ^ n16329 ^ n9076 ;
  assign n32194 = ( n5566 & n8849 ) | ( n5566 & ~n14731 ) | ( n8849 & ~n14731 ) ;
  assign n32195 = n32194 ^ n11468 ^ n6985 ;
  assign n32196 = n12411 ^ n1326 ^ n742 ;
  assign n32197 = n18832 | n32196 ;
  assign n32198 = n6398 & ~n32197 ;
  assign n32199 = ( n21309 & n25127 ) | ( n21309 & ~n32198 ) | ( n25127 & ~n32198 ) ;
  assign n32200 = n8172 & ~n11982 ;
  assign n32201 = n32200 ^ n26228 ^ 1'b0 ;
  assign n32202 = n32201 ^ n27111 ^ n26401 ;
  assign n32203 = n8914 & n26826 ;
  assign n32204 = n27248 & n32203 ;
  assign n32205 = n32204 ^ n24988 ^ n24944 ;
  assign n32206 = n12740 ^ n7586 ^ n706 ;
  assign n32207 = n1175 & n30617 ;
  assign n32208 = n27257 & n32207 ;
  assign n32209 = ( n4501 & n9131 ) | ( n4501 & n14955 ) | ( n9131 & n14955 ) ;
  assign n32210 = ( n4921 & n15497 ) | ( n4921 & ~n32209 ) | ( n15497 & ~n32209 ) ;
  assign n32213 = n21844 ^ n16428 ^ 1'b0 ;
  assign n32211 = n12749 ^ n11895 ^ n365 ;
  assign n32212 = ( x170 & n7764 ) | ( x170 & ~n32211 ) | ( n7764 & ~n32211 ) ;
  assign n32214 = n32213 ^ n32212 ^ n16146 ;
  assign n32215 = ( n2220 & n8093 ) | ( n2220 & n10744 ) | ( n8093 & n10744 ) ;
  assign n32216 = ( ~n6663 & n13795 ) | ( ~n6663 & n32215 ) | ( n13795 & n32215 ) ;
  assign n32217 = ( ~n9894 & n27372 ) | ( ~n9894 & n30044 ) | ( n27372 & n30044 ) ;
  assign n32218 = ( n1599 & ~n4953 ) | ( n1599 & n32217 ) | ( ~n4953 & n32217 ) ;
  assign n32219 = x193 & ~n4521 ;
  assign n32220 = ~n31713 & n32219 ;
  assign n32221 = n32220 ^ n17959 ^ 1'b0 ;
  assign n32222 = x188 & ~n24631 ;
  assign n32223 = n32221 & n32222 ;
  assign n32227 = n12035 ^ n9183 ^ n5377 ;
  assign n32224 = x244 & n9954 ;
  assign n32225 = n32224 ^ n26414 ^ 1'b0 ;
  assign n32226 = n32225 ^ n9422 ^ n5460 ;
  assign n32228 = n32227 ^ n32226 ^ 1'b0 ;
  assign n32229 = ( ~n2687 & n6852 ) | ( ~n2687 & n32228 ) | ( n6852 & n32228 ) ;
  assign n32230 = ( n5643 & n13081 ) | ( n5643 & n15315 ) | ( n13081 & n15315 ) ;
  assign n32231 = n25362 | n32230 ;
  assign n32243 = n13014 ^ n10560 ^ n4792 ;
  assign n32233 = n5972 ^ n4953 ^ n3134 ;
  assign n32232 = ( ~n7979 & n12371 ) | ( ~n7979 & n17938 ) | ( n12371 & n17938 ) ;
  assign n32234 = n32233 ^ n32232 ^ n24284 ;
  assign n32240 = n3205 ^ n1840 ^ 1'b0 ;
  assign n32239 = ( x234 & n2468 ) | ( x234 & ~n5069 ) | ( n2468 & ~n5069 ) ;
  assign n32235 = n8254 ^ n4985 ^ n2994 ;
  assign n32236 = n5751 | n20748 ;
  assign n32237 = n32235 | n32236 ;
  assign n32238 = ( n3227 & ~n4359 ) | ( n3227 & n32237 ) | ( ~n4359 & n32237 ) ;
  assign n32241 = n32240 ^ n32239 ^ n32238 ;
  assign n32242 = ~n32234 & n32241 ;
  assign n32244 = n32243 ^ n32242 ^ 1'b0 ;
  assign n32245 = n9375 & ~n32244 ;
  assign n32246 = n370 & n32245 ;
  assign n32247 = n32246 ^ n20238 ^ n4761 ;
  assign n32248 = ( n2256 & ~n4622 ) | ( n2256 & n17749 ) | ( ~n4622 & n17749 ) ;
  assign n32249 = n16004 ^ n7907 ^ n3762 ;
  assign n32250 = n16842 ^ n6106 ^ n1534 ;
  assign n32251 = n2780 & n32250 ;
  assign n32252 = ~n32249 & n32251 ;
  assign n32253 = ( ~n5203 & n31090 ) | ( ~n5203 & n32252 ) | ( n31090 & n32252 ) ;
  assign n32254 = n32248 & ~n32253 ;
  assign n32255 = n4199 & n32254 ;
  assign n32256 = n12162 ^ n5198 ^ 1'b0 ;
  assign n32257 = n5751 | n32256 ;
  assign n32258 = ( ~n15803 & n24038 ) | ( ~n15803 & n32257 ) | ( n24038 & n32257 ) ;
  assign n32259 = ( n4170 & n15824 ) | ( n4170 & ~n32258 ) | ( n15824 & ~n32258 ) ;
  assign n32260 = ~n17842 & n32259 ;
  assign n32261 = n12154 & n32260 ;
  assign n32263 = n28366 ^ n6600 ^ n5573 ;
  assign n32262 = n3667 & ~n7237 ;
  assign n32264 = n32263 ^ n32262 ^ 1'b0 ;
  assign n32265 = ( n16626 & n24474 ) | ( n16626 & n32264 ) | ( n24474 & n32264 ) ;
  assign n32266 = ( n696 & n23478 ) | ( n696 & n32265 ) | ( n23478 & n32265 ) ;
  assign n32267 = n12025 ^ n11239 ^ 1'b0 ;
  assign n32268 = n20988 | n32267 ;
  assign n32269 = ( n1007 & n3236 ) | ( n1007 & ~n10764 ) | ( n3236 & ~n10764 ) ;
  assign n32270 = ( n29014 & ~n32268 ) | ( n29014 & n32269 ) | ( ~n32268 & n32269 ) ;
  assign n32271 = ( n16876 & ~n26291 ) | ( n16876 & n31568 ) | ( ~n26291 & n31568 ) ;
  assign n32272 = ( n32266 & n32270 ) | ( n32266 & ~n32271 ) | ( n32270 & ~n32271 ) ;
  assign n32273 = n28222 ^ n8290 ^ n760 ;
  assign n32274 = n8460 & ~n32273 ;
  assign n32275 = ( n2764 & ~n4001 ) | ( n2764 & n24706 ) | ( ~n4001 & n24706 ) ;
  assign n32276 = n32275 ^ n23529 ^ n19023 ;
  assign n32277 = n17859 ^ n11234 ^ x138 ;
  assign n32278 = ( n25599 & ~n32276 ) | ( n25599 & n32277 ) | ( ~n32276 & n32277 ) ;
  assign n32279 = n25003 ^ n12613 ^ n4451 ;
  assign n32280 = n18439 | n27790 ;
  assign n32281 = ( ~n7136 & n8381 ) | ( ~n7136 & n19120 ) | ( n8381 & n19120 ) ;
  assign n32282 = ( n2514 & n12915 ) | ( n2514 & ~n14446 ) | ( n12915 & ~n14446 ) ;
  assign n32283 = ( n14387 & n32281 ) | ( n14387 & n32282 ) | ( n32281 & n32282 ) ;
  assign n32284 = ( n31677 & ~n32198 ) | ( n31677 & n32283 ) | ( ~n32198 & n32283 ) ;
  assign n32285 = ( n1326 & n2601 ) | ( n1326 & n6030 ) | ( n2601 & n6030 ) ;
  assign n32286 = n19493 ^ n12695 ^ 1'b0 ;
  assign n32287 = n20117 & ~n32286 ;
  assign n32288 = ( n18562 & n32285 ) | ( n18562 & n32287 ) | ( n32285 & n32287 ) ;
  assign n32289 = n32288 ^ n13280 ^ n3935 ;
  assign n32290 = ( n1295 & n3571 ) | ( n1295 & ~n12279 ) | ( n3571 & ~n12279 ) ;
  assign n32291 = ( n13169 & n23395 ) | ( n13169 & ~n32290 ) | ( n23395 & ~n32290 ) ;
  assign n32292 = n997 & ~n22235 ;
  assign n32293 = ( n9094 & n11650 ) | ( n9094 & ~n12420 ) | ( n11650 & ~n12420 ) ;
  assign n32294 = ( ~n3693 & n13575 ) | ( ~n3693 & n32293 ) | ( n13575 & n32293 ) ;
  assign n32295 = ( n17576 & ~n18987 ) | ( n17576 & n32294 ) | ( ~n18987 & n32294 ) ;
  assign n32296 = ( n3972 & n12281 ) | ( n3972 & n32295 ) | ( n12281 & n32295 ) ;
  assign n32297 = n32296 ^ n19031 ^ n8037 ;
  assign n32298 = ( n16223 & n18864 ) | ( n16223 & n21029 ) | ( n18864 & n21029 ) ;
  assign n32299 = n32298 ^ n28447 ^ n7899 ;
  assign n32300 = n17025 ^ n6890 ^ n6029 ;
  assign n32301 = n32300 ^ n17493 ^ 1'b0 ;
  assign n32302 = ( n5556 & ~n9689 ) | ( n5556 & n32301 ) | ( ~n9689 & n32301 ) ;
  assign n32303 = n12566 ^ n8127 ^ n3742 ;
  assign n32304 = n32303 ^ n26588 ^ n16061 ;
  assign n32305 = n26303 ^ n21898 ^ n4751 ;
  assign n32306 = ~n16207 & n32305 ;
  assign n32307 = n32306 ^ n18296 ^ 1'b0 ;
  assign n32308 = ( n7012 & n24963 ) | ( n7012 & n32307 ) | ( n24963 & n32307 ) ;
  assign n32309 = ~n2088 & n13140 ;
  assign n32310 = n19003 & n32309 ;
  assign n32311 = ( n7439 & ~n16695 ) | ( n7439 & n32310 ) | ( ~n16695 & n32310 ) ;
  assign n32312 = n10310 ^ n7051 ^ 1'b0 ;
  assign n32313 = ( n1980 & ~n7924 ) | ( n1980 & n32312 ) | ( ~n7924 & n32312 ) ;
  assign n32315 = n27612 ^ n10198 ^ n3244 ;
  assign n32314 = n2222 & ~n8760 ;
  assign n32316 = n32315 ^ n32314 ^ n23759 ;
  assign n32317 = ( n6735 & n19722 ) | ( n6735 & ~n21088 ) | ( n19722 & ~n21088 ) ;
  assign n32318 = ( n7764 & n26352 ) | ( n7764 & ~n30237 ) | ( n26352 & ~n30237 ) ;
  assign n32319 = ( ~n7045 & n29233 ) | ( ~n7045 & n30172 ) | ( n29233 & n30172 ) ;
  assign n32320 = n9021 ^ n266 ^ 1'b0 ;
  assign n32321 = ( n6956 & n14067 ) | ( n6956 & n32320 ) | ( n14067 & n32320 ) ;
  assign n32322 = ( n15921 & n23464 ) | ( n15921 & ~n32321 ) | ( n23464 & ~n32321 ) ;
  assign n32323 = ( n12849 & ~n26577 ) | ( n12849 & n32322 ) | ( ~n26577 & n32322 ) ;
  assign n32324 = n2118 & ~n10820 ;
  assign n32325 = n32324 ^ n1610 ^ 1'b0 ;
  assign n32326 = ( n18693 & n21408 ) | ( n18693 & ~n22695 ) | ( n21408 & ~n22695 ) ;
  assign n32327 = n32326 ^ n30906 ^ 1'b0 ;
  assign n32328 = n29629 ^ n8484 ^ n4465 ;
  assign n32329 = n26960 ^ n25709 ^ n17938 ;
  assign n32330 = ~n9665 & n32329 ;
  assign n32331 = n32330 ^ n8697 ^ 1'b0 ;
  assign n32332 = ( ~n14814 & n32328 ) | ( ~n14814 & n32331 ) | ( n32328 & n32331 ) ;
  assign n32335 = n3942 ^ n3414 ^ 1'b0 ;
  assign n32334 = n14090 ^ n6926 ^ 1'b0 ;
  assign n32336 = n32335 ^ n32334 ^ n20645 ;
  assign n32333 = ( n10273 & n17832 ) | ( n10273 & n23173 ) | ( n17832 & n23173 ) ;
  assign n32337 = n32336 ^ n32333 ^ n23090 ;
  assign n32338 = ( n12392 & ~n18048 ) | ( n12392 & n22372 ) | ( ~n18048 & n22372 ) ;
  assign n32339 = ( n1288 & ~n5866 ) | ( n1288 & n25424 ) | ( ~n5866 & n25424 ) ;
  assign n32340 = n32339 ^ n27206 ^ n19723 ;
  assign n32341 = ( ~n5417 & n12958 ) | ( ~n5417 & n32340 ) | ( n12958 & n32340 ) ;
  assign n32342 = ( n4986 & n11133 ) | ( n4986 & ~n25410 ) | ( n11133 & ~n25410 ) ;
  assign n32343 = n1758 | n32342 ;
  assign n32344 = ( n19063 & n25836 ) | ( n19063 & ~n32343 ) | ( n25836 & ~n32343 ) ;
  assign n32345 = n13741 ^ n9677 ^ n1114 ;
  assign n32346 = n32345 ^ n14997 ^ n2304 ;
  assign n32347 = n23161 ^ n11478 ^ n4638 ;
  assign n32348 = n32347 ^ n2804 ^ n297 ;
  assign n32349 = n14259 ^ n11797 ^ 1'b0 ;
  assign n32350 = n10065 & n32349 ;
  assign n32351 = n31649 & n32350 ;
  assign n32352 = ~n32348 & n32351 ;
  assign n32353 = n32352 ^ n31347 ^ n14913 ;
  assign n32354 = n6563 | n7368 ;
  assign n32355 = ( n4768 & ~n10753 ) | ( n4768 & n28583 ) | ( ~n10753 & n28583 ) ;
  assign n32356 = ~n14010 & n31773 ;
  assign n32357 = ~n6099 & n32356 ;
  assign n32358 = n15064 ^ n9219 ^ n1586 ;
  assign n32359 = n28162 ^ n4873 ^ 1'b0 ;
  assign n32360 = ~n32358 & n32359 ;
  assign n32361 = n5166 & ~n26935 ;
  assign n32362 = ~n7813 & n32361 ;
  assign n32363 = n32362 ^ n31753 ^ n16220 ;
  assign n32364 = n32360 & ~n32363 ;
  assign n32365 = n32364 ^ n27161 ^ 1'b0 ;
  assign n32366 = n30920 ^ n24586 ^ n2889 ;
  assign n32368 = n23631 ^ n14094 ^ n2638 ;
  assign n32369 = n32368 ^ n11818 ^ n7379 ;
  assign n32370 = ( n8680 & ~n9723 ) | ( n8680 & n32369 ) | ( ~n9723 & n32369 ) ;
  assign n32367 = n16271 ^ n15052 ^ n15045 ;
  assign n32371 = n32370 ^ n32367 ^ n18411 ;
  assign n32372 = n25683 ^ n25111 ^ n2890 ;
  assign n32373 = ( n1742 & n2644 ) | ( n1742 & ~n3480 ) | ( n2644 & ~n3480 ) ;
  assign n32374 = ( n7918 & ~n28093 ) | ( n7918 & n32373 ) | ( ~n28093 & n32373 ) ;
  assign n32375 = n18415 ^ n1900 ^ 1'b0 ;
  assign n32376 = n15267 & n32375 ;
  assign n32377 = n16141 ^ n16001 ^ 1'b0 ;
  assign n32378 = n23344 | n32377 ;
  assign n32380 = ( ~n5017 & n5464 ) | ( ~n5017 & n11965 ) | ( n5464 & n11965 ) ;
  assign n32379 = n32249 ^ n7675 ^ n1208 ;
  assign n32381 = n32380 ^ n32379 ^ n16392 ;
  assign n32382 = n32381 ^ n29512 ^ 1'b0 ;
  assign n32383 = n32378 | n32382 ;
  assign n32384 = n6940 ^ n4147 ^ n3797 ;
  assign n32385 = ~n11633 & n32384 ;
  assign n32386 = n2861 & n32385 ;
  assign n32387 = ( ~n6467 & n9961 ) | ( ~n6467 & n32386 ) | ( n9961 & n32386 ) ;
  assign n32388 = ~n1911 & n5729 ;
  assign n32389 = n32388 ^ n20491 ^ n8635 ;
  assign n32390 = n11219 ^ n837 ^ 1'b0 ;
  assign n32391 = ( n22020 & n32019 ) | ( n22020 & n32390 ) | ( n32019 & n32390 ) ;
  assign n32392 = n32391 ^ n23134 ^ n1602 ;
  assign n32393 = ( n21765 & n32038 ) | ( n21765 & n32392 ) | ( n32038 & n32392 ) ;
  assign n32394 = n32393 ^ n28863 ^ 1'b0 ;
  assign n32395 = n8651 & ~n32394 ;
  assign n32397 = ( n7779 & ~n8472 ) | ( n7779 & n10795 ) | ( ~n8472 & n10795 ) ;
  assign n32396 = n29881 ^ n11079 ^ n3762 ;
  assign n32398 = n32397 ^ n32396 ^ n8994 ;
  assign n32399 = n32398 ^ n21524 ^ 1'b0 ;
  assign n32403 = n21087 ^ n18906 ^ n1095 ;
  assign n32402 = n15836 ^ n9268 ^ 1'b0 ;
  assign n32404 = n32403 ^ n32402 ^ n18722 ;
  assign n32400 = n645 & ~n9626 ;
  assign n32401 = n32400 ^ n11148 ^ 1'b0 ;
  assign n32405 = n32404 ^ n32401 ^ n23896 ;
  assign n32406 = ( n14665 & ~n22412 ) | ( n14665 & n27922 ) | ( ~n22412 & n27922 ) ;
  assign n32407 = ( ~n6356 & n27238 ) | ( ~n6356 & n32402 ) | ( n27238 & n32402 ) ;
  assign n32408 = n24575 & ~n32407 ;
  assign n32409 = n7553 ^ n5491 ^ n1326 ;
  assign n32410 = n32409 ^ n22426 ^ n9705 ;
  assign n32411 = n15537 ^ n4152 ^ x53 ;
  assign n32412 = ( n11989 & ~n12142 ) | ( n11989 & n15819 ) | ( ~n12142 & n15819 ) ;
  assign n32413 = n32412 ^ n27839 ^ n18104 ;
  assign n32414 = n9154 ^ n7759 ^ n6369 ;
  assign n32415 = n13603 ^ n4354 ^ 1'b0 ;
  assign n32416 = n32415 ^ n22171 ^ n9783 ;
  assign n32417 = ( n3656 & n24407 ) | ( n3656 & ~n32416 ) | ( n24407 & ~n32416 ) ;
  assign n32418 = ( ~n19273 & n32414 ) | ( ~n19273 & n32417 ) | ( n32414 & n32417 ) ;
  assign n32419 = n8671 ^ n7212 ^ n346 ;
  assign n32420 = ( ~n11404 & n13661 ) | ( ~n11404 & n32419 ) | ( n13661 & n32419 ) ;
  assign n32421 = ( n8838 & n24041 ) | ( n8838 & ~n32420 ) | ( n24041 & ~n32420 ) ;
  assign n32422 = n12993 ^ n4468 ^ 1'b0 ;
  assign n32423 = n32421 & n32422 ;
  assign n32424 = ~n29992 & n30399 ;
  assign n32425 = ( n494 & n9739 ) | ( n494 & n32424 ) | ( n9739 & n32424 ) ;
  assign n32426 = x160 & n2236 ;
  assign n32427 = n32426 ^ n28492 ^ n11585 ;
  assign n32428 = ( n6717 & n6984 ) | ( n6717 & n23619 ) | ( n6984 & n23619 ) ;
  assign n32429 = ( ~n8029 & n14170 ) | ( ~n8029 & n32428 ) | ( n14170 & n32428 ) ;
  assign n32430 = ( n3401 & ~n12474 ) | ( n3401 & n32429 ) | ( ~n12474 & n32429 ) ;
  assign n32431 = n31959 ^ n17578 ^ n11905 ;
  assign n32432 = n1654 & ~n4112 ;
  assign n32435 = n31035 ^ n10070 ^ n6985 ;
  assign n32436 = ( n17382 & n26439 ) | ( n17382 & ~n32435 ) | ( n26439 & ~n32435 ) ;
  assign n32433 = n18926 ^ n1007 ^ 1'b0 ;
  assign n32434 = n6470 & ~n32433 ;
  assign n32437 = n32436 ^ n32434 ^ 1'b0 ;
  assign n32438 = n9283 ^ n5942 ^ n3911 ;
  assign n32439 = n32438 ^ n7505 ^ n7158 ;
  assign n32440 = ~n9898 & n32439 ;
  assign n32441 = n32440 ^ n12827 ^ 1'b0 ;
  assign n32445 = n30527 ^ n19756 ^ n18764 ;
  assign n32442 = n5078 ^ n1308 ^ 1'b0 ;
  assign n32443 = ~n2945 & n32442 ;
  assign n32444 = ( n5480 & n28121 ) | ( n5480 & n32443 ) | ( n28121 & n32443 ) ;
  assign n32446 = n32445 ^ n32444 ^ n18584 ;
  assign n32447 = n30944 ^ n10784 ^ n10608 ;
  assign n32448 = ( n4205 & n8831 ) | ( n4205 & n32447 ) | ( n8831 & n32447 ) ;
  assign n32449 = n18696 ^ n11739 ^ n1463 ;
  assign n32450 = ( n3960 & n5816 ) | ( n3960 & n32449 ) | ( n5816 & n32449 ) ;
  assign n32451 = n20347 ^ n19343 ^ n11643 ;
  assign n32452 = ( ~n6882 & n7661 ) | ( ~n6882 & n21140 ) | ( n7661 & n21140 ) ;
  assign n32453 = n14613 ^ n5409 ^ 1'b0 ;
  assign n32454 = n32452 & n32453 ;
  assign n32455 = ( n6699 & ~n8879 ) | ( n6699 & n15781 ) | ( ~n8879 & n15781 ) ;
  assign n32456 = ~n8944 & n32455 ;
  assign n32457 = n13664 ^ n10770 ^ n1215 ;
  assign n32458 = n28733 ^ n25320 ^ n22348 ;
  assign n32459 = n19846 ^ n4895 ^ 1'b0 ;
  assign n32460 = ( ~n10816 & n12915 ) | ( ~n10816 & n18123 ) | ( n12915 & n18123 ) ;
  assign n32461 = n32460 ^ n26666 ^ 1'b0 ;
  assign n32462 = n23583 & ~n32461 ;
  assign n32463 = n30441 ^ n26695 ^ n8617 ;
  assign n32464 = n32463 ^ n29131 ^ n10575 ;
  assign n32465 = n27198 ^ n6340 ^ n4115 ;
  assign n32466 = n6040 & n23933 ;
  assign n32467 = ( n19502 & n19519 ) | ( n19502 & ~n32466 ) | ( n19519 & ~n32466 ) ;
  assign n32468 = n19922 ^ n16227 ^ n3905 ;
  assign n32469 = ( ~n11958 & n23429 ) | ( ~n11958 & n32468 ) | ( n23429 & n32468 ) ;
  assign n32470 = ( n22980 & ~n24613 ) | ( n22980 & n24854 ) | ( ~n24613 & n24854 ) ;
  assign n32471 = n28689 ^ n10631 ^ n9896 ;
  assign n32472 = ( n13713 & n14410 ) | ( n13713 & n20106 ) | ( n14410 & n20106 ) ;
  assign n32473 = n32472 ^ n9994 ^ 1'b0 ;
  assign n32474 = n22255 & n32473 ;
  assign n32475 = ( n3011 & ~n13435 ) | ( n3011 & n18362 ) | ( ~n13435 & n18362 ) ;
  assign n32476 = n26152 ^ n25151 ^ n6109 ;
  assign n32477 = ( n4965 & n5981 ) | ( n4965 & n25612 ) | ( n5981 & n25612 ) ;
  assign n32478 = ( ~n5171 & n10846 ) | ( ~n5171 & n32477 ) | ( n10846 & n32477 ) ;
  assign n32479 = ( n20053 & n27971 ) | ( n20053 & n32478 ) | ( n27971 & n32478 ) ;
  assign n32480 = ( n32475 & n32476 ) | ( n32475 & ~n32479 ) | ( n32476 & ~n32479 ) ;
  assign n32481 = ( ~n2077 & n4903 ) | ( ~n2077 & n13206 ) | ( n4903 & n13206 ) ;
  assign n32482 = n32481 ^ n604 ^ 1'b0 ;
  assign n32483 = n6366 & n32482 ;
  assign n32484 = ( n2978 & n17236 ) | ( n2978 & ~n32483 ) | ( n17236 & ~n32483 ) ;
  assign n32485 = ( n3671 & ~n20524 ) | ( n3671 & n21006 ) | ( ~n20524 & n21006 ) ;
  assign n32486 = ( n16264 & n21636 ) | ( n16264 & ~n32485 ) | ( n21636 & ~n32485 ) ;
  assign n32489 = n22073 ^ n11350 ^ n9877 ;
  assign n32487 = n10209 ^ n9834 ^ n951 ;
  assign n32488 = n32487 ^ n14676 ^ n4068 ;
  assign n32490 = n32489 ^ n32488 ^ n13375 ;
  assign n32491 = ( n5282 & n14261 ) | ( n5282 & ~n32490 ) | ( n14261 & ~n32490 ) ;
  assign n32492 = ( ~n6423 & n32486 ) | ( ~n6423 & n32491 ) | ( n32486 & n32491 ) ;
  assign n32493 = n29996 ^ n21493 ^ n9926 ;
  assign n32494 = ( n2675 & ~n7655 ) | ( n2675 & n18251 ) | ( ~n7655 & n18251 ) ;
  assign n32495 = n3800 & ~n32494 ;
  assign n32496 = ( n10764 & ~n23059 ) | ( n10764 & n32495 ) | ( ~n23059 & n32495 ) ;
  assign n32497 = n32496 ^ n21651 ^ 1'b0 ;
  assign n32498 = ( n9786 & ~n27751 ) | ( n9786 & n32497 ) | ( ~n27751 & n32497 ) ;
  assign n32499 = n32498 ^ n8711 ^ n2557 ;
  assign n32500 = ( n18260 & n21076 ) | ( n18260 & n21250 ) | ( n21076 & n21250 ) ;
  assign n32501 = ( n1175 & ~n12933 ) | ( n1175 & n32500 ) | ( ~n12933 & n32500 ) ;
  assign n32502 = n22019 ^ n2512 ^ 1'b0 ;
  assign n32503 = ( n15085 & n21926 ) | ( n15085 & ~n32502 ) | ( n21926 & ~n32502 ) ;
  assign n32504 = ( ~n1403 & n25471 ) | ( ~n1403 & n32503 ) | ( n25471 & n32503 ) ;
  assign n32509 = ( n1900 & n4393 ) | ( n1900 & n26670 ) | ( n4393 & n26670 ) ;
  assign n32510 = ( n6369 & n14506 ) | ( n6369 & ~n30530 ) | ( n14506 & ~n30530 ) ;
  assign n32511 = ( n12993 & n32509 ) | ( n12993 & ~n32510 ) | ( n32509 & ~n32510 ) ;
  assign n32505 = n31376 ^ n17942 ^ n1821 ;
  assign n32506 = ( ~n4840 & n25355 ) | ( ~n4840 & n32505 ) | ( n25355 & n32505 ) ;
  assign n32507 = n21030 ^ n14922 ^ n3201 ;
  assign n32508 = ( n25570 & n32506 ) | ( n25570 & n32507 ) | ( n32506 & n32507 ) ;
  assign n32512 = n32511 ^ n32508 ^ n8076 ;
  assign n32513 = ( ~n14168 & n15402 ) | ( ~n14168 & n22828 ) | ( n15402 & n22828 ) ;
  assign n32514 = ( n6685 & n25083 ) | ( n6685 & n26702 ) | ( n25083 & n26702 ) ;
  assign n32515 = n32514 ^ n24537 ^ n21749 ;
  assign n32516 = ~n32513 & n32515 ;
  assign n32517 = n32516 ^ n6256 ^ 1'b0 ;
  assign n32518 = n18040 ^ n8978 ^ x17 ;
  assign n32519 = ( n23225 & n30012 ) | ( n23225 & ~n32518 ) | ( n30012 & ~n32518 ) ;
  assign n32526 = ( n3338 & ~n6138 ) | ( n3338 & n6573 ) | ( ~n6138 & n6573 ) ;
  assign n32527 = n4364 ^ n1248 ^ n438 ;
  assign n32528 = ( n7618 & n24429 ) | ( n7618 & ~n32527 ) | ( n24429 & ~n32527 ) ;
  assign n32529 = n32526 & n32528 ;
  assign n32530 = n32529 ^ n20113 ^ n14467 ;
  assign n32523 = ( n923 & n1325 ) | ( n923 & n5458 ) | ( n1325 & n5458 ) ;
  assign n32524 = ( ~n15782 & n15922 ) | ( ~n15782 & n22881 ) | ( n15922 & n22881 ) ;
  assign n32525 = ( ~n19991 & n32523 ) | ( ~n19991 & n32524 ) | ( n32523 & n32524 ) ;
  assign n32531 = n32530 ^ n32525 ^ n6013 ;
  assign n32521 = ~n10096 & n27510 ;
  assign n32522 = n11704 & n32521 ;
  assign n32532 = n32531 ^ n32522 ^ n11555 ;
  assign n32520 = ( n13422 & ~n15049 ) | ( n13422 & n25279 ) | ( ~n15049 & n25279 ) ;
  assign n32533 = n32532 ^ n32520 ^ 1'b0 ;
  assign n32534 = n9625 ^ n9132 ^ n7700 ;
  assign n32535 = n18333 ^ n7941 ^ 1'b0 ;
  assign n32536 = ~n1476 & n8642 ;
  assign n32537 = ~n32535 & n32536 ;
  assign n32538 = n29358 ^ n11759 ^ 1'b0 ;
  assign n32539 = n5877 & n32538 ;
  assign n32540 = ( ~n964 & n11585 ) | ( ~n964 & n32539 ) | ( n11585 & n32539 ) ;
  assign n32541 = n4776 | n9394 ;
  assign n32542 = n32541 ^ n15157 ^ 1'b0 ;
  assign n32543 = n16976 | n22548 ;
  assign n32544 = ( ~n1039 & n32542 ) | ( ~n1039 & n32543 ) | ( n32542 & n32543 ) ;
  assign n32546 = ( n3045 & n4477 ) | ( n3045 & ~n13742 ) | ( n4477 & ~n13742 ) ;
  assign n32547 = ( n14017 & ~n19290 ) | ( n14017 & n32546 ) | ( ~n19290 & n32546 ) ;
  assign n32545 = ~n5549 & n12008 ;
  assign n32548 = n32547 ^ n32545 ^ 1'b0 ;
  assign n32549 = ( n1572 & n5592 ) | ( n1572 & ~n16816 ) | ( n5592 & ~n16816 ) ;
  assign n32550 = n32549 ^ n18842 ^ n10558 ;
  assign n32551 = n32550 ^ n8310 ^ 1'b0 ;
  assign n32552 = n18132 & n32551 ;
  assign n32553 = ( n7831 & ~n22458 ) | ( n7831 & n32552 ) | ( ~n22458 & n32552 ) ;
  assign n32554 = ( n2299 & n13005 ) | ( n2299 & n32553 ) | ( n13005 & n32553 ) ;
  assign n32555 = n32554 ^ n8741 ^ n5310 ;
  assign n32556 = n26141 ^ n24090 ^ n23665 ;
  assign n32557 = ( n25523 & ~n32555 ) | ( n25523 & n32556 ) | ( ~n32555 & n32556 ) ;
  assign n32558 = ( ~n22693 & n32548 ) | ( ~n22693 & n32557 ) | ( n32548 & n32557 ) ;
  assign n32559 = n5790 ^ n2049 ^ n1108 ;
  assign n32560 = ( ~n10867 & n25317 ) | ( ~n10867 & n32559 ) | ( n25317 & n32559 ) ;
  assign n32561 = n21233 ^ n15656 ^ 1'b0 ;
  assign n32562 = n31916 ^ n9463 ^ n7390 ;
  assign n32563 = n15720 ^ n14784 ^ n3518 ;
  assign n32564 = n22870 ^ n18735 ^ n17939 ;
  assign n32567 = n3595 ^ n2964 ^ n2624 ;
  assign n32568 = ( n8721 & n16455 ) | ( n8721 & ~n32567 ) | ( n16455 & ~n32567 ) ;
  assign n32565 = n16814 ^ n6263 ^ n4472 ;
  assign n32566 = ( n2966 & n5459 ) | ( n2966 & n32565 ) | ( n5459 & n32565 ) ;
  assign n32569 = n32568 ^ n32566 ^ n1255 ;
  assign n32570 = n22047 ^ n7365 ^ 1'b0 ;
  assign n32571 = ( n1602 & n14022 ) | ( n1602 & ~n22458 ) | ( n14022 & ~n22458 ) ;
  assign n32572 = ( n12667 & ~n32570 ) | ( n12667 & n32571 ) | ( ~n32570 & n32571 ) ;
  assign n32573 = ( ~n1528 & n19406 ) | ( ~n1528 & n32572 ) | ( n19406 & n32572 ) ;
  assign n32575 = ( ~n7784 & n24404 ) | ( ~n7784 & n29523 ) | ( n24404 & n29523 ) ;
  assign n32576 = ( ~n1659 & n15302 ) | ( ~n1659 & n32575 ) | ( n15302 & n32575 ) ;
  assign n32574 = ~n21801 & n25766 ;
  assign n32577 = n32576 ^ n32574 ^ 1'b0 ;
  assign n32578 = n32577 ^ n21364 ^ n3417 ;
  assign n32579 = n8807 ^ n7968 ^ n3989 ;
  assign n32580 = n32579 ^ n28921 ^ n21431 ;
  assign n32581 = n32580 ^ n7743 ^ n3320 ;
  assign n32582 = n5802 & ~n31499 ;
  assign n32583 = n15800 ^ n8669 ^ n4168 ;
  assign n32584 = ( ~n10509 & n25212 ) | ( ~n10509 & n32583 ) | ( n25212 & n32583 ) ;
  assign n32585 = n32584 ^ n6855 ^ n5344 ;
  assign n32586 = ( n6638 & n27493 ) | ( n6638 & ~n32336 ) | ( n27493 & ~n32336 ) ;
  assign n32587 = ~n11249 & n23004 ;
  assign n32588 = ( n331 & n7774 ) | ( n331 & n14720 ) | ( n7774 & n14720 ) ;
  assign n32589 = ( n24872 & n30987 ) | ( n24872 & n32588 ) | ( n30987 & n32588 ) ;
  assign n32590 = n32589 ^ n22999 ^ n8664 ;
  assign n32591 = ( n11183 & n26774 ) | ( n11183 & ~n28356 ) | ( n26774 & ~n28356 ) ;
  assign n32592 = n32419 ^ n22313 ^ n9687 ;
  assign n32594 = n17139 ^ n13511 ^ 1'b0 ;
  assign n32593 = n27433 ^ n9587 ^ n4827 ;
  assign n32595 = n32594 ^ n32593 ^ n19803 ;
  assign n32596 = n32595 ^ n12499 ^ n4925 ;
  assign n32597 = n25022 ^ n6785 ^ 1'b0 ;
  assign n32598 = n17617 ^ n15289 ^ n1271 ;
  assign n32599 = ( n27393 & ~n32597 ) | ( n27393 & n32598 ) | ( ~n32597 & n32598 ) ;
  assign n32600 = n8654 ^ n2185 ^ 1'b0 ;
  assign n32601 = ( n12623 & n16260 ) | ( n12623 & ~n32600 ) | ( n16260 & ~n32600 ) ;
  assign n32602 = ( n411 & n19659 ) | ( n411 & n21233 ) | ( n19659 & n21233 ) ;
  assign n32603 = ( ~n1838 & n32601 ) | ( ~n1838 & n32602 ) | ( n32601 & n32602 ) ;
  assign n32604 = ( n2589 & n3070 ) | ( n2589 & ~n9260 ) | ( n3070 & ~n9260 ) ;
  assign n32605 = ( n4404 & n7212 ) | ( n4404 & ~n8975 ) | ( n7212 & ~n8975 ) ;
  assign n32609 = n14768 ^ n14366 ^ n6744 ;
  assign n32610 = n32609 ^ n28438 ^ n17207 ;
  assign n32611 = ( n6586 & ~n21017 ) | ( n6586 & n32610 ) | ( ~n21017 & n32610 ) ;
  assign n32608 = n24885 ^ n24155 ^ x108 ;
  assign n32606 = ( n5312 & n14267 ) | ( n5312 & n14617 ) | ( n14267 & n14617 ) ;
  assign n32607 = n32606 ^ n3800 ^ 1'b0 ;
  assign n32612 = n32611 ^ n32608 ^ n32607 ;
  assign n32615 = ( ~n11637 & n15515 ) | ( ~n11637 & n22019 ) | ( n15515 & n22019 ) ;
  assign n32613 = ( ~n684 & n11420 ) | ( ~n684 & n18868 ) | ( n11420 & n18868 ) ;
  assign n32614 = n32613 ^ n26713 ^ n13695 ;
  assign n32616 = n32615 ^ n32614 ^ n13065 ;
  assign n32620 = n1770 | n2373 ;
  assign n32621 = n32620 ^ n8412 ^ 1'b0 ;
  assign n32622 = ( n2995 & n3546 ) | ( n2995 & n32621 ) | ( n3546 & n32621 ) ;
  assign n32618 = n24869 ^ n24146 ^ 1'b0 ;
  assign n32617 = n5298 & n32265 ;
  assign n32619 = n32618 ^ n32617 ^ 1'b0 ;
  assign n32623 = n32622 ^ n32619 ^ n14359 ;
  assign n32624 = n21949 ^ n4087 ^ n909 ;
  assign n32625 = n32624 ^ n5121 ^ n4376 ;
  assign n32626 = n32625 ^ n11125 ^ x210 ;
  assign n32627 = n12432 & n32626 ;
  assign n32628 = n20935 ^ n11579 ^ n6638 ;
  assign n32629 = n32628 ^ n5376 ^ n1075 ;
  assign n32630 = ( n4291 & n21167 ) | ( n4291 & ~n32629 ) | ( n21167 & ~n32629 ) ;
  assign n32631 = ( n3465 & ~n13636 ) | ( n3465 & n32630 ) | ( ~n13636 & n32630 ) ;
  assign n32632 = n32631 ^ n14700 ^ 1'b0 ;
  assign n32633 = n32632 ^ n14317 ^ n13064 ;
  assign n32634 = ~n11588 & n14960 ;
  assign n32635 = n32634 ^ n4065 ^ 1'b0 ;
  assign n32636 = n19706 ^ n7993 ^ n1280 ;
  assign n32637 = n32636 ^ n17225 ^ n8029 ;
  assign n32638 = ( ~n909 & n32635 ) | ( ~n909 & n32637 ) | ( n32635 & n32637 ) ;
  assign n32639 = n26012 ^ n18975 ^ n3772 ;
  assign n32640 = n32639 ^ n21880 ^ n17623 ;
  assign n32641 = ( n1687 & n18315 ) | ( n1687 & ~n32640 ) | ( n18315 & ~n32640 ) ;
  assign n32642 = ( ~n4638 & n7622 ) | ( ~n4638 & n32641 ) | ( n7622 & n32641 ) ;
  assign n32643 = ( ~n7625 & n16213 ) | ( ~n7625 & n31483 ) | ( n16213 & n31483 ) ;
  assign n32644 = n17364 ^ n7754 ^ 1'b0 ;
  assign n32645 = ( n7428 & ~n10315 ) | ( n7428 & n32644 ) | ( ~n10315 & n32644 ) ;
  assign n32646 = n32645 ^ n14069 ^ n2213 ;
  assign n32647 = ( ~n2157 & n2661 ) | ( ~n2157 & n13719 ) | ( n2661 & n13719 ) ;
  assign n32648 = ( ~n1267 & n2218 ) | ( ~n1267 & n32647 ) | ( n2218 & n32647 ) ;
  assign n32649 = n2060 | n30116 ;
  assign n32650 = n24932 & ~n32649 ;
  assign n32651 = n32650 ^ n31958 ^ n18413 ;
  assign n32652 = ~n21912 & n32327 ;
  assign n32653 = n32652 ^ n10146 ^ 1'b0 ;
  assign n32658 = n15425 ^ n3172 ^ 1'b0 ;
  assign n32659 = n12964 & ~n32658 ;
  assign n32654 = ( n8603 & n14584 ) | ( n8603 & n28186 ) | ( n14584 & n28186 ) ;
  assign n32655 = ~n4501 & n32654 ;
  assign n32656 = ~n11922 & n32655 ;
  assign n32657 = n4213 & ~n32656 ;
  assign n32660 = n32659 ^ n32657 ^ 1'b0 ;
  assign n32664 = n6348 ^ n5639 ^ n4120 ;
  assign n32661 = ( ~n2916 & n8121 ) | ( ~n2916 & n15046 ) | ( n8121 & n15046 ) ;
  assign n32662 = n32661 ^ n31127 ^ n17829 ;
  assign n32663 = n32662 ^ n25580 ^ x66 ;
  assign n32665 = n32664 ^ n32663 ^ n17262 ;
  assign n32666 = ( ~n3307 & n3484 ) | ( ~n3307 & n7595 ) | ( n3484 & n7595 ) ;
  assign n32667 = n11099 ^ n10881 ^ n4013 ;
  assign n32668 = n32667 ^ n23839 ^ n18832 ;
  assign n32669 = n32668 ^ n28845 ^ n24191 ;
  assign n32670 = ( n30511 & ~n32666 ) | ( n30511 & n32669 ) | ( ~n32666 & n32669 ) ;
  assign n32671 = ( ~n3006 & n10263 ) | ( ~n3006 & n14564 ) | ( n10263 & n14564 ) ;
  assign n32672 = n20941 ^ n2247 ^ n1833 ;
  assign n32673 = n32672 ^ n32619 ^ n5348 ;
  assign n32674 = ~n2440 & n14863 ;
  assign n32675 = n32673 & n32674 ;
  assign n32676 = ( n5021 & ~n7960 ) | ( n5021 & n26854 ) | ( ~n7960 & n26854 ) ;
  assign n32677 = n32676 ^ n4957 ^ 1'b0 ;
  assign n32678 = n8230 | n32677 ;
  assign n32679 = ( n3232 & n3256 ) | ( n3232 & n6161 ) | ( n3256 & n6161 ) ;
  assign n32680 = n32679 ^ n32151 ^ n23219 ;
  assign n32681 = n32680 ^ n24114 ^ n12443 ;
  assign n32682 = n32678 | n32681 ;
  assign n32683 = n32682 ^ n14499 ^ 1'b0 ;
  assign n32684 = ~n7021 & n11814 ;
  assign n32685 = n32684 ^ n14835 ^ n3457 ;
  assign n32686 = n22311 ^ n16937 ^ n3439 ;
  assign n32687 = n23682 ^ n21278 ^ n10760 ;
  assign n32691 = n28277 ^ n13936 ^ n6922 ;
  assign n32689 = n32196 ^ n19709 ^ n16470 ;
  assign n32690 = n32689 ^ n19845 ^ n6770 ;
  assign n32688 = n22213 ^ n1172 ^ 1'b0 ;
  assign n32692 = n32691 ^ n32690 ^ n32688 ;
  assign n32693 = ( n32686 & n32687 ) | ( n32686 & n32692 ) | ( n32687 & n32692 ) ;
  assign n32694 = n30081 ^ n3268 ^ n2827 ;
  assign n32695 = n32694 ^ n14356 ^ 1'b0 ;
  assign n32696 = n25621 ^ n12447 ^ n11716 ;
  assign n32697 = n6605 & ~n31334 ;
  assign n32698 = n17824 & ~n21819 ;
  assign n32699 = n32697 & n32698 ;
  assign n32700 = n32111 ^ n20859 ^ n4842 ;
  assign n32701 = n32700 ^ n27183 ^ 1'b0 ;
  assign n32702 = n32701 ^ n16533 ^ n15097 ;
  assign n32705 = n9408 ^ n2181 ^ n1719 ;
  assign n32703 = n31445 ^ n26796 ^ 1'b0 ;
  assign n32704 = n917 & ~n32703 ;
  assign n32706 = n32705 ^ n32704 ^ n32018 ;
  assign n32707 = n10539 ^ n8386 ^ n5416 ;
  assign n32708 = n32707 ^ n23646 ^ n7890 ;
  assign n32709 = ( n3460 & n16140 ) | ( n3460 & ~n27245 ) | ( n16140 & ~n27245 ) ;
  assign n32710 = ( ~x248 & n2076 ) | ( ~x248 & n28283 ) | ( n2076 & n28283 ) ;
  assign n32711 = n24918 | n32710 ;
  assign n32712 = n32711 ^ n1910 ^ 1'b0 ;
  assign n32713 = n32712 ^ n19585 ^ n18311 ;
  assign n32714 = n26309 ^ n11818 ^ n3522 ;
  assign n32715 = n32714 ^ n19153 ^ n15996 ;
  assign n32716 = n21963 ^ n8204 ^ 1'b0 ;
  assign n32717 = n3558 | n32716 ;
  assign n32718 = ( n1445 & n12506 ) | ( n1445 & ~n18816 ) | ( n12506 & ~n18816 ) ;
  assign n32719 = n32718 ^ n11194 ^ n9928 ;
  assign n32720 = ( ~n28218 & n32717 ) | ( ~n28218 & n32719 ) | ( n32717 & n32719 ) ;
  assign n32721 = n19790 | n30475 ;
  assign n32722 = n32721 ^ n26134 ^ 1'b0 ;
  assign n32723 = n18613 ^ n367 ^ 1'b0 ;
  assign n32724 = ~n32722 & n32723 ;
  assign n32725 = n26149 ^ n11270 ^ n8522 ;
  assign n32726 = ( ~n15053 & n31343 ) | ( ~n15053 & n32725 ) | ( n31343 & n32725 ) ;
  assign n32727 = n28150 ^ n14293 ^ 1'b0 ;
  assign n32728 = ( ~n276 & n2433 ) | ( ~n276 & n9669 ) | ( n2433 & n9669 ) ;
  assign n32729 = n32728 ^ n856 ^ 1'b0 ;
  assign n32730 = ~n8385 & n32729 ;
  assign n32731 = n32730 ^ n31622 ^ n1734 ;
  assign n32732 = n20267 ^ n607 ^ 1'b0 ;
  assign n32733 = n6512 ^ n2551 ^ 1'b0 ;
  assign n32734 = ~n4133 & n32733 ;
  assign n32735 = ( x246 & n28866 ) | ( x246 & n32734 ) | ( n28866 & n32734 ) ;
  assign n32736 = n32735 ^ n29127 ^ n9254 ;
  assign n32737 = n24521 ^ n20453 ^ n1146 ;
  assign n32738 = ( n9591 & n11577 ) | ( n9591 & n32737 ) | ( n11577 & n32737 ) ;
  assign n32739 = ( ~n10919 & n31347 ) | ( ~n10919 & n32738 ) | ( n31347 & n32738 ) ;
  assign n32740 = n22036 ^ n7699 ^ n5932 ;
  assign n32741 = n13669 ^ n1356 ^ 1'b0 ;
  assign n32742 = n32741 ^ n9589 ^ n5234 ;
  assign n32743 = ( ~n940 & n32740 ) | ( ~n940 & n32742 ) | ( n32740 & n32742 ) ;
  assign n32744 = x223 & n2856 ;
  assign n32745 = n4788 & n32744 ;
  assign n32746 = n6957 & ~n32745 ;
  assign n32747 = n32746 ^ n12852 ^ 1'b0 ;
  assign n32748 = n18414 ^ n7554 ^ n5448 ;
  assign n32749 = n9964 ^ n5324 ^ 1'b0 ;
  assign n32750 = ~n11659 & n32749 ;
  assign n32751 = ( n32747 & n32748 ) | ( n32747 & ~n32750 ) | ( n32748 & ~n32750 ) ;
  assign n32755 = n22285 ^ n20088 ^ n6927 ;
  assign n32752 = n2009 & ~n2813 ;
  assign n32753 = n32752 ^ n25026 ^ 1'b0 ;
  assign n32754 = ( x228 & ~n15782 ) | ( x228 & n32753 ) | ( ~n15782 & n32753 ) ;
  assign n32756 = n32755 ^ n32754 ^ n3087 ;
  assign n32757 = n32756 ^ n24643 ^ n18016 ;
  assign n32758 = ( n12028 & n18158 ) | ( n12028 & n20409 ) | ( n18158 & n20409 ) ;
  assign n32759 = ( ~n4859 & n19292 ) | ( ~n4859 & n32758 ) | ( n19292 & n32758 ) ;
  assign n32760 = n15087 ^ n8923 ^ n5476 ;
  assign n32761 = ( n10134 & ~n11323 ) | ( n10134 & n23243 ) | ( ~n11323 & n23243 ) ;
  assign n32762 = ( x123 & ~n32760 ) | ( x123 & n32761 ) | ( ~n32760 & n32761 ) ;
  assign n32763 = ( n2984 & ~n27807 ) | ( n2984 & n32762 ) | ( ~n27807 & n32762 ) ;
  assign n32764 = n28487 ^ n20101 ^ 1'b0 ;
  assign n32765 = ( n4083 & ~n11436 ) | ( n4083 & n32764 ) | ( ~n11436 & n32764 ) ;
  assign n32766 = ( x66 & n14256 ) | ( x66 & n21698 ) | ( n14256 & n21698 ) ;
  assign n32767 = ( n11627 & ~n13281 ) | ( n11627 & n32766 ) | ( ~n13281 & n32766 ) ;
  assign n32768 = n5899 | n32767 ;
  assign n32769 = n32768 ^ n15136 ^ 1'b0 ;
  assign n32770 = ( n8180 & n12204 ) | ( n8180 & n14438 ) | ( n12204 & n14438 ) ;
  assign n32771 = n19204 ^ n3935 ^ n1340 ;
  assign n32772 = n26588 | n32771 ;
  assign n32773 = n32772 ^ n3237 ^ 1'b0 ;
  assign n32774 = ( n4338 & ~n18440 ) | ( n4338 & n32773 ) | ( ~n18440 & n32773 ) ;
  assign n32775 = n26200 ^ n22052 ^ n16961 ;
  assign n32776 = ( n8523 & ~n32774 ) | ( n8523 & n32775 ) | ( ~n32774 & n32775 ) ;
  assign n32777 = n32468 ^ n31211 ^ n11214 ;
  assign n32778 = ( n4395 & n7552 ) | ( n4395 & n15151 ) | ( n7552 & n15151 ) ;
  assign n32781 = ( ~n1816 & n15974 ) | ( ~n1816 & n17888 ) | ( n15974 & n17888 ) ;
  assign n32780 = n20415 ^ n13487 ^ n6905 ;
  assign n32779 = n26680 ^ n24824 ^ n3393 ;
  assign n32782 = n32781 ^ n32780 ^ n32779 ;
  assign n32783 = n31378 ^ n25629 ^ n20841 ;
  assign n32784 = ( n339 & n4760 ) | ( n339 & n29304 ) | ( n4760 & n29304 ) ;
  assign n32785 = n32488 ^ n26239 ^ 1'b0 ;
  assign n32786 = n12148 | n26741 ;
  assign n32787 = n7234 | n32786 ;
  assign n32788 = n2697 | n19907 ;
  assign n32789 = n32788 ^ n32472 ^ 1'b0 ;
  assign n32790 = n32789 ^ n12019 ^ n4164 ;
  assign n32791 = n21478 ^ x104 ^ 1'b0 ;
  assign n32792 = n12806 ^ n5012 ^ n2172 ;
  assign n32793 = n27388 & n32792 ;
  assign n32794 = n32793 ^ n16562 ^ 1'b0 ;
  assign n32795 = n32794 ^ n26103 ^ n16319 ;
  assign n32796 = n29875 ^ n1640 ^ n596 ;
  assign n32797 = ( n32380 & ~n32795 ) | ( n32380 & n32796 ) | ( ~n32795 & n32796 ) ;
  assign n32802 = ( n4632 & n14410 ) | ( n4632 & n17799 ) | ( n14410 & n17799 ) ;
  assign n32803 = ( n17201 & ~n17743 ) | ( n17201 & n32802 ) | ( ~n17743 & n32802 ) ;
  assign n32801 = ( ~n3857 & n10850 ) | ( ~n3857 & n10882 ) | ( n10850 & n10882 ) ;
  assign n32798 = ( n3437 & ~n3977 ) | ( n3437 & n19026 ) | ( ~n3977 & n19026 ) ;
  assign n32799 = n32798 ^ n10120 ^ n6098 ;
  assign n32800 = n32799 ^ n23725 ^ n7609 ;
  assign n32804 = n32803 ^ n32801 ^ n32800 ;
  assign n32805 = n4930 ^ n3005 ^ 1'b0 ;
  assign n32806 = n9692 ^ n7873 ^ n2967 ;
  assign n32807 = ~n20133 & n24363 ;
  assign n32808 = n32807 ^ n32548 ^ 1'b0 ;
  assign n32809 = n32808 ^ n17474 ^ n9355 ;
  assign n32810 = ( ~n20478 & n32806 ) | ( ~n20478 & n32809 ) | ( n32806 & n32809 ) ;
  assign n32811 = ( n6903 & n6915 ) | ( n6903 & n12099 ) | ( n6915 & n12099 ) ;
  assign n32812 = n12861 ^ n5399 ^ 1'b0 ;
  assign n32813 = ( n4223 & n29372 ) | ( n4223 & ~n32812 ) | ( n29372 & ~n32812 ) ;
  assign n32814 = n8707 ^ n4076 ^ 1'b0 ;
  assign n32815 = n1805 & n32814 ;
  assign n32816 = ( ~n11692 & n25111 ) | ( ~n11692 & n32815 ) | ( n25111 & n32815 ) ;
  assign n32817 = n32816 ^ n22502 ^ n1391 ;
  assign n32818 = ( n5461 & n11008 ) | ( n5461 & n20957 ) | ( n11008 & n20957 ) ;
  assign n32820 = n18947 ^ n5678 ^ n2103 ;
  assign n32819 = ( n1395 & n3850 ) | ( n1395 & n10287 ) | ( n3850 & n10287 ) ;
  assign n32821 = n32820 ^ n32819 ^ n1358 ;
  assign n32822 = ( n19377 & n32818 ) | ( n19377 & ~n32821 ) | ( n32818 & ~n32821 ) ;
  assign n32823 = ( ~n8527 & n29090 ) | ( ~n8527 & n32822 ) | ( n29090 & n32822 ) ;
  assign n32824 = ~x55 & n22830 ;
  assign n32825 = ~n16059 & n32824 ;
  assign n32826 = ( n9272 & ~n31016 ) | ( n9272 & n32825 ) | ( ~n31016 & n32825 ) ;
  assign n32827 = n32826 ^ n24904 ^ n11574 ;
  assign n32828 = ~n7886 & n32827 ;
  assign n32829 = n32828 ^ n24764 ^ 1'b0 ;
  assign n32830 = n1339 & n15101 ;
  assign n32831 = n8825 & n32830 ;
  assign n32832 = n32831 ^ n31388 ^ n14822 ;
  assign n32834 = ( n693 & n14446 ) | ( n693 & ~n22495 ) | ( n14446 & ~n22495 ) ;
  assign n32833 = n23713 ^ n5657 ^ n900 ;
  assign n32835 = n32834 ^ n32833 ^ n29973 ;
  assign n32836 = ( n1553 & ~n4900 ) | ( n1553 & n19199 ) | ( ~n4900 & n19199 ) ;
  assign n32837 = n6902 ^ n2018 ^ x188 ;
  assign n32838 = ( n2967 & n26184 ) | ( n2967 & n32837 ) | ( n26184 & n32837 ) ;
  assign n32839 = ( n6089 & ~n14987 ) | ( n6089 & n17696 ) | ( ~n14987 & n17696 ) ;
  assign n32840 = n32839 ^ n29100 ^ n9428 ;
  assign n32841 = n32840 ^ n26155 ^ n1562 ;
  assign n32842 = ( ~n2158 & n32838 ) | ( ~n2158 & n32841 ) | ( n32838 & n32841 ) ;
  assign n32843 = n13129 ^ n12657 ^ 1'b0 ;
  assign n32844 = n28232 ^ n14658 ^ n439 ;
  assign n32845 = ~n7764 & n32844 ;
  assign n32846 = n32845 ^ n30564 ^ 1'b0 ;
  assign n32848 = n29393 ^ n27351 ^ n5895 ;
  assign n32847 = n3950 & n18800 ;
  assign n32849 = n32848 ^ n32847 ^ 1'b0 ;
  assign n32850 = ( ~n13296 & n21952 ) | ( ~n13296 & n32849 ) | ( n21952 & n32849 ) ;
  assign n32852 = ( n8119 & n13809 ) | ( n8119 & n19356 ) | ( n13809 & n19356 ) ;
  assign n32853 = ( n1612 & ~n12552 ) | ( n1612 & n32852 ) | ( ~n12552 & n32852 ) ;
  assign n32851 = n30212 ^ n15436 ^ 1'b0 ;
  assign n32854 = n32853 ^ n32851 ^ n20259 ;
  assign n32855 = n25167 ^ n21724 ^ 1'b0 ;
  assign n32856 = n5762 & ~n26477 ;
  assign n32860 = ~n11850 & n19275 ;
  assign n32857 = ~n3123 & n11725 ;
  assign n32858 = ~n11912 & n32857 ;
  assign n32859 = n32858 ^ n11222 ^ n1120 ;
  assign n32861 = n32860 ^ n32859 ^ n16067 ;
  assign n32862 = n19272 ^ n7981 ^ n3851 ;
  assign n32863 = n32862 ^ n20397 ^ n6986 ;
  assign n32864 = n12269 ^ n6267 ^ n5204 ;
  assign n32865 = n32864 ^ n24988 ^ n7347 ;
  assign n32866 = ( ~n2455 & n12291 ) | ( ~n2455 & n32865 ) | ( n12291 & n32865 ) ;
  assign n32867 = n32863 | n32866 ;
  assign n32868 = n19504 | n32867 ;
  assign n32869 = n32868 ^ n5693 ^ n3584 ;
  assign n32870 = n5356 & ~n28532 ;
  assign n32871 = n32870 ^ n1411 ^ 1'b0 ;
  assign n32872 = n11666 ^ n3770 ^ n2457 ;
  assign n32873 = ( n938 & n2367 ) | ( n938 & n32872 ) | ( n2367 & n32872 ) ;
  assign n32875 = n4176 ^ n1726 ^ x195 ;
  assign n32876 = n26763 & ~n32875 ;
  assign n32874 = n5099 | n5757 ;
  assign n32877 = n32876 ^ n32874 ^ 1'b0 ;
  assign n32878 = n32877 ^ n30198 ^ n27257 ;
  assign n32879 = n28356 ^ n1227 ^ 1'b0 ;
  assign n32880 = ( n7052 & ~n20674 ) | ( n7052 & n29231 ) | ( ~n20674 & n29231 ) ;
  assign n32881 = ( ~n3564 & n7289 ) | ( ~n3564 & n27639 ) | ( n7289 & n27639 ) ;
  assign n32882 = n32881 ^ n31152 ^ n27871 ;
  assign n32884 = ( ~n12841 & n22124 ) | ( ~n12841 & n26010 ) | ( n22124 & n26010 ) ;
  assign n32883 = ( ~n9182 & n9789 ) | ( ~n9182 & n25712 ) | ( n9789 & n25712 ) ;
  assign n32885 = n32884 ^ n32883 ^ n18582 ;
  assign n32886 = n12810 ^ n7049 ^ 1'b0 ;
  assign n32887 = n3858 & ~n32886 ;
  assign n32888 = n29925 ^ n27963 ^ n23433 ;
  assign n32889 = ( n11669 & n21732 ) | ( n11669 & ~n32888 ) | ( n21732 & ~n32888 ) ;
  assign n32890 = ( n18309 & ~n21166 ) | ( n18309 & n32889 ) | ( ~n21166 & n32889 ) ;
  assign n32891 = n26042 ^ n22764 ^ n2062 ;
  assign n32892 = ( n32887 & ~n32890 ) | ( n32887 & n32891 ) | ( ~n32890 & n32891 ) ;
  assign n32893 = ( n469 & ~n4977 ) | ( n469 & n26278 ) | ( ~n4977 & n26278 ) ;
  assign n32894 = ( n26356 & n28991 ) | ( n26356 & n32893 ) | ( n28991 & n32893 ) ;
  assign n32895 = n9014 ^ x52 ^ 1'b0 ;
  assign n32896 = n32895 ^ n25937 ^ n12396 ;
  assign n32897 = n32896 ^ n20369 ^ n19804 ;
  assign n32898 = ( n7388 & ~n10556 ) | ( n7388 & n24370 ) | ( ~n10556 & n24370 ) ;
  assign n32899 = n32898 ^ n10144 ^ n9350 ;
  assign n32900 = n11466 | n17409 ;
  assign n32901 = n32900 ^ n13687 ^ 1'b0 ;
  assign n32902 = ( n15103 & n27373 ) | ( n15103 & n28285 ) | ( n27373 & n28285 ) ;
  assign n32903 = ( n809 & n22953 ) | ( n809 & n27990 ) | ( n22953 & n27990 ) ;
  assign n32904 = n6799 & n19888 ;
  assign n32905 = ( ~n16769 & n26611 ) | ( ~n16769 & n32904 ) | ( n26611 & n32904 ) ;
  assign n32906 = n16304 ^ n10865 ^ n9278 ;
  assign n32907 = ( n7103 & ~n26751 ) | ( n7103 & n30730 ) | ( ~n26751 & n30730 ) ;
  assign n32908 = ( ~n8782 & n12376 ) | ( ~n8782 & n32907 ) | ( n12376 & n32907 ) ;
  assign n32909 = ~n12623 & n23326 ;
  assign n32910 = n10570 & ~n26961 ;
  assign n32911 = n32910 ^ n3558 ^ 1'b0 ;
  assign n32912 = n32911 ^ n9787 ^ 1'b0 ;
  assign n32913 = ( ~n3273 & n11781 ) | ( ~n3273 & n21780 ) | ( n11781 & n21780 ) ;
  assign n32914 = n32913 ^ n32572 ^ n1269 ;
  assign n32915 = ~n9147 & n9886 ;
  assign n32916 = n21245 & n32915 ;
  assign n32917 = ( n11046 & n12621 ) | ( n11046 & n13714 ) | ( n12621 & n13714 ) ;
  assign n32918 = n32917 ^ n5990 ^ 1'b0 ;
  assign n32919 = ( n2713 & n13616 ) | ( n2713 & n32918 ) | ( n13616 & n32918 ) ;
  assign n32920 = ( n7216 & n32916 ) | ( n7216 & n32919 ) | ( n32916 & n32919 ) ;
  assign n32921 = ( x62 & n5263 ) | ( x62 & n32920 ) | ( n5263 & n32920 ) ;
  assign n32923 = ( n1195 & n3237 ) | ( n1195 & ~n5076 ) | ( n3237 & ~n5076 ) ;
  assign n32922 = n10838 ^ n7659 ^ x68 ;
  assign n32924 = n32923 ^ n32922 ^ n20002 ;
  assign n32925 = ( ~n15699 & n26693 ) | ( ~n15699 & n32180 ) | ( n26693 & n32180 ) ;
  assign n32926 = n3484 ^ n3037 ^ n1524 ;
  assign n32927 = n12659 | n32926 ;
  assign n32928 = ( n7208 & n14516 ) | ( n7208 & ~n25763 ) | ( n14516 & ~n25763 ) ;
  assign n32929 = ( n32925 & ~n32927 ) | ( n32925 & n32928 ) | ( ~n32927 & n32928 ) ;
  assign n32930 = n7430 ^ n5192 ^ 1'b0 ;
  assign n32931 = ( n4116 & n13596 ) | ( n4116 & ~n30627 ) | ( n13596 & ~n30627 ) ;
  assign n32932 = ( n7965 & n10380 ) | ( n7965 & ~n32931 ) | ( n10380 & ~n32931 ) ;
  assign n32933 = n32932 ^ n8228 ^ 1'b0 ;
  assign n32934 = ( n8699 & n11529 ) | ( n8699 & ~n32933 ) | ( n11529 & ~n32933 ) ;
  assign n32935 = n17110 ^ n3360 ^ n624 ;
  assign n32936 = n12556 | n27224 ;
  assign n32937 = n32936 ^ n18255 ^ n11460 ;
  assign n32938 = n32728 ^ n11704 ^ n7946 ;
  assign n32939 = ( n3564 & ~n5184 ) | ( n3564 & n8147 ) | ( ~n5184 & n8147 ) ;
  assign n32940 = ( n3448 & n32938 ) | ( n3448 & n32939 ) | ( n32938 & n32939 ) ;
  assign n32942 = n28720 ^ n27012 ^ n19453 ;
  assign n32941 = ( n3728 & n19393 ) | ( n3728 & n21022 ) | ( n19393 & n21022 ) ;
  assign n32943 = n32942 ^ n32941 ^ n25738 ;
  assign n32948 = n5097 & ~n16606 ;
  assign n32949 = n8524 & n32948 ;
  assign n32944 = ( n1127 & ~n18581 ) | ( n1127 & n20903 ) | ( ~n18581 & n20903 ) ;
  assign n32945 = n29270 ^ n6618 ^ 1'b0 ;
  assign n32946 = n22683 & ~n32945 ;
  assign n32947 = ( n17862 & n32944 ) | ( n17862 & ~n32946 ) | ( n32944 & ~n32946 ) ;
  assign n32950 = n32949 ^ n32947 ^ n20503 ;
  assign n32951 = ( n6919 & n8880 ) | ( n6919 & n23156 ) | ( n8880 & n23156 ) ;
  assign n32952 = n32951 ^ n25368 ^ n21333 ;
  assign n32953 = n32952 ^ n11281 ^ 1'b0 ;
  assign n32954 = n32953 ^ n30878 ^ n16310 ;
  assign n32955 = n8741 ^ n2271 ^ 1'b0 ;
  assign n32956 = n24074 ^ n12123 ^ x86 ;
  assign n32957 = n32956 ^ n16644 ^ n6076 ;
  assign n32958 = n10842 ^ n6724 ^ n3539 ;
  assign n32959 = ( n6113 & ~n7335 ) | ( n6113 & n32958 ) | ( ~n7335 & n32958 ) ;
  assign n32960 = n32959 ^ n30216 ^ n4784 ;
  assign n32961 = n32960 ^ n27506 ^ n21732 ;
  assign n32963 = ~n5090 & n17201 ;
  assign n32962 = n8897 ^ n6784 ^ 1'b0 ;
  assign n32964 = n32963 ^ n32962 ^ n7725 ;
  assign n32965 = ( n3147 & ~n32961 ) | ( n3147 & n32964 ) | ( ~n32961 & n32964 ) ;
  assign n32966 = n18284 ^ n11046 ^ n5393 ;
  assign n32967 = n3868 & n23688 ;
  assign n32968 = n32967 ^ n16416 ^ n12376 ;
  assign n32969 = ( x236 & n14592 ) | ( x236 & n16203 ) | ( n14592 & n16203 ) ;
  assign n32970 = ( n10455 & n22268 ) | ( n10455 & ~n32969 ) | ( n22268 & ~n32969 ) ;
  assign n32971 = n5571 & ~n9580 ;
  assign n32972 = ( n6667 & n30848 ) | ( n6667 & n32971 ) | ( n30848 & n32971 ) ;
  assign n32973 = ( n9202 & ~n15589 ) | ( n9202 & n32972 ) | ( ~n15589 & n32972 ) ;
  assign n32974 = n22970 | n32973 ;
  assign n32975 = n32970 | n32974 ;
  assign n32978 = n13594 & n24782 ;
  assign n32976 = n27850 ^ n2406 ^ 1'b0 ;
  assign n32977 = ( n11974 & ~n31385 ) | ( n11974 & n32976 ) | ( ~n31385 & n32976 ) ;
  assign n32979 = n32978 ^ n32977 ^ n6711 ;
  assign n32980 = ~n2948 & n9788 ;
  assign n32981 = n32979 & n32980 ;
  assign n32982 = n23825 ^ n20960 ^ n363 ;
  assign n32983 = n29622 ^ n21415 ^ n15159 ;
  assign n32984 = n32983 ^ n26593 ^ n7214 ;
  assign n32985 = ( n313 & n13218 ) | ( n313 & ~n18385 ) | ( n13218 & ~n18385 ) ;
  assign n32986 = ( ~n9395 & n18273 ) | ( ~n9395 & n32985 ) | ( n18273 & n32985 ) ;
  assign n32987 = n32986 ^ n13124 ^ n4248 ;
  assign n32988 = n18500 & ~n25436 ;
  assign n32989 = ( n7714 & ~n13160 ) | ( n7714 & n32988 ) | ( ~n13160 & n32988 ) ;
  assign n32990 = ( n1511 & n9519 ) | ( n1511 & n10010 ) | ( n9519 & n10010 ) ;
  assign n32991 = ( n1708 & ~n20414 ) | ( n1708 & n32990 ) | ( ~n20414 & n32990 ) ;
  assign n32992 = ( n5707 & n32989 ) | ( n5707 & n32991 ) | ( n32989 & n32991 ) ;
  assign n32993 = ( n11156 & n12195 ) | ( n11156 & ~n18780 ) | ( n12195 & ~n18780 ) ;
  assign n32994 = n1497 | n10775 ;
  assign n32995 = n2081 & ~n32994 ;
  assign n32996 = ( n832 & ~n7601 ) | ( n832 & n28954 ) | ( ~n7601 & n28954 ) ;
  assign n32997 = n17446 & ~n17480 ;
  assign n32998 = n32997 ^ n13744 ^ 1'b0 ;
  assign n32999 = n7103 | n32998 ;
  assign n33000 = n19135 & n32999 ;
  assign n33001 = ~n32996 & n33000 ;
  assign n33002 = n32995 | n33001 ;
  assign n33003 = n32993 | n33002 ;
  assign n33004 = n29296 ^ n27225 ^ n10167 ;
  assign n33005 = ( n26279 & ~n30398 ) | ( n26279 & n30710 ) | ( ~n30398 & n30710 ) ;
  assign n33006 = n11308 ^ n4724 ^ n449 ;
  assign n33007 = n9484 | n33006 ;
  assign n33008 = n33007 ^ n22446 ^ n13117 ;
  assign n33011 = ( n1905 & ~n2279 ) | ( n1905 & n2756 ) | ( ~n2279 & n2756 ) ;
  assign n33009 = n30642 ^ n21984 ^ n19914 ;
  assign n33010 = ( n3733 & n5013 ) | ( n3733 & ~n33009 ) | ( n5013 & ~n33009 ) ;
  assign n33012 = n33011 ^ n33010 ^ 1'b0 ;
  assign n33013 = n947 & ~n20133 ;
  assign n33014 = ~n9858 & n33013 ;
  assign n33016 = ( n3748 & ~n8065 ) | ( n3748 & n12627 ) | ( ~n8065 & n12627 ) ;
  assign n33015 = n14124 ^ n11220 ^ n7710 ;
  assign n33017 = n33016 ^ n33015 ^ n32463 ;
  assign n33018 = n27320 ^ n21106 ^ n20442 ;
  assign n33019 = n33018 ^ n19545 ^ n9925 ;
  assign n33021 = n13630 ^ n2022 ^ n544 ;
  assign n33022 = n33021 ^ n435 ^ n346 ;
  assign n33023 = n11187 & n25155 ;
  assign n33024 = n33023 ^ n31034 ^ 1'b0 ;
  assign n33025 = ( n22803 & ~n33022 ) | ( n22803 & n33024 ) | ( ~n33022 & n33024 ) ;
  assign n33020 = n18980 ^ n17765 ^ n15485 ;
  assign n33026 = n33025 ^ n33020 ^ n13634 ;
  assign n33027 = ( n1052 & n29117 ) | ( n1052 & n33026 ) | ( n29117 & n33026 ) ;
  assign n33028 = n21434 ^ n12793 ^ n8501 ;
  assign n33029 = n32839 ^ n24517 ^ n15333 ;
  assign n33030 = n33029 ^ n24821 ^ n8930 ;
  assign n33038 = n17449 ^ n11315 ^ n9524 ;
  assign n33031 = n12803 ^ n7037 ^ n579 ;
  assign n33032 = n33031 ^ n11809 ^ n11352 ;
  assign n33033 = n33032 ^ n9140 ^ 1'b0 ;
  assign n33034 = n9165 | n33033 ;
  assign n33035 = ( n2874 & n7451 ) | ( n2874 & ~n9613 ) | ( n7451 & ~n9613 ) ;
  assign n33036 = n33035 ^ n16969 ^ n8153 ;
  assign n33037 = n33034 & n33036 ;
  assign n33039 = n33038 ^ n33037 ^ 1'b0 ;
  assign n33040 = ~n12120 & n33039 ;
  assign n33042 = ( n4323 & n16558 ) | ( n4323 & n27941 ) | ( n16558 & n27941 ) ;
  assign n33041 = ( n11604 & ~n20180 ) | ( n11604 & n30950 ) | ( ~n20180 & n30950 ) ;
  assign n33043 = n33042 ^ n33041 ^ n14889 ;
  assign n33044 = n25054 ^ n24017 ^ n10484 ;
  assign n33046 = n8032 ^ n6450 ^ n3294 ;
  assign n33045 = ~n2517 & n9792 ;
  assign n33047 = n33046 ^ n33045 ^ n19339 ;
  assign n33048 = n28100 | n33047 ;
  assign n33049 = n33048 ^ n23841 ^ 1'b0 ;
  assign n33050 = n33049 ^ n10560 ^ 1'b0 ;
  assign n33053 = ( n2065 & n20140 ) | ( n2065 & ~n27256 ) | ( n20140 & ~n27256 ) ;
  assign n33051 = ( n2104 & n8576 ) | ( n2104 & n11674 ) | ( n8576 & n11674 ) ;
  assign n33052 = ( ~n22128 & n30312 ) | ( ~n22128 & n33051 ) | ( n30312 & n33051 ) ;
  assign n33054 = n33053 ^ n33052 ^ 1'b0 ;
  assign n33055 = n28233 ^ n27894 ^ n5521 ;
  assign n33056 = ( n9621 & n15494 ) | ( n9621 & n33055 ) | ( n15494 & n33055 ) ;
  assign n33057 = n30543 ^ n19424 ^ n17282 ;
  assign n33058 = n17454 | n33057 ;
  assign n33059 = n33056 & ~n33058 ;
  assign n33060 = n806 ^ n376 ^ 1'b0 ;
  assign n33061 = n622 & n33060 ;
  assign n33062 = n33061 ^ n3858 ^ 1'b0 ;
  assign n33063 = ~n4252 & n33062 ;
  assign n33064 = ( n12431 & ~n15471 ) | ( n12431 & n16371 ) | ( ~n15471 & n16371 ) ;
  assign n33065 = ( ~n21981 & n33063 ) | ( ~n21981 & n33064 ) | ( n33063 & n33064 ) ;
  assign n33066 = ( n2274 & ~n3149 ) | ( n2274 & n5231 ) | ( ~n3149 & n5231 ) ;
  assign n33067 = ( n10228 & n10866 ) | ( n10228 & n33066 ) | ( n10866 & n33066 ) ;
  assign n33068 = n33067 ^ n30740 ^ n13387 ;
  assign n33069 = ~n27768 & n33068 ;
  assign n33070 = ~n33065 & n33069 ;
  assign n33071 = ( n3228 & ~n8456 ) | ( n3228 & n9259 ) | ( ~n8456 & n9259 ) ;
  assign n33072 = ( ~n8788 & n13340 ) | ( ~n8788 & n14793 ) | ( n13340 & n14793 ) ;
  assign n33073 = ( n5006 & ~n33071 ) | ( n5006 & n33072 ) | ( ~n33071 & n33072 ) ;
  assign n33074 = n29915 ^ n16803 ^ 1'b0 ;
  assign n33076 = ( n8799 & ~n8931 ) | ( n8799 & n10291 ) | ( ~n8931 & n10291 ) ;
  assign n33077 = n33076 ^ n1519 ^ x0 ;
  assign n33075 = n8067 ^ x93 ^ 1'b0 ;
  assign n33078 = n33077 ^ n33075 ^ n13504 ;
  assign n33079 = ~n15715 & n18457 ;
  assign n33080 = n22930 ^ n10512 ^ n7654 ;
  assign n33081 = ( n5356 & n9428 ) | ( n5356 & n31741 ) | ( n9428 & n31741 ) ;
  assign n33082 = ( n3919 & ~n3939 ) | ( n3919 & n14769 ) | ( ~n3939 & n14769 ) ;
  assign n33083 = n26818 ^ n9359 ^ n835 ;
  assign n33084 = ( n33081 & n33082 ) | ( n33081 & ~n33083 ) | ( n33082 & ~n33083 ) ;
  assign n33085 = n10683 ^ n314 ^ 1'b0 ;
  assign n33086 = ~n8622 & n33085 ;
  assign n33087 = n3623 & ~n27980 ;
  assign n33088 = n33087 ^ n16087 ^ 1'b0 ;
  assign n33089 = n33088 ^ n19849 ^ n13283 ;
  assign n33090 = n18371 & ~n33089 ;
  assign n33091 = ~n28489 & n33090 ;
  assign n33092 = ( ~x248 & n1080 ) | ( ~x248 & n1348 ) | ( n1080 & n1348 ) ;
  assign n33093 = n33092 ^ n18414 ^ n18104 ;
  assign n33094 = ( ~n23807 & n33091 ) | ( ~n23807 & n33093 ) | ( n33091 & n33093 ) ;
  assign n33095 = n31690 ^ n18621 ^ n14818 ;
  assign n33096 = ( ~n10293 & n21902 ) | ( ~n10293 & n33095 ) | ( n21902 & n33095 ) ;
  assign n33097 = ( n31227 & n33094 ) | ( n31227 & ~n33096 ) | ( n33094 & ~n33096 ) ;
  assign n33099 = n11076 ^ n10378 ^ n5335 ;
  assign n33098 = n20181 ^ n7505 ^ n6961 ;
  assign n33100 = n33099 ^ n33098 ^ n26933 ;
  assign n33103 = n11398 ^ n9052 ^ n8070 ;
  assign n33104 = ( n12969 & n15872 ) | ( n12969 & n33103 ) | ( n15872 & n33103 ) ;
  assign n33101 = n9687 ^ n5407 ^ n1461 ;
  assign n33102 = n33101 ^ n20609 ^ n1189 ;
  assign n33105 = n33104 ^ n33102 ^ n16102 ;
  assign n33106 = ( n5607 & n16473 ) | ( n5607 & ~n33105 ) | ( n16473 & ~n33105 ) ;
  assign n33107 = ( n1499 & n4451 ) | ( n1499 & ~n14258 ) | ( n4451 & ~n14258 ) ;
  assign n33108 = n33107 ^ n26382 ^ 1'b0 ;
  assign n33109 = ( ~n5345 & n12841 ) | ( ~n5345 & n20212 ) | ( n12841 & n20212 ) ;
  assign n33110 = n19922 ^ n18119 ^ n18107 ;
  assign n33111 = n33110 ^ n25995 ^ n13718 ;
  assign n33112 = n16650 ^ n14887 ^ 1'b0 ;
  assign n33113 = n14190 ^ n865 ^ n747 ;
  assign n33114 = n33113 ^ n733 ^ x216 ;
  assign n33115 = ( ~n2392 & n28136 ) | ( ~n2392 & n31812 ) | ( n28136 & n31812 ) ;
  assign n33116 = n33115 ^ n9411 ^ 1'b0 ;
  assign n33117 = ( n33112 & n33114 ) | ( n33112 & n33116 ) | ( n33114 & n33116 ) ;
  assign n33118 = n17845 & ~n30901 ;
  assign n33119 = ( n4301 & n29660 ) | ( n4301 & n33118 ) | ( n29660 & n33118 ) ;
  assign n33120 = n20138 ^ n4652 ^ n2647 ;
  assign n33122 = n19091 ^ n1131 ^ n959 ;
  assign n33123 = n33122 ^ n21208 ^ n9730 ;
  assign n33121 = n26390 ^ n12056 ^ 1'b0 ;
  assign n33124 = n33123 ^ n33121 ^ n2286 ;
  assign n33125 = ( n7465 & n33120 ) | ( n7465 & n33124 ) | ( n33120 & n33124 ) ;
  assign n33126 = n26849 ^ n6686 ^ n2398 ;
  assign n33127 = n19849 ^ n8317 ^ n1532 ;
  assign n33128 = n27118 ^ n25410 ^ n17193 ;
  assign n33129 = ~n13009 & n33128 ;
  assign n33130 = ~n25416 & n33129 ;
  assign n33131 = ( n8959 & n33127 ) | ( n8959 & n33130 ) | ( n33127 & n33130 ) ;
  assign n33132 = n547 & n4645 ;
  assign n33133 = n33132 ^ n11539 ^ n7604 ;
  assign n33134 = n2719 & ~n15114 ;
  assign n33135 = n33134 ^ n11249 ^ 1'b0 ;
  assign n33136 = ~n5897 & n33135 ;
  assign n33137 = n3837 & n33136 ;
  assign n33138 = ( n6071 & ~n6197 ) | ( n6071 & n33137 ) | ( ~n6197 & n33137 ) ;
  assign n33139 = ( n2852 & n6259 ) | ( n2852 & n9886 ) | ( n6259 & n9886 ) ;
  assign n33140 = n33139 ^ n22433 ^ n4441 ;
  assign n33141 = n10386 ^ n10272 ^ n4913 ;
  assign n33142 = n33141 ^ n11001 ^ n2692 ;
  assign n33143 = n22731 ^ n7399 ^ n4648 ;
  assign n33144 = ( n18101 & n18268 ) | ( n18101 & ~n32248 ) | ( n18268 & ~n32248 ) ;
  assign n33145 = ( ~n26020 & n33143 ) | ( ~n26020 & n33144 ) | ( n33143 & n33144 ) ;
  assign n33146 = ( ~n3674 & n3923 ) | ( ~n3674 & n29556 ) | ( n3923 & n29556 ) ;
  assign n33147 = n12662 ^ n9950 ^ n476 ;
  assign n33148 = ( n20460 & n33146 ) | ( n20460 & ~n33147 ) | ( n33146 & ~n33147 ) ;
  assign n33150 = n17333 ^ n2751 ^ n1985 ;
  assign n33149 = n9630 ^ n8331 ^ n8188 ;
  assign n33151 = n33150 ^ n33149 ^ n11673 ;
  assign n33152 = n13938 | n28345 ;
  assign n33153 = n12731 | n33152 ;
  assign n33154 = n22599 ^ n19782 ^ n13175 ;
  assign n33155 = n33154 ^ n17233 ^ n10740 ;
  assign n33156 = n18831 ^ n9352 ^ n8611 ;
  assign n33157 = n4000 & ~n14854 ;
  assign n33158 = ( n30750 & n33156 ) | ( n30750 & n33157 ) | ( n33156 & n33157 ) ;
  assign n33162 = n17479 ^ n13803 ^ n10991 ;
  assign n33161 = n25366 ^ n15064 ^ 1'b0 ;
  assign n33159 = ( n2535 & n3739 ) | ( n2535 & n5960 ) | ( n3739 & n5960 ) ;
  assign n33160 = n33159 ^ n5882 ^ n3652 ;
  assign n33163 = n33162 ^ n33161 ^ n33160 ;
  assign n33164 = n12335 ^ n11855 ^ n9469 ;
  assign n33165 = n27917 & n31662 ;
  assign n33166 = ( n9102 & ~n31856 ) | ( n9102 & n33165 ) | ( ~n31856 & n33165 ) ;
  assign n33167 = n22554 ^ n4632 ^ n1618 ;
  assign n33168 = n33167 ^ n10430 ^ n7264 ;
  assign n33169 = n18900 ^ n8377 ^ 1'b0 ;
  assign n33170 = n25670 & ~n33169 ;
  assign n33171 = ( ~n11745 & n29883 ) | ( ~n11745 & n33170 ) | ( n29883 & n33170 ) ;
  assign n33172 = n7909 & n14047 ;
  assign n33173 = n7202 & n33172 ;
  assign n33174 = ( n5505 & n30194 ) | ( n5505 & ~n33173 ) | ( n30194 & ~n33173 ) ;
  assign n33175 = n25629 ^ n2703 ^ n520 ;
  assign n33176 = ( n4411 & ~n8667 ) | ( n4411 & n33175 ) | ( ~n8667 & n33175 ) ;
  assign n33177 = ( n8768 & n20377 ) | ( n8768 & ~n22329 ) | ( n20377 & ~n22329 ) ;
  assign n33183 = n19501 ^ n3048 ^ 1'b0 ;
  assign n33184 = ( ~n331 & n2760 ) | ( ~n331 & n3086 ) | ( n2760 & n3086 ) ;
  assign n33185 = ( x245 & n2666 ) | ( x245 & n33184 ) | ( n2666 & n33184 ) ;
  assign n33186 = n33185 ^ n15423 ^ n3793 ;
  assign n33187 = ( n4435 & n33183 ) | ( n4435 & n33186 ) | ( n33183 & n33186 ) ;
  assign n33178 = ( n293 & n2668 ) | ( n293 & ~n8005 ) | ( n2668 & ~n8005 ) ;
  assign n33179 = n33178 ^ n14010 ^ 1'b0 ;
  assign n33180 = n25224 & n33179 ;
  assign n33181 = ( ~n8236 & n10833 ) | ( ~n8236 & n33180 ) | ( n10833 & n33180 ) ;
  assign n33182 = ~n9238 & n33181 ;
  assign n33188 = n33187 ^ n33182 ^ 1'b0 ;
  assign n33189 = n1605 | n33188 ;
  assign n33190 = ( n3995 & n7719 ) | ( n3995 & n30445 ) | ( n7719 & n30445 ) ;
  assign n33191 = n26694 ^ n22626 ^ n6229 ;
  assign n33192 = ( n8849 & n26933 ) | ( n8849 & ~n33191 ) | ( n26933 & ~n33191 ) ;
  assign n33193 = n19206 ^ n4465 ^ n3586 ;
  assign n33194 = n33193 ^ n1783 ^ 1'b0 ;
  assign n33195 = n20142 & ~n33194 ;
  assign n33196 = n33195 ^ n3888 ^ 1'b0 ;
  assign n33197 = n1049 & ~n20661 ;
  assign n33198 = n33197 ^ n32567 ^ n14394 ;
  assign n33199 = n19386 ^ n11006 ^ n2575 ;
  assign n33200 = n807 & n33199 ;
  assign n33201 = ( n15181 & n24812 ) | ( n15181 & n29069 ) | ( n24812 & n29069 ) ;
  assign n33202 = n33201 ^ n19988 ^ n18589 ;
  assign n33203 = n14243 ^ n10698 ^ 1'b0 ;
  assign n33204 = n2230 | n33203 ;
  assign n33205 = n33204 ^ x16 ^ 1'b0 ;
  assign n33206 = n8448 & ~n33205 ;
  assign n33207 = n19623 ^ n11926 ^ n3496 ;
  assign n33208 = n33207 ^ n30706 ^ n19029 ;
  assign n33209 = n33208 ^ n27598 ^ n18774 ;
  assign n33210 = n18588 ^ n11097 ^ n6747 ;
  assign n33211 = ( n22973 & n26893 ) | ( n22973 & ~n33210 ) | ( n26893 & ~n33210 ) ;
  assign n33212 = n17678 & ~n33211 ;
  assign n33213 = n25668 ^ n14282 ^ 1'b0 ;
  assign n33214 = n10331 & n33213 ;
  assign n33215 = n33214 ^ n1812 ^ n1222 ;
  assign n33216 = ( n5806 & n17513 ) | ( n5806 & ~n31528 ) | ( n17513 & ~n31528 ) ;
  assign n33217 = n33216 ^ n16344 ^ n12948 ;
  assign n33218 = ( n5203 & n6514 ) | ( n5203 & ~n27116 ) | ( n6514 & ~n27116 ) ;
  assign n33219 = n33218 ^ n30741 ^ n30365 ;
  assign n33220 = ( n5492 & ~n33217 ) | ( n5492 & n33219 ) | ( ~n33217 & n33219 ) ;
  assign n33221 = n3511 | n7239 ;
  assign n33222 = n4406 | n10944 ;
  assign n33223 = n33221 & ~n33222 ;
  assign n33224 = n17373 | n24683 ;
  assign n33225 = n15076 | n33224 ;
  assign n33226 = n22966 ^ n22588 ^ n3541 ;
  assign n33227 = ( n3840 & n8289 ) | ( n3840 & n33226 ) | ( n8289 & n33226 ) ;
  assign n33228 = n15452 ^ n7783 ^ n5111 ;
  assign n33229 = n21854 ^ n14187 ^ n8101 ;
  assign n33230 = ( ~n5841 & n21770 ) | ( ~n5841 & n27706 ) | ( n21770 & n27706 ) ;
  assign n33231 = n33230 ^ n21743 ^ 1'b0 ;
  assign n33232 = x115 & ~n9623 ;
  assign n33233 = n33232 ^ n20130 ^ 1'b0 ;
  assign n33234 = ( n28512 & n33231 ) | ( n28512 & n33233 ) | ( n33231 & n33233 ) ;
  assign n33235 = n14280 & ~n19700 ;
  assign n33236 = ( n3349 & n9893 ) | ( n3349 & ~n18239 ) | ( n9893 & ~n18239 ) ;
  assign n33237 = ( ~n19782 & n33235 ) | ( ~n19782 & n33236 ) | ( n33235 & n33236 ) ;
  assign n33238 = ( n4240 & ~n14961 ) | ( n4240 & n26930 ) | ( ~n14961 & n26930 ) ;
  assign n33239 = n33238 ^ n13638 ^ n4148 ;
  assign n33240 = n9461 & ~n13932 ;
  assign n33241 = ( n2780 & ~n21820 ) | ( n2780 & n26455 ) | ( ~n21820 & n26455 ) ;
  assign n33242 = ( n29270 & n29318 ) | ( n29270 & n33241 ) | ( n29318 & n33241 ) ;
  assign n33243 = ( n19708 & ~n33240 ) | ( n19708 & n33242 ) | ( ~n33240 & n33242 ) ;
  assign n33244 = ~n3791 & n14604 ;
  assign n33245 = ( n6510 & n13501 ) | ( n6510 & ~n19658 ) | ( n13501 & ~n19658 ) ;
  assign n33246 = ( n27515 & n33244 ) | ( n27515 & ~n33245 ) | ( n33244 & ~n33245 ) ;
  assign n33249 = n4294 ^ n3264 ^ 1'b0 ;
  assign n33247 = ( n5858 & n11556 ) | ( n5858 & n19655 ) | ( n11556 & n19655 ) ;
  assign n33248 = n33247 ^ n4828 ^ n1447 ;
  assign n33250 = n33249 ^ n33248 ^ n16866 ;
  assign n33251 = n33250 ^ n11651 ^ n337 ;
  assign n33252 = n33251 ^ n21949 ^ n10763 ;
  assign n33259 = ~n6279 & n15321 ;
  assign n33260 = ~n9457 & n33259 ;
  assign n33257 = ( n8960 & n10080 ) | ( n8960 & n12478 ) | ( n10080 & n12478 ) ;
  assign n33258 = ( n6053 & n25844 ) | ( n6053 & n33257 ) | ( n25844 & n33257 ) ;
  assign n33253 = n15118 ^ n13936 ^ n3530 ;
  assign n33254 = ( n10763 & ~n23463 ) | ( n10763 & n33253 ) | ( ~n23463 & n33253 ) ;
  assign n33255 = n13052 | n33254 ;
  assign n33256 = ( n2105 & ~n19214 ) | ( n2105 & n33255 ) | ( ~n19214 & n33255 ) ;
  assign n33261 = n33260 ^ n33258 ^ n33256 ;
  assign n33262 = ( n1109 & ~n16135 ) | ( n1109 & n27230 ) | ( ~n16135 & n27230 ) ;
  assign n33263 = ( ~n2546 & n3478 ) | ( ~n2546 & n11169 ) | ( n3478 & n11169 ) ;
  assign n33264 = n33263 ^ n17362 ^ n16066 ;
  assign n33265 = n28348 ^ n7625 ^ n2506 ;
  assign n33266 = ( n24892 & ~n25818 ) | ( n24892 & n33265 ) | ( ~n25818 & n33265 ) ;
  assign n33267 = ( ~n11741 & n13834 ) | ( ~n11741 & n28437 ) | ( n13834 & n28437 ) ;
  assign n33268 = ( ~n12218 & n16495 ) | ( ~n12218 & n27562 ) | ( n16495 & n27562 ) ;
  assign n33269 = ( n9384 & ~n33267 ) | ( n9384 & n33268 ) | ( ~n33267 & n33268 ) ;
  assign n33272 = n5818 & n7686 ;
  assign n33270 = n10709 ^ n4558 ^ n283 ;
  assign n33271 = n33270 ^ n7423 ^ n4728 ;
  assign n33273 = n33272 ^ n33271 ^ n19874 ;
  assign n33274 = n33273 ^ n1142 ^ 1'b0 ;
  assign n33275 = ( n424 & n8025 ) | ( n424 & ~n8084 ) | ( n8025 & ~n8084 ) ;
  assign n33276 = ( n2145 & ~n27473 ) | ( n2145 & n33275 ) | ( ~n27473 & n33275 ) ;
  assign n33278 = n27865 ^ n23840 ^ 1'b0 ;
  assign n33277 = n27991 ^ n19121 ^ n3941 ;
  assign n33279 = n33278 ^ n33277 ^ n9848 ;
  assign n33280 = ( n17955 & ~n25028 ) | ( n17955 & n31001 ) | ( ~n25028 & n31001 ) ;
  assign n33281 = n6453 ^ n4976 ^ 1'b0 ;
  assign n33282 = ( n11361 & n33280 ) | ( n11361 & ~n33281 ) | ( n33280 & ~n33281 ) ;
  assign n33283 = n33282 ^ n9368 ^ n2758 ;
  assign n33284 = n21221 ^ n14814 ^ n14676 ;
  assign n33285 = ( n5668 & n8737 ) | ( n5668 & ~n33284 ) | ( n8737 & ~n33284 ) ;
  assign n33286 = ( n5926 & n16468 ) | ( n5926 & n33285 ) | ( n16468 & n33285 ) ;
  assign n33287 = ~n12350 & n25515 ;
  assign n33288 = n32904 ^ n15301 ^ n15219 ;
  assign n33289 = ( n20717 & n29099 ) | ( n20717 & ~n33288 ) | ( n29099 & ~n33288 ) ;
  assign n33291 = n19036 ^ n10103 ^ n8678 ;
  assign n33290 = ( n17762 & ~n24299 ) | ( n17762 & n32667 ) | ( ~n24299 & n32667 ) ;
  assign n33292 = n33291 ^ n33290 ^ n16941 ;
  assign n33293 = ( ~n16086 & n33289 ) | ( ~n16086 & n33292 ) | ( n33289 & n33292 ) ;
  assign n33294 = n7034 ^ n1143 ^ n694 ;
  assign n33295 = ( n3576 & n7252 ) | ( n3576 & ~n10995 ) | ( n7252 & ~n10995 ) ;
  assign n33296 = ( n304 & ~n14323 ) | ( n304 & n33295 ) | ( ~n14323 & n33295 ) ;
  assign n33302 = n29877 ^ n19757 ^ n15852 ;
  assign n33303 = ( n7479 & ~n9278 ) | ( n7479 & n33302 ) | ( ~n9278 & n33302 ) ;
  assign n33299 = n2624 & ~n7375 ;
  assign n33300 = n33299 ^ n21551 ^ 1'b0 ;
  assign n33297 = n28297 ^ n10154 ^ n6156 ;
  assign n33298 = ( ~n17097 & n26921 ) | ( ~n17097 & n33297 ) | ( n26921 & n33297 ) ;
  assign n33301 = n33300 ^ n33298 ^ n7255 ;
  assign n33304 = n33303 ^ n33301 ^ n11805 ;
  assign n33305 = ( n16887 & n32350 ) | ( n16887 & n33304 ) | ( n32350 & n33304 ) ;
  assign n33306 = n30181 ^ n23221 ^ 1'b0 ;
  assign n33307 = ~n30015 & n33306 ;
  assign n33309 = n21486 ^ n16255 ^ n5095 ;
  assign n33308 = n2156 & n26960 ;
  assign n33310 = n33309 ^ n33308 ^ 1'b0 ;
  assign n33311 = n23399 ^ n22932 ^ n19511 ;
  assign n33312 = ( n28948 & n29698 ) | ( n28948 & n33311 ) | ( n29698 & n33311 ) ;
  assign n33313 = ( n472 & ~n8760 ) | ( n472 & n10148 ) | ( ~n8760 & n10148 ) ;
  assign n33314 = n33313 ^ n9750 ^ 1'b0 ;
  assign n33315 = n30275 ^ n20939 ^ x206 ;
  assign n33316 = n19946 ^ n17836 ^ n1426 ;
  assign n33317 = n18104 ^ n17839 ^ 1'b0 ;
  assign n33318 = ( n33315 & n33316 ) | ( n33315 & n33317 ) | ( n33316 & n33317 ) ;
  assign n33319 = ~n1433 & n3039 ;
  assign n33320 = n33319 ^ n26568 ^ 1'b0 ;
  assign n33321 = ( n2054 & ~n4492 ) | ( n2054 & n9415 ) | ( ~n4492 & n9415 ) ;
  assign n33322 = ( x56 & ~n17198 ) | ( x56 & n26796 ) | ( ~n17198 & n26796 ) ;
  assign n33323 = n32748 ^ n31127 ^ n1940 ;
  assign n33324 = n33323 ^ n20071 ^ n12319 ;
  assign n33325 = ( n33321 & ~n33322 ) | ( n33321 & n33324 ) | ( ~n33322 & n33324 ) ;
  assign n33326 = ( ~n10202 & n25468 ) | ( ~n10202 & n27237 ) | ( n25468 & n27237 ) ;
  assign n33327 = ~n29061 & n33326 ;
  assign n33328 = n14602 ^ n12068 ^ 1'b0 ;
  assign n33329 = ~n26588 & n33328 ;
  assign n33330 = ( n4060 & n18730 ) | ( n4060 & n33329 ) | ( n18730 & n33329 ) ;
  assign n33331 = n25365 ^ n13319 ^ n9753 ;
  assign n33335 = ( ~n828 & n13824 ) | ( ~n828 & n13890 ) | ( n13824 & n13890 ) ;
  assign n33332 = n24143 ^ n14462 ^ n12257 ;
  assign n33333 = n33332 ^ n17795 ^ 1'b0 ;
  assign n33334 = n32496 & n33333 ;
  assign n33336 = n33335 ^ n33334 ^ n7533 ;
  assign n33337 = n33336 ^ n19215 ^ n10020 ;
  assign n33338 = ( n33330 & n33331 ) | ( n33330 & ~n33337 ) | ( n33331 & ~n33337 ) ;
  assign n33339 = n25975 ^ n13055 ^ n6683 ;
  assign n33340 = ~n13302 & n33339 ;
  assign n33341 = ( n5013 & n14334 ) | ( n5013 & ~n24815 ) | ( n14334 & ~n24815 ) ;
  assign n33342 = n16690 ^ n11247 ^ n5557 ;
  assign n33343 = ( ~n24682 & n33341 ) | ( ~n24682 & n33342 ) | ( n33341 & n33342 ) ;
  assign n33344 = n33100 ^ n9295 ^ 1'b0 ;
  assign n33345 = n22391 & n33344 ;
  assign n33349 = ( ~n10491 & n16654 ) | ( ~n10491 & n19203 ) | ( n16654 & n19203 ) ;
  assign n33350 = n33349 ^ n8033 ^ n4969 ;
  assign n33346 = n10522 ^ n593 ^ x135 ;
  assign n33347 = n33346 ^ n6287 ^ n1835 ;
  assign n33348 = ( n9441 & n22248 ) | ( n9441 & ~n33347 ) | ( n22248 & ~n33347 ) ;
  assign n33351 = n33350 ^ n33348 ^ n10291 ;
  assign n33356 = ( n826 & n1111 ) | ( n826 & n7021 ) | ( n1111 & n7021 ) ;
  assign n33352 = ( n7349 & n7788 ) | ( n7349 & ~n26696 ) | ( n7788 & ~n26696 ) ;
  assign n33353 = ( ~n2833 & n18038 ) | ( ~n2833 & n33253 ) | ( n18038 & n33253 ) ;
  assign n33354 = ( n16789 & ~n24742 ) | ( n16789 & n33353 ) | ( ~n24742 & n33353 ) ;
  assign n33355 = ( n30435 & n33352 ) | ( n30435 & n33354 ) | ( n33352 & n33354 ) ;
  assign n33357 = n33356 ^ n33355 ^ n31599 ;
  assign n33358 = n10311 ^ n5267 ^ 1'b0 ;
  assign n33359 = ~n9270 & n33358 ;
  assign n33360 = n22805 & n33359 ;
  assign n33361 = n33360 ^ n16986 ^ n4772 ;
  assign n33363 = n1049 & n20913 ;
  assign n33362 = n10429 ^ n8843 ^ n4293 ;
  assign n33364 = n33363 ^ n33362 ^ n17302 ;
  assign n33365 = n33364 ^ n20364 ^ n1521 ;
  assign n33366 = ( ~n1590 & n33361 ) | ( ~n1590 & n33365 ) | ( n33361 & n33365 ) ;
  assign n33367 = n9570 ^ n2742 ^ 1'b0 ;
  assign n33368 = n33367 ^ n22885 ^ 1'b0 ;
  assign n33369 = ( n2217 & n33366 ) | ( n2217 & n33368 ) | ( n33366 & n33368 ) ;
  assign n33375 = ( n6585 & ~n22641 ) | ( n6585 & n27260 ) | ( ~n22641 & n27260 ) ;
  assign n33370 = n13612 & ~n21224 ;
  assign n33371 = ~n4362 & n33370 ;
  assign n33372 = n3846 | n33082 ;
  assign n33373 = n33371 & ~n33372 ;
  assign n33374 = n33373 ^ n20830 ^ n12057 ;
  assign n33376 = n33375 ^ n33374 ^ n25920 ;
  assign n33377 = ( ~n1937 & n5026 ) | ( ~n1937 & n27427 ) | ( n5026 & n27427 ) ;
  assign n33378 = n26967 ^ n8910 ^ n7381 ;
  assign n33379 = ~n3666 & n33378 ;
  assign n33380 = n33379 ^ n12875 ^ 1'b0 ;
  assign n33381 = ( n15817 & ~n26588 ) | ( n15817 & n33380 ) | ( ~n26588 & n33380 ) ;
  assign n33382 = n4830 ^ n2298 ^ 1'b0 ;
  assign n33383 = n18495 | n33382 ;
  assign n33388 = n4542 ^ n1774 ^ 1'b0 ;
  assign n33389 = n33388 ^ n28744 ^ n25203 ;
  assign n33384 = ( ~x164 & n1656 ) | ( ~x164 & n3186 ) | ( n1656 & n3186 ) ;
  assign n33385 = n33384 ^ n29379 ^ n28605 ;
  assign n33386 = n33385 ^ n26453 ^ n22937 ;
  assign n33387 = ( n12376 & n16934 ) | ( n12376 & ~n33386 ) | ( n16934 & ~n33386 ) ;
  assign n33390 = n33389 ^ n33387 ^ n14134 ;
  assign n33391 = ( n547 & n705 ) | ( n547 & n2822 ) | ( n705 & n2822 ) ;
  assign n33392 = ( ~n9606 & n19329 ) | ( ~n9606 & n33391 ) | ( n19329 & n33391 ) ;
  assign n33393 = n33392 ^ n18876 ^ n15134 ;
  assign n33394 = ( n13636 & n20733 ) | ( n13636 & n33393 ) | ( n20733 & n33393 ) ;
  assign n33395 = ( x77 & n14723 ) | ( x77 & ~n16675 ) | ( n14723 & ~n16675 ) ;
  assign n33396 = ( n6082 & ~n10916 ) | ( n6082 & n13192 ) | ( ~n10916 & n13192 ) ;
  assign n33397 = n2273 & ~n33396 ;
  assign n33398 = n33397 ^ n1931 ^ 1'b0 ;
  assign n33399 = ( n12827 & n22481 ) | ( n12827 & ~n33398 ) | ( n22481 & ~n33398 ) ;
  assign n33400 = ( n5090 & ~n33395 ) | ( n5090 & n33399 ) | ( ~n33395 & n33399 ) ;
  assign n33401 = ( n7077 & ~n19438 ) | ( n7077 & n33400 ) | ( ~n19438 & n33400 ) ;
  assign n33402 = ( n8716 & ~n14555 ) | ( n8716 & n29568 ) | ( ~n14555 & n29568 ) ;
  assign n33403 = ( n15672 & n22051 ) | ( n15672 & n33402 ) | ( n22051 & n33402 ) ;
  assign n33404 = n33403 ^ n26409 ^ n8432 ;
  assign n33405 = n26139 & ~n33404 ;
  assign n33406 = n33405 ^ n1983 ^ 1'b0 ;
  assign n33407 = n8773 ^ n8288 ^ n6537 ;
  assign n33408 = ( n765 & n13233 ) | ( n765 & n15184 ) | ( n13233 & n15184 ) ;
  assign n33409 = n33408 ^ n21780 ^ n3415 ;
  assign n33410 = n25549 ^ n5718 ^ n862 ;
  assign n33411 = n33410 ^ n16072 ^ n2625 ;
  assign n33412 = ( n14826 & n33409 ) | ( n14826 & ~n33411 ) | ( n33409 & ~n33411 ) ;
  assign n33413 = n14952 ^ n367 ^ 1'b0 ;
  assign n33414 = n9334 & n33413 ;
  assign n33415 = ( n4954 & n10192 ) | ( n4954 & n33414 ) | ( n10192 & n33414 ) ;
  assign n33416 = n25086 ^ n4343 ^ 1'b0 ;
  assign n33417 = n20665 | n33416 ;
  assign n33418 = ( ~n23864 & n25225 ) | ( ~n23864 & n26522 ) | ( n25225 & n26522 ) ;
  assign n33419 = ( n4907 & n10970 ) | ( n4907 & ~n18273 ) | ( n10970 & ~n18273 ) ;
  assign n33420 = n29772 ^ n12893 ^ 1'b0 ;
  assign n33421 = n7974 & ~n33420 ;
  assign n33422 = n17567 ^ n2858 ^ n756 ;
  assign n33423 = ~n1579 & n16302 ;
  assign n33424 = ~n13182 & n33423 ;
  assign n33425 = ( n21047 & ~n33422 ) | ( n21047 & n33424 ) | ( ~n33422 & n33424 ) ;
  assign n33426 = ( ~n15082 & n17442 ) | ( ~n15082 & n33022 ) | ( n17442 & n33022 ) ;
  assign n33427 = n31660 ^ n12564 ^ n6540 ;
  assign n33428 = n6614 & n9336 ;
  assign n33429 = n654 & n33428 ;
  assign n33430 = n33429 ^ n19160 ^ n10801 ;
  assign n33431 = n33430 ^ n20844 ^ n6029 ;
  assign n33433 = n26115 ^ n17802 ^ n3150 ;
  assign n33434 = n33433 ^ n10257 ^ n7464 ;
  assign n33432 = n16076 & ~n31153 ;
  assign n33435 = n33434 ^ n33432 ^ 1'b0 ;
  assign n33436 = ( n4977 & n13899 ) | ( n4977 & ~n16997 ) | ( n13899 & ~n16997 ) ;
  assign n33437 = ~n2035 & n6335 ;
  assign n33438 = n33437 ^ n19086 ^ n4809 ;
  assign n33439 = n33438 ^ n23065 ^ 1'b0 ;
  assign n33440 = n11248 & ~n33439 ;
  assign n33441 = n2240 & n33440 ;
  assign n33442 = n33436 & n33441 ;
  assign n33443 = ( ~n263 & n8143 ) | ( ~n263 & n27983 ) | ( n8143 & n27983 ) ;
  assign n33444 = ( n13218 & n15752 ) | ( n13218 & n16500 ) | ( n15752 & n16500 ) ;
  assign n33445 = ( ~n6716 & n33443 ) | ( ~n6716 & n33444 ) | ( n33443 & n33444 ) ;
  assign n33446 = n6366 ^ n3264 ^ n2049 ;
  assign n33447 = ( ~n21938 & n31514 ) | ( ~n21938 & n33446 ) | ( n31514 & n33446 ) ;
  assign n33448 = n14819 | n30158 ;
  assign n33449 = n10763 & ~n33448 ;
  assign n33450 = ( n6124 & n29316 ) | ( n6124 & n33449 ) | ( n29316 & n33449 ) ;
  assign n33451 = ( ~n11104 & n28732 ) | ( ~n11104 & n32834 ) | ( n28732 & n32834 ) ;
  assign n33452 = n33451 ^ n33449 ^ 1'b0 ;
  assign n33453 = ( n21038 & ~n30281 ) | ( n21038 & n33452 ) | ( ~n30281 & n33452 ) ;
  assign n33454 = n11382 | n16334 ;
  assign n33455 = ( n12065 & ~n20346 ) | ( n12065 & n20674 ) | ( ~n20346 & n20674 ) ;
  assign n33456 = n26818 ^ x72 ^ 1'b0 ;
  assign n33461 = ( ~n14978 & n18223 ) | ( ~n14978 & n21082 ) | ( n18223 & n21082 ) ;
  assign n33459 = n24888 ^ n23914 ^ n14274 ;
  assign n33457 = n1828 & ~n9113 ;
  assign n33458 = n14861 & n33457 ;
  assign n33460 = n33459 ^ n33458 ^ n14566 ;
  assign n33462 = n33461 ^ n33460 ^ 1'b0 ;
  assign n33463 = ( n1124 & n2183 ) | ( n1124 & n14739 ) | ( n2183 & n14739 ) ;
  assign n33464 = ( n13711 & ~n29378 ) | ( n13711 & n33463 ) | ( ~n29378 & n33463 ) ;
  assign n33465 = n25182 ^ n17356 ^ n516 ;
  assign n33466 = n17028 ^ n16773 ^ n8079 ;
  assign n33467 = ( n14134 & n18493 ) | ( n14134 & ~n33466 ) | ( n18493 & ~n33466 ) ;
  assign n33468 = n18292 & ~n32766 ;
  assign n33469 = n33468 ^ n21559 ^ 1'b0 ;
  assign n33470 = ( n1236 & n6675 ) | ( n1236 & n9101 ) | ( n6675 & n9101 ) ;
  assign n33471 = n33470 ^ n30963 ^ 1'b0 ;
  assign n33472 = n19671 ^ n15506 ^ 1'b0 ;
  assign n33474 = n28373 ^ n25971 ^ n2484 ;
  assign n33473 = ( n6836 & n7238 ) | ( n6836 & ~n19935 ) | ( n7238 & ~n19935 ) ;
  assign n33475 = n33474 ^ n33473 ^ 1'b0 ;
  assign n33476 = n29217 ^ n17881 ^ n15566 ;
  assign n33479 = ( n13899 & ~n14647 ) | ( n13899 & n17476 ) | ( ~n14647 & n17476 ) ;
  assign n33477 = ( n16315 & ~n25408 ) | ( n16315 & n28283 ) | ( ~n25408 & n28283 ) ;
  assign n33478 = ( n7103 & n32397 ) | ( n7103 & n33477 ) | ( n32397 & n33477 ) ;
  assign n33480 = n33479 ^ n33478 ^ n19625 ;
  assign n33481 = n29114 ^ n12548 ^ 1'b0 ;
  assign n33482 = n33480 & n33481 ;
  assign n33486 = n8950 & n12728 ;
  assign n33487 = ( n18531 & ~n25283 ) | ( n18531 & n33486 ) | ( ~n25283 & n33486 ) ;
  assign n33484 = n15144 ^ n2267 ^ n850 ;
  assign n33483 = n33139 ^ n8577 ^ n6034 ;
  assign n33485 = n33484 ^ n33483 ^ n31141 ;
  assign n33488 = n33487 ^ n33485 ^ n4947 ;
  assign n33489 = ( n9986 & n13843 ) | ( n9986 & ~n22160 ) | ( n13843 & ~n22160 ) ;
  assign n33490 = n28864 ^ n6991 ^ n5402 ;
  assign n33491 = n15659 ^ x232 ^ 1'b0 ;
  assign n33492 = n33490 | n33491 ;
  assign n33493 = ( n11590 & ~n15150 ) | ( n11590 & n33492 ) | ( ~n15150 & n33492 ) ;
  assign n33494 = ( ~n13430 & n17044 ) | ( ~n13430 & n19681 ) | ( n17044 & n19681 ) ;
  assign n33495 = ( n11363 & ~n15211 ) | ( n11363 & n33494 ) | ( ~n15211 & n33494 ) ;
  assign n33496 = n33495 ^ n17304 ^ 1'b0 ;
  assign n33502 = ( n2515 & n10282 ) | ( n2515 & n29403 ) | ( n10282 & n29403 ) ;
  assign n33500 = n16879 ^ n8799 ^ n6976 ;
  assign n33501 = ( ~n5887 & n10986 ) | ( ~n5887 & n33500 ) | ( n10986 & n33500 ) ;
  assign n33503 = n33502 ^ n33501 ^ n11984 ;
  assign n33504 = ( n4620 & n14564 ) | ( n4620 & n33503 ) | ( n14564 & n33503 ) ;
  assign n33497 = ( n1393 & n2330 ) | ( n1393 & ~n3962 ) | ( n2330 & ~n3962 ) ;
  assign n33498 = n33497 ^ n13902 ^ n12919 ;
  assign n33499 = ( ~n419 & n12708 ) | ( ~n419 & n33498 ) | ( n12708 & n33498 ) ;
  assign n33505 = n33504 ^ n33499 ^ n21715 ;
  assign n33507 = ( n2697 & n16448 ) | ( n2697 & ~n19861 ) | ( n16448 & ~n19861 ) ;
  assign n33508 = n33507 ^ n14371 ^ n10906 ;
  assign n33506 = ( n3100 & ~n12029 ) | ( n3100 & n24921 ) | ( ~n12029 & n24921 ) ;
  assign n33509 = n33508 ^ n33506 ^ n2646 ;
  assign n33510 = ( n6444 & n17417 ) | ( n6444 & n28676 ) | ( n17417 & n28676 ) ;
  assign n33511 = ( n584 & ~n9447 ) | ( n584 & n26279 ) | ( ~n9447 & n26279 ) ;
  assign n33512 = ( x159 & ~n27921 ) | ( x159 & n33511 ) | ( ~n27921 & n33511 ) ;
  assign n33513 = ( n26674 & n27522 ) | ( n26674 & ~n33512 ) | ( n27522 & ~n33512 ) ;
  assign n33514 = n30421 ^ n25162 ^ n984 ;
  assign n33515 = ( n4415 & n19722 ) | ( n4415 & ~n33514 ) | ( n19722 & ~n33514 ) ;
  assign n33516 = n16861 ^ n15280 ^ n11450 ;
  assign n33517 = n13785 ^ n8400 ^ n2486 ;
  assign n33520 = ( ~n1164 & n9056 ) | ( ~n1164 & n27959 ) | ( n9056 & n27959 ) ;
  assign n33521 = ( ~n8349 & n11106 ) | ( ~n8349 & n33520 ) | ( n11106 & n33520 ) ;
  assign n33518 = n26424 ^ n7267 ^ n2097 ;
  assign n33519 = ( n6481 & n13841 ) | ( n6481 & n33518 ) | ( n13841 & n33518 ) ;
  assign n33522 = n33521 ^ n33519 ^ n11619 ;
  assign n33523 = n33522 ^ n6069 ^ n5219 ;
  assign n33524 = ( n33020 & n33517 ) | ( n33020 & ~n33523 ) | ( n33517 & ~n33523 ) ;
  assign n33525 = ( n5004 & ~n33516 ) | ( n5004 & n33524 ) | ( ~n33516 & n33524 ) ;
  assign n33526 = n21297 ^ n13807 ^ n8222 ;
  assign n33527 = n33526 ^ n29338 ^ n1164 ;
  assign n33528 = n33527 ^ n5665 ^ 1'b0 ;
  assign n33529 = n15016 ^ n1650 ^ 1'b0 ;
  assign n33533 = ( n21762 & n22372 ) | ( n21762 & n22713 ) | ( n22372 & n22713 ) ;
  assign n33530 = n9241 ^ n2353 ^ n1823 ;
  assign n33531 = n33530 ^ n22980 ^ n19377 ;
  assign n33532 = n33531 ^ n17705 ^ n12852 ;
  assign n33534 = n33533 ^ n33532 ^ n17780 ;
  assign n33535 = n26731 ^ n20986 ^ n18536 ;
  assign n33549 = ( n7188 & ~n16761 ) | ( n7188 & n26172 ) | ( ~n16761 & n26172 ) ;
  assign n33541 = ( n4230 & ~n13227 ) | ( n4230 & n25110 ) | ( ~n13227 & n25110 ) ;
  assign n33542 = ( ~n23968 & n30547 ) | ( ~n23968 & n33541 ) | ( n30547 & n33541 ) ;
  assign n33543 = n33542 ^ n25486 ^ 1'b0 ;
  assign n33544 = n13935 & n21134 ;
  assign n33545 = ~n3142 & n33544 ;
  assign n33546 = ( n27125 & n27807 ) | ( n27125 & n33545 ) | ( n27807 & n33545 ) ;
  assign n33547 = n33546 ^ n8333 ^ x142 ;
  assign n33548 = ( n22718 & ~n33543 ) | ( n22718 & n33547 ) | ( ~n33543 & n33547 ) ;
  assign n33536 = ( ~x144 & n1299 ) | ( ~x144 & n4060 ) | ( n1299 & n4060 ) ;
  assign n33537 = n22196 ^ n14672 ^ n1408 ;
  assign n33538 = ( n1370 & ~n33536 ) | ( n1370 & n33537 ) | ( ~n33536 & n33537 ) ;
  assign n33539 = n12803 ^ n8597 ^ n8270 ;
  assign n33540 = ( n15617 & ~n33538 ) | ( n15617 & n33539 ) | ( ~n33538 & n33539 ) ;
  assign n33550 = n33549 ^ n33548 ^ n33540 ;
  assign n33551 = ( ~n296 & n33535 ) | ( ~n296 & n33550 ) | ( n33535 & n33550 ) ;
  assign n33552 = n29806 ^ n26917 ^ n1526 ;
  assign n33553 = ( n1705 & ~n24018 ) | ( n1705 & n33552 ) | ( ~n24018 & n33552 ) ;
  assign n33554 = ( n7537 & n9108 ) | ( n7537 & ~n20254 ) | ( n9108 & ~n20254 ) ;
  assign n33555 = ( n462 & n10348 ) | ( n462 & n33554 ) | ( n10348 & n33554 ) ;
  assign n33556 = n33555 ^ n31844 ^ n25651 ;
  assign n33559 = n12395 ^ n8996 ^ n3385 ;
  assign n33560 = ( ~n2263 & n6312 ) | ( ~n2263 & n23494 ) | ( n6312 & n23494 ) ;
  assign n33561 = ( ~n5138 & n33559 ) | ( ~n5138 & n33560 ) | ( n33559 & n33560 ) ;
  assign n33557 = n10359 ^ n6761 ^ n4111 ;
  assign n33558 = n33557 ^ n22347 ^ n18674 ;
  assign n33562 = n33561 ^ n33558 ^ 1'b0 ;
  assign n33563 = ( n5192 & ~n19600 ) | ( n5192 & n21725 ) | ( ~n19600 & n21725 ) ;
  assign n33564 = n33563 ^ n18744 ^ n14753 ;
  assign n33565 = ( n6272 & n17328 ) | ( n6272 & n33564 ) | ( n17328 & n33564 ) ;
  assign n33567 = ( n3153 & n3792 ) | ( n3153 & n9686 ) | ( n3792 & n9686 ) ;
  assign n33568 = n33567 ^ n12787 ^ n5877 ;
  assign n33566 = n13424 ^ n6522 ^ 1'b0 ;
  assign n33569 = n33568 ^ n33566 ^ n9522 ;
  assign n33570 = ( n7089 & ~n21159 ) | ( n7089 & n30624 ) | ( ~n21159 & n30624 ) ;
  assign n33571 = n22947 ^ n16481 ^ 1'b0 ;
  assign n33572 = n33570 & n33571 ;
  assign n33573 = ( n1115 & ~n2597 ) | ( n1115 & n21073 ) | ( ~n2597 & n21073 ) ;
  assign n33574 = n32487 ^ n31424 ^ n10008 ;
  assign n33575 = ( n9440 & n33573 ) | ( n9440 & n33574 ) | ( n33573 & n33574 ) ;
  assign n33576 = n25791 ^ n11719 ^ n5946 ;
  assign n33577 = n7387 & n25224 ;
  assign n33578 = ~n1779 & n33577 ;
  assign n33579 = n292 & ~n33578 ;
  assign n33580 = n33579 ^ n21680 ^ 1'b0 ;
  assign n33581 = ( n1555 & ~n2833 ) | ( n1555 & n33580 ) | ( ~n2833 & n33580 ) ;
  assign n33582 = n30747 ^ n25603 ^ n5000 ;
  assign n33583 = n2055 | n33582 ;
  assign n33584 = n23454 ^ n20771 ^ n8672 ;
  assign n33585 = ( n6451 & ~n33583 ) | ( n6451 & n33584 ) | ( ~n33583 & n33584 ) ;
  assign n33586 = ( n7541 & n14015 ) | ( n7541 & ~n29407 ) | ( n14015 & ~n29407 ) ;
  assign n33587 = n31976 ^ n21404 ^ n7303 ;
  assign n33588 = ~n7128 & n33587 ;
  assign n33589 = n33588 ^ n9554 ^ 1'b0 ;
  assign n33590 = ( n1358 & ~n5647 ) | ( n1358 & n12094 ) | ( ~n5647 & n12094 ) ;
  assign n33591 = n8793 ^ n3401 ^ n2783 ;
  assign n33592 = n20343 ^ n18012 ^ n13040 ;
  assign n33593 = ( n12907 & n22024 ) | ( n12907 & n22870 ) | ( n22024 & n22870 ) ;
  assign n33594 = ( ~n5599 & n33592 ) | ( ~n5599 & n33593 ) | ( n33592 & n33593 ) ;
  assign n33595 = ( n33590 & ~n33591 ) | ( n33590 & n33594 ) | ( ~n33591 & n33594 ) ;
  assign n33596 = n9098 & ~n10450 ;
  assign n33597 = ~n33595 & n33596 ;
  assign n33598 = n33045 ^ n18738 ^ n14363 ;
  assign n33599 = ( n11943 & ~n21276 ) | ( n11943 & n33598 ) | ( ~n21276 & n33598 ) ;
  assign n33602 = n1539 & n12911 ;
  assign n33600 = ( x173 & n1485 ) | ( x173 & ~n26068 ) | ( n1485 & ~n26068 ) ;
  assign n33601 = n33600 ^ n13409 ^ n9544 ;
  assign n33603 = n33602 ^ n33601 ^ n2353 ;
  assign n33604 = n11640 ^ n7817 ^ n7511 ;
  assign n33605 = ( n11015 & ~n21301 ) | ( n11015 & n33604 ) | ( ~n21301 & n33604 ) ;
  assign n33606 = ( n10776 & n12804 ) | ( n10776 & ~n33605 ) | ( n12804 & ~n33605 ) ;
  assign n33607 = n29529 ^ n26319 ^ n25816 ;
  assign n33608 = n7516 ^ n3371 ^ x173 ;
  assign n33609 = ( n14001 & n16047 ) | ( n14001 & ~n33608 ) | ( n16047 & ~n33608 ) ;
  assign n33610 = n12843 & n14589 ;
  assign n33611 = n33609 & n33610 ;
  assign n33612 = ( x2 & n3728 ) | ( x2 & n4191 ) | ( n3728 & n4191 ) ;
  assign n33613 = ~n6270 & n33612 ;
  assign n33614 = n1781 & n33613 ;
  assign n33615 = n28103 ^ n24169 ^ 1'b0 ;
  assign n33616 = n33614 | n33615 ;
  assign n33617 = n29617 ^ n28514 ^ n13201 ;
  assign n33618 = ( n8065 & n33616 ) | ( n8065 & n33617 ) | ( n33616 & n33617 ) ;
  assign n33619 = ( n2591 & ~n5192 ) | ( n2591 & n21501 ) | ( ~n5192 & n21501 ) ;
  assign n33620 = ( n1118 & n25344 ) | ( n1118 & ~n33619 ) | ( n25344 & ~n33619 ) ;
  assign n33622 = n13263 ^ n5375 ^ n5368 ;
  assign n33623 = ( n387 & ~n17526 ) | ( n387 & n33622 ) | ( ~n17526 & n33622 ) ;
  assign n33624 = ( n1385 & n1427 ) | ( n1385 & ~n33623 ) | ( n1427 & ~n33623 ) ;
  assign n33621 = ( n6897 & ~n25176 ) | ( n6897 & n29451 ) | ( ~n25176 & n29451 ) ;
  assign n33625 = n33624 ^ n33621 ^ n25965 ;
  assign n33626 = n22024 ^ n13797 ^ n1868 ;
  assign n33627 = n33626 ^ n29715 ^ n11308 ;
  assign n33628 = ( n10816 & n29843 ) | ( n10816 & n30075 ) | ( n29843 & n30075 ) ;
  assign n33629 = n22545 ^ n4842 ^ 1'b0 ;
  assign n33630 = n33628 | n33629 ;
  assign n33631 = n29357 ^ n17963 ^ n10405 ;
  assign n33632 = n13972 ^ n11380 ^ 1'b0 ;
  assign n33633 = n2783 & n33632 ;
  assign n33634 = ~n27772 & n33633 ;
  assign n33635 = n33631 & n33634 ;
  assign n33636 = n7370 & ~n33635 ;
  assign n33637 = n25811 ^ n12536 ^ n3929 ;
  assign n33638 = n27865 ^ n26160 ^ n8752 ;
  assign n33639 = ( n12998 & ~n14669 ) | ( n12998 & n26168 ) | ( ~n14669 & n26168 ) ;
  assign n33641 = n8511 | n20488 ;
  assign n33640 = n30022 ^ n27046 ^ n23188 ;
  assign n33642 = n33641 ^ n33640 ^ n5074 ;
  assign n33643 = n16447 ^ n13996 ^ n8261 ;
  assign n33644 = n33643 ^ n13221 ^ n7579 ;
  assign n33645 = ( n1362 & n33316 ) | ( n1362 & n33644 ) | ( n33316 & n33644 ) ;
  assign n33646 = n33645 ^ n8522 ^ n6289 ;
  assign n33648 = n21932 ^ n5554 ^ n4316 ;
  assign n33647 = ( n15205 & n15730 ) | ( n15205 & ~n22084 ) | ( n15730 & ~n22084 ) ;
  assign n33649 = n33648 ^ n33647 ^ n7192 ;
  assign n33650 = ( n1233 & n30349 ) | ( n1233 & ~n33649 ) | ( n30349 & ~n33649 ) ;
  assign n33651 = ( n1062 & n2418 ) | ( n1062 & n22400 ) | ( n2418 & n22400 ) ;
  assign n33652 = n33651 ^ n24378 ^ n3074 ;
  assign n33653 = ( n8160 & ~n15852 ) | ( n8160 & n26618 ) | ( ~n15852 & n26618 ) ;
  assign n33654 = ( n2705 & n12489 ) | ( n2705 & ~n33653 ) | ( n12489 & ~n33653 ) ;
  assign n33655 = n33654 ^ n21883 ^ n9080 ;
  assign n33656 = ( ~n13337 & n25937 ) | ( ~n13337 & n33655 ) | ( n25937 & n33655 ) ;
  assign n33657 = ( n8274 & ~n10948 ) | ( n8274 & n11110 ) | ( ~n10948 & n11110 ) ;
  assign n33658 = ( n26097 & ~n33446 ) | ( n26097 & n33657 ) | ( ~n33446 & n33657 ) ;
  assign n33659 = n18119 ^ n14386 ^ 1'b0 ;
  assign n33660 = ~n33658 & n33659 ;
  assign n33661 = n15917 & ~n22100 ;
  assign n33662 = ~n4449 & n33661 ;
  assign n33668 = n27846 ^ n18945 ^ n1115 ;
  assign n33663 = ( n7195 & ~n9836 ) | ( n7195 & n28106 ) | ( ~n9836 & n28106 ) ;
  assign n33664 = ~n17791 & n28036 ;
  assign n33665 = ( x113 & ~n10279 ) | ( x113 & n33664 ) | ( ~n10279 & n33664 ) ;
  assign n33666 = ~n33663 & n33665 ;
  assign n33667 = n33666 ^ n21335 ^ 1'b0 ;
  assign n33669 = n33668 ^ n33667 ^ n14537 ;
  assign n33670 = ( n18360 & n30167 ) | ( n18360 & ~n30592 ) | ( n30167 & ~n30592 ) ;
  assign n33675 = n20783 ^ n2748 ^ n1965 ;
  assign n33676 = ( n14813 & ~n24565 ) | ( n14813 & n33675 ) | ( ~n24565 & n33675 ) ;
  assign n33673 = n9418 | n33403 ;
  assign n33674 = n33673 ^ n416 ^ 1'b0 ;
  assign n33671 = n27351 ^ n6588 ^ n3636 ;
  assign n33672 = ( n11688 & n13923 ) | ( n11688 & n33671 ) | ( n13923 & n33671 ) ;
  assign n33677 = n33676 ^ n33674 ^ n33672 ;
  assign n33679 = ( n5274 & n20938 ) | ( n5274 & n23231 ) | ( n20938 & n23231 ) ;
  assign n33678 = n25180 ^ n8843 ^ 1'b0 ;
  assign n33680 = n33679 ^ n33678 ^ n28768 ;
  assign n33681 = ( n8922 & ~n17313 ) | ( n8922 & n33361 ) | ( ~n17313 & n33361 ) ;
  assign n33682 = ( n4738 & ~n8843 ) | ( n4738 & n16643 ) | ( ~n8843 & n16643 ) ;
  assign n33683 = ( x160 & n4305 ) | ( x160 & n33682 ) | ( n4305 & n33682 ) ;
  assign n33684 = n18824 ^ n12440 ^ n1727 ;
  assign n33685 = ( n19721 & n19838 ) | ( n19721 & n25251 ) | ( n19838 & n25251 ) ;
  assign n33686 = n33685 ^ n12383 ^ 1'b0 ;
  assign n33687 = n33686 ^ n3189 ^ n2521 ;
  assign n33688 = ( n5091 & n9253 ) | ( n5091 & ~n20892 ) | ( n9253 & ~n20892 ) ;
  assign n33689 = ( n7828 & ~n16784 ) | ( n7828 & n30129 ) | ( ~n16784 & n30129 ) ;
  assign n33690 = n5968 & ~n11068 ;
  assign n33691 = n33690 ^ n9572 ^ 1'b0 ;
  assign n33692 = n33691 ^ n16511 ^ n12479 ;
  assign n33693 = n33692 ^ n9202 ^ 1'b0 ;
  assign n33694 = ~n33689 & n33693 ;
  assign n33695 = ( n15133 & n33688 ) | ( n15133 & ~n33694 ) | ( n33688 & ~n33694 ) ;
  assign n33696 = n33695 ^ n22574 ^ n14588 ;
  assign n33697 = n10345 & ~n26430 ;
  assign n33698 = n8231 & n33697 ;
  assign n33699 = n33698 ^ n29825 ^ n3871 ;
  assign n33700 = n33699 ^ n24192 ^ n2724 ;
  assign n33701 = n33700 ^ n27843 ^ n4780 ;
  assign n33702 = n9770 | n10660 ;
  assign n33703 = ~n25005 & n25669 ;
  assign n33704 = ~n2673 & n33703 ;
  assign n33705 = ( ~n5110 & n33702 ) | ( ~n5110 & n33704 ) | ( n33702 & n33704 ) ;
  assign n33706 = ( n24783 & n25245 ) | ( n24783 & n27691 ) | ( n25245 & n27691 ) ;
  assign n33707 = n33706 ^ n7188 ^ n6907 ;
  assign n33708 = n33538 ^ n3112 ^ 1'b0 ;
  assign n33709 = n19111 ^ n3219 ^ 1'b0 ;
  assign n33710 = ~n14752 & n33709 ;
  assign n33711 = n33710 ^ n22661 ^ n11631 ;
  assign n33712 = ( n9921 & n11453 ) | ( n9921 & n33711 ) | ( n11453 & n33711 ) ;
  assign n33713 = n33712 ^ n15640 ^ 1'b0 ;
  assign n33714 = ( n33707 & n33708 ) | ( n33707 & n33713 ) | ( n33708 & n33713 ) ;
  assign n33715 = n29516 ^ n16235 ^ n1240 ;
  assign n33719 = n17211 & n17479 ;
  assign n33720 = n33719 ^ n8514 ^ 1'b0 ;
  assign n33721 = n33720 ^ n15951 ^ n971 ;
  assign n33716 = n23617 ^ n22600 ^ 1'b0 ;
  assign n33717 = n15614 & ~n33716 ;
  assign n33718 = ( n5944 & n22740 ) | ( n5944 & n33717 ) | ( n22740 & n33717 ) ;
  assign n33722 = n33721 ^ n33718 ^ n27269 ;
  assign n33723 = ( n8129 & n11134 ) | ( n8129 & ~n28505 ) | ( n11134 & ~n28505 ) ;
  assign n33728 = n23214 ^ n2513 ^ n1064 ;
  assign n33725 = n7840 & ~n11254 ;
  assign n33726 = n33725 ^ n23696 ^ 1'b0 ;
  assign n33724 = ~n2692 & n27490 ;
  assign n33727 = n33726 ^ n33724 ^ n15516 ;
  assign n33729 = n33728 ^ n33727 ^ n17043 ;
  assign n33730 = n7862 ^ n6637 ^ n5616 ;
  assign n33731 = n26068 ^ n3773 ^ n2038 ;
  assign n33732 = n33731 ^ n21407 ^ n9918 ;
  assign n33733 = ( ~n12498 & n33730 ) | ( ~n12498 & n33732 ) | ( n33730 & n33732 ) ;
  assign n33734 = n27999 ^ n8756 ^ n1747 ;
  assign n33735 = ( ~n11148 & n19144 ) | ( ~n11148 & n33734 ) | ( n19144 & n33734 ) ;
  assign n33736 = n12392 ^ n2166 ^ 1'b0 ;
  assign n33737 = n10875 & n33736 ;
  assign n33738 = n20492 ^ n16072 ^ n2933 ;
  assign n33739 = n33738 ^ n4077 ^ 1'b0 ;
  assign n33740 = n4722 & ~n33739 ;
  assign n33741 = n23559 ^ n19188 ^ n14941 ;
  assign n33742 = ( n14708 & n16090 ) | ( n14708 & n33741 ) | ( n16090 & n33741 ) ;
  assign n33743 = n33742 ^ n24489 ^ n18586 ;
  assign n33744 = ( n2657 & ~n18546 ) | ( n2657 & n33743 ) | ( ~n18546 & n33743 ) ;
  assign n33745 = ( ~n6066 & n13419 ) | ( ~n6066 & n20744 ) | ( n13419 & n20744 ) ;
  assign n33746 = ( n11289 & n11620 ) | ( n11289 & ~n33745 ) | ( n11620 & ~n33745 ) ;
  assign n33747 = n31607 ^ n2127 ^ 1'b0 ;
  assign n33748 = n1254 & n6654 ;
  assign n33749 = ( n23191 & n30581 ) | ( n23191 & n31310 ) | ( n30581 & n31310 ) ;
  assign n33750 = n12324 ^ n10707 ^ n664 ;
  assign n33751 = ( n7667 & n25358 ) | ( n7667 & ~n33750 ) | ( n25358 & ~n33750 ) ;
  assign n33752 = n21232 & ~n29925 ;
  assign n33753 = n18595 ^ n8414 ^ n6368 ;
  assign n33754 = ( n13702 & ~n33752 ) | ( n13702 & n33753 ) | ( ~n33752 & n33753 ) ;
  assign n33755 = ( n457 & n7320 ) | ( n457 & ~n17248 ) | ( n7320 & ~n17248 ) ;
  assign n33756 = ( n2218 & ~n18562 ) | ( n2218 & n33755 ) | ( ~n18562 & n33755 ) ;
  assign n33757 = n19756 ^ n2835 ^ n693 ;
  assign n33758 = ( n19284 & ~n23974 ) | ( n19284 & n33757 ) | ( ~n23974 & n33757 ) ;
  assign n33759 = n26926 ^ n22238 ^ 1'b0 ;
  assign n33760 = n14824 & n22029 ;
  assign n33761 = ( n21828 & ~n33759 ) | ( n21828 & n33760 ) | ( ~n33759 & n33760 ) ;
  assign n33762 = n14966 & ~n33761 ;
  assign n33763 = n6389 & ~n24487 ;
  assign n33764 = ( n6803 & n12667 ) | ( n6803 & n12927 ) | ( n12667 & n12927 ) ;
  assign n33765 = n20167 ^ n10629 ^ n6884 ;
  assign n33766 = n33765 ^ n21397 ^ 1'b0 ;
  assign n33767 = n33764 & n33766 ;
  assign n33769 = ( n6695 & n9097 ) | ( n6695 & ~n24661 ) | ( n9097 & ~n24661 ) ;
  assign n33770 = ( ~n9437 & n12673 ) | ( ~n9437 & n33769 ) | ( n12673 & n33769 ) ;
  assign n33768 = n9200 & ~n33317 ;
  assign n33771 = n33770 ^ n33768 ^ 1'b0 ;
  assign n33772 = n3386 | n12586 ;
  assign n33773 = n24349 & ~n33772 ;
  assign n33774 = ( ~n4212 & n22538 ) | ( ~n4212 & n33773 ) | ( n22538 & n33773 ) ;
  assign n33775 = n33774 ^ n22330 ^ 1'b0 ;
  assign n33776 = n33771 & n33775 ;
  assign n33777 = n14183 ^ n8172 ^ n1606 ;
  assign n33778 = n3523 & n33777 ;
  assign n33779 = ( ~n4455 & n10706 ) | ( ~n4455 & n29176 ) | ( n10706 & n29176 ) ;
  assign n33783 = n23093 ^ n6741 ^ 1'b0 ;
  assign n33781 = ( n359 & n17697 ) | ( n359 & n22888 ) | ( n17697 & n22888 ) ;
  assign n33780 = ( n1900 & n2146 ) | ( n1900 & ~n13219 ) | ( n2146 & ~n13219 ) ;
  assign n33782 = n33781 ^ n33780 ^ n14740 ;
  assign n33784 = n33783 ^ n33782 ^ n30702 ;
  assign n33785 = n10633 ^ n2154 ^ n1509 ;
  assign n33786 = n33785 ^ n24460 ^ 1'b0 ;
  assign n33787 = n33786 ^ n26744 ^ n5336 ;
  assign n33788 = n3892 ^ n1730 ^ 1'b0 ;
  assign n33789 = ( n5727 & n25779 ) | ( n5727 & ~n28356 ) | ( n25779 & ~n28356 ) ;
  assign n33790 = ( n13799 & n29552 ) | ( n13799 & ~n33774 ) | ( n29552 & ~n33774 ) ;
  assign n33791 = n33790 ^ n28238 ^ n18963 ;
  assign n33792 = ( n1484 & n11637 ) | ( n1484 & ~n22548 ) | ( n11637 & ~n22548 ) ;
  assign n33793 = n33792 ^ n28814 ^ n15353 ;
  assign n33794 = n33793 ^ n30715 ^ n20848 ;
  assign n33795 = n26025 ^ n17840 ^ n17097 ;
  assign n33796 = n33795 ^ n19512 ^ 1'b0 ;
  assign n33797 = n15969 & ~n33796 ;
  assign n33798 = ~n3275 & n3885 ;
  assign n33799 = n33798 ^ n20556 ^ 1'b0 ;
  assign n33800 = ( n1497 & n5794 ) | ( n1497 & n29516 ) | ( n5794 & n29516 ) ;
  assign n33801 = n33800 ^ n13845 ^ n10395 ;
  assign n33803 = n16808 ^ n14451 ^ n941 ;
  assign n33802 = ( ~n4403 & n8736 ) | ( ~n4403 & n15574 ) | ( n8736 & n15574 ) ;
  assign n33804 = n33803 ^ n33802 ^ n17311 ;
  assign n33805 = n9005 | n19875 ;
  assign n33806 = ( ~n3449 & n27426 ) | ( ~n3449 & n33805 ) | ( n27426 & n33805 ) ;
  assign n33807 = n33806 ^ n8878 ^ x195 ;
  assign n33808 = ( n11945 & n14895 ) | ( n11945 & ~n33188 ) | ( n14895 & ~n33188 ) ;
  assign n33809 = ( n7057 & n8939 ) | ( n7057 & n14633 ) | ( n8939 & n14633 ) ;
  assign n33810 = n27251 ^ n10741 ^ n5782 ;
  assign n33811 = ( ~n29773 & n33809 ) | ( ~n29773 & n33810 ) | ( n33809 & n33810 ) ;
  assign n33812 = n14093 & ~n33811 ;
  assign n33813 = n33812 ^ n28250 ^ 1'b0 ;
  assign n33814 = n23453 ^ n5595 ^ n3819 ;
  assign n33815 = ( n9728 & n11560 ) | ( n9728 & n19060 ) | ( n11560 & n19060 ) ;
  assign n33816 = n33815 ^ n13970 ^ n7371 ;
  assign n33817 = n28748 ^ n16475 ^ n9550 ;
  assign n33818 = n5612 & n32629 ;
  assign n33819 = ~n7351 & n33818 ;
  assign n33820 = n1889 & ~n33819 ;
  assign n33821 = n33820 ^ n11655 ^ 1'b0 ;
  assign n33822 = n1469 | n7769 ;
  assign n33823 = n29488 & ~n33822 ;
  assign n33824 = ( n11582 & n33821 ) | ( n11582 & ~n33823 ) | ( n33821 & ~n33823 ) ;
  assign n33829 = n5796 | n23089 ;
  assign n33825 = ( ~n6667 & n7712 ) | ( ~n6667 & n8102 ) | ( n7712 & n8102 ) ;
  assign n33826 = n4048 ^ n3171 ^ n1340 ;
  assign n33827 = ( n16321 & n27583 ) | ( n16321 & ~n33826 ) | ( n27583 & ~n33826 ) ;
  assign n33828 = ( n5391 & n33825 ) | ( n5391 & n33827 ) | ( n33825 & n33827 ) ;
  assign n33830 = n33829 ^ n33828 ^ n23534 ;
  assign n33831 = n6701 & ~n27581 ;
  assign n33832 = n1522 & ~n18883 ;
  assign n33833 = n33832 ^ n33257 ^ 1'b0 ;
  assign n33834 = n24818 ^ n10230 ^ x157 ;
  assign n33835 = ( n26554 & n29714 ) | ( n26554 & ~n33834 ) | ( n29714 & ~n33834 ) ;
  assign n33836 = ( n20076 & n25653 ) | ( n20076 & ~n31578 ) | ( n25653 & ~n31578 ) ;
  assign n33837 = n18856 ^ n3332 ^ n632 ;
  assign n33838 = n27431 ^ n21770 ^ n8480 ;
  assign n33839 = n33838 ^ n16242 ^ n11059 ;
  assign n33841 = ( ~n23180 & n27230 ) | ( ~n23180 & n33720 ) | ( n27230 & n33720 ) ;
  assign n33840 = n11692 & n31653 ;
  assign n33842 = n33841 ^ n33840 ^ 1'b0 ;
  assign n33843 = ( n15576 & ~n20397 ) | ( n15576 & n25698 ) | ( ~n20397 & n25698 ) ;
  assign n33844 = n33843 ^ n14412 ^ n11924 ;
  assign n33845 = n22977 ^ n22075 ^ x22 ;
  assign n33851 = n3588 & n17100 ;
  assign n33847 = n22468 ^ n16451 ^ n7949 ;
  assign n33848 = n5070 & ~n5283 ;
  assign n33849 = n33537 & ~n33848 ;
  assign n33850 = n33847 & ~n33849 ;
  assign n33852 = n33851 ^ n33850 ^ 1'b0 ;
  assign n33846 = ( n3149 & n4907 ) | ( n3149 & ~n9952 ) | ( n4907 & ~n9952 ) ;
  assign n33853 = n33852 ^ n33846 ^ 1'b0 ;
  assign n33854 = n19731 & n33853 ;
  assign n33855 = ( ~n2541 & n6367 ) | ( ~n2541 & n6641 ) | ( n6367 & n6641 ) ;
  assign n33856 = n33855 ^ n30475 ^ n15147 ;
  assign n33857 = ( ~n1099 & n4070 ) | ( ~n1099 & n17359 ) | ( n4070 & n17359 ) ;
  assign n33860 = n6144 ^ n2841 ^ n2069 ;
  assign n33861 = n33860 ^ n8238 ^ n416 ;
  assign n33858 = ( n295 & n5321 ) | ( n295 & n13599 ) | ( n5321 & n13599 ) ;
  assign n33859 = n33858 ^ n30435 ^ n326 ;
  assign n33862 = n33861 ^ n33859 ^ n15944 ;
  assign n33863 = ( ~n3343 & n26382 ) | ( ~n3343 & n33862 ) | ( n26382 & n33862 ) ;
  assign n33864 = ( n6913 & n33857 ) | ( n6913 & ~n33863 ) | ( n33857 & ~n33863 ) ;
  assign n33866 = n2469 ^ n2053 ^ 1'b0 ;
  assign n33865 = ( n6292 & n15730 ) | ( n6292 & n33608 ) | ( n15730 & n33608 ) ;
  assign n33867 = n33866 ^ n33865 ^ n14653 ;
  assign n33868 = ( n33856 & n33864 ) | ( n33856 & ~n33867 ) | ( n33864 & ~n33867 ) ;
  assign n33871 = n17831 ^ n4909 ^ 1'b0 ;
  assign n33869 = n15735 | n19003 ;
  assign n33870 = n10095 | n33869 ;
  assign n33872 = n33871 ^ n33870 ^ n6995 ;
  assign n33873 = ( ~n20506 & n20988 ) | ( ~n20506 & n28210 ) | ( n20988 & n28210 ) ;
  assign n33874 = n33873 ^ n20697 ^ n12178 ;
  assign n33875 = ( ~n16167 & n22469 ) | ( ~n16167 & n31314 ) | ( n22469 & n31314 ) ;
  assign n33876 = n33875 ^ n21286 ^ n11493 ;
  assign n33877 = n28254 ^ n26158 ^ n22260 ;
  assign n33878 = ( n2774 & n33876 ) | ( n2774 & n33877 ) | ( n33876 & n33877 ) ;
  assign n33883 = ( n413 & n27414 ) | ( n413 & n32780 ) | ( n27414 & n32780 ) ;
  assign n33880 = ( n1481 & n6177 ) | ( n1481 & ~n14288 ) | ( n6177 & ~n14288 ) ;
  assign n33881 = ( ~n8603 & n18750 ) | ( ~n8603 & n33880 ) | ( n18750 & n33880 ) ;
  assign n33879 = ( n14327 & n17901 ) | ( n14327 & n31918 ) | ( n17901 & n31918 ) ;
  assign n33882 = n33881 ^ n33879 ^ n14718 ;
  assign n33884 = n33883 ^ n33882 ^ n22852 ;
  assign n33885 = ( ~n8973 & n18480 ) | ( ~n8973 & n32626 ) | ( n18480 & n32626 ) ;
  assign n33886 = n7766 | n12866 ;
  assign n33887 = ~n22917 & n33886 ;
  assign n33888 = n25867 ^ n15877 ^ n10257 ;
  assign n33889 = ( n3242 & n4235 ) | ( n3242 & n13064 ) | ( n4235 & n13064 ) ;
  assign n33890 = ( n12257 & n13487 ) | ( n12257 & n14520 ) | ( n13487 & n14520 ) ;
  assign n33891 = ( n3092 & n33889 ) | ( n3092 & n33890 ) | ( n33889 & n33890 ) ;
  assign n33892 = n17231 ^ n9663 ^ n763 ;
  assign n33893 = n33892 ^ n24893 ^ n7515 ;
  assign n33894 = n21100 ^ n16654 ^ n15439 ;
  assign n33895 = ( n2477 & n30333 ) | ( n2477 & n33894 ) | ( n30333 & n33894 ) ;
  assign n33896 = ~n957 & n18529 ;
  assign n33897 = n33896 ^ n28261 ^ n2195 ;
  assign n33899 = ( ~n8827 & n9688 ) | ( ~n8827 & n12458 ) | ( n9688 & n12458 ) ;
  assign n33898 = ~n30062 & n31709 ;
  assign n33900 = n33899 ^ n33898 ^ 1'b0 ;
  assign n33901 = n22140 ^ n14229 ^ n8329 ;
  assign n33902 = ( ~n3578 & n7977 ) | ( ~n3578 & n33901 ) | ( n7977 & n33901 ) ;
  assign n33903 = n33902 ^ n18580 ^ n13389 ;
  assign n33904 = n33903 ^ n27261 ^ n6327 ;
  assign n33906 = ~n2741 & n13114 ;
  assign n33907 = ( ~n4028 & n4935 ) | ( ~n4028 & n33906 ) | ( n4935 & n33906 ) ;
  assign n33905 = ( ~n537 & n2372 ) | ( ~n537 & n2483 ) | ( n2372 & n2483 ) ;
  assign n33908 = n33907 ^ n33905 ^ 1'b0 ;
  assign n33909 = n33908 ^ n8948 ^ n3969 ;
  assign n33910 = ( ~n26267 & n29813 ) | ( ~n26267 & n32978 ) | ( n29813 & n32978 ) ;
  assign n33911 = n23039 ^ n21008 ^ n2747 ;
  assign n33912 = n5099 | n10683 ;
  assign n33913 = n33911 | n33912 ;
  assign n33914 = ~n14389 & n24239 ;
  assign n33915 = n33914 ^ n24366 ^ n6055 ;
  assign n33916 = n8452 & ~n9677 ;
  assign n33917 = n33916 ^ n32641 ^ n16523 ;
  assign n33924 = ( n10869 & n13517 ) | ( n10869 & n32373 ) | ( n13517 & n32373 ) ;
  assign n33922 = n29826 ^ n24124 ^ 1'b0 ;
  assign n33918 = n11473 & ~n32502 ;
  assign n33919 = n28106 & n33918 ;
  assign n33920 = n33919 ^ n14868 ^ n8480 ;
  assign n33921 = n33920 ^ n27858 ^ n27480 ;
  assign n33923 = n33922 ^ n33921 ^ n10289 ;
  assign n33925 = n33924 ^ n33923 ^ n26701 ;
  assign n33926 = ( n4071 & ~n6592 ) | ( n4071 & n8891 ) | ( ~n6592 & n8891 ) ;
  assign n33927 = ( n18775 & n31979 ) | ( n18775 & n33926 ) | ( n31979 & n33926 ) ;
  assign n33928 = ( n7426 & n17438 ) | ( n7426 & ~n33927 ) | ( n17438 & ~n33927 ) ;
  assign n33930 = ( n4540 & ~n6433 ) | ( n4540 & n17364 ) | ( ~n6433 & n17364 ) ;
  assign n33929 = ( n6732 & n15970 ) | ( n6732 & n25042 ) | ( n15970 & n25042 ) ;
  assign n33931 = n33930 ^ n33929 ^ n12292 ;
  assign n33933 = n10647 ^ n7082 ^ n4217 ;
  assign n33934 = n19970 ^ n9683 ^ n6398 ;
  assign n33935 = ( n32495 & ~n33933 ) | ( n32495 & n33934 ) | ( ~n33933 & n33934 ) ;
  assign n33932 = n18883 ^ n11100 ^ n1067 ;
  assign n33936 = n33935 ^ n33932 ^ n16418 ;
  assign n33937 = n33936 ^ n23333 ^ n5505 ;
  assign n33938 = ( ~n14291 & n15141 ) | ( ~n14291 & n33937 ) | ( n15141 & n33937 ) ;
  assign n33939 = n28979 ^ n4302 ^ n3083 ;
  assign n33945 = ~n12099 & n13893 ;
  assign n33946 = n15875 & n33945 ;
  assign n33947 = n33946 ^ n9639 ^ n3177 ;
  assign n33942 = n18836 ^ n4595 ^ n3425 ;
  assign n33943 = n33942 ^ n16880 ^ n3225 ;
  assign n33944 = n33943 ^ n7046 ^ 1'b0 ;
  assign n33940 = n28475 ^ n18779 ^ n7568 ;
  assign n33941 = n33940 ^ n16875 ^ n8628 ;
  assign n33948 = n33947 ^ n33944 ^ n33941 ;
  assign n33951 = n11740 ^ n4292 ^ n2027 ;
  assign n33949 = n17500 | n32615 ;
  assign n33950 = n9147 & ~n33949 ;
  assign n33952 = n33951 ^ n33950 ^ n28192 ;
  assign n33953 = n28816 ^ n9196 ^ 1'b0 ;
  assign n33954 = n18480 & ~n33953 ;
  assign n33956 = n32895 ^ n13753 ^ n326 ;
  assign n33955 = ( n6513 & ~n29291 ) | ( n6513 & n29595 ) | ( ~n29291 & n29595 ) ;
  assign n33957 = n33956 ^ n33955 ^ n547 ;
  assign n33958 = ( n1356 & ~n4306 ) | ( n1356 & n4712 ) | ( ~n4306 & n4712 ) ;
  assign n33959 = ~n6128 & n33958 ;
  assign n33960 = n33959 ^ n12184 ^ n2016 ;
  assign n33961 = ( ~n1719 & n24123 ) | ( ~n1719 & n29305 ) | ( n24123 & n29305 ) ;
  assign n33962 = n33961 ^ n32766 ^ n11046 ;
  assign n33963 = n22612 ^ n21367 ^ n12152 ;
  assign n33964 = n33963 ^ n28712 ^ n5651 ;
  assign n33965 = n4781 & ~n19892 ;
  assign n33967 = n12245 ^ n10953 ^ n3680 ;
  assign n33968 = n33967 ^ n7653 ^ n4224 ;
  assign n33966 = n19566 ^ n8254 ^ n4235 ;
  assign n33969 = n33968 ^ n33966 ^ n11878 ;
  assign n33970 = n14883 ^ n9877 ^ n2710 ;
  assign n33971 = n33970 ^ n21871 ^ n9889 ;
  assign n33972 = n33971 ^ n13956 ^ n10709 ;
  assign n33973 = n33972 ^ n32143 ^ n7660 ;
  assign n33974 = n19952 | n33973 ;
  assign n33975 = n33974 ^ n30286 ^ 1'b0 ;
  assign n33976 = ( n11078 & n13488 ) | ( n11078 & n18994 ) | ( n13488 & n18994 ) ;
  assign n33977 = n33976 ^ n25460 ^ n5234 ;
  assign n33978 = n11002 ^ n2204 ^ 1'b0 ;
  assign n33979 = n33978 ^ n17151 ^ n5915 ;
  assign n33980 = n33979 ^ n30593 ^ n7779 ;
  assign n33981 = n4395 ^ n3254 ^ 1'b0 ;
  assign n33982 = n1323 | n1543 ;
  assign n33983 = n33982 ^ n27765 ^ n9327 ;
  assign n33984 = n33981 | n33983 ;
  assign n33985 = n33984 ^ n26426 ^ 1'b0 ;
  assign n33986 = n33985 ^ n31369 ^ n10914 ;
  assign n33987 = ( n3516 & n10633 ) | ( n3516 & ~n22574 ) | ( n10633 & ~n22574 ) ;
  assign n33988 = n32061 & ~n32275 ;
  assign n33989 = n33987 & n33988 ;
  assign n33990 = n8378 & ~n14233 ;
  assign n33991 = n7608 & n33990 ;
  assign n33992 = ( ~n1051 & n3539 ) | ( ~n1051 & n33991 ) | ( n3539 & n33991 ) ;
  assign n33993 = n19567 | n33992 ;
  assign n33994 = n4275 & ~n23851 ;
  assign n33995 = n3500 & n33994 ;
  assign n33996 = ( n8549 & ~n30963 ) | ( n8549 & n33995 ) | ( ~n30963 & n33995 ) ;
  assign n33997 = n28476 ^ n23896 ^ n18777 ;
  assign n33998 = ~n7573 & n24444 ;
  assign n33999 = ( n431 & n13971 ) | ( n431 & n26895 ) | ( n13971 & n26895 ) ;
  assign n34000 = n28295 ^ n19204 ^ n924 ;
  assign n34001 = ( n3630 & ~n18094 ) | ( n3630 & n34000 ) | ( ~n18094 & n34000 ) ;
  assign n34002 = n34001 ^ n32747 ^ n19921 ;
  assign n34003 = ( n5555 & ~n15694 ) | ( n5555 & n16466 ) | ( ~n15694 & n16466 ) ;
  assign n34004 = n34003 ^ n19835 ^ n13177 ;
  assign n34005 = n34004 ^ n24574 ^ 1'b0 ;
  assign n34006 = ( n18263 & ~n34002 ) | ( n18263 & n34005 ) | ( ~n34002 & n34005 ) ;
  assign n34007 = ( ~n8235 & n20004 ) | ( ~n8235 & n21842 ) | ( n20004 & n21842 ) ;
  assign n34008 = n2328 & ~n3727 ;
  assign n34009 = ~n14892 & n34008 ;
  assign n34010 = n34009 ^ n12630 ^ n1731 ;
  assign n34011 = ( n2732 & n6667 ) | ( n2732 & ~n34010 ) | ( n6667 & ~n34010 ) ;
  assign n34012 = ~n15808 & n34011 ;
  assign n34013 = n10053 & ~n17065 ;
  assign n34014 = n20302 ^ n14165 ^ n9629 ;
  assign n34015 = n34014 ^ n24400 ^ n14767 ;
  assign n34016 = ( x21 & n30906 ) | ( x21 & ~n34015 ) | ( n30906 & ~n34015 ) ;
  assign n34017 = ( n13962 & n14952 ) | ( n13962 & n18925 ) | ( n14952 & n18925 ) ;
  assign n34018 = n5351 & ~n25891 ;
  assign n34019 = n28805 | n34018 ;
  assign n34020 = n34017 | n34019 ;
  assign n34021 = ( ~n8978 & n22107 ) | ( ~n8978 & n23481 ) | ( n22107 & n23481 ) ;
  assign n34022 = n27253 ^ n4565 ^ 1'b0 ;
  assign n34023 = n34022 ^ n28270 ^ n10929 ;
  assign n34024 = n16321 ^ n12733 ^ 1'b0 ;
  assign n34025 = ( n5691 & n15393 ) | ( n5691 & n34024 ) | ( n15393 & n34024 ) ;
  assign n34026 = ~n22107 & n34025 ;
  assign n34027 = n22084 ^ n12157 ^ n7804 ;
  assign n34028 = ( ~n4757 & n5612 ) | ( ~n4757 & n9758 ) | ( n5612 & n9758 ) ;
  assign n34029 = ( n24158 & ~n28491 ) | ( n24158 & n34028 ) | ( ~n28491 & n34028 ) ;
  assign n34030 = ( n19289 & ~n32872 ) | ( n19289 & n34029 ) | ( ~n32872 & n34029 ) ;
  assign n34031 = n34030 ^ n18428 ^ n4345 ;
  assign n34032 = n14383 & ~n34031 ;
  assign n34033 = ~n28401 & n34032 ;
  assign n34034 = n5806 & ~n33207 ;
  assign n34035 = n24047 ^ n22186 ^ n2198 ;
  assign n34036 = n29536 & n34035 ;
  assign n34037 = ( ~x73 & n3243 ) | ( ~x73 & n18524 ) | ( n3243 & n18524 ) ;
  assign n34038 = n33067 & ~n34037 ;
  assign n34039 = ( x90 & ~n905 ) | ( x90 & n5623 ) | ( ~n905 & n5623 ) ;
  assign n34040 = ( n3965 & n6152 ) | ( n3965 & ~n33009 ) | ( n6152 & ~n33009 ) ;
  assign n34041 = ( n3219 & n8145 ) | ( n3219 & n13814 ) | ( n8145 & n13814 ) ;
  assign n34042 = n23277 ^ n20029 ^ n13750 ;
  assign n34043 = n30324 ^ n21901 ^ n2769 ;
  assign n34044 = ( ~n18509 & n26964 ) | ( ~n18509 & n34043 ) | ( n26964 & n34043 ) ;
  assign n34045 = ( n14931 & n34042 ) | ( n14931 & ~n34044 ) | ( n34042 & ~n34044 ) ;
  assign n34046 = ( ~n26803 & n34041 ) | ( ~n26803 & n34045 ) | ( n34041 & n34045 ) ;
  assign n34047 = ( n14551 & n34040 ) | ( n14551 & ~n34046 ) | ( n34040 & ~n34046 ) ;
  assign n34048 = ( n5680 & n34039 ) | ( n5680 & n34047 ) | ( n34039 & n34047 ) ;
  assign n34049 = n2829 | n25057 ;
  assign n34050 = n34049 ^ n30600 ^ 1'b0 ;
  assign n34051 = ( n7064 & n25843 ) | ( n7064 & ~n34050 ) | ( n25843 & ~n34050 ) ;
  assign n34052 = n25981 ^ n15356 ^ n1807 ;
  assign n34053 = ( n10248 & n34051 ) | ( n10248 & n34052 ) | ( n34051 & n34052 ) ;
  assign n34054 = n22900 ^ n16863 ^ n5019 ;
  assign n34055 = n4565 & n34054 ;
  assign n34056 = n34055 ^ n2888 ^ 1'b0 ;
  assign n34057 = n18847 ^ n1395 ^ 1'b0 ;
  assign n34058 = n33248 & n34057 ;
  assign n34059 = n11281 & n26366 ;
  assign n34060 = ( n10795 & n15769 ) | ( n10795 & ~n25196 ) | ( n15769 & ~n25196 ) ;
  assign n34061 = ~n3750 & n16757 ;
  assign n34062 = n34061 ^ n24661 ^ n2870 ;
  assign n34063 = n32360 ^ n16599 ^ n12294 ;
  assign n34064 = n14595 ^ n3221 ^ n292 ;
  assign n34065 = ( n12388 & n34063 ) | ( n12388 & ~n34064 ) | ( n34063 & ~n34064 ) ;
  assign n34066 = n14283 ^ n11801 ^ n1288 ;
  assign n34067 = ( n1459 & ~n6814 ) | ( n1459 & n34066 ) | ( ~n6814 & n34066 ) ;
  assign n34068 = n6553 & n8755 ;
  assign n34069 = n2625 & n34068 ;
  assign n34070 = n34069 ^ n19640 ^ 1'b0 ;
  assign n34071 = n27566 & ~n34070 ;
  assign n34072 = ~n5354 & n34071 ;
  assign n34073 = n33185 & n34072 ;
  assign n34074 = ( n20507 & ~n23499 ) | ( n20507 & n32606 ) | ( ~n23499 & n32606 ) ;
  assign n34075 = ( n18969 & ~n19440 ) | ( n18969 & n34074 ) | ( ~n19440 & n34074 ) ;
  assign n34076 = ( ~n12898 & n17429 ) | ( ~n12898 & n18994 ) | ( n17429 & n18994 ) ;
  assign n34077 = ( ~n18166 & n24275 ) | ( ~n18166 & n34076 ) | ( n24275 & n34076 ) ;
  assign n34078 = ( n4202 & n7343 ) | ( n4202 & ~n8378 ) | ( n7343 & ~n8378 ) ;
  assign n34079 = n34078 ^ n26247 ^ n17533 ;
  assign n34080 = n4455 ^ n3284 ^ x189 ;
  assign n34081 = ( n1235 & n3878 ) | ( n1235 & n7258 ) | ( n3878 & n7258 ) ;
  assign n34082 = ( n5790 & n34080 ) | ( n5790 & n34081 ) | ( n34080 & n34081 ) ;
  assign n34083 = ( n18746 & n25283 ) | ( n18746 & n34082 ) | ( n25283 & n34082 ) ;
  assign n34084 = ( n4474 & n11095 ) | ( n4474 & ~n21035 ) | ( n11095 & ~n21035 ) ;
  assign n34085 = ( n15426 & n29758 ) | ( n15426 & n34084 ) | ( n29758 & n34084 ) ;
  assign n34086 = ( n3954 & ~n20647 ) | ( n3954 & n34085 ) | ( ~n20647 & n34085 ) ;
  assign n34087 = ( n23128 & ~n31964 ) | ( n23128 & n32494 ) | ( ~n31964 & n32494 ) ;
  assign n34088 = n32584 ^ n25634 ^ n6192 ;
  assign n34089 = n1550 | n29491 ;
  assign n34090 = n34088 | n34089 ;
  assign n34091 = ( n18457 & ~n34087 ) | ( n18457 & n34090 ) | ( ~n34087 & n34090 ) ;
  assign n34092 = ( n14166 & n14185 ) | ( n14166 & ~n31907 ) | ( n14185 & ~n31907 ) ;
  assign n34093 = n34092 ^ n29074 ^ n3138 ;
  assign n34097 = n15955 ^ n7147 ^ x227 ;
  assign n34094 = ( x196 & n6433 ) | ( x196 & ~n25612 ) | ( n6433 & ~n25612 ) ;
  assign n34095 = n34094 ^ n23558 ^ n4967 ;
  assign n34096 = ( n25726 & ~n33926 ) | ( n25726 & n34095 ) | ( ~n33926 & n34095 ) ;
  assign n34098 = n34097 ^ n34096 ^ n2551 ;
  assign n34099 = ( x0 & n1447 ) | ( x0 & n30083 ) | ( n1447 & n30083 ) ;
  assign n34100 = n11089 ^ n10896 ^ 1'b0 ;
  assign n34101 = x36 & n3929 ;
  assign n34102 = n34101 ^ n20824 ^ 1'b0 ;
  assign n34104 = n24261 ^ n7289 ^ 1'b0 ;
  assign n34105 = n34104 ^ n10182 ^ n8820 ;
  assign n34103 = n10717 ^ n3607 ^ 1'b0 ;
  assign n34106 = n34105 ^ n34103 ^ n10429 ;
  assign n34107 = n26365 ^ n25099 ^ n10050 ;
  assign n34108 = ( x161 & ~n34106 ) | ( x161 & n34107 ) | ( ~n34106 & n34107 ) ;
  assign n34109 = n727 & ~n11121 ;
  assign n34110 = ( n761 & n4169 ) | ( n761 & ~n5069 ) | ( n4169 & ~n5069 ) ;
  assign n34111 = ( n11342 & n34109 ) | ( n11342 & ~n34110 ) | ( n34109 & ~n34110 ) ;
  assign n34112 = n34111 ^ n26848 ^ n11224 ;
  assign n34113 = n12663 ^ n7234 ^ n3798 ;
  assign n34114 = n34113 ^ n25528 ^ n24395 ;
  assign n34115 = n22056 ^ n18529 ^ n18527 ;
  assign n34116 = n34115 ^ n33958 ^ n24228 ;
  assign n34117 = n26604 ^ n8260 ^ n1886 ;
  assign n34118 = ( n13226 & ~n32815 ) | ( n13226 & n34117 ) | ( ~n32815 & n34117 ) ;
  assign n34119 = ( ~n7989 & n26539 ) | ( ~n7989 & n33536 ) | ( n26539 & n33536 ) ;
  assign n34120 = ~n1116 & n34119 ;
  assign n34121 = ~n29853 & n34120 ;
  assign n34122 = ( n6220 & n28157 ) | ( n6220 & n29500 ) | ( n28157 & n29500 ) ;
  assign n34123 = ( n1541 & n28574 ) | ( n1541 & ~n34122 ) | ( n28574 & ~n34122 ) ;
  assign n34124 = n10354 ^ n8403 ^ 1'b0 ;
  assign n34125 = n34124 ^ n22036 ^ n4345 ;
  assign n34126 = n25340 ^ n22615 ^ n16184 ;
  assign n34127 = ~n16478 & n19856 ;
  assign n34128 = n34127 ^ n17845 ^ n8084 ;
  assign n34129 = ( n15410 & ~n21483 ) | ( n15410 & n32671 ) | ( ~n21483 & n32671 ) ;
  assign n34130 = ( ~n6267 & n10105 ) | ( ~n6267 & n12795 ) | ( n10105 & n12795 ) ;
  assign n34131 = ( ~n6286 & n12897 ) | ( ~n6286 & n34130 ) | ( n12897 & n34130 ) ;
  assign n34132 = ( ~n16851 & n18253 ) | ( ~n16851 & n34131 ) | ( n18253 & n34131 ) ;
  assign n34133 = n13705 | n34132 ;
  assign n34134 = n29836 ^ n18637 ^ n2691 ;
  assign n34135 = ( n21687 & n23831 ) | ( n21687 & n26693 ) | ( n23831 & n26693 ) ;
  assign n34136 = n34135 ^ n26862 ^ n23948 ;
  assign n34137 = n5015 | n31187 ;
  assign n34138 = n1927 | n34137 ;
  assign n34139 = ( n8454 & n22641 ) | ( n8454 & n31326 ) | ( n22641 & n31326 ) ;
  assign n34140 = n1656 & n16260 ;
  assign n34141 = ( n3042 & ~n21168 ) | ( n3042 & n34140 ) | ( ~n21168 & n34140 ) ;
  assign n34142 = ( ~n23786 & n34139 ) | ( ~n23786 & n34141 ) | ( n34139 & n34141 ) ;
  assign n34143 = n4103 & ~n4521 ;
  assign n34144 = ( n8212 & ~n12694 ) | ( n8212 & n34143 ) | ( ~n12694 & n34143 ) ;
  assign n34145 = n27969 ^ n8381 ^ n5317 ;
  assign n34146 = ( n324 & ~n9752 ) | ( n324 & n9967 ) | ( ~n9752 & n9967 ) ;
  assign n34147 = ( n24943 & n34145 ) | ( n24943 & ~n34146 ) | ( n34145 & ~n34146 ) ;
  assign n34148 = n29523 ^ n6528 ^ n3924 ;
  assign n34149 = n34148 ^ n30743 ^ n27569 ;
  assign n34150 = ( ~n17386 & n34147 ) | ( ~n17386 & n34149 ) | ( n34147 & n34149 ) ;
  assign n34151 = n23309 ^ n19096 ^ n17194 ;
  assign n34152 = n34151 ^ n12625 ^ 1'b0 ;
  assign n34154 = n6844 | n15437 ;
  assign n34153 = n8034 ^ n6761 ^ n5136 ;
  assign n34155 = n34154 ^ n34153 ^ n7237 ;
  assign n34156 = n19844 ^ n16882 ^ n6783 ;
  assign n34157 = ( ~n11673 & n19672 ) | ( ~n11673 & n34156 ) | ( n19672 & n34156 ) ;
  assign n34158 = n34157 ^ n8983 ^ n6468 ;
  assign n34159 = ~n18519 & n26368 ;
  assign n34160 = n34159 ^ n12575 ^ n5934 ;
  assign n34161 = ( n34155 & n34158 ) | ( n34155 & n34160 ) | ( n34158 & n34160 ) ;
  assign n34163 = n3463 & ~n6625 ;
  assign n34164 = ~n3463 & n34163 ;
  assign n34162 = ( n4408 & n11953 ) | ( n4408 & n14142 ) | ( n11953 & n14142 ) ;
  assign n34165 = n34164 ^ n34162 ^ n21232 ;
  assign n34166 = n8865 ^ n8787 ^ n3368 ;
  assign n34167 = n25559 & n34166 ;
  assign n34168 = ( ~n12590 & n14300 ) | ( ~n12590 & n15199 ) | ( n14300 & n15199 ) ;
  assign n34169 = n34168 ^ n33598 ^ n20069 ;
  assign n34170 = x129 & n16311 ;
  assign n34171 = n34170 ^ n21190 ^ 1'b0 ;
  assign n34172 = ( ~n7422 & n17482 ) | ( ~n7422 & n34171 ) | ( n17482 & n34171 ) ;
  assign n34173 = n8065 ^ n7425 ^ 1'b0 ;
  assign n34174 = ( n5109 & n9847 ) | ( n5109 & n34173 ) | ( n9847 & n34173 ) ;
  assign n34175 = n34174 ^ n10449 ^ n7334 ;
  assign n34176 = ( n12698 & n24869 ) | ( n12698 & n34175 ) | ( n24869 & n34175 ) ;
  assign n34178 = n12831 ^ n11990 ^ 1'b0 ;
  assign n34177 = n19577 ^ n11924 ^ n8701 ;
  assign n34179 = n34178 ^ n34177 ^ n1007 ;
  assign n34180 = n34179 ^ n19534 ^ n17639 ;
  assign n34181 = n13407 ^ n6443 ^ n5636 ;
  assign n34182 = n30820 ^ n17159 ^ n3013 ;
  assign n34183 = n34182 ^ n23310 ^ n16619 ;
  assign n34184 = ( n22029 & n34181 ) | ( n22029 & n34183 ) | ( n34181 & n34183 ) ;
  assign n34185 = n29721 ^ n15718 ^ n12016 ;
  assign n34186 = n25882 ^ n21240 ^ n16258 ;
  assign n34187 = ( n8414 & ~n21091 ) | ( n8414 & n34186 ) | ( ~n21091 & n34186 ) ;
  assign n34188 = ( n19281 & ~n34185 ) | ( n19281 & n34187 ) | ( ~n34185 & n34187 ) ;
  assign n34189 = ( ~n8313 & n13952 ) | ( ~n8313 & n22146 ) | ( n13952 & n22146 ) ;
  assign n34190 = n3213 & n7984 ;
  assign n34191 = n34190 ^ n16117 ^ 1'b0 ;
  assign n34192 = ( n4779 & n28654 ) | ( n4779 & n34191 ) | ( n28654 & n34191 ) ;
  assign n34193 = ( n12116 & n23209 ) | ( n12116 & n34192 ) | ( n23209 & n34192 ) ;
  assign n34194 = n34193 ^ n17065 ^ n2078 ;
  assign n34195 = n28791 ^ n14581 ^ 1'b0 ;
  assign n34196 = n18741 ^ n2388 ^ n1380 ;
  assign n34197 = n34196 ^ n33653 ^ n25235 ;
  assign n34199 = ( n3562 & ~n14412 ) | ( n3562 & n23758 ) | ( ~n14412 & n23758 ) ;
  assign n34200 = n34199 ^ n12914 ^ n9083 ;
  assign n34201 = ( n288 & n5855 ) | ( n288 & ~n34200 ) | ( n5855 & ~n34200 ) ;
  assign n34198 = ~n522 & n13382 ;
  assign n34202 = n34201 ^ n34198 ^ 1'b0 ;
  assign n34203 = n34202 ^ n28940 ^ n25333 ;
  assign n34204 = n18837 ^ n14544 ^ n13531 ;
  assign n34205 = n34204 ^ n18750 ^ n7661 ;
  assign n34206 = n29849 ^ n16717 ^ n5972 ;
  assign n34207 = ~n22608 & n34206 ;
  assign n34208 = n34205 & n34207 ;
  assign n34209 = n32852 ^ n11398 ^ n2468 ;
  assign n34210 = ~n20060 & n22399 ;
  assign n34211 = ( n17394 & n26798 ) | ( n17394 & ~n34210 ) | ( n26798 & ~n34210 ) ;
  assign n34212 = ( n8353 & ~n33011 ) | ( n8353 & n34211 ) | ( ~n33011 & n34211 ) ;
  assign n34213 = ( n7682 & n11329 ) | ( n7682 & ~n14937 ) | ( n11329 & ~n14937 ) ;
  assign n34214 = n34213 ^ n18054 ^ n5931 ;
  assign n34215 = n34214 ^ n3971 ^ n2822 ;
  assign n34216 = ( n16300 & n23108 ) | ( n16300 & n34215 ) | ( n23108 & n34215 ) ;
  assign n34218 = n9187 ^ n1226 ^ 1'b0 ;
  assign n34219 = ~n6320 & n34218 ;
  assign n34217 = ( n3080 & n6751 ) | ( n3080 & ~n13473 ) | ( n6751 & ~n13473 ) ;
  assign n34220 = n34219 ^ n34217 ^ n5841 ;
  assign n34221 = n34220 ^ n29558 ^ n12873 ;
  assign n34222 = ( ~n2790 & n10017 ) | ( ~n2790 & n13383 ) | ( n10017 & n13383 ) ;
  assign n34223 = n34222 ^ n15394 ^ n12099 ;
  assign n34224 = n34221 & ~n34223 ;
  assign n34225 = n18267 ^ n17472 ^ n1907 ;
  assign n34228 = n18920 ^ n3776 ^ n1044 ;
  assign n34229 = n34228 ^ n9366 ^ n6950 ;
  assign n34226 = n15744 ^ n8073 ^ 1'b0 ;
  assign n34227 = ( n16325 & ~n31176 ) | ( n16325 & n34226 ) | ( ~n31176 & n34226 ) ;
  assign n34230 = n34229 ^ n34227 ^ n30628 ;
  assign n34231 = n34230 ^ n27360 ^ n10338 ;
  assign n34232 = ( ~n22320 & n32745 ) | ( ~n22320 & n33056 ) | ( n32745 & n33056 ) ;
  assign n34233 = ( n896 & n6389 ) | ( n896 & ~n28272 ) | ( n6389 & ~n28272 ) ;
  assign n34234 = ( ~n19749 & n29370 ) | ( ~n19749 & n34233 ) | ( n29370 & n34233 ) ;
  assign n34235 = n27974 & n34234 ;
  assign n34236 = n7299 & ~n11496 ;
  assign n34237 = ~n34235 & n34236 ;
  assign n34238 = n14718 | n18493 ;
  assign n34239 = n34238 ^ n16168 ^ 1'b0 ;
  assign n34240 = n33536 ^ n11894 ^ n6765 ;
  assign n34241 = ~n5981 & n34240 ;
  assign n34242 = ( ~n5339 & n13967 ) | ( ~n5339 & n16434 ) | ( n13967 & n16434 ) ;
  assign n34243 = n10880 & n25222 ;
  assign n34244 = n34242 & n34243 ;
  assign n34245 = n9482 & n34244 ;
  assign n34246 = ( n14838 & ~n34241 ) | ( n14838 & n34245 ) | ( ~n34241 & n34245 ) ;
  assign n34247 = n24168 ^ n19961 ^ n17209 ;
  assign n34248 = ( ~n30458 & n32953 ) | ( ~n30458 & n34247 ) | ( n32953 & n34247 ) ;
  assign n34249 = n26838 ^ n8133 ^ n1192 ;
  assign n34250 = ( n10479 & n15960 ) | ( n10479 & ~n34249 ) | ( n15960 & ~n34249 ) ;
  assign n34251 = ( n577 & n3781 ) | ( n577 & n11963 ) | ( n3781 & n11963 ) ;
  assign n34252 = n33876 ^ n12993 ^ n548 ;
  assign n34253 = ( n5835 & ~n11984 ) | ( n5835 & n15815 ) | ( ~n11984 & n15815 ) ;
  assign n34254 = n10678 ^ n2533 ^ n1411 ;
  assign n34255 = ( n32190 & n34253 ) | ( n32190 & ~n34254 ) | ( n34253 & ~n34254 ) ;
  assign n34256 = n792 | n23481 ;
  assign n34257 = n13743 & ~n34256 ;
  assign n34258 = ( n3612 & n8542 ) | ( n3612 & ~n20663 ) | ( n8542 & ~n20663 ) ;
  assign n34259 = ( n7612 & n34257 ) | ( n7612 & ~n34258 ) | ( n34257 & ~n34258 ) ;
  assign n34260 = n12513 ^ n3934 ^ n3414 ;
  assign n34261 = n34260 ^ n20653 ^ n3082 ;
  assign n34262 = n34261 ^ n15698 ^ n13593 ;
  assign n34263 = ( ~n7516 & n15798 ) | ( ~n7516 & n16031 ) | ( n15798 & n16031 ) ;
  assign n34264 = ( ~n6183 & n22698 ) | ( ~n6183 & n34263 ) | ( n22698 & n34263 ) ;
  assign n34265 = n34264 ^ n25694 ^ n22876 ;
  assign n34266 = n34265 ^ n31227 ^ n27654 ;
  assign n34267 = ( ~n842 & n3196 ) | ( ~n842 & n4850 ) | ( n3196 & n4850 ) ;
  assign n34268 = n34267 ^ n13661 ^ 1'b0 ;
  assign n34269 = n3827 ^ n3407 ^ 1'b0 ;
  assign n34270 = ~n34268 & n34269 ;
  assign n34271 = n33638 ^ n20844 ^ 1'b0 ;
  assign n34272 = n12495 & ~n34271 ;
  assign n34273 = n33922 ^ n2803 ^ n2206 ;
  assign n34275 = n21687 ^ n20166 ^ n14204 ;
  assign n34274 = ( n9269 & ~n15000 ) | ( n9269 & n30956 ) | ( ~n15000 & n30956 ) ;
  assign n34276 = n34275 ^ n34274 ^ n19612 ;
  assign n34277 = n9155 ^ n4074 ^ 1'b0 ;
  assign n34278 = n1153 | n34277 ;
  assign n34279 = ( ~n8013 & n12415 ) | ( ~n8013 & n16562 ) | ( n12415 & n16562 ) ;
  assign n34280 = n34279 ^ n6853 ^ 1'b0 ;
  assign n34281 = n34280 ^ n4686 ^ n1544 ;
  assign n34282 = ( n12850 & n34278 ) | ( n12850 & n34281 ) | ( n34278 & n34281 ) ;
  assign n34290 = n20625 ^ n9222 ^ n9097 ;
  assign n34291 = n34290 ^ n21431 ^ 1'b0 ;
  assign n34287 = n5533 ^ n3079 ^ n2695 ;
  assign n34288 = ~n1477 & n34287 ;
  assign n34284 = ( n680 & n5599 ) | ( n680 & n16866 ) | ( n5599 & n16866 ) ;
  assign n34283 = n17955 ^ n16414 ^ n4918 ;
  assign n34285 = n34284 ^ n34283 ^ n6320 ;
  assign n34286 = n34285 ^ n20015 ^ 1'b0 ;
  assign n34289 = n34288 ^ n34286 ^ n14333 ;
  assign n34292 = n34291 ^ n34289 ^ n32503 ;
  assign n34294 = n7621 | n19623 ;
  assign n34295 = ~n27830 & n29683 ;
  assign n34296 = ~n34294 & n34295 ;
  assign n34293 = ( x174 & n13600 ) | ( x174 & n16547 ) | ( n13600 & n16547 ) ;
  assign n34297 = n34296 ^ n34293 ^ n4312 ;
  assign n34298 = n2566 | n3300 ;
  assign n34299 = n3288 & ~n34298 ;
  assign n34301 = ( ~n3804 & n18808 ) | ( ~n3804 & n25678 ) | ( n18808 & n25678 ) ;
  assign n34300 = ~n13127 & n17101 ;
  assign n34302 = n34301 ^ n34300 ^ 1'b0 ;
  assign n34303 = n34302 ^ n26115 ^ n3614 ;
  assign n34304 = ( n2179 & n8203 ) | ( n2179 & ~n21938 ) | ( n8203 & ~n21938 ) ;
  assign n34305 = ~n15564 & n28764 ;
  assign n34306 = ~n6807 & n34305 ;
  assign n34307 = ( n310 & n785 ) | ( n310 & ~n16866 ) | ( n785 & ~n16866 ) ;
  assign n34308 = n34307 ^ n3694 ^ 1'b0 ;
  assign n34309 = n34308 ^ n6971 ^ n6073 ;
  assign n34310 = n34309 ^ n31997 ^ n6011 ;
  assign n34311 = ( ~n9853 & n29253 ) | ( ~n9853 & n34310 ) | ( n29253 & n34310 ) ;
  assign n34312 = n34311 ^ n33063 ^ n7117 ;
  assign n34313 = ( n9625 & n12399 ) | ( n9625 & ~n33550 ) | ( n12399 & ~n33550 ) ;
  assign n34314 = ( n3724 & n10773 ) | ( n3724 & n13939 ) | ( n10773 & n13939 ) ;
  assign n34315 = n34314 ^ n6546 ^ n2773 ;
  assign n34316 = n34315 ^ n29804 ^ 1'b0 ;
  assign n34317 = ( ~n5280 & n33322 ) | ( ~n5280 & n34316 ) | ( n33322 & n34316 ) ;
  assign n34318 = ( ~n3618 & n19146 ) | ( ~n3618 & n22412 ) | ( n19146 & n22412 ) ;
  assign n34319 = ( n12857 & ~n14412 ) | ( n12857 & n34318 ) | ( ~n14412 & n34318 ) ;
  assign n34320 = ( n6112 & ~n24482 ) | ( n6112 & n34035 ) | ( ~n24482 & n34035 ) ;
  assign n34321 = n10509 ^ n4002 ^ n262 ;
  assign n34322 = n14451 ^ n11664 ^ 1'b0 ;
  assign n34323 = n6256 & n34322 ;
  assign n34324 = ( ~n2991 & n4042 ) | ( ~n2991 & n16991 ) | ( n4042 & n16991 ) ;
  assign n34325 = ( n30490 & ~n34323 ) | ( n30490 & n34324 ) | ( ~n34323 & n34324 ) ;
  assign n34326 = n30445 ^ n3659 ^ 1'b0 ;
  assign n34327 = ~n34325 & n34326 ;
  assign n34328 = ( n5571 & n16060 ) | ( n5571 & n27347 ) | ( n16060 & n27347 ) ;
  assign n34331 = ~n4094 & n5084 ;
  assign n34329 = n16754 ^ n1718 ^ 1'b0 ;
  assign n34330 = n34329 ^ n9661 ^ n3759 ;
  assign n34332 = n34331 ^ n34330 ^ n13614 ;
  assign n34333 = n27064 ^ n25911 ^ n19213 ;
  assign n34337 = n8344 ^ n631 ^ 1'b0 ;
  assign n34338 = n6010 & n34337 ;
  assign n34339 = n34338 ^ n11820 ^ n2201 ;
  assign n34340 = ( n16708 & n26626 ) | ( n16708 & ~n34339 ) | ( n26626 & ~n34339 ) ;
  assign n34334 = n21097 ^ n19999 ^ n11328 ;
  assign n34335 = ( n3263 & ~n6829 ) | ( n3263 & n34334 ) | ( ~n6829 & n34334 ) ;
  assign n34336 = n34335 ^ n14976 ^ n13226 ;
  assign n34341 = n34340 ^ n34336 ^ n19685 ;
  assign n34345 = n15574 ^ n6646 ^ 1'b0 ;
  assign n34342 = ( ~n9510 & n11325 ) | ( ~n9510 & n25390 ) | ( n11325 & n25390 ) ;
  assign n34343 = ( ~n4927 & n24410 ) | ( ~n4927 & n34342 ) | ( n24410 & n34342 ) ;
  assign n34344 = n34343 ^ n14670 ^ n7085 ;
  assign n34346 = n34345 ^ n34344 ^ n12638 ;
  assign n34347 = ( ~x181 & n7646 ) | ( ~x181 & n9021 ) | ( n7646 & n9021 ) ;
  assign n34348 = ( ~n2045 & n14873 ) | ( ~n2045 & n27788 ) | ( n14873 & n27788 ) ;
  assign n34349 = n34348 ^ n20113 ^ 1'b0 ;
  assign n34350 = n34349 ^ n13288 ^ n511 ;
  assign n34351 = ( n11023 & ~n34347 ) | ( n11023 & n34350 ) | ( ~n34347 & n34350 ) ;
  assign n34359 = n19163 ^ n14030 ^ n6726 ;
  assign n34352 = n10515 ^ n9621 ^ n4610 ;
  assign n34353 = n25193 ^ n11288 ^ x235 ;
  assign n34354 = n25630 & n34353 ;
  assign n34355 = n34352 & n34354 ;
  assign n34356 = n14860 & ~n22932 ;
  assign n34357 = n34356 ^ n3235 ^ 1'b0 ;
  assign n34358 = ( n19313 & ~n34355 ) | ( n19313 & n34357 ) | ( ~n34355 & n34357 ) ;
  assign n34360 = n34359 ^ n34358 ^ n17722 ;
  assign n34361 = n34360 ^ n28918 ^ n28880 ;
  assign n34362 = n34361 ^ n11699 ^ n1770 ;
  assign n34363 = n10480 ^ n5995 ^ 1'b0 ;
  assign n34364 = ( n8045 & n18086 ) | ( n8045 & n22240 ) | ( n18086 & n22240 ) ;
  assign n34365 = n31005 ^ n17016 ^ n4726 ;
  assign n34366 = n27789 ^ n10598 ^ n2044 ;
  assign n34367 = ( n11001 & n21630 ) | ( n11001 & ~n34366 ) | ( n21630 & ~n34366 ) ;
  assign n34375 = ( n7345 & n8480 ) | ( n7345 & n12871 ) | ( n8480 & n12871 ) ;
  assign n34372 = n5784 | n13600 ;
  assign n34373 = n34372 ^ n26698 ^ 1'b0 ;
  assign n34374 = ( n8876 & n19767 ) | ( n8876 & ~n34373 ) | ( n19767 & ~n34373 ) ;
  assign n34368 = n15517 ^ n10887 ^ 1'b0 ;
  assign n34369 = n9381 & n34368 ;
  assign n34370 = ( n3205 & n23590 ) | ( n3205 & n33403 ) | ( n23590 & n33403 ) ;
  assign n34371 = ( n28787 & n34369 ) | ( n28787 & n34370 ) | ( n34369 & n34370 ) ;
  assign n34376 = n34375 ^ n34374 ^ n34371 ;
  assign n34377 = n13274 ^ n9836 ^ n4862 ;
  assign n34378 = ( n8744 & n19704 ) | ( n8744 & n34377 ) | ( n19704 & n34377 ) ;
  assign n34379 = ( ~n2015 & n17572 ) | ( ~n2015 & n20680 ) | ( n17572 & n20680 ) ;
  assign n34380 = ( n1341 & n21198 ) | ( n1341 & n26550 ) | ( n21198 & n26550 ) ;
  assign n34381 = ( ~n25487 & n34379 ) | ( ~n25487 & n34380 ) | ( n34379 & n34380 ) ;
  assign n34382 = n33483 ^ n25263 ^ n1231 ;
  assign n34383 = n27576 ^ n20405 ^ n3253 ;
  assign n34384 = n34383 ^ n17253 ^ n2061 ;
  assign n34385 = ( ~n7208 & n11611 ) | ( ~n7208 & n20796 ) | ( n11611 & n20796 ) ;
  assign n34386 = n20252 ^ n19358 ^ n7308 ;
  assign n34387 = n34386 ^ n31997 ^ 1'b0 ;
  assign n34389 = n6540 & ~n17379 ;
  assign n34390 = n34389 ^ n28979 ^ 1'b0 ;
  assign n34391 = n34390 ^ n16097 ^ n5261 ;
  assign n34392 = ( n8746 & ~n32911 ) | ( n8746 & n34391 ) | ( ~n32911 & n34391 ) ;
  assign n34388 = ( ~x83 & n2480 ) | ( ~x83 & n10179 ) | ( n2480 & n10179 ) ;
  assign n34393 = n34392 ^ n34388 ^ n5984 ;
  assign n34394 = n34393 ^ n33711 ^ n13093 ;
  assign n34395 = ( ~n422 & n14411 ) | ( ~n422 & n31703 ) | ( n14411 & n31703 ) ;
  assign n34396 = n34395 ^ n12207 ^ n4121 ;
  assign n34397 = ( n7173 & n8344 ) | ( n7173 & ~n26882 ) | ( n8344 & ~n26882 ) ;
  assign n34398 = n34397 ^ n27221 ^ n4283 ;
  assign n34402 = n24789 ^ n16689 ^ n3445 ;
  assign n34403 = n20576 ^ n18363 ^ n15849 ;
  assign n34404 = ( n7284 & ~n34402 ) | ( n7284 & n34403 ) | ( ~n34402 & n34403 ) ;
  assign n34405 = ( n4229 & ~n26437 ) | ( n4229 & n34404 ) | ( ~n26437 & n34404 ) ;
  assign n34400 = n13154 ^ n1198 ^ 1'b0 ;
  assign n34399 = ( n21449 & ~n28906 ) | ( n21449 & n33185 ) | ( ~n28906 & n33185 ) ;
  assign n34401 = n34400 ^ n34399 ^ x215 ;
  assign n34406 = n34405 ^ n34401 ^ n20988 ;
  assign n34407 = n5248 ^ n4509 ^ n3305 ;
  assign n34408 = n27913 | n34407 ;
  assign n34409 = n18857 & ~n34408 ;
  assign n34410 = ( n18963 & ~n32961 ) | ( n18963 & n34409 ) | ( ~n32961 & n34409 ) ;
  assign n34412 = ( x241 & ~n20842 ) | ( x241 & n22503 ) | ( ~n20842 & n22503 ) ;
  assign n34411 = ( n2741 & n6848 ) | ( n2741 & n10866 ) | ( n6848 & n10866 ) ;
  assign n34413 = n34412 ^ n34411 ^ n16253 ;
  assign n34414 = n21044 ^ n12435 ^ n3619 ;
  assign n34415 = n34414 ^ n13980 ^ n7668 ;
  assign n34416 = ( n2430 & ~n11633 ) | ( n2430 & n34415 ) | ( ~n11633 & n34415 ) ;
  assign n34417 = n4145 & ~n9611 ;
  assign n34418 = ~n20585 & n34417 ;
  assign n34419 = n19487 & ~n34418 ;
  assign n34420 = n8472 & n34419 ;
  assign n34422 = n12652 ^ n11716 ^ n8930 ;
  assign n34423 = n34422 ^ n13375 ^ n7943 ;
  assign n34421 = n26694 ^ n13448 ^ n3677 ;
  assign n34424 = n34423 ^ n34421 ^ n21394 ;
  assign n34425 = n26185 ^ n4877 ^ 1'b0 ;
  assign n34427 = ( n3202 & n16225 ) | ( n3202 & n21486 ) | ( n16225 & n21486 ) ;
  assign n34428 = ( ~n1380 & n25087 ) | ( ~n1380 & n34427 ) | ( n25087 & n34427 ) ;
  assign n34426 = n29420 ^ n13955 ^ n8761 ;
  assign n34429 = n34428 ^ n34426 ^ n27437 ;
  assign n34430 = n34429 ^ n33123 ^ n33091 ;
  assign n34432 = ( ~n5975 & n22871 ) | ( ~n5975 & n24590 ) | ( n22871 & n24590 ) ;
  assign n34431 = n26018 ^ n15213 ^ 1'b0 ;
  assign n34433 = n34432 ^ n34431 ^ n19085 ;
  assign n34434 = n18333 ^ n5769 ^ n5727 ;
  assign n34435 = n27882 ^ n20929 ^ n11613 ;
  assign n34436 = n10078 ^ n2840 ^ n368 ;
  assign n34437 = n34436 ^ n9296 ^ n1810 ;
  assign n34438 = n34437 ^ n17281 ^ n5360 ;
  assign n34439 = ( n21206 & n34435 ) | ( n21206 & ~n34438 ) | ( n34435 & ~n34438 ) ;
  assign n34440 = ( ~n14739 & n16640 ) | ( ~n14739 & n33530 ) | ( n16640 & n33530 ) ;
  assign n34441 = n11554 ^ n7908 ^ n6117 ;
  assign n34442 = ( n8054 & n8249 ) | ( n8054 & ~n34441 ) | ( n8249 & ~n34441 ) ;
  assign n34443 = ( ~n18181 & n32502 ) | ( ~n18181 & n34442 ) | ( n32502 & n34442 ) ;
  assign n34444 = ( ~n13993 & n29893 ) | ( ~n13993 & n34228 ) | ( n29893 & n34228 ) ;
  assign n34445 = ( ~n6261 & n18043 ) | ( ~n6261 & n34444 ) | ( n18043 & n34444 ) ;
  assign n34446 = n26654 ^ n20104 ^ 1'b0 ;
  assign n34447 = ( ~n6804 & n32570 ) | ( ~n6804 & n34446 ) | ( n32570 & n34446 ) ;
  assign n34448 = ( n7783 & n34104 ) | ( n7783 & n34447 ) | ( n34104 & n34447 ) ;
  assign n34449 = n31839 ^ n28791 ^ n26810 ;
  assign n34450 = ( n8564 & n28120 ) | ( n8564 & n28769 ) | ( n28120 & n28769 ) ;
  assign n34452 = n21256 ^ n4349 ^ 1'b0 ;
  assign n34453 = n26020 | n34452 ;
  assign n34454 = n34453 ^ n17467 ^ n5053 ;
  assign n34451 = ~n11823 & n17955 ;
  assign n34455 = n34454 ^ n34451 ^ 1'b0 ;
  assign n34456 = n8809 | n23231 ;
  assign n34457 = n34456 ^ n28845 ^ n8886 ;
  assign n34458 = n9364 & ~n18019 ;
  assign n34459 = n34458 ^ n32056 ^ 1'b0 ;
  assign n34460 = n24955 | n34459 ;
  assign n34461 = n34457 | n34460 ;
  assign n34462 = ( n741 & ~n5754 ) | ( n741 & n21450 ) | ( ~n5754 & n21450 ) ;
  assign n34463 = ( n3053 & ~n20384 ) | ( n3053 & n34462 ) | ( ~n20384 & n34462 ) ;
  assign n34464 = n10389 ^ n4344 ^ x72 ;
  assign n34465 = n34464 ^ n19509 ^ n14037 ;
  assign n34466 = ( n7094 & n17940 ) | ( n7094 & ~n20232 ) | ( n17940 & ~n20232 ) ;
  assign n34467 = n10203 ^ n6539 ^ 1'b0 ;
  assign n34468 = n8567 & ~n34467 ;
  assign n34469 = n22961 ^ n899 ^ 1'b0 ;
  assign n34470 = n34468 & ~n34469 ;
  assign n34471 = ~n4343 & n34470 ;
  assign n34472 = ~n29775 & n34471 ;
  assign n34473 = ( n14851 & ~n15292 ) | ( n14851 & n17075 ) | ( ~n15292 & n17075 ) ;
  assign n34474 = n9104 & n34473 ;
  assign n34475 = n7338 ^ n1864 ^ n502 ;
  assign n34476 = n34475 ^ n15333 ^ n5502 ;
  assign n34477 = n34476 ^ n33075 ^ n7908 ;
  assign n34478 = ( n26119 & n30209 ) | ( n26119 & ~n32860 ) | ( n30209 & ~n32860 ) ;
  assign n34479 = ( ~x63 & n4685 ) | ( ~x63 & n34478 ) | ( n4685 & n34478 ) ;
  assign n34484 = ( n3982 & n10602 ) | ( n3982 & n15114 ) | ( n10602 & n15114 ) ;
  assign n34483 = n17839 ^ n13478 ^ n2839 ;
  assign n34485 = n34484 ^ n34483 ^ n5314 ;
  assign n34480 = n11194 ^ n1143 ^ n444 ;
  assign n34481 = n575 & n34480 ;
  assign n34482 = n34481 ^ n23647 ^ n22656 ;
  assign n34486 = n34485 ^ n34482 ^ n30111 ;
  assign n34487 = n19493 ^ n7254 ^ 1'b0 ;
  assign n34488 = n33645 | n34487 ;
  assign n34489 = n34488 ^ n33624 ^ n3257 ;
  assign n34490 = n34489 ^ n28361 ^ n14866 ;
  assign n34491 = n1934 | n28639 ;
  assign n34492 = n19646 & ~n34491 ;
  assign n34493 = n4101 & n8034 ;
  assign n34494 = n8156 ^ n6142 ^ n1880 ;
  assign n34495 = n34494 ^ n18640 ^ n16295 ;
  assign n34496 = ( ~n2329 & n10810 ) | ( ~n2329 & n13210 ) | ( n10810 & n13210 ) ;
  assign n34497 = n8525 ^ n4839 ^ n3762 ;
  assign n34498 = n34497 ^ n31680 ^ n13113 ;
  assign n34504 = n14623 ^ n7191 ^ n5726 ;
  assign n34503 = n29478 ^ n9829 ^ x193 ;
  assign n34505 = n34504 ^ n34503 ^ n11758 ;
  assign n34501 = n18214 ^ n16438 ^ n9858 ;
  assign n34502 = n34501 ^ n31412 ^ n25148 ;
  assign n34506 = n34505 ^ n34502 ^ n6321 ;
  assign n34499 = n8716 ^ n5915 ^ n815 ;
  assign n34500 = n3274 & n34499 ;
  assign n34507 = n34506 ^ n34500 ^ 1'b0 ;
  assign n34508 = n16843 ^ n15317 ^ n3648 ;
  assign n34509 = ( ~n572 & n2433 ) | ( ~n572 & n34508 ) | ( n2433 & n34508 ) ;
  assign n34510 = ( x125 & n3645 ) | ( x125 & n15746 ) | ( n3645 & n15746 ) ;
  assign n34511 = n34510 ^ n18610 ^ n2029 ;
  assign n34512 = ( n28476 & ~n34509 ) | ( n28476 & n34511 ) | ( ~n34509 & n34511 ) ;
  assign n34513 = n33147 ^ n22591 ^ n21557 ;
  assign n34515 = ( x161 & n10433 ) | ( x161 & ~n10970 ) | ( n10433 & ~n10970 ) ;
  assign n34514 = ( ~n1586 & n13654 ) | ( ~n1586 & n18274 ) | ( n13654 & n18274 ) ;
  assign n34516 = n34515 ^ n34514 ^ n32000 ;
  assign n34517 = ( n2514 & n3467 ) | ( n2514 & ~n20524 ) | ( n3467 & ~n20524 ) ;
  assign n34518 = n34517 ^ n19736 ^ n8350 ;
  assign n34519 = n5315 | n17205 ;
  assign n34520 = n34519 ^ n23938 ^ 1'b0 ;
  assign n34521 = ( n19789 & n34518 ) | ( n19789 & n34520 ) | ( n34518 & n34520 ) ;
  assign n34522 = n31338 ^ n9487 ^ 1'b0 ;
  assign n34523 = ( ~n4802 & n8753 ) | ( ~n4802 & n21071 ) | ( n8753 & n21071 ) ;
  assign n34524 = n34523 ^ n27553 ^ n12673 ;
  assign n34525 = ( n2720 & n20033 ) | ( n2720 & ~n33358 ) | ( n20033 & ~n33358 ) ;
  assign n34526 = n33047 | n34525 ;
  assign n34527 = n5896 ^ n4181 ^ 1'b0 ;
  assign n34528 = n1748 & n34527 ;
  assign n34529 = ( ~n24843 & n33724 ) | ( ~n24843 & n34528 ) | ( n33724 & n34528 ) ;
  assign n34530 = n34529 ^ n25239 ^ n4835 ;
  assign n34531 = n5443 ^ n2957 ^ n1407 ;
  assign n34532 = n34531 ^ n31404 ^ n4544 ;
  assign n34533 = n34532 ^ n17184 ^ n10625 ;
  assign n34535 = n9111 ^ n8256 ^ n2415 ;
  assign n34534 = ~n21672 & n27862 ;
  assign n34536 = n34535 ^ n34534 ^ 1'b0 ;
  assign n34537 = n34536 ^ n29085 ^ n17683 ;
  assign n34538 = ( n6097 & ~n7576 ) | ( n6097 & n34537 ) | ( ~n7576 & n34537 ) ;
  assign n34539 = n17777 ^ n5730 ^ n890 ;
  assign n34540 = ( n5305 & ~n7321 ) | ( n5305 & n23059 ) | ( ~n7321 & n23059 ) ;
  assign n34541 = n10931 ^ n2968 ^ n1762 ;
  assign n34542 = ( n5805 & n34540 ) | ( n5805 & ~n34541 ) | ( n34540 & ~n34541 ) ;
  assign n34544 = n28432 ^ n15628 ^ n3234 ;
  assign n34545 = n34544 ^ n6444 ^ 1'b0 ;
  assign n34543 = n7070 & n9982 ;
  assign n34546 = n34545 ^ n34543 ^ 1'b0 ;
  assign n34547 = ( n5082 & n10832 ) | ( n5082 & ~n27106 ) | ( n10832 & ~n27106 ) ;
  assign n34548 = n20442 | n34547 ;
  assign n34549 = n34548 ^ n5934 ^ n1963 ;
  assign n34550 = ( n3404 & n7940 ) | ( n3404 & ~n32417 ) | ( n7940 & ~n32417 ) ;
  assign n34551 = x137 & n18126 ;
  assign n34552 = n34551 ^ n11364 ^ 1'b0 ;
  assign n34553 = n15421 ^ n12285 ^ 1'b0 ;
  assign n34554 = n34552 & ~n34553 ;
  assign n34555 = n9732 & n34554 ;
  assign n34556 = n25025 & n34555 ;
  assign n34557 = ( n6272 & n21388 ) | ( n6272 & ~n34556 ) | ( n21388 & ~n34556 ) ;
  assign n34558 = ( n14898 & n31437 ) | ( n14898 & ~n34557 ) | ( n31437 & ~n34557 ) ;
  assign n34559 = ( n7736 & ~n18527 ) | ( n7736 & n34558 ) | ( ~n18527 & n34558 ) ;
  assign n34560 = ( n3196 & n13874 ) | ( n3196 & ~n20027 ) | ( n13874 & ~n20027 ) ;
  assign n34561 = n2506 & n5629 ;
  assign n34562 = ~n33653 & n34561 ;
  assign n34563 = ( ~n27969 & n34560 ) | ( ~n27969 & n34562 ) | ( n34560 & n34562 ) ;
  assign n34564 = ( n2349 & n18620 ) | ( n2349 & ~n28631 ) | ( n18620 & ~n28631 ) ;
  assign n34565 = ( ~n858 & n2200 ) | ( ~n858 & n12403 ) | ( n2200 & n12403 ) ;
  assign n34566 = n24184 ^ n6748 ^ 1'b0 ;
  assign n34567 = n4551 | n34566 ;
  assign n34568 = n34567 ^ n30374 ^ n3119 ;
  assign n34569 = n34568 ^ n1515 ^ 1'b0 ;
  assign n34570 = ( n19965 & n33914 ) | ( n19965 & ~n34569 ) | ( n33914 & ~n34569 ) ;
  assign n34571 = ( n5767 & n8105 ) | ( n5767 & n24947 ) | ( n8105 & n24947 ) ;
  assign n34572 = n19351 ^ n4467 ^ n2443 ;
  assign n34573 = n34572 ^ n28048 ^ n12733 ;
  assign n34574 = n13090 ^ n4336 ^ 1'b0 ;
  assign n34575 = n10139 & ~n34574 ;
  assign n34576 = n34575 ^ n31989 ^ n30182 ;
  assign n34577 = n29617 ^ n9891 ^ n5975 ;
  assign n34578 = ( n713 & ~n21572 ) | ( n713 & n34577 ) | ( ~n21572 & n34577 ) ;
  assign n34579 = n16727 | n34578 ;
  assign n34580 = ( ~n2080 & n9500 ) | ( ~n2080 & n15587 ) | ( n9500 & n15587 ) ;
  assign n34581 = ( ~n6805 & n8270 ) | ( ~n6805 & n34580 ) | ( n8270 & n34580 ) ;
  assign n34582 = ~n30510 & n34581 ;
  assign n34583 = n34582 ^ n2267 ^ 1'b0 ;
  assign n34584 = n19448 ^ n10915 ^ 1'b0 ;
  assign n34585 = n34584 ^ n1029 ^ 1'b0 ;
  assign n34586 = n27518 & ~n34585 ;
  assign n34587 = n22838 ^ n19292 ^ n2181 ;
  assign n34588 = ~n11097 & n24018 ;
  assign n34589 = n34588 ^ n13713 ^ 1'b0 ;
  assign n34590 = n17747 ^ n17631 ^ 1'b0 ;
  assign n34591 = n3105 & ~n34590 ;
  assign n34592 = n34591 ^ n13797 ^ n1571 ;
  assign n34593 = ( n3640 & ~n34589 ) | ( n3640 & n34592 ) | ( ~n34589 & n34592 ) ;
  assign n34594 = n21825 & n22133 ;
  assign n34595 = n34594 ^ n34200 ^ 1'b0 ;
  assign n34596 = ~n14747 & n34595 ;
  assign n34597 = ~n25766 & n34596 ;
  assign n34598 = n2017 & n6585 ;
  assign n34599 = ~n2311 & n34598 ;
  assign n34600 = n23087 & ~n34599 ;
  assign n34601 = ( n12129 & n24135 ) | ( n12129 & ~n34600 ) | ( n24135 & ~n34600 ) ;
  assign n34602 = ( ~n13995 & n18300 ) | ( ~n13995 & n29660 ) | ( n18300 & n29660 ) ;
  assign n34603 = ( n1465 & ~n1681 ) | ( n1465 & n21393 ) | ( ~n1681 & n21393 ) ;
  assign n34604 = ( n21135 & n34602 ) | ( n21135 & ~n34603 ) | ( n34602 & ~n34603 ) ;
  assign n34605 = ( ~n16187 & n22993 ) | ( ~n16187 & n34604 ) | ( n22993 & n34604 ) ;
  assign n34606 = ( n2426 & ~n12458 ) | ( n2426 & n17931 ) | ( ~n12458 & n17931 ) ;
  assign n34607 = n34606 ^ n15113 ^ n14225 ;
  assign n34609 = n23473 ^ n18701 ^ n17120 ;
  assign n34608 = ( n848 & ~n11457 ) | ( n848 & n14491 ) | ( ~n11457 & n14491 ) ;
  assign n34610 = n34609 ^ n34608 ^ n5093 ;
  assign n34611 = n34610 ^ n17020 ^ n7160 ;
  assign n34612 = ( n3223 & n5338 ) | ( n3223 & n7365 ) | ( n5338 & n7365 ) ;
  assign n34613 = n34612 ^ n20945 ^ n11929 ;
  assign n34614 = n20151 ^ n5383 ^ n1181 ;
  assign n34615 = n12914 | n34614 ;
  assign n34616 = n18640 | n34615 ;
  assign n34617 = ( n1569 & n4009 ) | ( n1569 & ~n6501 ) | ( n4009 & ~n6501 ) ;
  assign n34618 = n34617 ^ n6296 ^ n327 ;
  assign n34619 = n34618 ^ n22917 ^ 1'b0 ;
  assign n34620 = n6959 ^ n6341 ^ n3338 ;
  assign n34621 = ( n466 & ~n8365 ) | ( n466 & n21765 ) | ( ~n8365 & n21765 ) ;
  assign n34622 = n34621 ^ n31899 ^ x7 ;
  assign n34623 = ( n2493 & n3407 ) | ( n2493 & ~n25553 ) | ( n3407 & ~n25553 ) ;
  assign n34625 = ( ~n5752 & n10215 ) | ( ~n5752 & n12871 ) | ( n10215 & n12871 ) ;
  assign n34626 = n34625 ^ n20865 ^ 1'b0 ;
  assign n34624 = ~n27830 & n28269 ;
  assign n34627 = n34626 ^ n34624 ^ 1'b0 ;
  assign n34628 = n23017 ^ n10634 ^ n4442 ;
  assign n34629 = n26236 ^ n22109 ^ n8934 ;
  assign n34630 = n14158 ^ n7808 ^ n6491 ;
  assign n34631 = n34630 ^ n7252 ^ n3797 ;
  assign n34632 = ( ~n2052 & n34629 ) | ( ~n2052 & n34631 ) | ( n34629 & n34631 ) ;
  assign n34633 = n34632 ^ n31173 ^ n7700 ;
  assign n34634 = n34633 ^ n27356 ^ n12579 ;
  assign n34635 = ( n14467 & n34628 ) | ( n14467 & ~n34634 ) | ( n34628 & ~n34634 ) ;
  assign n34636 = n24865 ^ n11688 ^ n612 ;
  assign n34637 = n28301 ^ n27751 ^ n18620 ;
  assign n34638 = ( n6150 & ~n34636 ) | ( n6150 & n34637 ) | ( ~n34636 & n34637 ) ;
  assign n34639 = n34638 ^ n31483 ^ n15937 ;
  assign n34640 = n29226 ^ n22326 ^ n4292 ;
  assign n34641 = n9700 ^ n4608 ^ n2644 ;
  assign n34642 = ( n18526 & ~n25404 ) | ( n18526 & n34641 ) | ( ~n25404 & n34641 ) ;
  assign n34646 = ( n9703 & n16963 ) | ( n9703 & ~n16976 ) | ( n16963 & ~n16976 ) ;
  assign n34644 = n16267 ^ n3441 ^ 1'b0 ;
  assign n34645 = n34644 ^ n22987 ^ n16505 ;
  assign n34647 = n34646 ^ n34645 ^ n11866 ;
  assign n34643 = n1117 & n5710 ;
  assign n34648 = n34647 ^ n34643 ^ 1'b0 ;
  assign n34649 = n34648 ^ n27625 ^ n3804 ;
  assign n34650 = n7962 ^ n6761 ^ n5384 ;
  assign n34651 = n3040 & ~n34650 ;
  assign n34652 = n34651 ^ n33385 ^ 1'b0 ;
  assign n34653 = ( n22176 & n31219 ) | ( n22176 & ~n34652 ) | ( n31219 & ~n34652 ) ;
  assign n34654 = n9600 & n20945 ;
  assign n34655 = ~n5442 & n34654 ;
  assign n34656 = ( n1000 & n18064 ) | ( n1000 & n30881 ) | ( n18064 & n30881 ) ;
  assign n34657 = ( ~n1540 & n2750 ) | ( ~n1540 & n34656 ) | ( n2750 & n34656 ) ;
  assign n34658 = ( ~n7373 & n9030 ) | ( ~n7373 & n9182 ) | ( n9030 & n9182 ) ;
  assign n34659 = ( n12048 & n30014 ) | ( n12048 & n34658 ) | ( n30014 & n34658 ) ;
  assign n34660 = n34659 ^ n21824 ^ n11473 ;
  assign n34661 = n922 | n17047 ;
  assign n34662 = n34660 | n34661 ;
  assign n34663 = n34662 ^ n6703 ^ 1'b0 ;
  assign n34664 = n8209 ^ n1550 ^ 1'b0 ;
  assign n34665 = ( x77 & n27046 ) | ( x77 & ~n34664 ) | ( n27046 & ~n34664 ) ;
  assign n34666 = n12520 ^ n11499 ^ n4658 ;
  assign n34667 = n7703 ^ n5800 ^ n2222 ;
  assign n34668 = ( n4435 & n34666 ) | ( n4435 & ~n34667 ) | ( n34666 & ~n34667 ) ;
  assign n34669 = n34668 ^ n8329 ^ n8196 ;
  assign n34670 = n34665 | n34669 ;
  assign n34671 = ( n6594 & ~n15541 ) | ( n6594 & n34670 ) | ( ~n15541 & n34670 ) ;
  assign n34672 = n20913 ^ n7207 ^ n4034 ;
  assign n34673 = n34672 ^ n27206 ^ n12724 ;
  assign n34674 = ( n6822 & n26419 ) | ( n6822 & ~n34673 ) | ( n26419 & ~n34673 ) ;
  assign n34675 = n2556 & ~n27401 ;
  assign n34676 = n34675 ^ n352 ^ 1'b0 ;
  assign n34677 = n34676 ^ n33914 ^ n3772 ;
  assign n34678 = ~n2535 & n15022 ;
  assign n34679 = n22992 & n34678 ;
  assign n34680 = ( ~n17383 & n26927 ) | ( ~n17383 & n28424 ) | ( n26927 & n28424 ) ;
  assign n34681 = n18689 & n25594 ;
  assign n34682 = ( n3374 & n3468 ) | ( n3374 & ~n34634 ) | ( n3468 & ~n34634 ) ;
  assign n34683 = ( n21196 & ~n34681 ) | ( n21196 & n34682 ) | ( ~n34681 & n34682 ) ;
  assign n34684 = n32497 ^ n24013 ^ n22627 ;
  assign n34685 = ( n480 & n1442 ) | ( n480 & ~n9200 ) | ( n1442 & ~n9200 ) ;
  assign n34686 = n34685 ^ n22717 ^ n11915 ;
  assign n34687 = ( ~n3652 & n34684 ) | ( ~n3652 & n34686 ) | ( n34684 & n34686 ) ;
  assign n34688 = n30225 ^ n21183 ^ n19121 ;
  assign n34689 = n8467 ^ n5068 ^ 1'b0 ;
  assign n34690 = n34688 | n34689 ;
  assign n34691 = ( n6513 & ~n7802 ) | ( n6513 & n8915 ) | ( ~n7802 & n8915 ) ;
  assign n34692 = n16913 ^ n11446 ^ n11142 ;
  assign n34693 = n28250 ^ n12552 ^ n4677 ;
  assign n34694 = ( n34691 & ~n34692 ) | ( n34691 & n34693 ) | ( ~n34692 & n34693 ) ;
  assign n34695 = n7011 ^ n2774 ^ 1'b0 ;
  assign n34696 = n21341 ^ n11415 ^ 1'b0 ;
  assign n34697 = ( n2033 & n34695 ) | ( n2033 & ~n34696 ) | ( n34695 & ~n34696 ) ;
  assign n34699 = n19860 ^ n17524 ^ n5249 ;
  assign n34698 = n17832 ^ n14771 ^ n5467 ;
  assign n34700 = n34699 ^ n34698 ^ n17710 ;
  assign n34701 = n30918 ^ n29437 ^ n16911 ;
  assign n34702 = ( n1684 & n3746 ) | ( n1684 & n18008 ) | ( n3746 & n18008 ) ;
  assign n34703 = ( ~n9420 & n14467 ) | ( ~n9420 & n29908 ) | ( n14467 & n29908 ) ;
  assign n34704 = n34703 ^ n20040 ^ 1'b0 ;
  assign n34705 = n8083 | n27606 ;
  assign n34706 = n34705 ^ n19978 ^ 1'b0 ;
  assign n34707 = ( n1150 & ~n17947 ) | ( n1150 & n24386 ) | ( ~n17947 & n24386 ) ;
  assign n34708 = ( n17154 & n25965 ) | ( n17154 & n28770 ) | ( n25965 & n28770 ) ;
  assign n34709 = ( n1088 & n2661 ) | ( n1088 & n13360 ) | ( n2661 & n13360 ) ;
  assign n34710 = n21938 ^ n9742 ^ 1'b0 ;
  assign n34711 = ~n34709 & n34710 ;
  assign n34712 = n32530 ^ n28801 ^ n10939 ;
  assign n34713 = n34712 ^ n27982 ^ 1'b0 ;
  assign n34714 = ~n17377 & n25977 ;
  assign n34716 = n10887 | n28006 ;
  assign n34717 = n5931 | n34716 ;
  assign n34715 = n13572 ^ n9626 ^ n6643 ;
  assign n34718 = n34717 ^ n34715 ^ n14748 ;
  assign n34719 = ~n12136 & n17281 ;
  assign n34720 = n34719 ^ n15129 ^ 1'b0 ;
  assign n34721 = ( n371 & ~n13396 ) | ( n371 & n34720 ) | ( ~n13396 & n34720 ) ;
  assign n34722 = ( ~n9523 & n21356 ) | ( ~n9523 & n34721 ) | ( n21356 & n34721 ) ;
  assign n34723 = n34722 ^ n28409 ^ n27313 ;
  assign n34724 = n8542 | n33584 ;
  assign n34725 = n14894 & ~n34724 ;
  assign n34726 = n32600 ^ n4776 ^ 1'b0 ;
  assign n34727 = ( n24466 & n34352 ) | ( n24466 & ~n34726 ) | ( n34352 & ~n34726 ) ;
  assign n34728 = n9967 ^ n3469 ^ n1361 ;
  assign n34729 = n34728 ^ n17564 ^ n3097 ;
  assign n34730 = ( ~n4321 & n12493 ) | ( ~n4321 & n34729 ) | ( n12493 & n34729 ) ;
  assign n34731 = n32303 ^ n31110 ^ n461 ;
  assign n34734 = n10764 ^ n3544 ^ 1'b0 ;
  assign n34732 = n20443 ^ n1505 ^ 1'b0 ;
  assign n34733 = n8351 & ~n34732 ;
  assign n34735 = n34734 ^ n34733 ^ n19988 ;
  assign n34736 = n30801 ^ n22757 ^ n3404 ;
  assign n34737 = ( ~n643 & n33595 ) | ( ~n643 & n34736 ) | ( n33595 & n34736 ) ;
  assign n34738 = n22360 ^ n6398 ^ n6392 ;
  assign n34742 = x149 & n2745 ;
  assign n34739 = ~n11342 & n21446 ;
  assign n34740 = n34739 ^ n20728 ^ n17777 ;
  assign n34741 = ~n6973 & n34740 ;
  assign n34743 = n34742 ^ n34741 ^ n16762 ;
  assign n34744 = n15773 ^ n15171 ^ 1'b0 ;
  assign n34745 = ~n2399 & n34744 ;
  assign n34746 = n34745 ^ n2061 ^ 1'b0 ;
  assign n34747 = n34743 & n34746 ;
  assign n34748 = n24492 ^ n13096 ^ n1754 ;
  assign n34749 = ( n1892 & n20466 ) | ( n1892 & n33731 ) | ( n20466 & n33731 ) ;
  assign n34750 = n5522 & ~n34749 ;
  assign n34751 = n19631 & n34750 ;
  assign n34752 = n34748 | n34751 ;
  assign n34753 = x205 & n3508 ;
  assign n34754 = n9728 & n34753 ;
  assign n34755 = n34754 ^ n5663 ^ n4381 ;
  assign n34756 = ( n17653 & n32742 ) | ( n17653 & ~n34755 ) | ( n32742 & ~n34755 ) ;
  assign n34757 = n14064 ^ n5502 ^ n5160 ;
  assign n34758 = n34757 ^ n884 ^ n490 ;
  assign n34759 = n32548 ^ n23500 ^ n3872 ;
  assign n34760 = n28948 ^ n26273 ^ n24184 ;
  assign n34761 = ( n18125 & n34759 ) | ( n18125 & ~n34760 ) | ( n34759 & ~n34760 ) ;
  assign n34762 = ( n31115 & n34758 ) | ( n31115 & n34761 ) | ( n34758 & n34761 ) ;
  assign n34763 = n7439 & n7892 ;
  assign n34764 = n13017 & n34763 ;
  assign n34765 = ( n2690 & n4965 ) | ( n2690 & n29665 ) | ( n4965 & n29665 ) ;
  assign n34766 = n3916 & n34765 ;
  assign n34767 = n34766 ^ n2785 ^ 1'b0 ;
  assign n34768 = n3007 ^ n2725 ^ n1197 ;
  assign n34769 = ( n24904 & n27360 ) | ( n24904 & ~n34768 ) | ( n27360 & ~n34768 ) ;
  assign n34770 = n21670 ^ n10034 ^ n2020 ;
  assign n34771 = n27744 ^ n20532 ^ n1818 ;
  assign n34772 = ( n5870 & n34770 ) | ( n5870 & ~n34771 ) | ( n34770 & ~n34771 ) ;
  assign n34773 = n9134 ^ n1883 ^ n1537 ;
  assign n34774 = n13905 ^ n8141 ^ 1'b0 ;
  assign n34775 = n34773 & ~n34774 ;
  assign n34776 = ( n7906 & n18217 ) | ( n7906 & ~n34775 ) | ( n18217 & ~n34775 ) ;
  assign n34777 = ( n851 & ~n26539 ) | ( n851 & n34776 ) | ( ~n26539 & n34776 ) ;
  assign n34778 = n19625 ^ n9710 ^ n1175 ;
  assign n34779 = n30262 & ~n34778 ;
  assign n34780 = n34779 ^ n22580 ^ 1'b0 ;
  assign n34781 = n8300 & n18621 ;
  assign n34782 = n21017 ^ n16094 ^ n2814 ;
  assign n34784 = ( n11492 & n16448 ) | ( n11492 & ~n22554 ) | ( n16448 & ~n22554 ) ;
  assign n34785 = n34784 ^ n22753 ^ n12747 ;
  assign n34786 = n34785 ^ n16619 ^ n2925 ;
  assign n34787 = n13061 ^ n4717 ^ 1'b0 ;
  assign n34788 = n34786 | n34787 ;
  assign n34783 = n7984 & n31626 ;
  assign n34789 = n34788 ^ n34783 ^ 1'b0 ;
  assign n34790 = n29100 ^ n19121 ^ n3490 ;
  assign n34791 = n26192 ^ n11689 ^ n4986 ;
  assign n34792 = ( n4275 & n6099 ) | ( n4275 & ~n34791 ) | ( n6099 & ~n34791 ) ;
  assign n34793 = ( n28235 & n34790 ) | ( n28235 & n34792 ) | ( n34790 & n34792 ) ;
  assign n34794 = n19977 ^ n11225 ^ n6288 ;
  assign n34795 = ( ~n31253 & n33214 ) | ( ~n31253 & n34794 ) | ( n33214 & n34794 ) ;
  assign n34798 = ( n2842 & n8107 ) | ( n2842 & ~n11180 ) | ( n8107 & ~n11180 ) ;
  assign n34797 = n19540 ^ n704 ^ x162 ;
  assign n34796 = ( n10605 & n13762 ) | ( n10605 & ~n23526 ) | ( n13762 & ~n23526 ) ;
  assign n34799 = n34798 ^ n34797 ^ n34796 ;
  assign n34800 = ( n379 & ~n8530 ) | ( n379 & n21150 ) | ( ~n8530 & n21150 ) ;
  assign n34801 = n6243 & n34800 ;
  assign n34802 = n6162 & n34801 ;
  assign n34803 = ( n19065 & n24178 ) | ( n19065 & n34802 ) | ( n24178 & n34802 ) ;
  assign n34804 = n1917 & ~n23080 ;
  assign n34805 = ~n7447 & n34804 ;
  assign n34806 = n5115 | n34805 ;
  assign n34807 = n24270 | n34806 ;
  assign n34808 = ( n5927 & ~n9707 ) | ( n5927 & n34807 ) | ( ~n9707 & n34807 ) ;
  assign n34809 = ( ~n3768 & n27349 ) | ( ~n3768 & n30368 ) | ( n27349 & n30368 ) ;
  assign n34810 = n5573 ^ n3768 ^ n3762 ;
  assign n34811 = ~n16020 & n34810 ;
  assign n34812 = ( n2395 & n10738 ) | ( n2395 & n21243 ) | ( n10738 & n21243 ) ;
  assign n34813 = n11503 ^ n5932 ^ n3901 ;
  assign n34814 = ( n1784 & ~n34812 ) | ( n1784 & n34813 ) | ( ~n34812 & n34813 ) ;
  assign n34815 = n26239 ^ n10566 ^ 1'b0 ;
  assign n34816 = n28740 ^ n22275 ^ n10190 ;
  assign n34817 = n34816 ^ n25391 ^ 1'b0 ;
  assign n34818 = ~n34815 & n34817 ;
  assign n34819 = n8246 ^ n8220 ^ 1'b0 ;
  assign n34820 = n19340 ^ n7582 ^ n7404 ;
  assign n34821 = n1319 | n13078 ;
  assign n34822 = n33932 ^ n31229 ^ n10302 ;
  assign n34825 = n12009 ^ n6292 ^ n2535 ;
  assign n34826 = n34825 ^ n21808 ^ n21179 ;
  assign n34823 = n13760 & n28057 ;
  assign n34824 = ~n25549 & n34823 ;
  assign n34827 = n34826 ^ n34824 ^ n717 ;
  assign n34828 = n34827 ^ n2978 ^ 1'b0 ;
  assign n34829 = n28196 ^ n17564 ^ n2714 ;
  assign n34830 = n34829 ^ n15726 ^ 1'b0 ;
  assign n34831 = n287 & ~n34830 ;
  assign n34832 = n13435 ^ n12394 ^ n8784 ;
  assign n34833 = n34832 ^ n8084 ^ 1'b0 ;
  assign n34834 = n9263 ^ n5164 ^ n3375 ;
  assign n34835 = n34834 ^ n22802 ^ n9134 ;
  assign n34836 = n8914 ^ n7252 ^ n5168 ;
  assign n34837 = ( n559 & n33038 ) | ( n559 & ~n34836 ) | ( n33038 & ~n34836 ) ;
  assign n34838 = ( ~n1433 & n16548 ) | ( ~n1433 & n23682 ) | ( n16548 & n23682 ) ;
  assign n34839 = ( ~n12616 & n22132 ) | ( ~n12616 & n34838 ) | ( n22132 & n34838 ) ;
  assign n34840 = n8605 | n34839 ;
  assign n34841 = ( n17026 & n20563 ) | ( n17026 & n25425 ) | ( n20563 & n25425 ) ;
  assign n34842 = n25866 ^ n7748 ^ 1'b0 ;
  assign n34843 = n34841 | n34842 ;
  assign n34844 = ( ~n4740 & n16658 ) | ( ~n4740 & n34843 ) | ( n16658 & n34843 ) ;
  assign n34848 = ( n334 & n19514 ) | ( n334 & ~n20924 ) | ( n19514 & ~n20924 ) ;
  assign n34849 = n5344 & ~n34848 ;
  assign n34850 = ~n17829 & n34849 ;
  assign n34845 = n10782 ^ n10535 ^ n5064 ;
  assign n34846 = n7212 | n34845 ;
  assign n34847 = n4350 | n34846 ;
  assign n34851 = n34850 ^ n34847 ^ 1'b0 ;
  assign n34852 = n34844 & ~n34851 ;
  assign n34854 = n18637 | n20532 ;
  assign n34855 = n34854 ^ n33695 ^ n12277 ;
  assign n34853 = n20535 ^ n4113 ^ x223 ;
  assign n34856 = n34855 ^ n34853 ^ n6770 ;
  assign n34857 = ( ~n4142 & n12577 ) | ( ~n4142 & n13469 ) | ( n12577 & n13469 ) ;
  assign n34858 = n24468 ^ n22790 ^ 1'b0 ;
  assign n34859 = n34858 ^ n23178 ^ n511 ;
  assign n34860 = ( n6013 & ~n19782 ) | ( n6013 & n27574 ) | ( ~n19782 & n27574 ) ;
  assign n34861 = n34860 ^ n19131 ^ n18221 ;
  assign n34862 = n25893 ^ n14989 ^ n11163 ;
  assign n34863 = ( ~n10049 & n34861 ) | ( ~n10049 & n34862 ) | ( n34861 & n34862 ) ;
  assign n34864 = ( ~n819 & n7637 ) | ( ~n819 & n31683 ) | ( n7637 & n31683 ) ;
  assign n34865 = n34444 ^ n332 ^ 1'b0 ;
  assign n34866 = n24288 & n34865 ;
  assign n34867 = n1615 & n6887 ;
  assign n34868 = n34867 ^ n28538 ^ 1'b0 ;
  assign n34869 = n13957 ^ n13765 ^ n9542 ;
  assign n34870 = ( n2270 & n13124 ) | ( n2270 & ~n34869 ) | ( n13124 & ~n34869 ) ;
  assign n34871 = ( ~n3950 & n4585 ) | ( ~n3950 & n27494 ) | ( n4585 & n27494 ) ;
  assign n34872 = ( n13229 & n25558 ) | ( n13229 & ~n27293 ) | ( n25558 & ~n27293 ) ;
  assign n34873 = ( n24953 & ~n31120 ) | ( n24953 & n34872 ) | ( ~n31120 & n34872 ) ;
  assign n34874 = ( n7770 & n8701 ) | ( n7770 & ~n28208 ) | ( n8701 & ~n28208 ) ;
  assign n34875 = n34874 ^ n31746 ^ n31280 ;
  assign n34876 = n34875 ^ n20837 ^ 1'b0 ;
  assign n34877 = n18734 ^ n11657 ^ n10085 ;
  assign n34878 = ( n27135 & n29453 ) | ( n27135 & ~n34877 ) | ( n29453 & ~n34877 ) ;
  assign n34879 = n22290 ^ n18373 ^ n11510 ;
  assign n34880 = n34879 ^ n11365 ^ n3717 ;
  assign n34889 = n22560 ^ n10075 ^ n5306 ;
  assign n34886 = n7040 ^ n2795 ^ 1'b0 ;
  assign n34887 = n1612 & ~n34886 ;
  assign n34888 = ( n21465 & ~n32476 ) | ( n21465 & n34887 ) | ( ~n32476 & n34887 ) ;
  assign n34884 = n22941 ^ n21809 ^ n10347 ;
  assign n34881 = n21105 ^ n5715 ^ 1'b0 ;
  assign n34882 = ( ~n8673 & n17278 ) | ( ~n8673 & n34881 ) | ( n17278 & n34881 ) ;
  assign n34883 = n34882 ^ n26874 ^ n9074 ;
  assign n34885 = n34884 ^ n34883 ^ n21856 ;
  assign n34890 = n34889 ^ n34888 ^ n34885 ;
  assign n34891 = n27240 ^ n23026 ^ n11245 ;
  assign n34894 = ( n8261 & ~n16571 ) | ( n8261 & n22380 ) | ( ~n16571 & n22380 ) ;
  assign n34892 = n33218 ^ n19621 ^ 1'b0 ;
  assign n34893 = n10337 & n34892 ;
  assign n34895 = n34894 ^ n34893 ^ n8868 ;
  assign n34896 = n23292 ^ n7531 ^ n6106 ;
  assign n34897 = n34896 ^ n33546 ^ n7751 ;
  assign n34898 = ( n7397 & n7807 ) | ( n7397 & n12558 ) | ( n7807 & n12558 ) ;
  assign n34899 = ( n4140 & n11005 ) | ( n4140 & ~n12871 ) | ( n11005 & ~n12871 ) ;
  assign n34900 = n4154 & ~n6637 ;
  assign n34901 = n6769 & n34900 ;
  assign n34902 = n7262 | n34901 ;
  assign n34903 = n23480 ^ n7611 ^ x103 ;
  assign n34904 = ( ~n1963 & n34399 ) | ( ~n1963 & n34903 ) | ( n34399 & n34903 ) ;
  assign n34905 = n20418 ^ n17260 ^ n12585 ;
  assign n34906 = n499 & ~n34905 ;
  assign n34907 = n18760 ^ n10977 ^ 1'b0 ;
  assign n34908 = ( n19836 & n22363 ) | ( n19836 & n34907 ) | ( n22363 & n34907 ) ;
  assign n34909 = ~n16043 & n17371 ;
  assign n34910 = n34909 ^ n23399 ^ n9894 ;
  assign n34911 = n34910 ^ n9787 ^ n3091 ;
  assign n34912 = n34441 ^ n9823 ^ n5093 ;
  assign n34913 = ( n4649 & n7947 ) | ( n4649 & n14961 ) | ( n7947 & n14961 ) ;
  assign n34914 = n34913 ^ n15811 ^ n4791 ;
  assign n34915 = n34914 ^ n7447 ^ 1'b0 ;
  assign n34916 = ~n16299 & n34915 ;
  assign n34917 = n34916 ^ n23514 ^ n7680 ;
  assign n34918 = n34917 ^ n29176 ^ n3900 ;
  assign n34919 = ( n11764 & n34912 ) | ( n11764 & ~n34918 ) | ( n34912 & ~n34918 ) ;
  assign n34921 = n30921 ^ n27690 ^ n300 ;
  assign n34920 = n16512 & ~n18015 ;
  assign n34922 = n34921 ^ n34920 ^ 1'b0 ;
  assign n34923 = ( x164 & n987 ) | ( x164 & ~n19501 ) | ( n987 & ~n19501 ) ;
  assign n34924 = ~n1094 & n13928 ;
  assign n34925 = ~n34923 & n34924 ;
  assign n34926 = n11566 ^ n11354 ^ n10878 ;
  assign n34930 = ( ~n1710 & n18457 ) | ( ~n1710 & n21131 ) | ( n18457 & n21131 ) ;
  assign n34928 = n32679 ^ n27857 ^ n20106 ;
  assign n34927 = n2174 & ~n6686 ;
  assign n34929 = n34928 ^ n34927 ^ 1'b0 ;
  assign n34931 = n34930 ^ n34929 ^ n33331 ;
  assign n34932 = n18854 ^ n11734 ^ n5411 ;
  assign n34933 = ( n17054 & n21138 ) | ( n17054 & n23552 ) | ( n21138 & n23552 ) ;
  assign n34934 = ( ~n18464 & n23703 ) | ( ~n18464 & n34933 ) | ( n23703 & n34933 ) ;
  assign n34935 = ( ~n4444 & n9180 ) | ( ~n4444 & n10263 ) | ( n9180 & n10263 ) ;
  assign n34936 = n34022 ^ n31347 ^ n9233 ;
  assign n34937 = n20562 ^ n5912 ^ n4334 ;
  assign n34938 = ( n34935 & ~n34936 ) | ( n34935 & n34937 ) | ( ~n34936 & n34937 ) ;
  assign n34939 = n33902 ^ n29056 ^ n21314 ;
  assign n34940 = n34939 ^ n32641 ^ n6690 ;
  assign n34943 = ( ~n964 & n7733 ) | ( ~n964 & n10070 ) | ( n7733 & n10070 ) ;
  assign n34944 = n34943 ^ n32265 ^ n8808 ;
  assign n34941 = n5165 | n8767 ;
  assign n34942 = ( ~n2534 & n20576 ) | ( ~n2534 & n34941 ) | ( n20576 & n34941 ) ;
  assign n34945 = n34944 ^ n34942 ^ n3888 ;
  assign n34948 = ( ~n2536 & n6187 ) | ( ~n2536 & n28877 ) | ( n6187 & n28877 ) ;
  assign n34946 = n16208 ^ n4258 ^ n3180 ;
  assign n34947 = ( ~n8829 & n32969 ) | ( ~n8829 & n34946 ) | ( n32969 & n34946 ) ;
  assign n34949 = n34948 ^ n34947 ^ n12980 ;
  assign n34950 = n34949 ^ n17723 ^ 1'b0 ;
  assign n34951 = n30075 ^ n26263 ^ n8882 ;
  assign n34952 = n20347 ^ n15878 ^ n4709 ;
  assign n34953 = ( n19952 & n21076 ) | ( n19952 & n34952 ) | ( n21076 & n34952 ) ;
  assign n34956 = n17077 ^ n15581 ^ n5916 ;
  assign n34957 = n34956 ^ n21646 ^ 1'b0 ;
  assign n34954 = n16915 | n29666 ;
  assign n34955 = n9723 & ~n34954 ;
  assign n34958 = n34957 ^ n34955 ^ 1'b0 ;
  assign n34959 = n23187 ^ n22891 ^ n6479 ;
  assign n34960 = n27860 ^ n12086 ^ n2826 ;
  assign n34961 = ( ~n2278 & n30956 ) | ( ~n2278 & n34960 ) | ( n30956 & n34960 ) ;
  assign n34963 = n27975 ^ n15395 ^ n13330 ;
  assign n34962 = ( n5644 & n23215 ) | ( n5644 & n27357 ) | ( n23215 & n27357 ) ;
  assign n34964 = n34963 ^ n34962 ^ n14245 ;
  assign n34965 = ~n20105 & n27383 ;
  assign n34966 = ( n8363 & n23603 ) | ( n8363 & n34965 ) | ( n23603 & n34965 ) ;
  assign n34967 = n27637 ^ n16035 ^ n6851 ;
  assign n34968 = ( n5512 & n7667 ) | ( n5512 & n17710 ) | ( n7667 & n17710 ) ;
  assign n34969 = n34968 ^ n12001 ^ 1'b0 ;
  assign n34970 = ( n17541 & n18439 ) | ( n17541 & n34969 ) | ( n18439 & n34969 ) ;
  assign n34971 = n27759 ^ n7253 ^ n4839 ;
  assign n34972 = ( ~n2272 & n3037 ) | ( ~n2272 & n34971 ) | ( n3037 & n34971 ) ;
  assign n34973 = ( n23259 & n26072 ) | ( n23259 & ~n34972 ) | ( n26072 & ~n34972 ) ;
  assign n34974 = n34973 ^ n27308 ^ n2420 ;
  assign n34975 = ( n3424 & ~n4693 ) | ( n3424 & n16161 ) | ( ~n4693 & n16161 ) ;
  assign n34976 = n34975 ^ n11177 ^ n6363 ;
  assign n34977 = n23875 ^ n18218 ^ 1'b0 ;
  assign n34978 = n1489 & ~n34977 ;
  assign n34979 = ( n8161 & n9006 ) | ( n8161 & n26726 ) | ( n9006 & n26726 ) ;
  assign n34980 = n13548 | n34979 ;
  assign n34981 = ( ~n6061 & n11259 ) | ( ~n6061 & n18561 ) | ( n11259 & n18561 ) ;
  assign n34982 = n34981 ^ n25638 ^ n17567 ;
  assign n34983 = n20542 ^ n7815 ^ n1947 ;
  assign n34990 = ( n2850 & n4600 ) | ( n2850 & ~n17530 ) | ( n4600 & ~n17530 ) ;
  assign n34987 = ~n1247 & n1927 ;
  assign n34988 = n8716 & n34987 ;
  assign n34984 = n5956 ^ n5147 ^ n2375 ;
  assign n34985 = n20533 ^ n10381 ^ n3279 ;
  assign n34986 = ( n3173 & n34984 ) | ( n3173 & ~n34985 ) | ( n34984 & ~n34985 ) ;
  assign n34989 = n34988 ^ n34986 ^ n33123 ;
  assign n34991 = n34990 ^ n34989 ^ n27328 ;
  assign n34992 = n34991 ^ n25458 ^ n12213 ;
  assign n34996 = n922 | n2049 ;
  assign n34997 = n9233 & ~n34996 ;
  assign n34998 = n34997 ^ n17710 ^ 1'b0 ;
  assign n34994 = n13736 ^ n3561 ^ n1511 ;
  assign n34993 = ( ~n9927 & n19858 ) | ( ~n9927 & n22974 ) | ( n19858 & n22974 ) ;
  assign n34995 = n34994 ^ n34993 ^ n6643 ;
  assign n34999 = n34998 ^ n34995 ^ n22912 ;
  assign n35000 = n32941 ^ n21553 ^ n6136 ;
  assign n35001 = ( ~n21132 & n21589 ) | ( ~n21132 & n22731 ) | ( n21589 & n22731 ) ;
  assign n35002 = n1337 & n15555 ;
  assign n35003 = ~n35001 & n35002 ;
  assign n35004 = ( n464 & n3969 ) | ( n464 & n35003 ) | ( n3969 & n35003 ) ;
  assign n35005 = ( ~n4794 & n35000 ) | ( ~n4794 & n35004 ) | ( n35000 & n35004 ) ;
  assign n35006 = n28639 ^ n2730 ^ n606 ;
  assign n35007 = ( n1428 & n3409 ) | ( n1428 & n35006 ) | ( n3409 & n35006 ) ;
  assign n35008 = n22414 ^ n16258 ^ x64 ;
  assign n35009 = ( x216 & n22649 ) | ( x216 & n27117 ) | ( n22649 & n27117 ) ;
  assign n35010 = ( n16216 & n31151 ) | ( n16216 & ~n32237 ) | ( n31151 & ~n32237 ) ;
  assign n35011 = ( n3044 & n30895 ) | ( n3044 & n35010 ) | ( n30895 & n35010 ) ;
  assign n35012 = ( ~n2801 & n3591 ) | ( ~n2801 & n4464 ) | ( n3591 & n4464 ) ;
  assign n35013 = n28137 ^ n982 ^ 1'b0 ;
  assign n35014 = n35012 & n35013 ;
  assign n35016 = n16219 ^ n16066 ^ n9806 ;
  assign n35015 = n5713 & n28326 ;
  assign n35017 = n35016 ^ n35015 ^ 1'b0 ;
  assign n35018 = ( n9716 & ~n23512 ) | ( n9716 & n28522 ) | ( ~n23512 & n28522 ) ;
  assign n35019 = n25222 ^ n4720 ^ 1'b0 ;
  assign n35020 = ( n2113 & ~n3072 ) | ( n2113 & n15800 ) | ( ~n3072 & n15800 ) ;
  assign n35021 = ( n5774 & n35019 ) | ( n5774 & ~n35020 ) | ( n35019 & ~n35020 ) ;
  assign n35022 = n35021 ^ n23752 ^ n12946 ;
  assign n35023 = ( n991 & n28536 ) | ( n991 & ~n31853 ) | ( n28536 & ~n31853 ) ;
  assign n35024 = n31368 ^ n29587 ^ n4096 ;
  assign n35025 = ( n4096 & n10098 ) | ( n4096 & ~n16712 ) | ( n10098 & ~n16712 ) ;
  assign n35031 = ( n6356 & n13831 ) | ( n6356 & ~n33371 ) | ( n13831 & ~n33371 ) ;
  assign n35026 = n19031 ^ n6756 ^ n6702 ;
  assign n35027 = n11154 ^ n8053 ^ n5738 ;
  assign n35028 = ( n1246 & n17551 ) | ( n1246 & n35027 ) | ( n17551 & n35027 ) ;
  assign n35029 = ( n14134 & ~n35026 ) | ( n14134 & n35028 ) | ( ~n35026 & n35028 ) ;
  assign n35030 = ~n8194 & n35029 ;
  assign n35032 = n35031 ^ n35030 ^ n18150 ;
  assign n35033 = n18143 ^ n14096 ^ n12594 ;
  assign n35034 = ( n3607 & n18524 ) | ( n3607 & ~n23475 ) | ( n18524 & ~n23475 ) ;
  assign n35035 = ( n34263 & ~n35033 ) | ( n34263 & n35034 ) | ( ~n35033 & n35034 ) ;
  assign n35036 = n26409 & ~n31445 ;
  assign n35037 = ( n5783 & n32745 ) | ( n5783 & ~n35036 ) | ( n32745 & ~n35036 ) ;
  assign n35038 = n18084 ^ n16320 ^ 1'b0 ;
  assign n35039 = n11985 | n35038 ;
  assign n35040 = n35039 ^ n16418 ^ n6776 ;
  assign n35041 = n35040 ^ n31690 ^ n17237 ;
  assign n35044 = n7870 ^ n6605 ^ n3693 ;
  assign n35042 = n32926 ^ n18749 ^ 1'b0 ;
  assign n35043 = n28107 | n35042 ;
  assign n35045 = n35044 ^ n35043 ^ n1418 ;
  assign n35046 = n35045 ^ n22476 ^ n2634 ;
  assign n35047 = n12535 ^ n11606 ^ n10147 ;
  assign n35048 = n35047 ^ n2954 ^ 1'b0 ;
  assign n35049 = n24418 & ~n35048 ;
  assign n35050 = n31424 ^ n30590 ^ n5997 ;
  assign n35051 = n9978 ^ n6924 ^ 1'b0 ;
  assign n35052 = ~n3125 & n26064 ;
  assign n35053 = n35052 ^ n14558 ^ 1'b0 ;
  assign n35054 = ( n4056 & ~n4700 ) | ( n4056 & n11716 ) | ( ~n4700 & n11716 ) ;
  assign n35055 = ( ~n17168 & n22649 ) | ( ~n17168 & n35054 ) | ( n22649 & n35054 ) ;
  assign n35056 = n19321 ^ n10903 ^ n8903 ;
  assign n35057 = n30503 ^ n13477 ^ 1'b0 ;
  assign n35058 = n26245 & ~n35057 ;
  assign n35059 = n4184 | n8554 ;
  assign n35060 = ( ~n5631 & n31985 ) | ( ~n5631 & n35059 ) | ( n31985 & n35059 ) ;
  assign n35061 = ( ~n3976 & n19381 ) | ( ~n3976 & n35060 ) | ( n19381 & n35060 ) ;
  assign n35062 = n7790 & n30895 ;
  assign n35063 = ( n589 & n12662 ) | ( n589 & n35062 ) | ( n12662 & n35062 ) ;
  assign n35064 = ( n6952 & ~n31642 ) | ( n6952 & n35063 ) | ( ~n31642 & n35063 ) ;
  assign n35065 = n10781 ^ n8665 ^ n400 ;
  assign n35066 = ( n9655 & n23225 ) | ( n9655 & ~n33981 ) | ( n23225 & ~n33981 ) ;
  assign n35067 = ( n31617 & ~n35065 ) | ( n31617 & n35066 ) | ( ~n35065 & n35066 ) ;
  assign n35068 = n28432 ^ n17333 ^ n2778 ;
  assign n35069 = ( ~n9493 & n13429 ) | ( ~n9493 & n23353 ) | ( n13429 & n23353 ) ;
  assign n35070 = n35069 ^ n22142 ^ n15917 ;
  assign n35071 = n35070 ^ n8369 ^ n7333 ;
  assign n35072 = ( n1205 & n7320 ) | ( n1205 & ~n35071 ) | ( n7320 & ~n35071 ) ;
  assign n35073 = ( n14776 & n15779 ) | ( n14776 & ~n17715 ) | ( n15779 & ~n17715 ) ;
  assign n35074 = ( n11014 & n13868 ) | ( n11014 & ~n35073 ) | ( n13868 & ~n35073 ) ;
  assign n35075 = n16726 & n29612 ;
  assign n35076 = n35075 ^ n14695 ^ n12268 ;
  assign n35077 = ( n15376 & ~n22618 ) | ( n15376 & n27437 ) | ( ~n22618 & n27437 ) ;
  assign n35078 = n35077 ^ n31070 ^ n4344 ;
  assign n35079 = ( n4633 & n6385 ) | ( n4633 & ~n22415 ) | ( n6385 & ~n22415 ) ;
  assign n35080 = n35079 ^ n27110 ^ n5795 ;
  assign n35081 = ( n261 & ~n3018 ) | ( n261 & n34802 ) | ( ~n3018 & n34802 ) ;
  assign n35082 = n16801 | n23446 ;
  assign n35083 = n35082 ^ n12708 ^ 1'b0 ;
  assign n35084 = n5740 & ~n31256 ;
  assign n35085 = n4483 ^ n898 ^ 1'b0 ;
  assign n35086 = n35085 ^ n21374 ^ n6067 ;
  assign n35087 = n6390 | n35086 ;
  assign n35088 = n35084 & ~n35087 ;
  assign n35089 = n19635 ^ n9650 ^ n1950 ;
  assign n35090 = n5494 ^ n1313 ^ 1'b0 ;
  assign n35091 = ( n30469 & n32147 ) | ( n30469 & n35090 ) | ( n32147 & n35090 ) ;
  assign n35094 = ( n12673 & n14046 ) | ( n12673 & ~n22568 ) | ( n14046 & ~n22568 ) ;
  assign n35092 = n4928 & ~n10409 ;
  assign n35093 = n35092 ^ n4123 ^ 1'b0 ;
  assign n35095 = n35094 ^ n35093 ^ n34963 ;
  assign n35096 = n34155 ^ n20865 ^ 1'b0 ;
  assign n35097 = ~n31374 & n35096 ;
  assign n35098 = ( n4222 & ~n29368 ) | ( n4222 & n35097 ) | ( ~n29368 & n35097 ) ;
  assign n35099 = ( n5452 & ~n15391 ) | ( n5452 & n23178 ) | ( ~n15391 & n23178 ) ;
  assign n35100 = n35099 ^ n20542 ^ n1504 ;
  assign n35101 = n35100 ^ n4780 ^ 1'b0 ;
  assign n35102 = n13189 ^ n9360 ^ 1'b0 ;
  assign n35103 = n20877 & n35102 ;
  assign n35104 = ( n15330 & n18438 ) | ( n15330 & n23477 ) | ( n18438 & n23477 ) ;
  assign n35105 = ( n5596 & ~n14654 ) | ( n5596 & n22498 ) | ( ~n14654 & n22498 ) ;
  assign n35106 = n24865 ^ n21805 ^ n17484 ;
  assign n35107 = n35106 ^ n5688 ^ 1'b0 ;
  assign n35108 = n25597 & n35107 ;
  assign n35109 = n35108 ^ n20578 ^ n3131 ;
  assign n35110 = ( n35104 & n35105 ) | ( n35104 & n35109 ) | ( n35105 & n35109 ) ;
  assign n35111 = n13574 ^ n9523 ^ n1150 ;
  assign n35112 = n35111 ^ n10667 ^ n7434 ;
  assign n35113 = n35112 ^ n14032 ^ x127 ;
  assign n35114 = n25563 ^ n21154 ^ n7552 ;
  assign n35115 = ~n9668 & n12499 ;
  assign n35116 = ~n5739 & n35115 ;
  assign n35117 = n35116 ^ n11411 ^ n690 ;
  assign n35118 = n1073 | n9998 ;
  assign n35119 = n19263 ^ n3493 ^ 1'b0 ;
  assign n35120 = n27408 | n35119 ;
  assign n35121 = ( ~n15792 & n17682 ) | ( ~n15792 & n24613 ) | ( n17682 & n24613 ) ;
  assign n35122 = ( ~n12179 & n28445 ) | ( ~n12179 & n35121 ) | ( n28445 & n35121 ) ;
  assign n35123 = n35122 ^ n7715 ^ n4571 ;
  assign n35124 = n35123 ^ n24983 ^ n10220 ;
  assign n35125 = ( n854 & ~n2397 ) | ( n854 & n22113 ) | ( ~n2397 & n22113 ) ;
  assign n35126 = n24528 ^ n6559 ^ 1'b0 ;
  assign n35127 = n35126 ^ n5594 ^ n4288 ;
  assign n35128 = ( x93 & n7805 ) | ( x93 & ~n10187 ) | ( n7805 & ~n10187 ) ;
  assign n35129 = n35128 ^ n33022 ^ n8050 ;
  assign n35130 = n2563 & n3049 ;
  assign n35131 = n35130 ^ n17781 ^ n2922 ;
  assign n35132 = n21142 ^ n20286 ^ n11233 ;
  assign n35133 = ( ~n1165 & n24074 ) | ( ~n1165 & n35132 ) | ( n24074 & n35132 ) ;
  assign n35134 = ( x88 & ~n21535 ) | ( x88 & n34039 ) | ( ~n21535 & n34039 ) ;
  assign n35135 = ( n2199 & n15475 ) | ( n2199 & n35134 ) | ( n15475 & n35134 ) ;
  assign n35136 = n35135 ^ n17611 ^ 1'b0 ;
  assign n35137 = n35136 ^ n32295 ^ n4638 ;
  assign n35138 = n35137 ^ n30306 ^ n6327 ;
  assign n35139 = ( n10848 & ~n16359 ) | ( n10848 & n35138 ) | ( ~n16359 & n35138 ) ;
  assign n35140 = n7067 & ~n21357 ;
  assign n35141 = n35140 ^ n23326 ^ 1'b0 ;
  assign n35142 = n30730 ^ n18608 ^ 1'b0 ;
  assign n35143 = n35142 ^ n22446 ^ n12355 ;
  assign n35144 = ( n4197 & n7892 ) | ( n4197 & ~n8995 ) | ( n7892 & ~n8995 ) ;
  assign n35145 = ( n1869 & n4248 ) | ( n1869 & n10267 ) | ( n4248 & n10267 ) ;
  assign n35146 = ( n4637 & ~n5900 ) | ( n4637 & n35145 ) | ( ~n5900 & n35145 ) ;
  assign n35147 = ( n31751 & ~n35144 ) | ( n31751 & n35146 ) | ( ~n35144 & n35146 ) ;
  assign n35148 = n4586 ^ x128 ^ 1'b0 ;
  assign n35149 = n34807 ^ n23113 ^ n20700 ;
  assign n35150 = ( ~n5647 & n16514 ) | ( ~n5647 & n19530 ) | ( n16514 & n19530 ) ;
  assign n35151 = n1094 | n1158 ;
  assign n35152 = n17899 | n35151 ;
  assign n35153 = ( n2220 & n5782 ) | ( n2220 & ~n12816 ) | ( n5782 & ~n12816 ) ;
  assign n35154 = n35153 ^ n33064 ^ n3449 ;
  assign n35155 = n15765 ^ n10643 ^ 1'b0 ;
  assign n35156 = n1287 & ~n35155 ;
  assign n35157 = n35156 ^ n22554 ^ n16286 ;
  assign n35158 = n35157 ^ n30820 ^ n26326 ;
  assign n35159 = n15221 ^ n11703 ^ n8106 ;
  assign n35160 = ~n12677 & n24301 ;
  assign n35161 = n35160 ^ n14193 ^ 1'b0 ;
  assign n35162 = n35161 ^ n28331 ^ 1'b0 ;
  assign n35163 = ( n2433 & n5990 ) | ( n2433 & ~n6897 ) | ( n5990 & ~n6897 ) ;
  assign n35164 = ( n4587 & n17697 ) | ( n4587 & ~n21790 ) | ( n17697 & ~n21790 ) ;
  assign n35165 = n19565 ^ n11346 ^ n6118 ;
  assign n35166 = n4777 ^ n4553 ^ 1'b0 ;
  assign n35167 = n14233 | n35166 ;
  assign n35168 = ( ~n22431 & n35165 ) | ( ~n22431 & n35167 ) | ( n35165 & n35167 ) ;
  assign n35169 = n35168 ^ n28478 ^ 1'b0 ;
  assign n35170 = n35164 & ~n35169 ;
  assign n35171 = ( n23003 & n35163 ) | ( n23003 & n35170 ) | ( n35163 & n35170 ) ;
  assign n35172 = n26414 ^ n24711 ^ n5609 ;
  assign n35173 = ( n16034 & n29333 ) | ( n16034 & n30593 ) | ( n29333 & n30593 ) ;
  assign n35174 = n23692 ^ n21753 ^ 1'b0 ;
  assign n35175 = ~n20820 & n23884 ;
  assign n35176 = ~x31 & n35175 ;
  assign n35177 = n3369 & ~n4265 ;
  assign n35178 = ( n4600 & ~n8067 ) | ( n4600 & n35177 ) | ( ~n8067 & n35177 ) ;
  assign n35179 = n30340 | n33284 ;
  assign n35180 = n35179 ^ n1220 ^ 1'b0 ;
  assign n35181 = ( n20756 & ~n25750 ) | ( n20756 & n35180 ) | ( ~n25750 & n35180 ) ;
  assign n35182 = n34080 ^ n31495 ^ n12561 ;
  assign n35183 = n4894 ^ x40 ^ 1'b0 ;
  assign n35184 = ~n15279 & n35183 ;
  assign n35185 = ( n10835 & ~n35182 ) | ( n10835 & n35184 ) | ( ~n35182 & n35184 ) ;
  assign n35188 = n5685 ^ n1577 ^ 1'b0 ;
  assign n35186 = ( n1738 & ~n6462 ) | ( n1738 & n22972 ) | ( ~n6462 & n22972 ) ;
  assign n35187 = n35186 ^ n23121 ^ n13827 ;
  assign n35189 = n35188 ^ n35187 ^ n9534 ;
  assign n35190 = ( n16256 & n21315 ) | ( n16256 & n25747 ) | ( n21315 & n25747 ) ;
  assign n35191 = n35190 ^ n4633 ^ x155 ;
  assign n35192 = n18166 ^ n6784 ^ n981 ;
  assign n35193 = ~n18424 & n35192 ;
  assign n35194 = n35193 ^ n7181 ^ 1'b0 ;
  assign n35195 = n32069 ^ n7532 ^ n3357 ;
  assign n35196 = n35195 ^ n7385 ^ n2284 ;
  assign n35197 = n17355 ^ n16213 ^ n7540 ;
  assign n35198 = ( n16909 & ~n27660 ) | ( n16909 & n31576 ) | ( ~n27660 & n31576 ) ;
  assign n35199 = n13088 ^ n5495 ^ 1'b0 ;
  assign n35200 = n10415 & ~n35199 ;
  assign n35201 = n18974 ^ n10326 ^ n8878 ;
  assign n35202 = ( ~n16544 & n30378 ) | ( ~n16544 & n35201 ) | ( n30378 & n35201 ) ;
  assign n35203 = n12093 & n35202 ;
  assign n35204 = n5253 & n35203 ;
  assign n35205 = n32339 ^ n22617 ^ n14902 ;
  assign n35206 = ( n12121 & ~n17605 ) | ( n12121 & n35205 ) | ( ~n17605 & n35205 ) ;
  assign n35207 = n23005 ^ n8765 ^ n3180 ;
  assign n35208 = n23149 ^ n16748 ^ 1'b0 ;
  assign n35209 = ( n6848 & n23082 ) | ( n6848 & ~n35208 ) | ( n23082 & ~n35208 ) ;
  assign n35211 = ~n1093 & n11853 ;
  assign n35212 = ( n5780 & n14422 ) | ( n5780 & ~n35211 ) | ( n14422 & ~n35211 ) ;
  assign n35210 = n4125 | n18432 ;
  assign n35213 = n35212 ^ n35210 ^ 1'b0 ;
  assign n35214 = ( n35207 & ~n35209 ) | ( n35207 & n35213 ) | ( ~n35209 & n35213 ) ;
  assign n35215 = n28219 ^ n12179 ^ n5468 ;
  assign n35216 = ( n1148 & ~n2795 ) | ( n1148 & n3269 ) | ( ~n2795 & n3269 ) ;
  assign n35217 = ~n28849 & n35216 ;
  assign n35218 = n11353 | n22097 ;
  assign n35219 = ( n24197 & n28582 ) | ( n24197 & n35218 ) | ( n28582 & n35218 ) ;
  assign n35220 = ( ~n2091 & n22142 ) | ( ~n2091 & n35219 ) | ( n22142 & n35219 ) ;
  assign n35223 = ( ~n2590 & n18511 ) | ( ~n2590 & n19478 ) | ( n18511 & n19478 ) ;
  assign n35221 = ( ~x249 & n8031 ) | ( ~x249 & n29941 ) | ( n8031 & n29941 ) ;
  assign n35222 = n10796 & n35221 ;
  assign n35224 = n35223 ^ n35222 ^ 1'b0 ;
  assign n35225 = n18888 ^ n9633 ^ n4384 ;
  assign n35226 = ( n5226 & ~n28048 ) | ( n5226 & n35225 ) | ( ~n28048 & n35225 ) ;
  assign n35227 = ( ~n2337 & n8083 ) | ( ~n2337 & n21754 ) | ( n8083 & n21754 ) ;
  assign n35228 = ( x146 & n2537 ) | ( x146 & n6824 ) | ( n2537 & n6824 ) ;
  assign n35229 = ( n23250 & ~n35227 ) | ( n23250 & n35228 ) | ( ~n35227 & n35228 ) ;
  assign n35230 = n15115 ^ n13140 ^ 1'b0 ;
  assign n35231 = ( n19950 & n34494 ) | ( n19950 & n35230 ) | ( n34494 & n35230 ) ;
  assign n35232 = n35231 ^ n13827 ^ n9721 ;
  assign n35233 = ( n12570 & n33815 ) | ( n12570 & ~n35232 ) | ( n33815 & ~n35232 ) ;
  assign n35234 = ( n2717 & n19665 ) | ( n2717 & n24638 ) | ( n19665 & n24638 ) ;
  assign n35235 = ( n2933 & n6770 ) | ( n2933 & n27896 ) | ( n6770 & n27896 ) ;
  assign n35236 = n35235 ^ n5287 ^ n4213 ;
  assign n35237 = n23956 | n30692 ;
  assign n35238 = n35236 & ~n35237 ;
  assign n35239 = ~n22087 & n25882 ;
  assign n35240 = ~n15754 & n35239 ;
  assign n35241 = n19415 ^ n17505 ^ n11599 ;
  assign n35242 = ( ~n8627 & n10040 ) | ( ~n8627 & n35241 ) | ( n10040 & n35241 ) ;
  assign n35243 = n30754 ^ n27854 ^ n11913 ;
  assign n35244 = ( n1358 & n1377 ) | ( n1358 & ~n3886 ) | ( n1377 & ~n3886 ) ;
  assign n35245 = n35244 ^ n23893 ^ n7740 ;
  assign n35246 = n4247 & ~n35245 ;
  assign n35247 = ( n2314 & n2373 ) | ( n2314 & n29955 ) | ( n2373 & n29955 ) ;
  assign n35248 = n35247 ^ n31087 ^ 1'b0 ;
  assign n35249 = ( n31297 & n31603 ) | ( n31297 & ~n32379 ) | ( n31603 & ~n32379 ) ;
  assign n35250 = n35249 ^ n29008 ^ n9754 ;
  assign n35251 = n22136 | n35250 ;
  assign n35252 = n30935 & ~n35251 ;
  assign n35253 = n19183 ^ n12094 ^ n6789 ;
  assign n35254 = ( ~n3009 & n12097 ) | ( ~n3009 & n35253 ) | ( n12097 & n35253 ) ;
  assign n35255 = n35254 ^ n13252 ^ n5491 ;
  assign n35256 = n35255 ^ n19098 ^ n1548 ;
  assign n35257 = n35256 ^ n7870 ^ 1'b0 ;
  assign n35258 = ( n9619 & n25626 ) | ( n9619 & ~n34577 ) | ( n25626 & ~n34577 ) ;
  assign n35259 = ( ~n4041 & n9797 ) | ( ~n4041 & n25931 ) | ( n9797 & n25931 ) ;
  assign n35260 = n9107 & n18827 ;
  assign n35261 = n22143 & n35260 ;
  assign n35262 = ( n4899 & n21808 ) | ( n4899 & n35261 ) | ( n21808 & n35261 ) ;
  assign n35263 = x209 ^ x130 ^ 1'b0 ;
  assign n35264 = ~n1925 & n35263 ;
  assign n35265 = ( n3927 & n22233 ) | ( n3927 & ~n35264 ) | ( n22233 & ~n35264 ) ;
  assign n35266 = ( n11084 & ~n13484 ) | ( n11084 & n35265 ) | ( ~n13484 & n35265 ) ;
  assign n35268 = ( n1065 & n25636 ) | ( n1065 & n25770 ) | ( n25636 & n25770 ) ;
  assign n35267 = n23791 ^ n12418 ^ n4395 ;
  assign n35269 = n35268 ^ n35267 ^ n34645 ;
  assign n35270 = ( n6641 & n35266 ) | ( n6641 & n35269 ) | ( n35266 & n35269 ) ;
  assign n35273 = n12172 ^ n2938 ^ n1737 ;
  assign n35271 = n23589 ^ n9141 ^ n2712 ;
  assign n35272 = n7034 & ~n35271 ;
  assign n35274 = n35273 ^ n35272 ^ n32263 ;
  assign n35275 = n34692 ^ n30044 ^ n24803 ;
  assign n35276 = ( ~n28076 & n28657 ) | ( ~n28076 & n35275 ) | ( n28657 & n35275 ) ;
  assign n35277 = ( n6645 & n28172 ) | ( n6645 & n35276 ) | ( n28172 & n35276 ) ;
  assign n35278 = ( n11171 & n12326 ) | ( n11171 & n16101 ) | ( n12326 & n16101 ) ;
  assign n35279 = ( n277 & n365 ) | ( n277 & n11898 ) | ( n365 & n11898 ) ;
  assign n35280 = ( ~n9566 & n9721 ) | ( ~n9566 & n35279 ) | ( n9721 & n35279 ) ;
  assign n35281 = ( n288 & ~n8161 ) | ( n288 & n16504 ) | ( ~n8161 & n16504 ) ;
  assign n35282 = n35281 ^ n21591 ^ n15067 ;
  assign n35283 = ( n10810 & n11498 ) | ( n10810 & n35282 ) | ( n11498 & n35282 ) ;
  assign n35284 = ( n22809 & n35280 ) | ( n22809 & ~n35283 ) | ( n35280 & ~n35283 ) ;
  assign n35285 = n11146 & n21820 ;
  assign n35286 = n7888 ^ n7231 ^ n1218 ;
  assign n35287 = n35286 ^ n34874 ^ n24091 ;
  assign n35291 = n24562 ^ n3387 ^ n580 ;
  assign n35292 = n6694 & n35291 ;
  assign n35293 = n35292 ^ n22453 ^ 1'b0 ;
  assign n35290 = n17753 ^ n8654 ^ 1'b0 ;
  assign n35288 = n26175 ^ n22613 ^ n11007 ;
  assign n35289 = n35288 ^ n28285 ^ n12393 ;
  assign n35294 = n35293 ^ n35290 ^ n35289 ;
  assign n35295 = ( n2606 & n6606 ) | ( n2606 & ~n19287 ) | ( n6606 & ~n19287 ) ;
  assign n35296 = n35295 ^ n27858 ^ n2615 ;
  assign n35297 = n28532 ^ n16443 ^ n2759 ;
  assign n35298 = ( n13926 & ~n29331 ) | ( n13926 & n35297 ) | ( ~n29331 & n35297 ) ;
  assign n35299 = n17615 ^ n10386 ^ 1'b0 ;
  assign n35300 = n35298 & n35299 ;
  assign n35301 = ( n5784 & n23265 ) | ( n5784 & n35300 ) | ( n23265 & n35300 ) ;
  assign n35302 = ( n7177 & n22312 ) | ( n7177 & ~n28037 ) | ( n22312 & ~n28037 ) ;
  assign n35303 = n35302 ^ n27990 ^ n27410 ;
  assign n35304 = n3343 & n35303 ;
  assign n35305 = n35304 ^ n18206 ^ 1'b0 ;
  assign n35306 = ( ~n10940 & n19823 ) | ( ~n10940 & n21505 ) | ( n19823 & n21505 ) ;
  assign n35307 = ( ~n4487 & n17937 ) | ( ~n4487 & n35306 ) | ( n17937 & n35306 ) ;
  assign n35308 = ( n9905 & n11989 ) | ( n9905 & ~n35307 ) | ( n11989 & ~n35307 ) ;
  assign n35309 = n4925 ^ n3390 ^ n280 ;
  assign n35310 = n4384 ^ n2803 ^ n2704 ;
  assign n35311 = ( n4299 & n35309 ) | ( n4299 & ~n35310 ) | ( n35309 & ~n35310 ) ;
  assign n35312 = n16067 ^ n11477 ^ n4738 ;
  assign n35313 = ( n2204 & n5809 ) | ( n2204 & n9054 ) | ( n5809 & n9054 ) ;
  assign n35314 = ( n5766 & ~n8226 ) | ( n5766 & n35313 ) | ( ~n8226 & n35313 ) ;
  assign n35315 = ( n19047 & n24551 ) | ( n19047 & ~n35314 ) | ( n24551 & ~n35314 ) ;
  assign n35316 = ( n20344 & n35312 ) | ( n20344 & n35315 ) | ( n35312 & n35315 ) ;
  assign n35317 = n18068 ^ n4785 ^ 1'b0 ;
  assign n35318 = n27982 & ~n35317 ;
  assign n35319 = ( n34540 & ~n35316 ) | ( n34540 & n35318 ) | ( ~n35316 & n35318 ) ;
  assign n35320 = ( n27221 & n35311 ) | ( n27221 & ~n35319 ) | ( n35311 & ~n35319 ) ;
  assign n35321 = n35031 ^ n6144 ^ n2087 ;
  assign n35322 = n35321 ^ n14283 ^ n4787 ;
  assign n35323 = n7657 & ~n13937 ;
  assign n35324 = n22476 & n35323 ;
  assign n35326 = ( n9801 & n11918 ) | ( n9801 & ~n16415 ) | ( n11918 & ~n16415 ) ;
  assign n35325 = ( ~n2255 & n13307 ) | ( ~n2255 & n17328 ) | ( n13307 & n17328 ) ;
  assign n35327 = n35326 ^ n35325 ^ n3727 ;
  assign n35328 = n35327 ^ n13258 ^ 1'b0 ;
  assign n35333 = n16202 ^ n12735 ^ 1'b0 ;
  assign n35334 = n17576 ^ n11126 ^ n4556 ;
  assign n35335 = ( n28013 & n35333 ) | ( n28013 & ~n35334 ) | ( n35333 & ~n35334 ) ;
  assign n35329 = ( n23711 & n24744 ) | ( n23711 & n26769 ) | ( n24744 & n26769 ) ;
  assign n35330 = ( n2695 & n17689 ) | ( n2695 & ~n35329 ) | ( n17689 & ~n35329 ) ;
  assign n35331 = ( ~n6644 & n10408 ) | ( ~n6644 & n35330 ) | ( n10408 & n35330 ) ;
  assign n35332 = n10266 | n35331 ;
  assign n35336 = n35335 ^ n35332 ^ n23166 ;
  assign n35337 = ( ~n415 & n17816 ) | ( ~n415 & n19349 ) | ( n17816 & n19349 ) ;
  assign n35338 = ( n6652 & n10311 ) | ( n6652 & ~n35337 ) | ( n10311 & ~n35337 ) ;
  assign n35341 = ( n314 & n3008 ) | ( n314 & ~n12949 ) | ( n3008 & ~n12949 ) ;
  assign n35339 = n23080 ^ n15486 ^ 1'b0 ;
  assign n35340 = ~n3030 & n35339 ;
  assign n35342 = n35341 ^ n35340 ^ n29181 ;
  assign n35343 = n25876 ^ n5647 ^ n459 ;
  assign n35344 = ( n4329 & n23918 ) | ( n4329 & ~n35343 ) | ( n23918 & ~n35343 ) ;
  assign n35345 = n35344 ^ n32089 ^ n2894 ;
  assign n35346 = n7191 ^ n3404 ^ 1'b0 ;
  assign n35347 = n8040 ^ n6646 ^ n5459 ;
  assign n35348 = ( n14727 & n31220 ) | ( n14727 & ~n35347 ) | ( n31220 & ~n35347 ) ;
  assign n35349 = n3284 | n9991 ;
  assign n35350 = n35349 ^ n15803 ^ 1'b0 ;
  assign n35351 = n35350 ^ n24674 ^ n18345 ;
  assign n35352 = ( n2894 & n3809 ) | ( n2894 & ~n29256 ) | ( n3809 & ~n29256 ) ;
  assign n35353 = n18822 ^ n16538 ^ n16492 ;
  assign n35354 = ( n2345 & n4886 ) | ( n2345 & n25853 ) | ( n4886 & n25853 ) ;
  assign n35355 = n7933 & n30864 ;
  assign n35356 = n35355 ^ n14397 ^ 1'b0 ;
  assign n35357 = ( ~n7038 & n14323 ) | ( ~n7038 & n35356 ) | ( n14323 & n35356 ) ;
  assign n35359 = n21679 ^ n6513 ^ n3986 ;
  assign n35358 = ( n10253 & ~n28162 ) | ( n10253 & n29333 ) | ( ~n28162 & n29333 ) ;
  assign n35360 = n35359 ^ n35358 ^ n24360 ;
  assign n35361 = n9536 ^ n7259 ^ n6746 ;
  assign n35362 = n4021 | n26473 ;
  assign n35363 = n18440 & ~n35362 ;
  assign n35364 = ( n3595 & n9507 ) | ( n3595 & ~n12823 ) | ( n9507 & ~n12823 ) ;
  assign n35365 = n35364 ^ n26987 ^ n13206 ;
  assign n35366 = n27885 ^ n19804 ^ x240 ;
  assign n35367 = ( ~n10173 & n29055 ) | ( ~n10173 & n33446 ) | ( n29055 & n33446 ) ;
  assign n35372 = ( n428 & n895 ) | ( n428 & ~n947 ) | ( n895 & ~n947 ) ;
  assign n35371 = n17054 ^ n13294 ^ n7566 ;
  assign n35373 = n35372 ^ n35371 ^ 1'b0 ;
  assign n35368 = n22615 ^ n16130 ^ n5694 ;
  assign n35369 = n35368 ^ n20150 ^ n2823 ;
  assign n35370 = n35369 ^ n20073 ^ n1895 ;
  assign n35374 = n35373 ^ n35370 ^ n8921 ;
  assign n35375 = ~n21828 & n33250 ;
  assign n35376 = ~n14685 & n35375 ;
  assign n35377 = ( n1278 & n17237 ) | ( n1278 & ~n19849 ) | ( n17237 & ~n19849 ) ;
  assign n35383 = ( n4271 & n12901 ) | ( n4271 & n34528 ) | ( n12901 & n34528 ) ;
  assign n35381 = ( ~n4762 & n8268 ) | ( ~n4762 & n25448 ) | ( n8268 & n25448 ) ;
  assign n35379 = ( n5060 & ~n15976 ) | ( n5060 & n17510 ) | ( ~n15976 & n17510 ) ;
  assign n35378 = n17312 ^ n7046 ^ n1035 ;
  assign n35380 = n35379 ^ n35378 ^ n3286 ;
  assign n35382 = n35381 ^ n35380 ^ n12117 ;
  assign n35384 = n35383 ^ n35382 ^ 1'b0 ;
  assign n35385 = n35377 | n35384 ;
  assign n35386 = n25725 ^ n19314 ^ n3158 ;
  assign n35387 = n35386 ^ n26020 ^ n2612 ;
  assign n35388 = n23413 ^ n8542 ^ n1644 ;
  assign n35391 = n20632 ^ n10994 ^ n5343 ;
  assign n35389 = n8783 & ~n12814 ;
  assign n35390 = n7055 & n35389 ;
  assign n35392 = n35391 ^ n35390 ^ n19425 ;
  assign n35393 = n11803 ^ n4473 ^ x12 ;
  assign n35394 = n6830 ^ n1028 ^ 1'b0 ;
  assign n35395 = ( n5292 & ~n35393 ) | ( n5292 & n35394 ) | ( ~n35393 & n35394 ) ;
  assign n35396 = n7560 ^ n6073 ^ 1'b0 ;
  assign n35397 = ~n28175 & n35396 ;
  assign n35398 = n11814 ^ n6652 ^ n878 ;
  assign n35399 = n1545 & ~n11056 ;
  assign n35400 = ~n22908 & n35399 ;
  assign n35401 = n35400 ^ n15551 ^ 1'b0 ;
  assign n35402 = n35398 & n35401 ;
  assign n35403 = n17853 ^ n1708 ^ 1'b0 ;
  assign n35404 = ~n29211 & n35403 ;
  assign n35405 = ( n7703 & ~n28771 ) | ( n7703 & n35404 ) | ( ~n28771 & n35404 ) ;
  assign n35406 = n25570 ^ n18004 ^ n8539 ;
  assign n35407 = n35406 ^ n26795 ^ n14533 ;
  assign n35408 = n16934 ^ n9986 ^ 1'b0 ;
  assign n35409 = ~n918 & n35408 ;
  assign n35410 = n23594 ^ n19400 ^ n10760 ;
  assign n35411 = ( n9565 & n28960 ) | ( n9565 & n35410 ) | ( n28960 & n35410 ) ;
  assign n35412 = ( n1852 & n35409 ) | ( n1852 & ~n35411 ) | ( n35409 & ~n35411 ) ;
  assign n35413 = n22542 ^ n20340 ^ n17386 ;
  assign n35414 = ( n2523 & n33902 ) | ( n2523 & ~n35413 ) | ( n33902 & ~n35413 ) ;
  assign n35415 = ( ~n22629 & n23740 ) | ( ~n22629 & n28384 ) | ( n23740 & n28384 ) ;
  assign n35416 = ( ~n2248 & n24184 ) | ( ~n2248 & n35415 ) | ( n24184 & n35415 ) ;
  assign n35417 = n6685 ^ n5179 ^ n3498 ;
  assign n35418 = n35417 ^ n18946 ^ n558 ;
  assign n35420 = ( ~n6001 & n13904 ) | ( ~n6001 & n20026 ) | ( n13904 & n20026 ) ;
  assign n35419 = n22463 ^ n18469 ^ n8955 ;
  assign n35421 = n35420 ^ n35419 ^ 1'b0 ;
  assign n35422 = n14817 ^ n11039 ^ n8178 ;
  assign n35423 = ( n2895 & n3124 ) | ( n2895 & n4013 ) | ( n3124 & n4013 ) ;
  assign n35424 = n35423 ^ n5814 ^ n4057 ;
  assign n35425 = n35424 ^ n16417 ^ 1'b0 ;
  assign n35426 = ~n35422 & n35425 ;
  assign n35427 = ( n11976 & n19639 ) | ( n11976 & ~n35426 ) | ( n19639 & ~n35426 ) ;
  assign n35428 = n18474 ^ n10560 ^ n2777 ;
  assign n35429 = n25049 & ~n35428 ;
  assign n35430 = ( ~n4731 & n6484 ) | ( ~n4731 & n18058 ) | ( n6484 & n18058 ) ;
  assign n35431 = ( n17540 & ~n23575 ) | ( n17540 & n35430 ) | ( ~n23575 & n35430 ) ;
  assign n35432 = ( n5769 & ~n14659 ) | ( n5769 & n16001 ) | ( ~n14659 & n16001 ) ;
  assign n35433 = ( n8671 & ~n33363 ) | ( n8671 & n35432 ) | ( ~n33363 & n35432 ) ;
  assign n35434 = n14935 & n35433 ;
  assign n35435 = ( n16975 & ~n19373 ) | ( n16975 & n35434 ) | ( ~n19373 & n35434 ) ;
  assign n35436 = ( n29978 & n35431 ) | ( n29978 & n35435 ) | ( n35431 & n35435 ) ;
  assign n35437 = ( n2345 & n4568 ) | ( n2345 & ~n21187 ) | ( n4568 & ~n21187 ) ;
  assign n35438 = n35437 ^ n4575 ^ n3532 ;
  assign n35439 = n35438 ^ n16676 ^ x9 ;
  assign n35440 = n6964 & n35439 ;
  assign n35441 = ~n19863 & n35440 ;
  assign n35443 = ( n22132 & n23353 ) | ( n22132 & n35165 ) | ( n23353 & n35165 ) ;
  assign n35442 = n3805 & n12221 ;
  assign n35444 = n35443 ^ n35442 ^ 1'b0 ;
  assign n35445 = ( n14346 & n32773 ) | ( n14346 & ~n35444 ) | ( n32773 & ~n35444 ) ;
  assign n35446 = n35445 ^ n18703 ^ 1'b0 ;
  assign n35448 = n20314 ^ n6895 ^ n6580 ;
  assign n35449 = n35448 ^ n12266 ^ n3790 ;
  assign n35447 = n34692 ^ n15406 ^ n1210 ;
  assign n35450 = n35449 ^ n35447 ^ n16701 ;
  assign n35451 = n11733 & ~n27612 ;
  assign n35452 = ( ~n2366 & n10551 ) | ( ~n2366 & n35451 ) | ( n10551 & n35451 ) ;
  assign n35453 = n35452 ^ n32252 ^ 1'b0 ;
  assign n35460 = n15849 ^ n8484 ^ n2546 ;
  assign n35461 = n35460 ^ n18974 ^ x66 ;
  assign n35462 = ( n940 & n7250 ) | ( n940 & ~n35461 ) | ( n7250 & ~n35461 ) ;
  assign n35458 = n32315 ^ n9746 ^ n3650 ;
  assign n35459 = ( ~n7241 & n12406 ) | ( ~n7241 & n35458 ) | ( n12406 & n35458 ) ;
  assign n35454 = ( n1409 & ~n4970 ) | ( n1409 & n11473 ) | ( ~n4970 & n11473 ) ;
  assign n35455 = ( n22047 & n30592 ) | ( n22047 & n35454 ) | ( n30592 & n35454 ) ;
  assign n35456 = ( n3815 & n5172 ) | ( n3815 & ~n35455 ) | ( n5172 & ~n35455 ) ;
  assign n35457 = n35456 ^ n16481 ^ n10242 ;
  assign n35463 = n35462 ^ n35459 ^ n35457 ;
  assign n35464 = ( n2618 & n5495 ) | ( n2618 & ~n9905 ) | ( n5495 & ~n9905 ) ;
  assign n35465 = n24287 ^ n11771 ^ 1'b0 ;
  assign n35466 = ( n16273 & ~n35464 ) | ( n16273 & n35465 ) | ( ~n35464 & n35465 ) ;
  assign n35469 = n29456 ^ n16933 ^ 1'b0 ;
  assign n35467 = n6836 & n35144 ;
  assign n35468 = ~n15135 & n35467 ;
  assign n35470 = n35469 ^ n35468 ^ n20241 ;
  assign n35471 = n28517 ^ n26695 ^ n24891 ;
  assign n35472 = ( n5429 & n6483 ) | ( n5429 & n10426 ) | ( n6483 & n10426 ) ;
  assign n35473 = ( n702 & n6279 ) | ( n702 & ~n35472 ) | ( n6279 & ~n35472 ) ;
  assign n35478 = n7283 ^ n7160 ^ n6818 ;
  assign n35474 = ( n1103 & ~n7875 ) | ( n1103 & n22939 ) | ( ~n7875 & n22939 ) ;
  assign n35475 = n33521 ^ n10649 ^ n6631 ;
  assign n35476 = ( n20788 & n35474 ) | ( n20788 & n35475 ) | ( n35474 & n35475 ) ;
  assign n35477 = n35476 ^ n30906 ^ n13795 ;
  assign n35479 = n35478 ^ n35477 ^ n3004 ;
  assign n35480 = n19999 ^ n16047 ^ 1'b0 ;
  assign n35481 = n335 & ~n35480 ;
  assign n35482 = n7946 ^ n2450 ^ 1'b0 ;
  assign n35483 = n35481 & ~n35482 ;
  assign n35485 = n16291 ^ n13508 ^ n10737 ;
  assign n35484 = n25656 & n30909 ;
  assign n35486 = n35485 ^ n35484 ^ n28447 ;
  assign n35487 = n13710 ^ n9726 ^ n4355 ;
  assign n35488 = n16128 & ~n29167 ;
  assign n35489 = ~n13169 & n35488 ;
  assign n35490 = n35489 ^ n15924 ^ n11315 ;
  assign n35492 = ( ~n1326 & n2551 ) | ( ~n1326 & n3677 ) | ( n2551 & n3677 ) ;
  assign n35491 = n27330 ^ n17591 ^ n414 ;
  assign n35493 = n35492 ^ n35491 ^ n19815 ;
  assign n35494 = n18892 ^ n13584 ^ n13118 ;
  assign n35495 = n35494 ^ n27045 ^ n14205 ;
  assign n35496 = n28927 ^ n21133 ^ n18820 ;
  assign n35497 = n35496 ^ n33066 ^ 1'b0 ;
  assign n35498 = n30148 ^ n15856 ^ n14682 ;
  assign n35499 = n11640 ^ n5001 ^ 1'b0 ;
  assign n35500 = ( n4420 & ~n6148 ) | ( n4420 & n18908 ) | ( ~n6148 & n18908 ) ;
  assign n35501 = ~n2059 & n2252 ;
  assign n35502 = n35501 ^ n13980 ^ 1'b0 ;
  assign n35503 = ( n5832 & ~n33160 ) | ( n5832 & n35502 ) | ( ~n33160 & n35502 ) ;
  assign n35504 = ( n17868 & n35500 ) | ( n17868 & n35503 ) | ( n35500 & n35503 ) ;
  assign n35505 = ( n26874 & n35499 ) | ( n26874 & ~n35504 ) | ( n35499 & ~n35504 ) ;
  assign n35506 = ~n10578 & n30281 ;
  assign n35507 = n35505 & n35506 ;
  assign n35508 = ( n681 & n13847 ) | ( n681 & n14089 ) | ( n13847 & n14089 ) ;
  assign n35509 = ~n14756 & n35508 ;
  assign n35510 = n35509 ^ n23569 ^ n9855 ;
  assign n35511 = n18904 ^ n14242 ^ n4163 ;
  assign n35512 = n23639 ^ n15100 ^ n11530 ;
  assign n35513 = ( n35510 & n35511 ) | ( n35510 & ~n35512 ) | ( n35511 & ~n35512 ) ;
  assign n35514 = ( ~n2118 & n14751 ) | ( ~n2118 & n25997 ) | ( n14751 & n25997 ) ;
  assign n35515 = ( n27948 & n35513 ) | ( n27948 & ~n35514 ) | ( n35513 & ~n35514 ) ;
  assign n35516 = n11098 ^ n8716 ^ n2491 ;
  assign n35517 = n24200 ^ n22585 ^ n7076 ;
  assign n35518 = ( n4694 & ~n21424 ) | ( n4694 & n21862 ) | ( ~n21424 & n21862 ) ;
  assign n35519 = ( n3278 & n8335 ) | ( n3278 & ~n35518 ) | ( n8335 & ~n35518 ) ;
  assign n35520 = n35519 ^ n32320 ^ n1904 ;
  assign n35521 = ( ~n30901 & n31187 ) | ( ~n30901 & n35520 ) | ( n31187 & n35520 ) ;
  assign n35522 = ( ~n3373 & n19394 ) | ( ~n3373 & n20917 ) | ( n19394 & n20917 ) ;
  assign n35529 = ( n4934 & n5351 ) | ( n4934 & n17697 ) | ( n5351 & n17697 ) ;
  assign n35523 = ( ~n8294 & n8460 ) | ( ~n8294 & n13337 ) | ( n8460 & n13337 ) ;
  assign n35524 = n35523 ^ x225 ^ 1'b0 ;
  assign n35525 = n35524 ^ n21553 ^ n14252 ;
  assign n35526 = ( ~n3495 & n7748 ) | ( ~n3495 & n10719 ) | ( n7748 & n10719 ) ;
  assign n35527 = ( n2415 & n8938 ) | ( n2415 & ~n35526 ) | ( n8938 & ~n35526 ) ;
  assign n35528 = ( n4144 & ~n35525 ) | ( n4144 & n35527 ) | ( ~n35525 & n35527 ) ;
  assign n35530 = n35529 ^ n35528 ^ 1'b0 ;
  assign n35531 = n14998 & ~n35530 ;
  assign n35532 = ( n15141 & n35522 ) | ( n15141 & ~n35531 ) | ( n35522 & ~n35531 ) ;
  assign n35533 = ~n1822 & n25894 ;
  assign n35534 = n35533 ^ n15109 ^ n12330 ;
  assign n35535 = n35534 ^ n23958 ^ n18587 ;
  assign n35537 = n13214 ^ n3649 ^ n3302 ;
  assign n35536 = n1562 & ~n14925 ;
  assign n35538 = n35537 ^ n35536 ^ 1'b0 ;
  assign n35539 = ( ~n13300 & n14835 ) | ( ~n13300 & n35538 ) | ( n14835 & n35538 ) ;
  assign n35540 = ( ~n18100 & n21397 ) | ( ~n18100 & n34309 ) | ( n21397 & n34309 ) ;
  assign n35541 = n29392 ^ n18934 ^ n5489 ;
  assign n35542 = ( n7714 & n20015 ) | ( n7714 & ~n35541 ) | ( n20015 & ~n35541 ) ;
  assign n35543 = n31075 | n35542 ;
  assign n35544 = n34321 & n35543 ;
  assign n35545 = ~n35540 & n35544 ;
  assign n35546 = n7606 ^ x184 ^ 1'b0 ;
  assign n35547 = ~n10278 & n35546 ;
  assign n35548 = n35547 ^ n13837 ^ n13360 ;
  assign n35549 = ( n15791 & n16612 ) | ( n15791 & ~n23232 ) | ( n16612 & ~n23232 ) ;
  assign n35550 = ( n5962 & n18068 ) | ( n5962 & ~n35549 ) | ( n18068 & ~n35549 ) ;
  assign n35551 = n11600 ^ n2811 ^ 1'b0 ;
  assign n35552 = n35551 ^ n29168 ^ n2994 ;
  assign n35554 = ~n2938 & n5540 ;
  assign n35555 = n35554 ^ n10031 ^ n4283 ;
  assign n35553 = n11898 & n24868 ;
  assign n35556 = n35555 ^ n35553 ^ 1'b0 ;
  assign n35557 = ( n6573 & n7183 ) | ( n6573 & n35556 ) | ( n7183 & n35556 ) ;
  assign n35559 = n8508 & n30403 ;
  assign n35560 = n35559 ^ n8793 ^ 1'b0 ;
  assign n35558 = n3462 & n35028 ;
  assign n35561 = n35560 ^ n35558 ^ n16244 ;
  assign n35562 = n26027 ^ n10205 ^ n9069 ;
  assign n35563 = ( n15329 & n20062 ) | ( n15329 & n35562 ) | ( n20062 & n35562 ) ;
  assign n35564 = ( n22020 & n33295 ) | ( n22020 & n35563 ) | ( n33295 & n35563 ) ;
  assign n35565 = ( n272 & ~n10299 ) | ( n272 & n26249 ) | ( ~n10299 & n26249 ) ;
  assign n35566 = ~n22112 & n35565 ;
  assign n35567 = n35566 ^ n30616 ^ 1'b0 ;
  assign n35571 = ( n6008 & n11152 ) | ( n6008 & n34054 ) | ( n11152 & n34054 ) ;
  assign n35568 = ( x131 & n5197 ) | ( x131 & ~n6587 ) | ( n5197 & ~n6587 ) ;
  assign n35569 = ( n2515 & ~n21438 ) | ( n2515 & n35568 ) | ( ~n21438 & n35568 ) ;
  assign n35570 = n35569 ^ n9541 ^ n5648 ;
  assign n35572 = n35571 ^ n35570 ^ n34633 ;
  assign n35573 = n5663 & ~n14398 ;
  assign n35574 = ( n18679 & n27914 ) | ( n18679 & n35573 ) | ( n27914 & n35573 ) ;
  assign n35576 = n18976 ^ n8835 ^ n4651 ;
  assign n35577 = n35576 ^ n18058 ^ n9661 ;
  assign n35575 = n28684 ^ n17818 ^ n5919 ;
  assign n35578 = n35577 ^ n35575 ^ n32916 ;
  assign n35579 = n33479 ^ n8249 ^ n5344 ;
  assign n35580 = ( n33517 & ~n34745 ) | ( n33517 & n35579 ) | ( ~n34745 & n35579 ) ;
  assign n35581 = ( n282 & ~n808 ) | ( n282 & n35580 ) | ( ~n808 & n35580 ) ;
  assign n35582 = n25049 ^ n18656 ^ n5689 ;
  assign n35583 = ~n1787 & n3170 ;
  assign n35584 = ( n12651 & n16375 ) | ( n12651 & ~n16619 ) | ( n16375 & ~n16619 ) ;
  assign n35585 = n9504 & n31211 ;
  assign n35586 = n35585 ^ n9685 ^ 1'b0 ;
  assign n35587 = n16816 ^ n3367 ^ n1789 ;
  assign n35588 = n35587 ^ n24586 ^ n4039 ;
  assign n35589 = ( n10976 & n16342 ) | ( n10976 & ~n25739 ) | ( n16342 & ~n25739 ) ;
  assign n35590 = n35589 ^ n30963 ^ n8639 ;
  assign n35591 = ( n12220 & n35588 ) | ( n12220 & n35590 ) | ( n35588 & n35590 ) ;
  assign n35592 = ( n35584 & ~n35586 ) | ( n35584 & n35591 ) | ( ~n35586 & n35591 ) ;
  assign n35593 = n20059 ^ n7293 ^ 1'b0 ;
  assign n35594 = ~n2380 & n35593 ;
  assign n35595 = n4516 & ~n35594 ;
  assign n35596 = n35595 ^ n28779 ^ n6202 ;
  assign n35597 = ( ~n35583 & n35592 ) | ( ~n35583 & n35596 ) | ( n35592 & n35596 ) ;
  assign n35598 = ( n2288 & ~n12286 ) | ( n2288 & n30706 ) | ( ~n12286 & n30706 ) ;
  assign n35599 = ( n2612 & n4855 ) | ( n2612 & n28986 ) | ( n4855 & n28986 ) ;
  assign n35600 = n11332 & ~n34267 ;
  assign n35601 = n35600 ^ n22081 ^ n15685 ;
  assign n35602 = ( n20268 & n34206 ) | ( n20268 & ~n35601 ) | ( n34206 & ~n35601 ) ;
  assign n35603 = ( n12545 & n20582 ) | ( n12545 & n29953 ) | ( n20582 & n29953 ) ;
  assign n35604 = n22620 & n35603 ;
  assign n35605 = ( n1648 & ~n4519 ) | ( n1648 & n8087 ) | ( ~n4519 & n8087 ) ;
  assign n35606 = n20497 | n35605 ;
  assign n35607 = ( ~n11619 & n27299 ) | ( ~n11619 & n35606 ) | ( n27299 & n35606 ) ;
  assign n35608 = n7407 & n35607 ;
  assign n35609 = ~n34111 & n35608 ;
  assign n35610 = n35609 ^ n29539 ^ n19888 ;
  assign n35611 = ( n25372 & ~n35604 ) | ( n25372 & n35610 ) | ( ~n35604 & n35610 ) ;
  assign n35612 = n13412 ^ n7968 ^ n4340 ;
  assign n35613 = ( n461 & n1365 ) | ( n461 & ~n10810 ) | ( n1365 & ~n10810 ) ;
  assign n35614 = n11699 & ~n14656 ;
  assign n35615 = ( n4141 & n35613 ) | ( n4141 & ~n35614 ) | ( n35613 & ~n35614 ) ;
  assign n35616 = n23722 ^ n18151 ^ n4074 ;
  assign n35617 = ( n3831 & n22330 ) | ( n3831 & n35616 ) | ( n22330 & n35616 ) ;
  assign n35618 = n23169 | n30291 ;
  assign n35620 = ( n931 & ~n21970 ) | ( n931 & n25806 ) | ( ~n21970 & n25806 ) ;
  assign n35619 = ( n9082 & n27807 ) | ( n9082 & n31460 ) | ( n27807 & n31460 ) ;
  assign n35621 = n35620 ^ n35619 ^ n32780 ;
  assign n35622 = n9776 ^ n3815 ^ 1'b0 ;
  assign n35623 = ( n4825 & n9517 ) | ( n4825 & n24327 ) | ( n9517 & n24327 ) ;
  assign n35624 = ( n35484 & n35622 ) | ( n35484 & n35623 ) | ( n35622 & n35623 ) ;
  assign n35625 = ( n1484 & n18810 ) | ( n1484 & ~n24533 ) | ( n18810 & ~n24533 ) ;
  assign n35626 = ~n21024 & n29323 ;
  assign n35627 = n1852 & ~n33924 ;
  assign n35628 = n35627 ^ n23032 ^ 1'b0 ;
  assign n35629 = ( ~n24182 & n26726 ) | ( ~n24182 & n35529 ) | ( n26726 & n35529 ) ;
  assign n35630 = ( n12547 & ~n19487 ) | ( n12547 & n20954 ) | ( ~n19487 & n20954 ) ;
  assign n35631 = n35630 ^ n28834 ^ n872 ;
  assign n35632 = n35631 ^ n18643 ^ n15064 ;
  assign n35633 = n20815 ^ n15863 ^ n4043 ;
  assign n35634 = n23846 ^ n11117 ^ n2493 ;
  assign n35635 = n35634 ^ n13392 ^ n7257 ;
  assign n35636 = ( n22138 & n35633 ) | ( n22138 & ~n35635 ) | ( n35633 & ~n35635 ) ;
  assign n35637 = n5235 ^ n3382 ^ n823 ;
  assign n35638 = n35637 ^ n15321 ^ n8403 ;
  assign n35639 = n34473 | n35638 ;
  assign n35640 = n18663 & ~n35639 ;
  assign n35641 = n35640 ^ n14132 ^ n5477 ;
  assign n35642 = ( ~n671 & n8219 ) | ( ~n671 & n25257 ) | ( n8219 & n25257 ) ;
  assign n35643 = ( ~n704 & n8870 ) | ( ~n704 & n35642 ) | ( n8870 & n35642 ) ;
  assign n35644 = ( n15553 & ~n23014 ) | ( n15553 & n35643 ) | ( ~n23014 & n35643 ) ;
  assign n35645 = ( n4830 & ~n21648 ) | ( n4830 & n27983 ) | ( ~n21648 & n27983 ) ;
  assign n35646 = n34667 ^ n618 ^ x85 ;
  assign n35647 = ( n5061 & n35645 ) | ( n5061 & ~n35646 ) | ( n35645 & ~n35646 ) ;
  assign n35649 = n10689 ^ n9177 ^ 1'b0 ;
  assign n35650 = n10710 & ~n35649 ;
  assign n35651 = ( n4945 & ~n13998 ) | ( n4945 & n35650 ) | ( ~n13998 & n35650 ) ;
  assign n35652 = n35651 ^ n28222 ^ 1'b0 ;
  assign n35653 = n8683 & ~n35652 ;
  assign n35648 = n3568 & n27317 ;
  assign n35654 = n35653 ^ n35648 ^ 1'b0 ;
  assign n35655 = n12506 ^ n8056 ^ 1'b0 ;
  assign n35656 = n9715 ^ n4436 ^ n3396 ;
  assign n35657 = ( ~n1301 & n3763 ) | ( ~n1301 & n35656 ) | ( n3763 & n35656 ) ;
  assign n35658 = n35657 ^ n33021 ^ n18437 ;
  assign n35659 = n35658 ^ n20657 ^ n1934 ;
  assign n35660 = ( n9806 & n35655 ) | ( n9806 & n35659 ) | ( n35655 & n35659 ) ;
  assign n35661 = ( n3584 & n5995 ) | ( n3584 & n35660 ) | ( n5995 & n35660 ) ;
  assign n35665 = n5439 ^ n1752 ^ 1'b0 ;
  assign n35666 = n9591 & n35665 ;
  assign n35662 = n12748 ^ n1702 ^ 1'b0 ;
  assign n35663 = n16595 | n35662 ;
  assign n35664 = n35663 ^ n28425 ^ n257 ;
  assign n35667 = n35666 ^ n35664 ^ n35412 ;
  assign n35668 = ( ~n4947 & n6830 ) | ( ~n4947 & n12545 ) | ( n6830 & n12545 ) ;
  assign n35669 = n26574 ^ n13730 ^ n1410 ;
  assign n35670 = ( ~n11821 & n35668 ) | ( ~n11821 & n35669 ) | ( n35668 & n35669 ) ;
  assign n35671 = ( n5889 & ~n13907 ) | ( n5889 & n35670 ) | ( ~n13907 & n35670 ) ;
  assign n35672 = n19023 ^ n3435 ^ n2173 ;
  assign n35673 = n35672 ^ n34475 ^ n26538 ;
  assign n35674 = n31875 ^ n20168 ^ n8536 ;
  assign n35675 = ( n4950 & ~n11080 ) | ( n4950 & n18132 ) | ( ~n11080 & n18132 ) ;
  assign n35676 = n11181 & n35675 ;
  assign n35678 = n19667 ^ n7516 ^ n3148 ;
  assign n35679 = n9772 & ~n35678 ;
  assign n35677 = n11679 ^ n6584 ^ n2710 ;
  assign n35680 = n35679 ^ n35677 ^ n33774 ;
  assign n35681 = n18487 ^ n15788 ^ n13803 ;
  assign n35682 = n35681 ^ n20728 ^ n18602 ;
  assign n35683 = n35682 ^ n11266 ^ n9767 ;
  assign n35684 = n1094 | n31969 ;
  assign n35685 = n35684 ^ n24080 ^ 1'b0 ;
  assign n35686 = n35685 ^ n18603 ^ n625 ;
  assign n35687 = n12067 ^ n11614 ^ n5253 ;
  assign n35688 = ( n2362 & n26963 ) | ( n2362 & n28007 ) | ( n26963 & n28007 ) ;
  assign n35689 = ( n25536 & n31633 ) | ( n25536 & ~n35688 ) | ( n31633 & ~n35688 ) ;
  assign n35690 = n17294 ^ n13251 ^ 1'b0 ;
  assign n35691 = n23028 | n35690 ;
  assign n35692 = ( ~n3247 & n15794 ) | ( ~n3247 & n35691 ) | ( n15794 & n35691 ) ;
  assign n35697 = n18656 ^ n10042 ^ n6861 ;
  assign n35693 = n5174 & n7418 ;
  assign n35694 = n3116 & n35693 ;
  assign n35695 = n17421 ^ n10462 ^ 1'b0 ;
  assign n35696 = ( n28983 & ~n35694 ) | ( n28983 & n35695 ) | ( ~n35694 & n35695 ) ;
  assign n35698 = n35697 ^ n35696 ^ n21599 ;
  assign n35699 = ( ~n12836 & n15317 ) | ( ~n12836 & n35698 ) | ( n15317 & n35698 ) ;
  assign n35700 = ( ~n12893 & n16314 ) | ( ~n12893 & n21045 ) | ( n16314 & n21045 ) ;
  assign n35701 = ( n2138 & n23377 ) | ( n2138 & ~n35700 ) | ( n23377 & ~n35700 ) ;
  assign n35702 = n35701 ^ n20168 ^ n16473 ;
  assign n35703 = n35702 ^ n10342 ^ 1'b0 ;
  assign n35704 = ~n1390 & n35703 ;
  assign n35705 = n34242 ^ n27650 ^ n12708 ;
  assign n35707 = n7051 | n22163 ;
  assign n35706 = n11837 & ~n28468 ;
  assign n35708 = n35707 ^ n35706 ^ 1'b0 ;
  assign n35709 = ( n7839 & ~n28993 ) | ( n7839 & n35708 ) | ( ~n28993 & n35708 ) ;
  assign n35710 = n35709 ^ n18521 ^ 1'b0 ;
  assign n35711 = ( ~n2918 & n10985 ) | ( ~n2918 & n28370 ) | ( n10985 & n28370 ) ;
  assign n35712 = n35711 ^ n9572 ^ n649 ;
  assign n35713 = n35712 ^ n3601 ^ x175 ;
  assign n35714 = ( n4241 & n7572 ) | ( n4241 & ~n12954 ) | ( n7572 & ~n12954 ) ;
  assign n35715 = n31036 ^ n10078 ^ n5185 ;
  assign n35716 = ( ~n5230 & n10016 ) | ( ~n5230 & n35715 ) | ( n10016 & n35715 ) ;
  assign n35717 = n35716 ^ n31235 ^ n19553 ;
  assign n35718 = ( n27913 & n35714 ) | ( n27913 & n35717 ) | ( n35714 & n35717 ) ;
  assign n35719 = n17512 ^ n5534 ^ n3877 ;
  assign n35720 = ( ~n30049 & n30695 ) | ( ~n30049 & n35719 ) | ( n30695 & n35719 ) ;
  assign n35721 = ( n6073 & n11769 ) | ( n6073 & n35513 ) | ( n11769 & n35513 ) ;
  assign n35722 = n19080 | n29588 ;
  assign n35723 = n35721 | n35722 ;
  assign n35724 = n12085 ^ n10889 ^ n5030 ;
  assign n35725 = n35724 ^ n6921 ^ 1'b0 ;
  assign n35726 = ~n4375 & n35725 ;
  assign n35727 = n35726 ^ n20028 ^ n9905 ;
  assign n35728 = ( n9289 & n28473 ) | ( n9289 & n32403 ) | ( n28473 & n32403 ) ;
  assign n35729 = n35728 ^ n10374 ^ n8721 ;
  assign n35730 = ( n10839 & n35727 ) | ( n10839 & n35729 ) | ( n35727 & n35729 ) ;
  assign n35731 = n3887 & ~n13506 ;
  assign n35732 = n972 & n35731 ;
  assign n35733 = n35732 ^ n32566 ^ n2898 ;
  assign n35734 = n35733 ^ n22561 ^ n21005 ;
  assign n35735 = ( n3720 & n7712 ) | ( n3720 & n10099 ) | ( n7712 & n10099 ) ;
  assign n35736 = n21932 ^ n14859 ^ n6698 ;
  assign n35737 = ( ~n15818 & n35735 ) | ( ~n15818 & n35736 ) | ( n35735 & n35736 ) ;
  assign n35740 = ( n555 & n10256 ) | ( n555 & n18532 ) | ( n10256 & n18532 ) ;
  assign n35739 = ( n10348 & n18467 ) | ( n10348 & n30044 ) | ( n18467 & n30044 ) ;
  assign n35738 = n33181 ^ n11374 ^ n5352 ;
  assign n35741 = n35740 ^ n35739 ^ n35738 ;
  assign n35742 = n375 & ~n35741 ;
  assign n35743 = n35742 ^ n9748 ^ 1'b0 ;
  assign n35744 = n23926 ^ n8178 ^ n4470 ;
  assign n35745 = n35744 ^ n17994 ^ n13493 ;
  assign n35746 = ( n4558 & ~n4874 ) | ( n4558 & n9042 ) | ( ~n4874 & n9042 ) ;
  assign n35747 = n28720 ^ n17172 ^ n8323 ;
  assign n35748 = ( n35745 & ~n35746 ) | ( n35745 & n35747 ) | ( ~n35746 & n35747 ) ;
  assign n35749 = n8281 ^ n8256 ^ n7528 ;
  assign n35751 = n17642 ^ n15848 ^ n1749 ;
  assign n35750 = ~n6503 & n34727 ;
  assign n35752 = n35751 ^ n35750 ^ 1'b0 ;
  assign n35753 = n21233 ^ n8772 ^ 1'b0 ;
  assign n35754 = n24261 & n35753 ;
  assign n35755 = ( n7232 & n12019 ) | ( n7232 & ~n28580 ) | ( n12019 & ~n28580 ) ;
  assign n35756 = n35755 ^ n20644 ^ 1'b0 ;
  assign n35757 = ~n4320 & n35756 ;
  assign n35758 = ( ~n4122 & n8153 ) | ( ~n4122 & n24474 ) | ( n8153 & n24474 ) ;
  assign n35759 = ( n11612 & n25905 ) | ( n11612 & n35758 ) | ( n25905 & n35758 ) ;
  assign n35760 = n4770 | n11315 ;
  assign n35761 = n19356 ^ n9190 ^ n6900 ;
  assign n35762 = ( n9481 & ~n35760 ) | ( n9481 & n35761 ) | ( ~n35760 & n35761 ) ;
  assign n35763 = ( n18831 & n27223 ) | ( n18831 & n35762 ) | ( n27223 & n35762 ) ;
  assign n35764 = n23933 ^ n11562 ^ n8145 ;
  assign n35765 = ( n2439 & ~n11139 ) | ( n2439 & n35764 ) | ( ~n11139 & n35764 ) ;
  assign n35766 = ( n16591 & n19843 ) | ( n16591 & ~n34092 ) | ( n19843 & ~n34092 ) ;
  assign n35767 = ( n16758 & n27786 ) | ( n16758 & ~n35766 ) | ( n27786 & ~n35766 ) ;
  assign n35768 = n22431 ^ n794 ^ 1'b0 ;
  assign n35769 = n7418 & n35768 ;
  assign n35770 = x177 & n35769 ;
  assign n35771 = n6060 & n35770 ;
  assign n35772 = ( n4875 & n6008 ) | ( n4875 & ~n12170 ) | ( n6008 & ~n12170 ) ;
  assign n35773 = ( n23175 & n27907 ) | ( n23175 & n35772 ) | ( n27907 & n35772 ) ;
  assign n35774 = ( n3828 & n35771 ) | ( n3828 & ~n35773 ) | ( n35771 & ~n35773 ) ;
  assign n35775 = ( n28579 & n31107 ) | ( n28579 & n35774 ) | ( n31107 & n35774 ) ;
  assign n35776 = n35775 ^ n28613 ^ n8171 ;
  assign n35782 = ( ~n6346 & n19905 ) | ( ~n6346 & n23784 ) | ( n19905 & n23784 ) ;
  assign n35777 = ( n2101 & ~n8385 ) | ( n2101 & n12110 ) | ( ~n8385 & n12110 ) ;
  assign n35778 = n35777 ^ n7276 ^ n3450 ;
  assign n35779 = n10993 & ~n35778 ;
  assign n35780 = ~n30264 & n35779 ;
  assign n35781 = n35780 ^ n4037 ^ n2635 ;
  assign n35783 = n35782 ^ n35781 ^ n30384 ;
  assign n35784 = n21805 ^ n6136 ^ n4521 ;
  assign n35785 = n35784 ^ n24628 ^ n7239 ;
  assign n35786 = n28175 ^ n4702 ^ 1'b0 ;
  assign n35787 = n19868 ^ n11153 ^ 1'b0 ;
  assign n35788 = ( n29741 & n35786 ) | ( n29741 & n35787 ) | ( n35786 & n35787 ) ;
  assign n35789 = n7362 ^ x122 ^ 1'b0 ;
  assign n35790 = ( n2336 & ~n10391 ) | ( n2336 & n35789 ) | ( ~n10391 & n35789 ) ;
  assign n35791 = n24363 ^ n14048 ^ n7708 ;
  assign n35792 = ( ~x227 & n2016 ) | ( ~x227 & n35791 ) | ( n2016 & n35791 ) ;
  assign n35793 = ( n11245 & n34656 ) | ( n11245 & ~n35792 ) | ( n34656 & ~n35792 ) ;
  assign n35794 = n35793 ^ n30252 ^ n5201 ;
  assign n35795 = n32440 ^ n16216 ^ n880 ;
  assign n35796 = n35795 ^ n34494 ^ n1527 ;
  assign n35797 = ( n2023 & n5867 ) | ( n2023 & ~n20367 ) | ( n5867 & ~n20367 ) ;
  assign n35798 = n20488 | n35797 ;
  assign n35799 = n35798 ^ n18675 ^ 1'b0 ;
  assign n35800 = ( n12904 & n23376 ) | ( n12904 & n29550 ) | ( n23376 & n29550 ) ;
  assign n35801 = n35800 ^ n24800 ^ n6099 ;
  assign n35802 = n11668 ^ n414 ^ 1'b0 ;
  assign n35803 = ~n1960 & n35802 ;
  assign n35804 = ~n12971 & n35803 ;
  assign n35805 = ( n1195 & n24835 ) | ( n1195 & ~n35804 ) | ( n24835 & ~n35804 ) ;
  assign n35809 = n365 & ~n4010 ;
  assign n35807 = ( n9032 & n31406 ) | ( n9032 & ~n34069 ) | ( n31406 & ~n34069 ) ;
  assign n35806 = ( n10511 & n28210 ) | ( n10511 & n31271 ) | ( n28210 & n31271 ) ;
  assign n35808 = n35807 ^ n35806 ^ n33356 ;
  assign n35810 = n35809 ^ n35808 ^ n32606 ;
  assign n35811 = n6118 ^ n3881 ^ 1'b0 ;
  assign n35812 = ~n7548 & n35811 ;
  assign n35813 = n35812 ^ n30189 ^ n15333 ;
  assign n35814 = n34791 ^ n8932 ^ n4054 ;
  assign n35815 = n35814 ^ n6001 ^ n4442 ;
  assign n35816 = n3121 & n35815 ;
  assign n35817 = n35816 ^ n4159 ^ 1'b0 ;
  assign n35818 = ( n3807 & n7048 ) | ( n3807 & ~n18758 ) | ( n7048 & ~n18758 ) ;
  assign n35819 = n35818 ^ n24416 ^ 1'b0 ;
  assign n35820 = n28966 | n35819 ;
  assign n35821 = n23797 ^ n22101 ^ n14180 ;
  assign n35822 = n20375 ^ n18103 ^ n11212 ;
  assign n35830 = n27939 ^ n16246 ^ n7466 ;
  assign n35828 = ( n4625 & n5710 ) | ( n4625 & n15109 ) | ( n5710 & n15109 ) ;
  assign n35823 = ( n12131 & ~n13309 ) | ( n12131 & n23706 ) | ( ~n13309 & n23706 ) ;
  assign n35824 = ( ~n2767 & n24873 ) | ( ~n2767 & n35823 ) | ( n24873 & n35823 ) ;
  assign n35825 = ( n1817 & n2219 ) | ( n1817 & ~n16202 ) | ( n2219 & ~n16202 ) ;
  assign n35826 = n19786 & n35825 ;
  assign n35827 = ( ~n9482 & n35824 ) | ( ~n9482 & n35826 ) | ( n35824 & n35826 ) ;
  assign n35829 = n35828 ^ n35827 ^ n13477 ;
  assign n35831 = n35830 ^ n35829 ^ n25605 ;
  assign n35832 = n24244 ^ n23699 ^ n5923 ;
  assign n35833 = ( x17 & ~n35077 ) | ( x17 & n35832 ) | ( ~n35077 & n35832 ) ;
  assign n35834 = n3998 & n11048 ;
  assign n35835 = n35834 ^ n26949 ^ 1'b0 ;
  assign n35836 = n35835 ^ n27119 ^ n19660 ;
  assign n35837 = n27317 ^ n27251 ^ n25194 ;
  assign n35838 = ( n4093 & ~n5287 ) | ( n4093 & n9729 ) | ( ~n5287 & n9729 ) ;
  assign n35839 = n35838 ^ n18561 ^ n7998 ;
  assign n35840 = n35839 ^ n26792 ^ n8281 ;
  assign n35841 = n18184 & n35840 ;
  assign n35842 = n35841 ^ n9927 ^ 1'b0 ;
  assign n35843 = n35842 ^ n24536 ^ 1'b0 ;
  assign n35844 = ( n3949 & n28781 ) | ( n3949 & ~n35843 ) | ( n28781 & ~n35843 ) ;
  assign n35845 = n21973 ^ n19244 ^ n4668 ;
  assign n35853 = ~n25816 & n30985 ;
  assign n35854 = ~n17833 & n35853 ;
  assign n35855 = n35854 ^ n7492 ^ n3233 ;
  assign n35846 = n13762 ^ n9624 ^ 1'b0 ;
  assign n35847 = n35846 ^ n16937 ^ n13477 ;
  assign n35848 = n35847 ^ n1053 ^ 1'b0 ;
  assign n35849 = n19353 ^ n16622 ^ 1'b0 ;
  assign n35850 = n8030 & ~n35849 ;
  assign n35851 = n35850 ^ n29119 ^ n6758 ;
  assign n35852 = ( n12386 & ~n35848 ) | ( n12386 & n35851 ) | ( ~n35848 & n35851 ) ;
  assign n35856 = n35855 ^ n35852 ^ n31329 ;
  assign n35857 = ( n2370 & n3374 ) | ( n2370 & ~n25025 ) | ( n3374 & ~n25025 ) ;
  assign n35858 = n35857 ^ n28984 ^ n28948 ;
  assign n35859 = n7793 & n9164 ;
  assign n35860 = ( n1530 & ~n7861 ) | ( n1530 & n16592 ) | ( ~n7861 & n16592 ) ;
  assign n35861 = ( ~n2174 & n10122 ) | ( ~n2174 & n11438 ) | ( n10122 & n11438 ) ;
  assign n35862 = n35860 & ~n35861 ;
  assign n35863 = ( n3135 & n10535 ) | ( n3135 & n15501 ) | ( n10535 & n15501 ) ;
  assign n35864 = ~n4679 & n28026 ;
  assign n35865 = n22075 ^ n13874 ^ n13204 ;
  assign n35866 = n17917 ^ n14919 ^ n9372 ;
  assign n35867 = n18382 & n35866 ;
  assign n35868 = ( n14878 & n35865 ) | ( n14878 & n35867 ) | ( n35865 & n35867 ) ;
  assign n35869 = ( n5480 & n5901 ) | ( n5480 & n35868 ) | ( n5901 & n35868 ) ;
  assign n35870 = ~n6645 & n14489 ;
  assign n35872 = n6496 ^ n3592 ^ x218 ;
  assign n35873 = n35872 ^ n17560 ^ 1'b0 ;
  assign n35874 = n3552 | n35873 ;
  assign n35871 = n9649 ^ n6662 ^ n3886 ;
  assign n35875 = n35874 ^ n35871 ^ n24819 ;
  assign n35876 = n35875 ^ n22746 ^ n10908 ;
  assign n35877 = n35876 ^ n16288 ^ 1'b0 ;
  assign n35878 = ~n35870 & n35877 ;
  assign n35879 = ( n5997 & ~n13972 ) | ( n5997 & n30148 ) | ( ~n13972 & n30148 ) ;
  assign n35880 = n14861 ^ n13958 ^ n11353 ;
  assign n35881 = n35880 ^ n7120 ^ n801 ;
  assign n35882 = n5574 & n35881 ;
  assign n35883 = n12654 ^ n11791 ^ n10279 ;
  assign n35884 = n35883 ^ n35293 ^ n21635 ;
  assign n35885 = ( n14243 & n27526 ) | ( n14243 & n35884 ) | ( n27526 & n35884 ) ;
  assign n35886 = n24699 ^ n13299 ^ n9523 ;
  assign n35887 = n29117 ^ n28982 ^ n2403 ;
  assign n35891 = ( n681 & n8095 ) | ( n681 & n15960 ) | ( n8095 & n15960 ) ;
  assign n35890 = ( n1643 & n6381 ) | ( n1643 & n17684 ) | ( n6381 & n17684 ) ;
  assign n35888 = n12205 ^ n7417 ^ n3486 ;
  assign n35889 = ( ~n2593 & n16271 ) | ( ~n2593 & n35888 ) | ( n16271 & n35888 ) ;
  assign n35892 = n35891 ^ n35890 ^ n35889 ;
  assign n35893 = ( n2970 & ~n9056 ) | ( n2970 & n35892 ) | ( ~n9056 & n35892 ) ;
  assign n35894 = ( n2815 & ~n3283 ) | ( n2815 & n11827 ) | ( ~n3283 & n11827 ) ;
  assign n35895 = n35894 ^ n31369 ^ n4378 ;
  assign n35896 = ( n10192 & n12715 ) | ( n10192 & n33724 ) | ( n12715 & n33724 ) ;
  assign n35897 = ( n2415 & n29313 ) | ( n2415 & ~n35896 ) | ( n29313 & ~n35896 ) ;
  assign n35898 = n20490 ^ n9969 ^ n2728 ;
  assign n35899 = n35898 ^ n23645 ^ 1'b0 ;
  assign n35900 = n35664 ^ n10530 ^ n881 ;
  assign n35901 = n19314 & ~n34545 ;
  assign n35902 = n30437 ^ n9594 ^ 1'b0 ;
  assign n35903 = n34000 | n35902 ;
  assign n35904 = n35903 ^ n26370 ^ n3248 ;
  assign n35905 = n18055 ^ n2664 ^ n2316 ;
  assign n35908 = ~n3768 & n8370 ;
  assign n35906 = n31972 ^ n5908 ^ n5907 ;
  assign n35907 = n35906 ^ n13638 ^ n9358 ;
  assign n35909 = n35908 ^ n35907 ^ n24242 ;
  assign n35910 = ( n14766 & ~n16288 ) | ( n14766 & n19541 ) | ( ~n16288 & n19541 ) ;
  assign n35911 = n23394 ^ n19009 ^ n14869 ;
  assign n35912 = n13045 ^ n8852 ^ n4067 ;
  assign n35913 = n1083 & n35912 ;
  assign n35914 = n35913 ^ n22582 ^ 1'b0 ;
  assign n35915 = ( n35910 & n35911 ) | ( n35910 & n35914 ) | ( n35911 & n35914 ) ;
  assign n35916 = n35915 ^ n11061 ^ n3350 ;
  assign n35917 = n34993 ^ n17829 ^ n3899 ;
  assign n35918 = ( n1686 & n30961 ) | ( n1686 & ~n35917 ) | ( n30961 & ~n35917 ) ;
  assign n35919 = ( ~n20554 & n26803 ) | ( ~n20554 & n35918 ) | ( n26803 & n35918 ) ;
  assign n35920 = n11083 ^ n4656 ^ x36 ;
  assign n35921 = n35920 ^ n24391 ^ n2389 ;
  assign n35922 = n21521 ^ n13200 ^ 1'b0 ;
  assign n35923 = ~n6969 & n35922 ;
  assign n35924 = n26803 & n29009 ;
  assign n35925 = n18679 & n35924 ;
  assign n35926 = ( ~n11531 & n12720 ) | ( ~n11531 & n17737 ) | ( n12720 & n17737 ) ;
  assign n35927 = n35926 ^ n15118 ^ n11613 ;
  assign n35928 = n8334 & n22313 ;
  assign n35929 = n35928 ^ n5283 ^ 1'b0 ;
  assign n35930 = n35929 ^ n13484 ^ n2233 ;
  assign n35931 = ( n16076 & n25895 ) | ( n16076 & n35930 ) | ( n25895 & n35930 ) ;
  assign n35932 = ~n22901 & n28247 ;
  assign n35933 = ~n1446 & n35932 ;
  assign n35934 = n35933 ^ n11181 ^ n2883 ;
  assign n35935 = n3457 & n12815 ;
  assign n35945 = n26287 ^ n16376 ^ n1304 ;
  assign n35946 = n35945 ^ n2966 ^ 1'b0 ;
  assign n35943 = n22718 ^ n16984 ^ 1'b0 ;
  assign n35944 = n15698 | n35943 ;
  assign n35938 = ( n5339 & n8757 ) | ( n5339 & ~n13293 ) | ( n8757 & ~n13293 ) ;
  assign n35937 = n9298 ^ n3848 ^ n2470 ;
  assign n35939 = n35938 ^ n35937 ^ 1'b0 ;
  assign n35936 = n6785 ^ n6623 ^ 1'b0 ;
  assign n35940 = n35939 ^ n35936 ^ n1155 ;
  assign n35941 = ~n8942 & n35940 ;
  assign n35942 = n35941 ^ n31583 ^ 1'b0 ;
  assign n35947 = n35946 ^ n35944 ^ n35942 ;
  assign n35948 = n35947 ^ n34153 ^ n6991 ;
  assign n35949 = n19250 ^ n7519 ^ n7378 ;
  assign n35950 = n35949 ^ n14450 ^ 1'b0 ;
  assign n35951 = n35950 ^ n21222 ^ n14057 ;
  assign n35952 = n22796 ^ n18008 ^ 1'b0 ;
  assign n35953 = n32506 ^ n27811 ^ n2271 ;
  assign n35954 = n34200 ^ n29388 ^ n760 ;
  assign n35955 = ( n812 & n24133 ) | ( n812 & n30691 ) | ( n24133 & n30691 ) ;
  assign n35956 = n14982 & n16327 ;
  assign n35957 = ( ~n35954 & n35955 ) | ( ~n35954 & n35956 ) | ( n35955 & n35956 ) ;
  assign n35960 = n22059 ^ n14114 ^ n8727 ;
  assign n35958 = n19459 ^ n16452 ^ n6037 ;
  assign n35959 = n35958 ^ n6709 ^ n4070 ;
  assign n35961 = n35960 ^ n35959 ^ n8768 ;
  assign n35962 = n25647 ^ n2770 ^ 1'b0 ;
  assign n35963 = n35962 ^ n19625 ^ n2015 ;
  assign n35964 = n27026 ^ n2923 ^ 1'b0 ;
  assign n35965 = n35963 & ~n35964 ;
  assign n35967 = ( n6728 & ~n14187 ) | ( n6728 & n20545 ) | ( ~n14187 & n20545 ) ;
  assign n35966 = n9063 ^ n4374 ^ n806 ;
  assign n35968 = n35967 ^ n35966 ^ n3244 ;
  assign n35969 = n17290 ^ n870 ^ 1'b0 ;
  assign n35970 = n14803 | n35969 ;
  assign n35971 = ( n1089 & ~n3019 ) | ( n1089 & n12559 ) | ( ~n3019 & n12559 ) ;
  assign n35972 = ~n15452 & n16637 ;
  assign n35973 = ( n3749 & n21518 ) | ( n3749 & n35972 ) | ( n21518 & n35972 ) ;
  assign n35974 = ( n15022 & n18578 ) | ( n15022 & ~n35973 ) | ( n18578 & ~n35973 ) ;
  assign n35975 = ( n35970 & n35971 ) | ( n35970 & n35974 ) | ( n35971 & n35974 ) ;
  assign n35976 = n16785 ^ n16034 ^ n715 ;
  assign n35977 = ( n5562 & n17316 ) | ( n5562 & ~n35976 ) | ( n17316 & ~n35976 ) ;
  assign n35978 = n14952 ^ n8661 ^ n4229 ;
  assign n35979 = ( ~n6737 & n7205 ) | ( ~n6737 & n35978 ) | ( n7205 & n35978 ) ;
  assign n35980 = n35979 ^ n27413 ^ n21260 ;
  assign n35981 = ( n4326 & n24592 ) | ( n4326 & ~n35980 ) | ( n24592 & ~n35980 ) ;
  assign n35982 = n7991 & n29445 ;
  assign n35983 = n35982 ^ n10493 ^ n295 ;
  assign n35984 = ( ~n2572 & n7738 ) | ( ~n2572 & n8584 ) | ( n7738 & n8584 ) ;
  assign n35988 = n23149 ^ n15817 ^ n8078 ;
  assign n35989 = n25570 & n35988 ;
  assign n35990 = n35989 ^ n10937 ^ 1'b0 ;
  assign n35985 = ~n7217 & n22400 ;
  assign n35986 = ~n21691 & n35985 ;
  assign n35987 = n16252 | n35986 ;
  assign n35991 = n35990 ^ n35987 ^ 1'b0 ;
  assign n35992 = n35991 ^ n29792 ^ n6502 ;
  assign n35993 = ~n3334 & n24986 ;
  assign n35994 = n35993 ^ n11413 ^ 1'b0 ;
  assign n35995 = ( n8561 & n19445 ) | ( n8561 & ~n35994 ) | ( n19445 & ~n35994 ) ;
  assign n35996 = n35995 ^ n21631 ^ n296 ;
  assign n35997 = ( n6303 & ~n6461 ) | ( n6303 & n9591 ) | ( ~n6461 & n9591 ) ;
  assign n35998 = ( n4905 & n15941 ) | ( n4905 & n35997 ) | ( n15941 & n35997 ) ;
  assign n35999 = ( n16092 & ~n35996 ) | ( n16092 & n35998 ) | ( ~n35996 & n35998 ) ;
  assign n36001 = ~n6437 & n7984 ;
  assign n36002 = n36001 ^ n17641 ^ 1'b0 ;
  assign n36000 = n21478 ^ n18702 ^ n6382 ;
  assign n36003 = n36002 ^ n36000 ^ 1'b0 ;
  assign n36004 = ( n6007 & n6202 ) | ( n6007 & ~n11822 ) | ( n6202 & ~n11822 ) ;
  assign n36005 = ( n5805 & ~n15668 ) | ( n5805 & n20597 ) | ( ~n15668 & n20597 ) ;
  assign n36006 = ~n36004 & n36005 ;
  assign n36007 = ~n5184 & n36006 ;
  assign n36008 = n30848 ^ n30038 ^ n2292 ;
  assign n36009 = ( n3483 & n20308 ) | ( n3483 & n22665 ) | ( n20308 & n22665 ) ;
  assign n36010 = n36009 ^ n21485 ^ 1'b0 ;
  assign n36011 = n20104 ^ n6600 ^ n2250 ;
  assign n36012 = n36011 ^ n12524 ^ 1'b0 ;
  assign n36013 = n5946 & n14227 ;
  assign n36014 = ~n10135 & n36013 ;
  assign n36015 = n36014 ^ n775 ^ 1'b0 ;
  assign n36016 = ( ~n5910 & n9907 ) | ( ~n5910 & n14336 ) | ( n9907 & n14336 ) ;
  assign n36017 = ( n8431 & ~n15242 ) | ( n8431 & n17844 ) | ( ~n15242 & n17844 ) ;
  assign n36018 = ( n14979 & ~n36016 ) | ( n14979 & n36017 ) | ( ~n36016 & n36017 ) ;
  assign n36019 = ( n25815 & n36015 ) | ( n25815 & n36018 ) | ( n36015 & n36018 ) ;
  assign n36020 = ( n9554 & n22097 ) | ( n9554 & n36019 ) | ( n22097 & n36019 ) ;
  assign n36021 = ( n3251 & n19979 ) | ( n3251 & ~n25301 ) | ( n19979 & ~n25301 ) ;
  assign n36022 = n33826 ^ n21083 ^ n15760 ;
  assign n36023 = n21291 & n36022 ;
  assign n36024 = ~n36021 & n36023 ;
  assign n36025 = ( n507 & ~n32312 ) | ( n507 & n34633 ) | ( ~n32312 & n34633 ) ;
  assign n36028 = n2512 ^ n1834 ^ n648 ;
  assign n36027 = ( n1783 & n2968 ) | ( n1783 & n30806 ) | ( n2968 & n30806 ) ;
  assign n36029 = n36028 ^ n36027 ^ n13365 ;
  assign n36026 = n975 & n4213 ;
  assign n36030 = n36029 ^ n36026 ^ 1'b0 ;
  assign n36031 = ( n12916 & ~n23647 ) | ( n12916 & n36030 ) | ( ~n23647 & n36030 ) ;
  assign n36032 = n9133 & ~n14056 ;
  assign n36033 = ~n953 & n36032 ;
  assign n36034 = n23366 ^ n9197 ^ 1'b0 ;
  assign n36035 = n6538 & n36034 ;
  assign n36036 = n36035 ^ n22662 ^ n18195 ;
  assign n36037 = ( n657 & n36033 ) | ( n657 & n36036 ) | ( n36033 & n36036 ) ;
  assign n36038 = ( n1932 & n6072 ) | ( n1932 & n11117 ) | ( n6072 & n11117 ) ;
  assign n36039 = ( ~n22179 & n26456 ) | ( ~n22179 & n28664 ) | ( n26456 & n28664 ) ;
  assign n36040 = n36039 ^ n17389 ^ n8833 ;
  assign n36041 = ( n24123 & n36038 ) | ( n24123 & n36040 ) | ( n36038 & n36040 ) ;
  assign n36042 = n10924 ^ n4859 ^ n2245 ;
  assign n36043 = n9398 | n21793 ;
  assign n36045 = ~n6340 & n6560 ;
  assign n36046 = n36045 ^ n12965 ^ 1'b0 ;
  assign n36044 = ( ~n2298 & n4823 ) | ( ~n2298 & n24733 ) | ( n4823 & n24733 ) ;
  assign n36047 = n36046 ^ n36044 ^ n8910 ;
  assign n36048 = n27667 ^ n15399 ^ n8070 ;
  assign n36049 = ( n5841 & ~n28455 ) | ( n5841 & n36048 ) | ( ~n28455 & n36048 ) ;
  assign n36050 = ( n9999 & n14887 ) | ( n9999 & ~n29193 ) | ( n14887 & ~n29193 ) ;
  assign n36051 = ~n8556 & n16744 ;
  assign n36052 = ( n18160 & ~n19671 ) | ( n18160 & n36051 ) | ( ~n19671 & n36051 ) ;
  assign n36053 = ( ~n1632 & n2822 ) | ( ~n1632 & n16272 ) | ( n2822 & n16272 ) ;
  assign n36054 = n6837 & n24990 ;
  assign n36055 = n36054 ^ n35857 ^ 1'b0 ;
  assign n36056 = n20714 | n24951 ;
  assign n36057 = n10230 | n36056 ;
  assign n36058 = n36057 ^ n32917 ^ n30849 ;
  assign n36059 = n23458 ^ n21356 ^ n18868 ;
  assign n36060 = ( n22624 & ~n36058 ) | ( n22624 & n36059 ) | ( ~n36058 & n36059 ) ;
  assign n36062 = ~n2181 & n20724 ;
  assign n36063 = n10744 & n36062 ;
  assign n36061 = ( n5844 & n15056 ) | ( n5844 & ~n20020 ) | ( n15056 & ~n20020 ) ;
  assign n36064 = n36063 ^ n36061 ^ n10415 ;
  assign n36065 = ( ~n898 & n7135 ) | ( ~n898 & n11159 ) | ( n7135 & n11159 ) ;
  assign n36066 = n14085 ^ n11084 ^ 1'b0 ;
  assign n36067 = ~n36065 & n36066 ;
  assign n36068 = ( n5652 & n16930 ) | ( n5652 & n36067 ) | ( n16930 & n36067 ) ;
  assign n36069 = ( n26439 & n31720 ) | ( n26439 & ~n36068 ) | ( n31720 & ~n36068 ) ;
  assign n36070 = n16071 ^ n11159 ^ n2959 ;
  assign n36071 = n18007 ^ n15333 ^ n6405 ;
  assign n36072 = n29465 ^ n13719 ^ n5965 ;
  assign n36073 = n4458 ^ n4287 ^ 1'b0 ;
  assign n36074 = n8078 ^ n7619 ^ n5272 ;
  assign n36075 = ( n10003 & ~n21502 ) | ( n10003 & n26279 ) | ( ~n21502 & n26279 ) ;
  assign n36076 = ( n1559 & n36074 ) | ( n1559 & n36075 ) | ( n36074 & n36075 ) ;
  assign n36077 = ( n17288 & n17475 ) | ( n17288 & ~n25552 ) | ( n17475 & ~n25552 ) ;
  assign n36078 = n34438 ^ n26477 ^ n17415 ;
  assign n36079 = n23611 | n26532 ;
  assign n36080 = n36079 ^ n18516 ^ 1'b0 ;
  assign n36081 = ( ~n2336 & n19170 ) | ( ~n2336 & n36080 ) | ( n19170 & n36080 ) ;
  assign n36082 = n31397 ^ n31236 ^ n21018 ;
  assign n36083 = ( n10158 & n28498 ) | ( n10158 & n36082 ) | ( n28498 & n36082 ) ;
  assign n36084 = n36083 ^ n27745 ^ n16128 ;
  assign n36085 = n28483 ^ n23912 ^ n4584 ;
  assign n36086 = ( n15749 & n24133 ) | ( n15749 & n35212 ) | ( n24133 & n35212 ) ;
  assign n36087 = ( n2156 & ~n34029 ) | ( n2156 & n36086 ) | ( ~n34029 & n36086 ) ;
  assign n36088 = ( n8747 & n36085 ) | ( n8747 & ~n36087 ) | ( n36085 & ~n36087 ) ;
  assign n36089 = n36088 ^ n16449 ^ n7649 ;
  assign n36091 = n23083 ^ n20037 ^ n8913 ;
  assign n36090 = ( x236 & ~n9587 ) | ( x236 & n19320 ) | ( ~n9587 & n19320 ) ;
  assign n36092 = n36091 ^ n36090 ^ n12457 ;
  assign n36093 = ( n1911 & n29932 ) | ( n1911 & n36092 ) | ( n29932 & n36092 ) ;
  assign n36094 = n36093 ^ n35738 ^ n4502 ;
  assign n36095 = n28853 ^ n17378 ^ n7814 ;
  assign n36096 = n12585 ^ n11683 ^ n8607 ;
  assign n36097 = ( n14594 & n30897 ) | ( n14594 & n36096 ) | ( n30897 & n36096 ) ;
  assign n36098 = ( n20041 & n36095 ) | ( n20041 & ~n36097 ) | ( n36095 & ~n36097 ) ;
  assign n36099 = ( ~n2572 & n27141 ) | ( ~n2572 & n29996 ) | ( n27141 & n29996 ) ;
  assign n36100 = n36099 ^ n33143 ^ n8308 ;
  assign n36101 = ( n21072 & n30393 ) | ( n21072 & ~n36100 ) | ( n30393 & ~n36100 ) ;
  assign n36102 = n24042 ^ n9719 ^ n8495 ;
  assign n36103 = ( n13432 & n14485 ) | ( n13432 & ~n36102 ) | ( n14485 & ~n36102 ) ;
  assign n36104 = ( n11824 & n23529 ) | ( n11824 & n27637 ) | ( n23529 & n27637 ) ;
  assign n36105 = n36104 ^ n16082 ^ 1'b0 ;
  assign n36106 = n36105 ^ n27612 ^ n25709 ;
  assign n36107 = n35106 ^ n13239 ^ 1'b0 ;
  assign n36108 = ( n5411 & ~n36106 ) | ( n5411 & n36107 ) | ( ~n36106 & n36107 ) ;
  assign n36110 = n19952 ^ n6857 ^ n6680 ;
  assign n36109 = n11906 ^ n11404 ^ n1489 ;
  assign n36111 = n36110 ^ n36109 ^ n6013 ;
  assign n36112 = n7783 ^ n7100 ^ n2711 ;
  assign n36113 = ( n1991 & ~n30486 ) | ( n1991 & n36112 ) | ( ~n30486 & n36112 ) ;
  assign n36114 = ( n3115 & n25113 ) | ( n3115 & ~n30528 ) | ( n25113 & ~n30528 ) ;
  assign n36115 = n19980 ^ n10985 ^ 1'b0 ;
  assign n36116 = x119 & n36115 ;
  assign n36117 = n24480 ^ n20628 ^ n5314 ;
  assign n36118 = n25496 ^ n24493 ^ 1'b0 ;
  assign n36119 = ( n7014 & n14933 ) | ( n7014 & ~n25110 ) | ( n14933 & ~n25110 ) ;
  assign n36120 = n11433 ^ n6829 ^ n1384 ;
  assign n36121 = n36120 ^ n32666 ^ x0 ;
  assign n36123 = n22022 ^ n12281 ^ n8669 ;
  assign n36124 = ~n8318 & n13259 ;
  assign n36125 = n36124 ^ n3898 ^ 1'b0 ;
  assign n36126 = n28548 & ~n36125 ;
  assign n36127 = ~n36123 & n36126 ;
  assign n36122 = n2278 & ~n3304 ;
  assign n36128 = n36127 ^ n36122 ^ 1'b0 ;
  assign n36129 = ( n5172 & ~n22047 ) | ( n5172 & n27142 ) | ( ~n22047 & n27142 ) ;
  assign n36130 = n36129 ^ n12652 ^ n1101 ;
  assign n36131 = n32570 ^ n23467 ^ 1'b0 ;
  assign n36132 = n13248 & ~n36131 ;
  assign n36133 = ( n11170 & ~n11992 ) | ( n11170 & n36132 ) | ( ~n11992 & n36132 ) ;
  assign n36134 = ( n11198 & ~n15196 ) | ( n11198 & n17739 ) | ( ~n15196 & n17739 ) ;
  assign n36135 = ( n27282 & ~n36133 ) | ( n27282 & n36134 ) | ( ~n36133 & n36134 ) ;
  assign n36136 = ~n4117 & n9520 ;
  assign n36137 = ( n8531 & ~n9800 ) | ( n8531 & n36136 ) | ( ~n9800 & n36136 ) ;
  assign n36138 = n36137 ^ n29020 ^ n12313 ;
  assign n36139 = n10588 & ~n25488 ;
  assign n36140 = ~n36138 & n36139 ;
  assign n36141 = ( n34929 & ~n36135 ) | ( n34929 & n36140 ) | ( ~n36135 & n36140 ) ;
  assign n36142 = n327 & ~n24370 ;
  assign n36143 = n36142 ^ n15690 ^ 1'b0 ;
  assign n36144 = n14515 & ~n15085 ;
  assign n36145 = n36144 ^ n21367 ^ 1'b0 ;
  assign n36146 = ~n14931 & n36145 ;
  assign n36147 = n567 | n28090 ;
  assign n36148 = n15943 & ~n36147 ;
  assign n36149 = n11770 ^ n2356 ^ n1586 ;
  assign n36150 = n36149 ^ n21116 ^ n14764 ;
  assign n36151 = ( ~n9821 & n36148 ) | ( ~n9821 & n36150 ) | ( n36148 & n36150 ) ;
  assign n36152 = ( ~n4939 & n8238 ) | ( ~n4939 & n8995 ) | ( n8238 & n8995 ) ;
  assign n36153 = ( n15220 & n33981 ) | ( n15220 & ~n36152 ) | ( n33981 & ~n36152 ) ;
  assign n36154 = n13960 ^ n7993 ^ n1442 ;
  assign n36155 = ( n4886 & n5013 ) | ( n4886 & ~n36154 ) | ( n5013 & ~n36154 ) ;
  assign n36156 = ( n22030 & n36153 ) | ( n22030 & n36155 ) | ( n36153 & n36155 ) ;
  assign n36157 = ( n1393 & n12373 ) | ( n1393 & ~n16015 ) | ( n12373 & ~n16015 ) ;
  assign n36158 = ( ~n9630 & n28531 ) | ( ~n9630 & n35995 ) | ( n28531 & n35995 ) ;
  assign n36159 = n36158 ^ n30636 ^ n23176 ;
  assign n36160 = n36159 ^ n24691 ^ n21407 ;
  assign n36161 = n4187 | n15878 ;
  assign n36162 = n7972 & ~n36161 ;
  assign n36163 = n3281 | n36162 ;
  assign n36164 = n32095 | n36163 ;
  assign n36165 = ( n2636 & n10646 ) | ( n2636 & n21168 ) | ( n10646 & n21168 ) ;
  assign n36166 = ( n12890 & n36164 ) | ( n12890 & n36165 ) | ( n36164 & n36165 ) ;
  assign n36167 = n36166 ^ n5820 ^ n1064 ;
  assign n36168 = n20662 ^ n10915 ^ n669 ;
  assign n36169 = n36168 ^ n17747 ^ n17456 ;
  assign n36170 = n17402 ^ n11195 ^ n341 ;
  assign n36171 = ( n3796 & n18437 ) | ( n3796 & n36170 ) | ( n18437 & n36170 ) ;
  assign n36172 = n18569 ^ n14439 ^ n3323 ;
  assign n36173 = n32565 & n36172 ;
  assign n36174 = n17595 | n36173 ;
  assign n36175 = ( ~n5060 & n10717 ) | ( ~n5060 & n31038 ) | ( n10717 & n31038 ) ;
  assign n36176 = ( n5781 & ~n7303 ) | ( n5781 & n8129 ) | ( ~n7303 & n8129 ) ;
  assign n36177 = ( n5801 & n36175 ) | ( n5801 & ~n36176 ) | ( n36175 & ~n36176 ) ;
  assign n36178 = ( n36171 & ~n36174 ) | ( n36171 & n36177 ) | ( ~n36174 & n36177 ) ;
  assign n36182 = n23899 ^ n17271 ^ n1165 ;
  assign n36179 = n27654 ^ n23377 ^ n1115 ;
  assign n36180 = n17418 | n36179 ;
  assign n36181 = n20162 & ~n36180 ;
  assign n36183 = n36182 ^ n36181 ^ n15125 ;
  assign n36184 = n23734 ^ n14859 ^ n12809 ;
  assign n36185 = n15410 & n34560 ;
  assign n36186 = ( n22728 & n23684 ) | ( n22728 & n23905 ) | ( n23684 & n23905 ) ;
  assign n36187 = ( n612 & n25220 ) | ( n612 & n30706 ) | ( n25220 & n30706 ) ;
  assign n36188 = ( n9865 & n24953 ) | ( n9865 & n30861 ) | ( n24953 & n30861 ) ;
  assign n36189 = n31551 | n36188 ;
  assign n36190 = n33026 ^ n8212 ^ n1187 ;
  assign n36191 = n29142 ^ n17785 ^ 1'b0 ;
  assign n36192 = ~n10448 & n36191 ;
  assign n36193 = n1772 & n36192 ;
  assign n36194 = ( ~n2801 & n20843 ) | ( ~n2801 & n36193 ) | ( n20843 & n36193 ) ;
  assign n36195 = n6840 | n16875 ;
  assign n36196 = ( n275 & n13893 ) | ( n275 & ~n21341 ) | ( n13893 & ~n21341 ) ;
  assign n36197 = n36196 ^ n8922 ^ n7994 ;
  assign n36198 = n36197 ^ n22755 ^ n15685 ;
  assign n36199 = ( n12165 & ~n36195 ) | ( n12165 & n36198 ) | ( ~n36195 & n36198 ) ;
  assign n36200 = ( ~n17172 & n20109 ) | ( ~n17172 & n33594 ) | ( n20109 & n33594 ) ;
  assign n36203 = n33356 ^ n21842 ^ n4585 ;
  assign n36201 = n31787 ^ n21013 ^ 1'b0 ;
  assign n36202 = n27528 | n36201 ;
  assign n36204 = n36203 ^ n36202 ^ n6118 ;
  assign n36205 = n22769 ^ n15262 ^ n5760 ;
  assign n36207 = ( n5480 & ~n8178 ) | ( n5480 & n18529 ) | ( ~n8178 & n18529 ) ;
  assign n36206 = n8066 ^ n1790 ^ 1'b0 ;
  assign n36208 = n36207 ^ n36206 ^ n3038 ;
  assign n36209 = ( ~n14943 & n34217 ) | ( ~n14943 & n36208 ) | ( n34217 & n36208 ) ;
  assign n36210 = ( n4850 & ~n32947 ) | ( n4850 & n36209 ) | ( ~n32947 & n36209 ) ;
  assign n36211 = ( n20876 & ~n26528 ) | ( n20876 & n29828 ) | ( ~n26528 & n29828 ) ;
  assign n36212 = n19231 ^ n11564 ^ 1'b0 ;
  assign n36213 = ~n24950 & n36212 ;
  assign n36214 = n5287 & n10680 ;
  assign n36215 = n874 & ~n36214 ;
  assign n36216 = n23784 ^ n10267 ^ 1'b0 ;
  assign n36217 = ( ~n16288 & n19514 ) | ( ~n16288 & n32895 ) | ( n19514 & n32895 ) ;
  assign n36218 = ( n14070 & ~n18886 ) | ( n14070 & n23091 ) | ( ~n18886 & n23091 ) ;
  assign n36219 = n36218 ^ n33424 ^ n7842 ;
  assign n36220 = ( ~n20588 & n29425 ) | ( ~n20588 & n36219 ) | ( n29425 & n36219 ) ;
  assign n36221 = ( ~n5461 & n16942 ) | ( ~n5461 & n35228 ) | ( n16942 & n35228 ) ;
  assign n36222 = ( n494 & ~n13952 ) | ( n494 & n36221 ) | ( ~n13952 & n36221 ) ;
  assign n36223 = ( ~n3464 & n28748 ) | ( ~n3464 & n36222 ) | ( n28748 & n36222 ) ;
  assign n36224 = ( n4789 & n11217 ) | ( n4789 & n13198 ) | ( n11217 & n13198 ) ;
  assign n36225 = n14989 & n36224 ;
  assign n36226 = n873 & n36225 ;
  assign n36227 = n11895 ^ n10033 ^ n1328 ;
  assign n36228 = ( n19432 & ~n19904 ) | ( n19432 & n36227 ) | ( ~n19904 & n36227 ) ;
  assign n36229 = n19876 ^ n12667 ^ n8843 ;
  assign n36230 = n36229 ^ n28716 ^ n24513 ;
  assign n36231 = ( n5471 & n13369 ) | ( n5471 & ~n27189 ) | ( n13369 & ~n27189 ) ;
  assign n36234 = n19728 ^ n11136 ^ n2198 ;
  assign n36235 = n36234 ^ n20964 ^ n11093 ;
  assign n36232 = ( n2869 & n11181 ) | ( n2869 & n23226 ) | ( n11181 & n23226 ) ;
  assign n36233 = ( n33461 & ~n36224 ) | ( n33461 & n36232 ) | ( ~n36224 & n36232 ) ;
  assign n36236 = n36235 ^ n36233 ^ n4174 ;
  assign n36237 = n31326 ^ n5386 ^ n2438 ;
  assign n36241 = ( ~n2236 & n2922 ) | ( ~n2236 & n2966 ) | ( n2922 & n2966 ) ;
  assign n36240 = n25888 ^ n11673 ^ n4494 ;
  assign n36238 = n14172 ^ n3066 ^ 1'b0 ;
  assign n36239 = ( n2364 & n11045 ) | ( n2364 & ~n36238 ) | ( n11045 & ~n36238 ) ;
  assign n36242 = n36241 ^ n36240 ^ n36239 ;
  assign n36243 = ( x1 & n22394 ) | ( x1 & ~n34464 ) | ( n22394 & ~n34464 ) ;
  assign n36244 = n29964 ^ n7573 ^ n6626 ;
  assign n36246 = n14965 ^ n6512 ^ n2678 ;
  assign n36245 = n14045 ^ n10765 ^ n4224 ;
  assign n36247 = n36246 ^ n36245 ^ n741 ;
  assign n36248 = n34103 ^ n20996 ^ n19314 ;
  assign n36249 = ~n14643 & n20189 ;
  assign n36250 = ( n2226 & n9681 ) | ( n2226 & ~n36249 ) | ( n9681 & ~n36249 ) ;
  assign n36251 = n36250 ^ n13121 ^ n9919 ;
  assign n36252 = n21545 ^ n4445 ^ n652 ;
  assign n36253 = n36252 ^ n29857 ^ n8353 ;
  assign n36254 = n36253 ^ n24150 ^ n8012 ;
  assign n36255 = n9214 & ~n30379 ;
  assign n36256 = n36255 ^ n419 ^ 1'b0 ;
  assign n36257 = n23049 ^ n10878 ^ n8418 ;
  assign n36258 = n31613 & ~n36257 ;
  assign n36259 = ( ~n6698 & n11298 ) | ( ~n6698 & n12310 ) | ( n11298 & n12310 ) ;
  assign n36260 = ( n13729 & n23236 ) | ( n13729 & ~n27317 ) | ( n23236 & ~n27317 ) ;
  assign n36261 = n16950 ^ n9373 ^ n3311 ;
  assign n36262 = n19545 ^ n5614 ^ 1'b0 ;
  assign n36263 = ~n14752 & n36262 ;
  assign n36264 = n36263 ^ n5980 ^ 1'b0 ;
  assign n36265 = n29214 ^ n20431 ^ 1'b0 ;
  assign n36266 = n36264 | n36265 ;
  assign n36267 = ( ~n5655 & n5681 ) | ( ~n5655 & n17331 ) | ( n5681 & n17331 ) ;
  assign n36268 = n36267 ^ n24253 ^ n4927 ;
  assign n36269 = n13857 ^ n539 ^ 1'b0 ;
  assign n36270 = n2567 & ~n36269 ;
  assign n36271 = ( n8482 & n12942 ) | ( n8482 & ~n36270 ) | ( n12942 & ~n36270 ) ;
  assign n36272 = ( n14501 & n36268 ) | ( n14501 & n36271 ) | ( n36268 & n36271 ) ;
  assign n36273 = ( n10675 & n13373 ) | ( n10675 & n23753 ) | ( n13373 & n23753 ) ;
  assign n36274 = n33254 ^ n14998 ^ n5729 ;
  assign n36275 = n36274 ^ n17022 ^ n1747 ;
  assign n36276 = n36275 ^ n14324 ^ n5145 ;
  assign n36280 = ( n2827 & n5231 ) | ( n2827 & n11618 ) | ( n5231 & n11618 ) ;
  assign n36277 = n13376 ^ n13365 ^ n3483 ;
  assign n36278 = n13282 ^ x182 ^ 1'b0 ;
  assign n36279 = n36277 & n36278 ;
  assign n36281 = n36280 ^ n36279 ^ n6121 ;
  assign n36285 = ( ~n5877 & n15244 ) | ( ~n5877 & n24089 ) | ( n15244 & n24089 ) ;
  assign n36282 = ( n11012 & n19108 ) | ( n11012 & n21970 ) | ( n19108 & n21970 ) ;
  assign n36283 = n27399 ^ n17412 ^ 1'b0 ;
  assign n36284 = n36282 & ~n36283 ;
  assign n36286 = n36285 ^ n36284 ^ 1'b0 ;
  assign n36287 = ( n12861 & n21857 ) | ( n12861 & n36286 ) | ( n21857 & n36286 ) ;
  assign n36288 = n23091 ^ n9382 ^ 1'b0 ;
  assign n36289 = n36288 ^ n19242 ^ n1118 ;
  assign n36290 = ( n2879 & ~n28461 ) | ( n2879 & n29850 ) | ( ~n28461 & n29850 ) ;
  assign n36291 = n36290 ^ n8009 ^ n4460 ;
  assign n36292 = ( n478 & n11745 ) | ( n478 & n36291 ) | ( n11745 & n36291 ) ;
  assign n36293 = n26901 ^ n10694 ^ 1'b0 ;
  assign n36294 = n19450 ^ n3843 ^ x183 ;
  assign n36295 = n27518 ^ n15672 ^ n11912 ;
  assign n36296 = n36295 ^ n23843 ^ n11231 ;
  assign n36297 = ( n31719 & n33360 ) | ( n31719 & n36296 ) | ( n33360 & n36296 ) ;
  assign n36298 = n27519 ^ n25005 ^ n10275 ;
  assign n36299 = n18791 ^ n4137 ^ 1'b0 ;
  assign n36300 = n16389 & n36299 ;
  assign n36301 = ( ~n10319 & n22081 ) | ( ~n10319 & n33973 ) | ( n22081 & n33973 ) ;
  assign n36302 = ( n3440 & n3591 ) | ( n3440 & ~n18752 ) | ( n3591 & ~n18752 ) ;
  assign n36303 = n27410 ^ n9763 ^ n2345 ;
  assign n36304 = ( n8527 & n10517 ) | ( n8527 & ~n36303 ) | ( n10517 & ~n36303 ) ;
  assign n36305 = n36304 ^ n17092 ^ n13151 ;
  assign n36306 = ( n800 & ~n877 ) | ( n800 & n10239 ) | ( ~n877 & n10239 ) ;
  assign n36307 = ( n22847 & n36305 ) | ( n22847 & ~n36306 ) | ( n36305 & ~n36306 ) ;
  assign n36308 = ( n24506 & n36302 ) | ( n24506 & n36307 ) | ( n36302 & n36307 ) ;
  assign n36309 = n2098 & ~n27166 ;
  assign n36310 = n36309 ^ n1014 ^ 1'b0 ;
  assign n36311 = n15053 ^ n9222 ^ n6414 ;
  assign n36312 = n36311 ^ n26573 ^ n14117 ;
  assign n36313 = ( n2151 & n18897 ) | ( n2151 & n20945 ) | ( n18897 & n20945 ) ;
  assign n36314 = ( n36310 & n36312 ) | ( n36310 & n36313 ) | ( n36312 & n36313 ) ;
  assign n36315 = n11267 ^ n6874 ^ n3012 ;
  assign n36316 = n36315 ^ n5672 ^ n1211 ;
  assign n36317 = n36316 ^ n23042 ^ n15793 ;
  assign n36318 = ( ~n1537 & n20338 ) | ( ~n1537 & n24536 ) | ( n20338 & n24536 ) ;
  assign n36319 = ~n11771 & n33104 ;
  assign n36320 = n15288 & n36319 ;
  assign n36321 = n36320 ^ n20061 ^ n5600 ;
  assign n36322 = ( n11758 & n36318 ) | ( n11758 & n36321 ) | ( n36318 & n36321 ) ;
  assign n36323 = n22215 ^ n14026 ^ n11343 ;
  assign n36324 = n31446 ^ n29620 ^ 1'b0 ;
  assign n36325 = ( n23644 & n24348 ) | ( n23644 & n36324 ) | ( n24348 & n36324 ) ;
  assign n36326 = ( x1 & n16501 ) | ( x1 & n31909 ) | ( n16501 & n31909 ) ;
  assign n36327 = n20903 ^ n18299 ^ 1'b0 ;
  assign n36328 = ( n16122 & ~n20654 ) | ( n16122 & n36327 ) | ( ~n20654 & n36327 ) ;
  assign n36329 = n29169 ^ n16172 ^ n12323 ;
  assign n36330 = ( n4707 & n23028 ) | ( n4707 & ~n36329 ) | ( n23028 & ~n36329 ) ;
  assign n36331 = n14193 ^ n13688 ^ n3508 ;
  assign n36332 = ( n14422 & ~n36330 ) | ( n14422 & n36331 ) | ( ~n36330 & n36331 ) ;
  assign n36340 = ( n2700 & n7078 ) | ( n2700 & n10718 ) | ( n7078 & n10718 ) ;
  assign n36333 = n3212 & n13141 ;
  assign n36334 = ( n4977 & n17738 ) | ( n4977 & ~n31940 ) | ( n17738 & ~n31940 ) ;
  assign n36335 = ( ~n20400 & n27041 ) | ( ~n20400 & n36334 ) | ( n27041 & n36334 ) ;
  assign n36336 = n36335 ^ n17526 ^ n17423 ;
  assign n36337 = ( n18462 & n23122 ) | ( n18462 & ~n36336 ) | ( n23122 & ~n36336 ) ;
  assign n36338 = ( ~n4784 & n36333 ) | ( ~n4784 & n36337 ) | ( n36333 & n36337 ) ;
  assign n36339 = n36338 ^ n17301 ^ n11014 ;
  assign n36341 = n36340 ^ n36339 ^ n19324 ;
  assign n36342 = n15397 ^ n5445 ^ n5038 ;
  assign n36343 = n36342 ^ n17580 ^ n13438 ;
  assign n36345 = ( n6901 & ~n23282 ) | ( n6901 & n31479 ) | ( ~n23282 & n31479 ) ;
  assign n36344 = ~n11867 & n12976 ;
  assign n36346 = n36345 ^ n36344 ^ 1'b0 ;
  assign n36347 = ( n10680 & ~n19847 ) | ( n10680 & n27771 ) | ( ~n19847 & n27771 ) ;
  assign n36348 = n36347 ^ n32419 ^ n28543 ;
  assign n36349 = n31350 ^ n29451 ^ n11821 ;
  assign n36350 = n7978 ^ n5694 ^ n2133 ;
  assign n36351 = ( n1862 & n16008 ) | ( n1862 & n36350 ) | ( n16008 & n36350 ) ;
  assign n36352 = ( ~n2203 & n15429 ) | ( ~n2203 & n29273 ) | ( n15429 & n29273 ) ;
  assign n36353 = ( n15699 & ~n36351 ) | ( n15699 & n36352 ) | ( ~n36351 & n36352 ) ;
  assign n36359 = ( n699 & ~n2250 ) | ( n699 & n30170 ) | ( ~n2250 & n30170 ) ;
  assign n36356 = n25235 ^ n18116 ^ n7886 ;
  assign n36354 = n3642 & ~n25477 ;
  assign n36355 = n16144 & n36354 ;
  assign n36357 = n36356 ^ n36355 ^ n3425 ;
  assign n36358 = n36357 ^ n24447 ^ n21986 ;
  assign n36360 = n36359 ^ n36358 ^ n2845 ;
  assign n36361 = n36360 ^ n31477 ^ n29298 ;
  assign n36362 = n10676 | n30170 ;
  assign n36363 = ( ~n9143 & n14926 ) | ( ~n9143 & n35153 ) | ( n14926 & n35153 ) ;
  assign n36367 = ( n1105 & ~n15103 ) | ( n1105 & n18310 ) | ( ~n15103 & n18310 ) ;
  assign n36364 = n26234 ^ n18583 ^ n7754 ;
  assign n36365 = ( ~n2029 & n11292 ) | ( ~n2029 & n18428 ) | ( n11292 & n18428 ) ;
  assign n36366 = ~n36364 & n36365 ;
  assign n36368 = n36367 ^ n36366 ^ 1'b0 ;
  assign n36369 = n36368 ^ n15880 ^ 1'b0 ;
  assign n36370 = n36363 | n36369 ;
  assign n36371 = ( n3861 & n22714 ) | ( n3861 & n34037 ) | ( n22714 & n34037 ) ;
  assign n36374 = n12988 ^ n995 ^ x194 ;
  assign n36375 = n36374 ^ n5239 ^ n4676 ;
  assign n36372 = n15593 ^ n9052 ^ n8692 ;
  assign n36373 = n36372 ^ n32211 ^ n1824 ;
  assign n36376 = n36375 ^ n36373 ^ n33066 ;
  assign n36377 = ( n7397 & n25664 ) | ( n7397 & n36376 ) | ( n25664 & n36376 ) ;
  assign n36378 = ( n10579 & n20697 ) | ( n10579 & ~n36377 ) | ( n20697 & ~n36377 ) ;
  assign n36379 = ( ~n7525 & n10197 ) | ( ~n7525 & n36378 ) | ( n10197 & n36378 ) ;
  assign n36384 = n17440 ^ n8386 ^ n1166 ;
  assign n36382 = n2996 ^ n2699 ^ n858 ;
  assign n36380 = n14410 ^ n10779 ^ n1397 ;
  assign n36381 = ( n21262 & n31219 ) | ( n21262 & n36380 ) | ( n31219 & n36380 ) ;
  assign n36383 = n36382 ^ n36381 ^ n15363 ;
  assign n36385 = n36384 ^ n36383 ^ n6650 ;
  assign n36386 = n11540 & ~n26343 ;
  assign n36387 = n23216 & n36386 ;
  assign n36388 = ( n3790 & ~n21468 ) | ( n3790 & n24074 ) | ( ~n21468 & n24074 ) ;
  assign n36389 = ( n2256 & n6827 ) | ( n2256 & n36388 ) | ( n6827 & n36388 ) ;
  assign n36390 = n36389 ^ n9287 ^ 1'b0 ;
  assign n36391 = n2553 & ~n36390 ;
  assign n36393 = n14502 ^ n8890 ^ n5441 ;
  assign n36392 = n9771 ^ n6327 ^ 1'b0 ;
  assign n36394 = n36393 ^ n36392 ^ n26007 ;
  assign n36395 = ( ~n2171 & n7661 ) | ( ~n2171 & n7800 ) | ( n7661 & n7800 ) ;
  assign n36396 = n35167 ^ n22941 ^ n12927 ;
  assign n36397 = ( n750 & ~n36395 ) | ( n750 & n36396 ) | ( ~n36395 & n36396 ) ;
  assign n36398 = n36397 ^ n20260 ^ n11327 ;
  assign n36399 = ~n7080 & n17563 ;
  assign n36400 = ( ~n19961 & n20299 ) | ( ~n19961 & n36399 ) | ( n20299 & n36399 ) ;
  assign n36401 = n36400 ^ n36137 ^ n31864 ;
  assign n36402 = ( ~n5300 & n6695 ) | ( ~n5300 & n19073 ) | ( n6695 & n19073 ) ;
  assign n36403 = n3860 & n20114 ;
  assign n36404 = n36403 ^ n7785 ^ 1'b0 ;
  assign n36405 = ( n32667 & n36402 ) | ( n32667 & ~n36404 ) | ( n36402 & ~n36404 ) ;
  assign n36406 = ( n26117 & n29778 ) | ( n26117 & ~n36405 ) | ( n29778 & ~n36405 ) ;
  assign n36407 = n25714 ^ n20347 ^ n5766 ;
  assign n36408 = ( n26759 & ~n36406 ) | ( n26759 & n36407 ) | ( ~n36406 & n36407 ) ;
  assign n36409 = ( n7552 & ~n11066 ) | ( n7552 & n29074 ) | ( ~n11066 & n29074 ) ;
  assign n36410 = n31938 ^ n20298 ^ n2483 ;
  assign n36411 = ( n14357 & n17327 ) | ( n14357 & ~n23167 ) | ( n17327 & ~n23167 ) ;
  assign n36412 = ( n11363 & n16236 ) | ( n11363 & n36411 ) | ( n16236 & n36411 ) ;
  assign n36414 = ( n2602 & ~n2998 ) | ( n2602 & n19429 ) | ( ~n2998 & n19429 ) ;
  assign n36415 = ( ~n11580 & n26286 ) | ( ~n11580 & n36414 ) | ( n26286 & n36414 ) ;
  assign n36413 = n21293 ^ n13791 ^ 1'b0 ;
  assign n36416 = n36415 ^ n36413 ^ n6929 ;
  assign n36417 = ( ~n22730 & n22979 ) | ( ~n22730 & n34001 ) | ( n22979 & n34001 ) ;
  assign n36418 = n3181 & ~n6359 ;
  assign n36419 = ( n2598 & n13731 ) | ( n2598 & ~n36418 ) | ( n13731 & ~n36418 ) ;
  assign n36420 = ~n24243 & n26763 ;
  assign n36421 = n30013 & n36420 ;
  assign n36423 = ( n5355 & n7443 ) | ( n5355 & n24990 ) | ( n7443 & n24990 ) ;
  assign n36422 = n19235 & n23558 ;
  assign n36424 = n36423 ^ n36422 ^ n7559 ;
  assign n36425 = n23598 ^ n16125 ^ n12849 ;
  assign n36426 = n36425 ^ n29999 ^ n12345 ;
  assign n36427 = n36426 ^ n6138 ^ n4271 ;
  assign n36428 = n18307 ^ n10046 ^ 1'b0 ;
  assign n36429 = n20033 | n36428 ;
  assign n36430 = n36429 ^ n26494 ^ n23783 ;
  assign n36432 = n15970 ^ n6302 ^ n4674 ;
  assign n36433 = n36432 ^ n24895 ^ n15217 ;
  assign n36431 = n18543 ^ n14371 ^ n7960 ;
  assign n36434 = n36433 ^ n36431 ^ n15260 ;
  assign n36435 = ( ~n13954 & n17411 ) | ( ~n13954 & n36434 ) | ( n17411 & n36434 ) ;
  assign n36436 = ( n4649 & ~n12798 ) | ( n4649 & n13245 ) | ( ~n12798 & n13245 ) ;
  assign n36437 = ( n397 & n36357 ) | ( n397 & n36436 ) | ( n36357 & n36436 ) ;
  assign n36441 = n19243 ^ n7267 ^ 1'b0 ;
  assign n36439 = ( n6454 & ~n8124 ) | ( n6454 & n16899 ) | ( ~n8124 & n16899 ) ;
  assign n36440 = n36439 ^ n31110 ^ 1'b0 ;
  assign n36442 = n36441 ^ n36440 ^ n18659 ;
  assign n36438 = n18402 & ~n25359 ;
  assign n36443 = n36442 ^ n36438 ^ 1'b0 ;
  assign n36444 = ( n18003 & ~n20212 ) | ( n18003 & n34784 ) | ( ~n20212 & n34784 ) ;
  assign n36446 = ( x46 & n5778 ) | ( x46 & ~n9200 ) | ( n5778 & ~n9200 ) ;
  assign n36447 = ~n15833 & n36446 ;
  assign n36445 = n18244 ^ n11137 ^ n10062 ;
  assign n36448 = n36447 ^ n36445 ^ n1371 ;
  assign n36449 = n30606 ^ n23991 ^ n8353 ;
  assign n36450 = ( ~n832 & n2257 ) | ( ~n832 & n5675 ) | ( n2257 & n5675 ) ;
  assign n36451 = n11320 & n36450 ;
  assign n36452 = n36451 ^ n3744 ^ 1'b0 ;
  assign n36453 = n1060 & n4420 ;
  assign n36454 = ~n6725 & n36453 ;
  assign n36455 = ~n6939 & n36454 ;
  assign n36456 = ~n2608 & n25940 ;
  assign n36457 = ( n22618 & ~n23334 ) | ( n22618 & n36456 ) | ( ~n23334 & n36456 ) ;
  assign n36459 = ( n4556 & ~n7623 ) | ( n4556 & n12235 ) | ( ~n7623 & n12235 ) ;
  assign n36458 = ( x179 & ~n13162 ) | ( x179 & n21338 ) | ( ~n13162 & n21338 ) ;
  assign n36460 = n36459 ^ n36458 ^ n30282 ;
  assign n36462 = n3108 & n3181 ;
  assign n36463 = n36462 ^ n1345 ^ 1'b0 ;
  assign n36461 = n35806 ^ n15805 ^ n2674 ;
  assign n36464 = n36463 ^ n36461 ^ n16104 ;
  assign n36465 = n21747 ^ n2324 ^ 1'b0 ;
  assign n36466 = n24380 | n36465 ;
  assign n36468 = ( n9988 & ~n11958 ) | ( n9988 & n21011 ) | ( ~n11958 & n21011 ) ;
  assign n36467 = ( x211 & n18439 ) | ( x211 & ~n27034 ) | ( n18439 & ~n27034 ) ;
  assign n36469 = n36468 ^ n36467 ^ n22214 ;
  assign n36470 = ( n338 & n9989 ) | ( n338 & ~n22037 ) | ( n9989 & ~n22037 ) ;
  assign n36471 = n33378 ^ n27770 ^ n2061 ;
  assign n36472 = n36471 ^ n4690 ^ 1'b0 ;
  assign n36473 = n36470 | n36472 ;
  assign n36475 = ( n1269 & n21591 ) | ( n1269 & ~n24864 ) | ( n21591 & ~n24864 ) ;
  assign n36474 = n1335 & n21521 ;
  assign n36476 = n36475 ^ n36474 ^ 1'b0 ;
  assign n36477 = n34591 ^ n33092 ^ n27858 ;
  assign n36481 = ( n9973 & ~n11160 ) | ( n9973 & n23371 ) | ( ~n11160 & n23371 ) ;
  assign n36478 = n18423 & n24220 ;
  assign n36479 = n36478 ^ n5562 ^ 1'b0 ;
  assign n36480 = n36479 ^ n13827 ^ n4588 ;
  assign n36482 = n36481 ^ n36480 ^ n2247 ;
  assign n36483 = n28591 ^ n17395 ^ n2706 ;
  assign n36484 = n6473 & ~n7601 ;
  assign n36485 = n36484 ^ n16327 ^ 1'b0 ;
  assign n36486 = n15128 ^ n13367 ^ n11590 ;
  assign n36487 = ( n1990 & ~n4985 ) | ( n1990 & n36486 ) | ( ~n4985 & n36486 ) ;
  assign n36488 = n10988 ^ n6198 ^ n5485 ;
  assign n36489 = n20340 & ~n36488 ;
  assign n36490 = n3498 & n24803 ;
  assign n36491 = ~n10634 & n36490 ;
  assign n36492 = ( n3558 & n36489 ) | ( n3558 & ~n36491 ) | ( n36489 & ~n36491 ) ;
  assign n36493 = ( n6683 & n31969 ) | ( n6683 & ~n36492 ) | ( n31969 & ~n36492 ) ;
  assign n36494 = n16304 ^ n10793 ^ n7552 ;
  assign n36495 = ( n1254 & n4445 ) | ( n1254 & n19212 ) | ( n4445 & n19212 ) ;
  assign n36496 = n36495 ^ n18569 ^ n4885 ;
  assign n36497 = n23756 & ~n25236 ;
  assign n36498 = ( n13496 & n36496 ) | ( n13496 & ~n36497 ) | ( n36496 & ~n36497 ) ;
  assign n36499 = ( n30080 & ~n36494 ) | ( n30080 & n36498 ) | ( ~n36494 & n36498 ) ;
  assign n36500 = ( n10640 & ~n20324 ) | ( n10640 & n27655 ) | ( ~n20324 & n27655 ) ;
  assign n36501 = ( n295 & n1314 ) | ( n295 & n6360 ) | ( n1314 & n6360 ) ;
  assign n36502 = ( n12808 & ~n19454 ) | ( n12808 & n36501 ) | ( ~n19454 & n36501 ) ;
  assign n36503 = n36502 ^ n34629 ^ 1'b0 ;
  assign n36505 = ( n10730 & ~n10820 ) | ( n10730 & n29596 ) | ( ~n10820 & n29596 ) ;
  assign n36504 = ( n2469 & ~n3384 ) | ( n2469 & n6686 ) | ( ~n3384 & n6686 ) ;
  assign n36506 = n36505 ^ n36504 ^ n6539 ;
  assign n36507 = n14647 ^ n9948 ^ n611 ;
  assign n36508 = ( n2147 & n21334 ) | ( n2147 & n35633 ) | ( n21334 & n35633 ) ;
  assign n36509 = n26175 ^ n10310 ^ 1'b0 ;
  assign n36510 = n29362 & ~n36509 ;
  assign n36511 = ( n10224 & n22664 ) | ( n10224 & ~n33032 ) | ( n22664 & ~n33032 ) ;
  assign n36512 = ( ~n834 & n36510 ) | ( ~n834 & n36511 ) | ( n36510 & n36511 ) ;
  assign n36513 = ( n15778 & n18392 ) | ( n15778 & ~n36512 ) | ( n18392 & ~n36512 ) ;
  assign n36514 = ( ~n4029 & n8258 ) | ( ~n4029 & n36513 ) | ( n8258 & n36513 ) ;
  assign n36515 = ( ~n9165 & n36508 ) | ( ~n9165 & n36514 ) | ( n36508 & n36514 ) ;
  assign n36516 = n17098 & n35571 ;
  assign n36517 = n36516 ^ n31735 ^ 1'b0 ;
  assign n36518 = n32654 ^ n25175 ^ n5251 ;
  assign n36519 = n15524 ^ n1413 ^ 1'b0 ;
  assign n36520 = ( n5382 & ~n27545 ) | ( n5382 & n36519 ) | ( ~n27545 & n36519 ) ;
  assign n36521 = n10677 & n20473 ;
  assign n36522 = n25523 ^ n20150 ^ n4869 ;
  assign n36523 = n36522 ^ n8964 ^ 1'b0 ;
  assign n36524 = n36523 ^ n9749 ^ n730 ;
  assign n36525 = ( n3825 & n20377 ) | ( n3825 & ~n36524 ) | ( n20377 & ~n36524 ) ;
  assign n36526 = n29358 ^ n12330 ^ n4538 ;
  assign n36527 = ~n36525 & n36526 ;
  assign n36528 = ( ~n1837 & n19830 ) | ( ~n1837 & n31422 ) | ( n19830 & n31422 ) ;
  assign n36529 = n36528 ^ n3860 ^ n3216 ;
  assign n36530 = n28139 ^ n10194 ^ n774 ;
  assign n36531 = ( ~n6151 & n32803 ) | ( ~n6151 & n36530 ) | ( n32803 & n36530 ) ;
  assign n36532 = n36531 ^ n2691 ^ 1'b0 ;
  assign n36533 = n1338 & n36532 ;
  assign n36534 = n30398 ^ n28298 ^ n10415 ;
  assign n36535 = n36534 ^ n27344 ^ n17821 ;
  assign n36536 = ( n13464 & n19056 ) | ( n13464 & n22042 ) | ( n19056 & n22042 ) ;
  assign n36537 = ( n2484 & n21005 ) | ( n2484 & n30697 ) | ( n21005 & n30697 ) ;
  assign n36538 = ( n2793 & ~n22503 ) | ( n2793 & n24407 ) | ( ~n22503 & n24407 ) ;
  assign n36539 = ( ~n36536 & n36537 ) | ( ~n36536 & n36538 ) | ( n36537 & n36538 ) ;
  assign n36540 = n17736 ^ n10649 ^ n4077 ;
  assign n36541 = ~n12222 & n13103 ;
  assign n36542 = n36541 ^ n33396 ^ 1'b0 ;
  assign n36544 = ( n14060 & n16629 ) | ( n14060 & ~n30134 ) | ( n16629 & ~n30134 ) ;
  assign n36543 = n8080 & n9034 ;
  assign n36545 = n36544 ^ n36543 ^ 1'b0 ;
  assign n36546 = ( x172 & n8035 ) | ( x172 & ~n10626 ) | ( n8035 & ~n10626 ) ;
  assign n36547 = ( n478 & n3699 ) | ( n478 & ~n10520 ) | ( n3699 & ~n10520 ) ;
  assign n36548 = ( ~n20443 & n36546 ) | ( ~n20443 & n36547 ) | ( n36546 & n36547 ) ;
  assign n36549 = n36548 ^ n23091 ^ n3492 ;
  assign n36552 = n18610 ^ n14882 ^ n12449 ;
  assign n36550 = n16796 ^ n11543 ^ 1'b0 ;
  assign n36551 = ~n8542 & n36550 ;
  assign n36553 = n36552 ^ n36551 ^ n16189 ;
  assign n36554 = n36553 ^ n22350 ^ n18563 ;
  assign n36555 = n2949 & ~n19173 ;
  assign n36556 = n9934 ^ n2153 ^ x147 ;
  assign n36557 = ( n4783 & n18360 ) | ( n4783 & ~n36556 ) | ( n18360 & ~n36556 ) ;
  assign n36558 = n36557 ^ n29543 ^ n6516 ;
  assign n36559 = ( ~n3378 & n5930 ) | ( ~n3378 & n22876 ) | ( n5930 & n22876 ) ;
  assign n36560 = n36559 ^ n36149 ^ 1'b0 ;
  assign n36561 = n16945 ^ n9437 ^ 1'b0 ;
  assign n36562 = ~n15518 & n36561 ;
  assign n36563 = ( ~n12446 & n28024 ) | ( ~n12446 & n36562 ) | ( n28024 & n36562 ) ;
  assign n36564 = ( ~n1580 & n12248 ) | ( ~n1580 & n23329 ) | ( n12248 & n23329 ) ;
  assign n36565 = ( n4877 & n7246 ) | ( n4877 & n30409 ) | ( n7246 & n30409 ) ;
  assign n36566 = ( ~n5998 & n25359 ) | ( ~n5998 & n35153 ) | ( n25359 & n35153 ) ;
  assign n36567 = ( n18159 & n29101 ) | ( n18159 & ~n36566 ) | ( n29101 & ~n36566 ) ;
  assign n36568 = n36567 ^ n4543 ^ x133 ;
  assign n36569 = n12116 | n27215 ;
  assign n36570 = n3132 & ~n36569 ;
  assign n36571 = n36570 ^ n5341 ^ 1'b0 ;
  assign n36572 = n1829 & n5390 ;
  assign n36573 = ( n9000 & n15116 ) | ( n9000 & n17672 ) | ( n15116 & n17672 ) ;
  assign n36574 = ~n5175 & n31217 ;
  assign n36575 = n36574 ^ n18230 ^ 1'b0 ;
  assign n36576 = ( n33360 & ~n36573 ) | ( n33360 & n36575 ) | ( ~n36573 & n36575 ) ;
  assign n36579 = n21778 ^ n16477 ^ n10840 ;
  assign n36580 = n13461 & n36579 ;
  assign n36581 = n11796 & n36580 ;
  assign n36577 = n9364 ^ n6805 ^ 1'b0 ;
  assign n36578 = n14400 | n36577 ;
  assign n36582 = n36581 ^ n36578 ^ n6552 ;
  assign n36583 = ( x162 & ~n15100 ) | ( x162 & n26325 ) | ( ~n15100 & n26325 ) ;
  assign n36584 = n36583 ^ n10132 ^ 1'b0 ;
  assign n36585 = ( n24574 & n26072 ) | ( n24574 & ~n35773 ) | ( n26072 & ~n35773 ) ;
  assign n36586 = ( ~n12467 & n17073 ) | ( ~n12467 & n25385 ) | ( n17073 & n25385 ) ;
  assign n36589 = n23708 ^ n22740 ^ n9693 ;
  assign n36590 = n36589 ^ n30329 ^ n6660 ;
  assign n36591 = n36590 ^ n8867 ^ n3192 ;
  assign n36587 = n25540 ^ n6323 ^ 1'b0 ;
  assign n36588 = ~n8867 & n36587 ;
  assign n36592 = n36591 ^ n36588 ^ n26369 ;
  assign n36593 = ( n1376 & ~n6550 ) | ( n1376 & n36592 ) | ( ~n6550 & n36592 ) ;
  assign n36594 = ( n3585 & n6318 ) | ( n3585 & n11124 ) | ( n6318 & n11124 ) ;
  assign n36595 = n21393 ^ n2398 ^ n1496 ;
  assign n36596 = n11412 ^ n7188 ^ 1'b0 ;
  assign n36597 = n9083 & ~n36596 ;
  assign n36598 = ( n378 & n36595 ) | ( n378 & n36597 ) | ( n36595 & n36597 ) ;
  assign n36599 = ( n24952 & n36594 ) | ( n24952 & n36598 ) | ( n36594 & n36598 ) ;
  assign n36600 = ( n20055 & n22917 ) | ( n20055 & ~n32584 ) | ( n22917 & ~n32584 ) ;
  assign n36601 = n36600 ^ n11873 ^ n4245 ;
  assign n36602 = ~n18736 & n32515 ;
  assign n36603 = n36602 ^ n1284 ^ 1'b0 ;
  assign n36604 = n14264 ^ n3903 ^ n2786 ;
  assign n36605 = ( n5730 & n18033 ) | ( n5730 & ~n32766 ) | ( n18033 & ~n32766 ) ;
  assign n36606 = n36605 ^ n20459 ^ n19937 ;
  assign n36607 = ( n12158 & ~n36604 ) | ( n12158 & n36606 ) | ( ~n36604 & n36606 ) ;
  assign n36610 = ( ~n3294 & n17726 ) | ( ~n3294 & n28465 ) | ( n17726 & n28465 ) ;
  assign n36611 = n36610 ^ n27846 ^ n10635 ;
  assign n36608 = ( n3357 & n3376 ) | ( n3357 & ~n4761 ) | ( n3376 & ~n4761 ) ;
  assign n36609 = ( ~n6762 & n34411 ) | ( ~n6762 & n36608 ) | ( n34411 & n36608 ) ;
  assign n36612 = n36611 ^ n36609 ^ n9335 ;
  assign n36613 = n14998 ^ n13301 ^ n6399 ;
  assign n36617 = ( n399 & n8775 ) | ( n399 & n19167 ) | ( n8775 & n19167 ) ;
  assign n36614 = ( n3379 & ~n13671 ) | ( n3379 & n22142 ) | ( ~n13671 & n22142 ) ;
  assign n36615 = n36614 ^ n17943 ^ 1'b0 ;
  assign n36616 = n3541 & ~n36615 ;
  assign n36618 = n36617 ^ n36616 ^ n21674 ;
  assign n36619 = n20189 ^ n18086 ^ n966 ;
  assign n36620 = ~n10126 & n23332 ;
  assign n36621 = n14868 ^ n10253 ^ 1'b0 ;
  assign n36622 = n36621 ^ n16325 ^ n2326 ;
  assign n36623 = n36622 ^ n33519 ^ n10350 ;
  assign n36624 = ( n8766 & n14600 ) | ( n8766 & n36623 ) | ( n14600 & n36623 ) ;
  assign n36626 = n11982 ^ n8682 ^ n2926 ;
  assign n36625 = n27285 ^ n17058 ^ n15785 ;
  assign n36627 = n36626 ^ n36625 ^ n484 ;
  assign n36628 = ~n15637 & n28925 ;
  assign n36629 = ( ~n23389 & n28979 ) | ( ~n23389 & n35211 ) | ( n28979 & n35211 ) ;
  assign n36630 = n36629 ^ n26944 ^ n22158 ;
  assign n36631 = n18419 & ~n36630 ;
  assign n36632 = ( n4760 & n16545 ) | ( n4760 & ~n26814 ) | ( n16545 & ~n26814 ) ;
  assign n36633 = ( n5106 & n13425 ) | ( n5106 & ~n36632 ) | ( n13425 & ~n36632 ) ;
  assign n36634 = ( n9550 & n10608 ) | ( n9550 & n17753 ) | ( n10608 & n17753 ) ;
  assign n36635 = ~n10607 & n36530 ;
  assign n36636 = ( x71 & n15576 ) | ( x71 & n27332 ) | ( n15576 & n27332 ) ;
  assign n36637 = ( n31296 & n36635 ) | ( n31296 & ~n36636 ) | ( n36635 & ~n36636 ) ;
  assign n36638 = ( n16930 & ~n24045 ) | ( n16930 & n36637 ) | ( ~n24045 & n36637 ) ;
  assign n36639 = n36311 ^ n34541 ^ n6537 ;
  assign n36640 = ( n6875 & ~n16098 ) | ( n6875 & n29541 ) | ( ~n16098 & n29541 ) ;
  assign n36641 = n36640 ^ n10485 ^ n9664 ;
  assign n36642 = ( n24871 & n31239 ) | ( n24871 & n36641 ) | ( n31239 & n36641 ) ;
  assign n36643 = n7977 | n21436 ;
  assign n36644 = n36643 ^ n3259 ^ 1'b0 ;
  assign n36645 = ( n11855 & n21472 ) | ( n11855 & ~n36644 ) | ( n21472 & ~n36644 ) ;
  assign n36648 = n19548 ^ n12021 ^ n9377 ;
  assign n36646 = n34798 ^ n19081 ^ n12285 ;
  assign n36647 = ( n10493 & ~n20055 ) | ( n10493 & n36646 ) | ( ~n20055 & n36646 ) ;
  assign n36649 = n36648 ^ n36647 ^ n22820 ;
  assign n36650 = n19248 & ~n32096 ;
  assign n36651 = n28124 & n36650 ;
  assign n36652 = ( n13357 & n13427 ) | ( n13357 & n22766 ) | ( n13427 & n22766 ) ;
  assign n36653 = n32907 ^ n2847 ^ n1706 ;
  assign n36654 = ( n14618 & n28400 ) | ( n14618 & n36653 ) | ( n28400 & n36653 ) ;
  assign n36655 = n24541 ^ n22691 ^ n17595 ;
  assign n36657 = n25081 & n29666 ;
  assign n36656 = n31775 ^ n11439 ^ n3776 ;
  assign n36658 = n36657 ^ n36656 ^ n6288 ;
  assign n36659 = n36658 ^ n7622 ^ n1819 ;
  assign n36660 = n33590 ^ n18123 ^ 1'b0 ;
  assign n36661 = n36660 ^ n27854 ^ n25038 ;
  assign n36662 = n31897 ^ n8544 ^ n3318 ;
  assign n36663 = n36662 ^ n19067 ^ n9744 ;
  assign n36664 = n36663 ^ n9215 ^ n8751 ;
  assign n36666 = n21207 ^ n18267 ^ 1'b0 ;
  assign n36665 = ( n7077 & ~n16815 ) | ( n7077 & n30298 ) | ( ~n16815 & n30298 ) ;
  assign n36667 = n36666 ^ n36665 ^ n318 ;
  assign n36670 = n23691 ^ n17790 ^ n14328 ;
  assign n36671 = ( n1783 & n19386 ) | ( n1783 & n36670 ) | ( n19386 & n36670 ) ;
  assign n36672 = n36671 ^ n27576 ^ n15511 ;
  assign n36668 = n3558 | n25530 ;
  assign n36669 = n36668 ^ n36657 ^ 1'b0 ;
  assign n36673 = n36672 ^ n36669 ^ n3696 ;
  assign n36674 = ( n8171 & ~n25988 ) | ( n8171 & n26845 ) | ( ~n25988 & n26845 ) ;
  assign n36675 = n5400 & ~n36674 ;
  assign n36676 = n36675 ^ n9499 ^ 1'b0 ;
  assign n36677 = ~n17052 & n36676 ;
  assign n36678 = ( ~n12372 & n16676 ) | ( ~n12372 & n22604 ) | ( n16676 & n22604 ) ;
  assign n36679 = n6967 & n31440 ;
  assign n36680 = n14159 | n36679 ;
  assign n36681 = n19821 & ~n36680 ;
  assign n36682 = n36681 ^ n21666 ^ n9547 ;
  assign n36683 = n30545 ^ n22211 ^ n13117 ;
  assign n36684 = n21713 & ~n36683 ;
  assign n36685 = n33769 & n36684 ;
  assign n36687 = n22814 ^ n19861 ^ n9760 ;
  assign n36686 = n25975 ^ n25611 ^ n8754 ;
  assign n36688 = n36687 ^ n36686 ^ n23552 ;
  assign n36689 = ( ~n7789 & n9098 ) | ( ~n7789 & n22380 ) | ( n9098 & n22380 ) ;
  assign n36690 = ( n3988 & n8676 ) | ( n3988 & n10165 ) | ( n8676 & n10165 ) ;
  assign n36691 = n36690 ^ n15698 ^ 1'b0 ;
  assign n36692 = n36691 ^ n24853 ^ n22137 ;
  assign n36693 = ( n5494 & n15313 ) | ( n5494 & ~n32812 ) | ( n15313 & ~n32812 ) ;
  assign n36694 = n7877 & ~n23043 ;
  assign n36695 = n23854 ^ n18609 ^ n3391 ;
  assign n36696 = n1824 | n2926 ;
  assign n36697 = n21262 | n36696 ;
  assign n36698 = ( n16937 & ~n35610 ) | ( n16937 & n36697 ) | ( ~n35610 & n36697 ) ;
  assign n36699 = n22452 ^ n17593 ^ n10264 ;
  assign n36700 = n36699 ^ n17974 ^ n13330 ;
  assign n36701 = n17068 ^ n11498 ^ n10827 ;
  assign n36702 = n36701 ^ n31159 ^ n20767 ;
  assign n36703 = n15714 ^ n6053 ^ n5445 ;
  assign n36704 = ( n13663 & n26745 ) | ( n13663 & ~n36703 ) | ( n26745 & ~n36703 ) ;
  assign n36705 = ( ~n9233 & n22196 ) | ( ~n9233 & n36704 ) | ( n22196 & n36704 ) ;
  assign n36706 = ~n9787 & n36705 ;
  assign n36707 = n36706 ^ n2350 ^ 1'b0 ;
  assign n36708 = ( n4764 & n4842 ) | ( n4764 & ~n6799 ) | ( n4842 & ~n6799 ) ;
  assign n36709 = ( n883 & n14380 ) | ( n883 & n16306 ) | ( n14380 & n16306 ) ;
  assign n36710 = n36709 ^ n17010 ^ n1080 ;
  assign n36711 = n1790 & ~n36710 ;
  assign n36712 = ( n4651 & n15423 ) | ( n4651 & n29243 ) | ( n15423 & n29243 ) ;
  assign n36713 = ( ~n9438 & n10292 ) | ( ~n9438 & n22598 ) | ( n10292 & n22598 ) ;
  assign n36714 = ~n22236 & n36713 ;
  assign n36715 = n36714 ^ n32712 ^ 1'b0 ;
  assign n36716 = ( ~n2171 & n36712 ) | ( ~n2171 & n36715 ) | ( n36712 & n36715 ) ;
  assign n36717 = n28727 | n36716 ;
  assign n36718 = n36717 ^ n9972 ^ 1'b0 ;
  assign n36719 = n15332 ^ n11006 ^ n4228 ;
  assign n36720 = ( n1440 & n14466 ) | ( n1440 & ~n20122 ) | ( n14466 & ~n20122 ) ;
  assign n36721 = n16158 ^ n5831 ^ n1349 ;
  assign n36722 = ( n15087 & ~n36720 ) | ( n15087 & n36721 ) | ( ~n36720 & n36721 ) ;
  assign n36723 = ( ~n16259 & n36719 ) | ( ~n16259 & n36722 ) | ( n36719 & n36722 ) ;
  assign n36724 = n36723 ^ n19285 ^ 1'b0 ;
  assign n36725 = ~n7304 & n36724 ;
  assign n36726 = n31477 ^ n14401 ^ n7538 ;
  assign n36727 = ( n29445 & n30530 ) | ( n29445 & ~n31642 ) | ( n30530 & ~n31642 ) ;
  assign n36728 = ( n8901 & n19955 ) | ( n8901 & n28566 ) | ( n19955 & n28566 ) ;
  assign n36729 = n36728 ^ n27431 ^ n10809 ;
  assign n36730 = n25136 ^ n24717 ^ n8174 ;
  assign n36731 = ( n3632 & n8227 ) | ( n3632 & n36730 ) | ( n8227 & n36730 ) ;
  assign n36732 = n32741 ^ n12294 ^ 1'b0 ;
  assign n36733 = n35912 & n36732 ;
  assign n36734 = n6297 & n36459 ;
  assign n36735 = n36734 ^ n7031 ^ 1'b0 ;
  assign n36736 = n29517 ^ n2137 ^ 1'b0 ;
  assign n36741 = ( n9515 & ~n21019 ) | ( n9515 & n32380 ) | ( ~n21019 & n32380 ) ;
  assign n36742 = ( n5672 & n26963 ) | ( n5672 & ~n36741 ) | ( n26963 & ~n36741 ) ;
  assign n36740 = ( n15368 & ~n18345 ) | ( n15368 & n28239 ) | ( ~n18345 & n28239 ) ;
  assign n36737 = n2635 & n25629 ;
  assign n36738 = n3581 & n36737 ;
  assign n36739 = ( n6171 & n6570 ) | ( n6171 & ~n36738 ) | ( n6570 & ~n36738 ) ;
  assign n36743 = n36742 ^ n36740 ^ n36739 ;
  assign n36744 = n27407 ^ n14463 ^ n8178 ;
  assign n36745 = n25530 ^ n8212 ^ n4617 ;
  assign n36746 = ( ~n3951 & n11889 ) | ( ~n3951 & n36745 ) | ( n11889 & n36745 ) ;
  assign n36747 = ( n5851 & n21190 ) | ( n5851 & n32978 ) | ( n21190 & n32978 ) ;
  assign n36748 = n27130 ^ n12162 ^ n1309 ;
  assign n36749 = n36748 ^ n28090 ^ n20647 ;
  assign n36751 = n19440 ^ n8872 ^ n4258 ;
  assign n36750 = n18783 | n29500 ;
  assign n36752 = n36751 ^ n36750 ^ 1'b0 ;
  assign n36753 = n36752 ^ n24233 ^ 1'b0 ;
  assign n36754 = n36749 & n36753 ;
  assign n36755 = n36754 ^ n11443 ^ n3834 ;
  assign n36756 = ( n6742 & n17222 ) | ( n6742 & n17874 ) | ( n17222 & n17874 ) ;
  assign n36757 = n32303 ^ n4679 ^ n1716 ;
  assign n36758 = n24744 ^ n19906 ^ n1259 ;
  assign n36759 = n15133 ^ n12089 ^ n7143 ;
  assign n36760 = ( n36757 & ~n36758 ) | ( n36757 & n36759 ) | ( ~n36758 & n36759 ) ;
  assign n36761 = ( ~n26167 & n36756 ) | ( ~n26167 & n36760 ) | ( n36756 & n36760 ) ;
  assign n36762 = ( n2365 & n16570 ) | ( n2365 & ~n36761 ) | ( n16570 & ~n36761 ) ;
  assign n36763 = n31135 ^ n18570 ^ n5605 ;
  assign n36764 = n24319 ^ n14286 ^ n1543 ;
  assign n36765 = n36764 ^ n15487 ^ x143 ;
  assign n36766 = n19668 & n36765 ;
  assign n36767 = n12799 & n36766 ;
  assign n36768 = n6291 ^ n2620 ^ n2580 ;
  assign n36769 = ( n13472 & n19455 ) | ( n13472 & ~n36768 ) | ( n19455 & ~n36768 ) ;
  assign n36770 = ( n2006 & ~n28815 ) | ( n2006 & n36769 ) | ( ~n28815 & n36769 ) ;
  assign n36771 = n23662 ^ n1936 ^ n1351 ;
  assign n36772 = n3562 | n6183 ;
  assign n36773 = n6791 | n36772 ;
  assign n36774 = ( ~n23560 & n36771 ) | ( ~n23560 & n36773 ) | ( n36771 & n36773 ) ;
  assign n36775 = n36774 ^ n12783 ^ n6124 ;
  assign n36776 = n13530 & ~n14141 ;
  assign n36777 = ( ~n5450 & n14344 ) | ( ~n5450 & n36776 ) | ( n14344 & n36776 ) ;
  assign n36778 = ( n5925 & n11311 ) | ( n5925 & n36777 ) | ( n11311 & n36777 ) ;
  assign n36780 = ( ~n5024 & n6780 ) | ( ~n5024 & n24192 ) | ( n6780 & n24192 ) ;
  assign n36781 = ( ~n24819 & n24852 ) | ( ~n24819 & n36780 ) | ( n24852 & n36780 ) ;
  assign n36782 = n14365 ^ n11934 ^ n6605 ;
  assign n36783 = n36782 ^ n21428 ^ n6401 ;
  assign n36784 = ( n31441 & n36781 ) | ( n31441 & ~n36783 ) | ( n36781 & ~n36783 ) ;
  assign n36779 = n8196 ^ n3181 ^ n2621 ;
  assign n36785 = n36784 ^ n36779 ^ n1319 ;
  assign n36786 = ( n14085 & n18827 ) | ( n14085 & n33460 ) | ( n18827 & n33460 ) ;
  assign n36787 = n36786 ^ n14368 ^ n8446 ;
  assign n36788 = n15326 ^ n15265 ^ n5626 ;
  assign n36789 = ( n1196 & ~n11154 ) | ( n1196 & n11358 ) | ( ~n11154 & n11358 ) ;
  assign n36790 = n8472 ^ n3194 ^ n1546 ;
  assign n36791 = ( ~x179 & n10909 ) | ( ~x179 & n12045 ) | ( n10909 & n12045 ) ;
  assign n36792 = ( n2675 & n36790 ) | ( n2675 & ~n36791 ) | ( n36790 & ~n36791 ) ;
  assign n36793 = n36792 ^ n703 ^ 1'b0 ;
  assign n36794 = ~n36789 & n36793 ;
  assign n36795 = n16628 ^ n13748 ^ n13322 ;
  assign n36796 = ( n9951 & ~n14039 ) | ( n9951 & n36795 ) | ( ~n14039 & n36795 ) ;
  assign n36797 = ( ~n9361 & n17531 ) | ( ~n9361 & n23846 ) | ( n17531 & n23846 ) ;
  assign n36798 = ( ~x168 & n7202 ) | ( ~x168 & n17864 ) | ( n7202 & n17864 ) ;
  assign n36799 = n2792 & n16723 ;
  assign n36800 = n32310 ^ n15104 ^ 1'b0 ;
  assign n36801 = n36799 | n36800 ;
  assign n36802 = ( n10054 & ~n32953 ) | ( n10054 & n36801 ) | ( ~n32953 & n36801 ) ;
  assign n36803 = n16095 ^ n15612 ^ n6886 ;
  assign n36804 = n30084 ^ n8731 ^ n465 ;
  assign n36805 = ( n9248 & n36803 ) | ( n9248 & ~n36804 ) | ( n36803 & ~n36804 ) ;
  assign n36806 = ( n2865 & n4385 ) | ( n2865 & ~n6286 ) | ( n4385 & ~n6286 ) ;
  assign n36807 = n36806 ^ n25848 ^ n20671 ;
  assign n36808 = ( ~n22196 & n34962 ) | ( ~n22196 & n36807 ) | ( n34962 & n36807 ) ;
  assign n36809 = n10261 & n34041 ;
  assign n36810 = n2968 & n36809 ;
  assign n36811 = ( n19255 & ~n23115 ) | ( n19255 & n26402 ) | ( ~n23115 & n26402 ) ;
  assign n36812 = ( n21135 & n25114 ) | ( n21135 & ~n34427 ) | ( n25114 & ~n34427 ) ;
  assign n36813 = n24936 ^ n17663 ^ n4950 ;
  assign n36814 = n36813 ^ n36235 ^ n21134 ;
  assign n36815 = n6103 & ~n36814 ;
  assign n36816 = n13548 ^ n12884 ^ n4012 ;
  assign n36817 = n36816 ^ n10180 ^ 1'b0 ;
  assign n36818 = n34839 & n36817 ;
  assign n36819 = ( n8867 & ~n17895 ) | ( n8867 & n24739 ) | ( ~n17895 & n24739 ) ;
  assign n36821 = n15561 & ~n33720 ;
  assign n36822 = ( n1042 & ~n15256 ) | ( n1042 & n36821 ) | ( ~n15256 & n36821 ) ;
  assign n36820 = ~n4133 & n8772 ;
  assign n36823 = n36822 ^ n36820 ^ 1'b0 ;
  assign n36824 = n36823 ^ n28339 ^ n14044 ;
  assign n36825 = n36824 ^ n1263 ^ n359 ;
  assign n36826 = ( n19219 & n24009 ) | ( n19219 & n35286 ) | ( n24009 & n35286 ) ;
  assign n36833 = ( n5947 & ~n13227 ) | ( n5947 & n16382 ) | ( ~n13227 & n16382 ) ;
  assign n36827 = ( n891 & n1034 ) | ( n891 & n15552 ) | ( n1034 & n15552 ) ;
  assign n36828 = ( n8538 & ~n10341 ) | ( n8538 & n11673 ) | ( ~n10341 & n11673 ) ;
  assign n36829 = ( n554 & n1605 ) | ( n554 & n36828 ) | ( n1605 & n36828 ) ;
  assign n36830 = ( ~n12112 & n17476 ) | ( ~n12112 & n17903 ) | ( n17476 & n17903 ) ;
  assign n36831 = ( ~n6695 & n36829 ) | ( ~n6695 & n36830 ) | ( n36829 & n36830 ) ;
  assign n36832 = ( n10001 & n36827 ) | ( n10001 & n36831 ) | ( n36827 & n36831 ) ;
  assign n36834 = n36833 ^ n36832 ^ n9643 ;
  assign n36835 = n22702 ^ n18381 ^ n1532 ;
  assign n36836 = n36835 ^ n12927 ^ n6509 ;
  assign n36837 = n36836 ^ n19446 ^ n10258 ;
  assign n36838 = ( n5461 & ~n13768 ) | ( n5461 & n17320 ) | ( ~n13768 & n17320 ) ;
  assign n36839 = n20875 & n36838 ;
  assign n36840 = n29244 ^ n20517 ^ n4598 ;
  assign n36841 = ( n19406 & n35435 ) | ( n19406 & n36840 ) | ( n35435 & n36840 ) ;
  assign n36842 = n26646 ^ n23634 ^ n12153 ;
  assign n36843 = ( n1545 & n18393 ) | ( n1545 & ~n18427 ) | ( n18393 & ~n18427 ) ;
  assign n36844 = n36843 ^ n11714 ^ n9008 ;
  assign n36845 = n19572 ^ n13737 ^ 1'b0 ;
  assign n36846 = ~n21833 & n36845 ;
  assign n36847 = n32872 ^ n5626 ^ n799 ;
  assign n36848 = ( ~n20765 & n36846 ) | ( ~n20765 & n36847 ) | ( n36846 & n36847 ) ;
  assign n36849 = n36848 ^ n25981 ^ n23016 ;
  assign n36850 = n4223 ^ n4057 ^ 1'b0 ;
  assign n36851 = ( n572 & n21792 ) | ( n572 & n36850 ) | ( n21792 & n36850 ) ;
  assign n36852 = ( n7692 & n18178 ) | ( n7692 & ~n18592 ) | ( n18178 & ~n18592 ) ;
  assign n36853 = ~n9479 & n36852 ;
  assign n36854 = ~n2822 & n36853 ;
  assign n36855 = ~n21973 & n33254 ;
  assign n36856 = n6318 & ~n10795 ;
  assign n36857 = n36856 ^ n17754 ^ 1'b0 ;
  assign n36858 = n36857 ^ n20162 ^ n13998 ;
  assign n36859 = ( ~n8841 & n13436 ) | ( ~n8841 & n23087 ) | ( n13436 & n23087 ) ;
  assign n36860 = n36859 ^ n32263 ^ n384 ;
  assign n36861 = n36860 ^ n6269 ^ n1757 ;
  assign n36862 = ( ~n22175 & n31897 ) | ( ~n22175 & n36861 ) | ( n31897 & n36861 ) ;
  assign n36863 = ~n2668 & n22004 ;
  assign n36864 = n36863 ^ n30853 ^ 1'b0 ;
  assign n36865 = ~n9656 & n36864 ;
  assign n36866 = n35090 ^ n18383 ^ 1'b0 ;
  assign n36867 = n36865 & n36866 ;
  assign n36868 = n36867 ^ n26225 ^ n22715 ;
  assign n36869 = n36868 ^ n20276 ^ n3854 ;
  assign n36872 = n4417 | n5103 ;
  assign n36870 = n5711 ^ n3994 ^ n3861 ;
  assign n36871 = n36870 ^ n33970 ^ n1532 ;
  assign n36873 = n36872 ^ n36871 ^ n17005 ;
  assign n36874 = n24145 | n25034 ;
  assign n36875 = n19043 & ~n36874 ;
  assign n36876 = ( n21325 & n27307 ) | ( n21325 & ~n33554 ) | ( n27307 & ~n33554 ) ;
  assign n36877 = n36875 | n36876 ;
  assign n36878 = ( ~n2350 & n8128 ) | ( ~n2350 & n9621 ) | ( n8128 & n9621 ) ;
  assign n36879 = n36878 ^ n22907 ^ n2346 ;
  assign n36880 = n28226 ^ n23953 ^ n8256 ;
  assign n36881 = ( n2317 & ~n2831 ) | ( n2317 & n30678 ) | ( ~n2831 & n30678 ) ;
  assign n36882 = ( n5741 & ~n17315 ) | ( n5741 & n36881 ) | ( ~n17315 & n36881 ) ;
  assign n36883 = ( ~n389 & n2529 ) | ( ~n389 & n5884 ) | ( n2529 & n5884 ) ;
  assign n36884 = ( ~n7279 & n31150 ) | ( ~n7279 & n36883 ) | ( n31150 & n36883 ) ;
  assign n36885 = ( n19509 & ~n25798 ) | ( n19509 & n36884 ) | ( ~n25798 & n36884 ) ;
  assign n36886 = ~n313 & n25506 ;
  assign n36887 = n36885 & n36886 ;
  assign n36888 = ~n5983 & n9869 ;
  assign n36889 = n19220 ^ n4649 ^ 1'b0 ;
  assign n36890 = ( n3101 & n6854 ) | ( n3101 & ~n26711 ) | ( n6854 & ~n26711 ) ;
  assign n36891 = n16275 ^ n8042 ^ n2758 ;
  assign n36892 = n36891 ^ n17273 ^ n624 ;
  assign n36893 = n36892 ^ n23340 ^ n17900 ;
  assign n36894 = n7649 ^ n5659 ^ n4984 ;
  assign n36895 = n20930 ^ n17123 ^ n12662 ;
  assign n36896 = ( ~n4283 & n29992 ) | ( ~n4283 & n36895 ) | ( n29992 & n36895 ) ;
  assign n36897 = ( n18159 & n36894 ) | ( n18159 & ~n36896 ) | ( n36894 & ~n36896 ) ;
  assign n36898 = n22111 | n36897 ;
  assign n36899 = n1868 & ~n36898 ;
  assign n36900 = n29243 ^ n20229 ^ n3173 ;
  assign n36901 = n12094 ^ n4001 ^ n694 ;
  assign n36902 = ( n5658 & n36525 ) | ( n5658 & n36901 ) | ( n36525 & n36901 ) ;
  assign n36903 = n22238 ^ n605 ^ 1'b0 ;
  assign n36907 = n1358 & ~n12669 ;
  assign n36908 = ~n26360 & n36907 ;
  assign n36909 = n36908 ^ n25412 ^ n23740 ;
  assign n36904 = ( ~n23121 & n24060 ) | ( ~n23121 & n25371 ) | ( n24060 & n25371 ) ;
  assign n36905 = n16160 & n36904 ;
  assign n36906 = n36905 ^ n14603 ^ n8303 ;
  assign n36910 = n36909 ^ n36906 ^ n8115 ;
  assign n36911 = n13143 ^ n11353 ^ n4344 ;
  assign n36912 = ( n26626 & n29230 ) | ( n26626 & n36911 ) | ( n29230 & n36911 ) ;
  assign n36913 = n5505 ^ n4758 ^ n1287 ;
  assign n36914 = ( n1244 & ~n3013 ) | ( n1244 & n21432 ) | ( ~n3013 & n21432 ) ;
  assign n36915 = ( n9989 & n36913 ) | ( n9989 & n36914 ) | ( n36913 & n36914 ) ;
  assign n36916 = ( ~n6873 & n11106 ) | ( ~n6873 & n19147 ) | ( n11106 & n19147 ) ;
  assign n36917 = ( n4286 & ~n19646 ) | ( n4286 & n35398 ) | ( ~n19646 & n35398 ) ;
  assign n36918 = n23452 ^ n7672 ^ n5511 ;
  assign n36919 = n36917 & n36918 ;
  assign n36920 = n36916 & n36919 ;
  assign n36921 = n32445 ^ n30426 ^ 1'b0 ;
  assign n36922 = ( n23841 & ~n36920 ) | ( n23841 & n36921 ) | ( ~n36920 & n36921 ) ;
  assign n36923 = ( n17067 & n33857 ) | ( n17067 & ~n36922 ) | ( n33857 & ~n36922 ) ;
  assign n36925 = ( n5922 & ~n13067 ) | ( n5922 & n17651 ) | ( ~n13067 & n17651 ) ;
  assign n36926 = ( ~n1543 & n20667 ) | ( ~n1543 & n36925 ) | ( n20667 & n36925 ) ;
  assign n36924 = ( n3214 & n3945 ) | ( n3214 & n24115 ) | ( n3945 & n24115 ) ;
  assign n36927 = n36926 ^ n36924 ^ n16223 ;
  assign n36929 = n4394 & n8508 ;
  assign n36930 = ~n5947 & n36929 ;
  assign n36928 = n9913 & ~n17406 ;
  assign n36931 = n36930 ^ n36928 ^ 1'b0 ;
  assign n36932 = n27071 ^ n26548 ^ n23340 ;
  assign n36933 = ( n769 & n36931 ) | ( n769 & ~n36932 ) | ( n36931 & ~n36932 ) ;
  assign n36934 = n13872 ^ n11279 ^ n2754 ;
  assign n36935 = ( n9268 & ~n19161 ) | ( n9268 & n36934 ) | ( ~n19161 & n36934 ) ;
  assign n36937 = ( n645 & n1841 ) | ( n645 & n10763 ) | ( n1841 & n10763 ) ;
  assign n36938 = n36937 ^ n25831 ^ n15952 ;
  assign n36936 = ( ~n18318 & n36239 ) | ( ~n18318 & n36514 ) | ( n36239 & n36514 ) ;
  assign n36939 = n36938 ^ n36936 ^ n20052 ;
  assign n36940 = n30160 | n35990 ;
  assign n36943 = n4784 ^ n4723 ^ n3100 ;
  assign n36941 = n19720 ^ n6798 ^ n2737 ;
  assign n36942 = n36941 ^ n11267 ^ n1314 ;
  assign n36944 = n36943 ^ n36942 ^ n16515 ;
  assign n36945 = n19210 ^ n8821 ^ 1'b0 ;
  assign n36946 = n36944 & n36945 ;
  assign n36947 = n25952 ^ n19071 ^ n14470 ;
  assign n36949 = n33815 ^ n6805 ^ n3363 ;
  assign n36948 = n21821 & n23372 ;
  assign n36950 = n36949 ^ n36948 ^ 1'b0 ;
  assign n36951 = n16640 ^ n14742 ^ n718 ;
  assign n36952 = ( ~n13643 & n18966 ) | ( ~n13643 & n36951 ) | ( n18966 & n36951 ) ;
  assign n36953 = ( n12898 & n18818 ) | ( n12898 & n36952 ) | ( n18818 & n36952 ) ;
  assign n36954 = ( ~n28870 & n36636 ) | ( ~n28870 & n36953 ) | ( n36636 & n36953 ) ;
  assign n36955 = ( n36947 & ~n36950 ) | ( n36947 & n36954 ) | ( ~n36950 & n36954 ) ;
  assign n36958 = n15551 | n34785 ;
  assign n36959 = n36958 ^ n11242 ^ 1'b0 ;
  assign n36956 = n30592 ^ n28098 ^ n5880 ;
  assign n36957 = ( n29389 & n29925 ) | ( n29389 & ~n36956 ) | ( n29925 & ~n36956 ) ;
  assign n36960 = n36959 ^ n36957 ^ n33522 ;
  assign n36961 = n1109 & n18842 ;
  assign n36962 = n36961 ^ n2183 ^ 1'b0 ;
  assign n36963 = n33614 | n36962 ;
  assign n36964 = n16659 & ~n29142 ;
  assign n36965 = n36964 ^ n14936 ^ 1'b0 ;
  assign n36966 = ( n14338 & ~n31958 ) | ( n14338 & n36965 ) | ( ~n31958 & n36965 ) ;
  assign n36967 = n22125 & n31651 ;
  assign n36968 = ( ~n5218 & n6357 ) | ( ~n5218 & n20632 ) | ( n6357 & n20632 ) ;
  assign n36969 = ( x158 & n36941 ) | ( x158 & n36968 ) | ( n36941 & n36968 ) ;
  assign n36970 = n19504 ^ n12169 ^ n5534 ;
  assign n36971 = n36970 ^ n13476 ^ 1'b0 ;
  assign n36972 = n13182 & ~n36971 ;
  assign n36973 = n36972 ^ n22074 ^ n4987 ;
  assign n36974 = ( n5929 & ~n24827 ) | ( n5929 & n25772 ) | ( ~n24827 & n25772 ) ;
  assign n36975 = n36974 ^ n17503 ^ n1395 ;
  assign n36976 = ( n906 & n12249 ) | ( n906 & ~n28085 ) | ( n12249 & ~n28085 ) ;
  assign n36977 = ( ~n2180 & n2224 ) | ( ~n2180 & n20094 ) | ( n2224 & n20094 ) ;
  assign n36978 = ( ~n1935 & n6095 ) | ( ~n1935 & n36604 ) | ( n6095 & n36604 ) ;
  assign n36979 = n30292 ^ n1213 ^ 1'b0 ;
  assign n36980 = ~n11696 & n36979 ;
  assign n36981 = n9375 & ~n12781 ;
  assign n36982 = ~n4602 & n36981 ;
  assign n36983 = n24067 & n36982 ;
  assign n36984 = ( ~n1146 & n1440 ) | ( ~n1146 & n35407 ) | ( n1440 & n35407 ) ;
  assign n36989 = n2521 ^ n411 ^ x30 ;
  assign n36985 = n22618 & ~n27456 ;
  assign n36986 = n36985 ^ n5816 ^ 1'b0 ;
  assign n36987 = n36986 ^ n10326 ^ n8413 ;
  assign n36988 = ( ~n6248 & n19759 ) | ( ~n6248 & n36987 ) | ( n19759 & n36987 ) ;
  assign n36990 = n36989 ^ n36988 ^ n24161 ;
  assign n36996 = ~n2271 & n26696 ;
  assign n36997 = n19541 | n36996 ;
  assign n36993 = n18659 & ~n26217 ;
  assign n36994 = n21445 & n36993 ;
  assign n36991 = ( n2599 & ~n10286 ) | ( n2599 & n30346 ) | ( ~n10286 & n30346 ) ;
  assign n36992 = n36991 ^ n33934 ^ n1182 ;
  assign n36995 = n36994 ^ n36992 ^ n23862 ;
  assign n36998 = n36997 ^ n36995 ^ n6639 ;
  assign n36999 = ( n3580 & ~n9338 ) | ( n3580 & n27774 ) | ( ~n9338 & n27774 ) ;
  assign n37000 = ( n4823 & n35020 ) | ( n4823 & n36999 ) | ( n35020 & n36999 ) ;
  assign n37001 = n27533 ^ n27046 ^ n25484 ;
  assign n37002 = ( n12021 & n17185 ) | ( n12021 & ~n25840 ) | ( n17185 & ~n25840 ) ;
  assign n37003 = ( n1477 & ~n8299 ) | ( n1477 & n37002 ) | ( ~n8299 & n37002 ) ;
  assign n37004 = ( n23567 & n37001 ) | ( n23567 & n37003 ) | ( n37001 & n37003 ) ;
  assign n37005 = n33861 & ~n37004 ;
  assign n37006 = n1884 & n37005 ;
  assign n37007 = n29419 ^ n21271 ^ n1143 ;
  assign n37008 = n5070 | n22429 ;
  assign n37009 = n37008 ^ n1158 ^ 1'b0 ;
  assign n37010 = n37009 ^ n16698 ^ n2719 ;
  assign n37011 = n37010 ^ n22256 ^ n8993 ;
  assign n37012 = ( n12085 & n13684 ) | ( n12085 & n37011 ) | ( n13684 & n37011 ) ;
  assign n37013 = ( n356 & n1078 ) | ( n356 & n3558 ) | ( n1078 & n3558 ) ;
  assign n37014 = n26385 ^ n1247 ^ 1'b0 ;
  assign n37015 = ~n30045 & n37014 ;
  assign n37016 = n37015 ^ n14684 ^ n8317 ;
  assign n37017 = n4852 | n18499 ;
  assign n37018 = n37017 ^ n31057 ^ 1'b0 ;
  assign n37019 = n14942 ^ n10631 ^ n2279 ;
  assign n37020 = n16970 ^ n15306 ^ n6710 ;
  assign n37021 = ( n16429 & n27916 ) | ( n16429 & ~n37020 ) | ( n27916 & ~n37020 ) ;
  assign n37022 = ( n15800 & n37019 ) | ( n15800 & ~n37021 ) | ( n37019 & ~n37021 ) ;
  assign n37023 = ~n2089 & n37022 ;
  assign n37024 = n37023 ^ n5388 ^ 1'b0 ;
  assign n37025 = ( n448 & n10607 ) | ( n448 & n15826 ) | ( n10607 & n15826 ) ;
  assign n37026 = ( ~n679 & n3048 ) | ( ~n679 & n37025 ) | ( n3048 & n37025 ) ;
  assign n37027 = x57 & n37026 ;
  assign n37028 = ( n3049 & n5386 ) | ( n3049 & ~n11986 ) | ( n5386 & ~n11986 ) ;
  assign n37029 = ( x201 & n1612 ) | ( x201 & n37028 ) | ( n1612 & n37028 ) ;
  assign n37030 = n37029 ^ n34228 ^ n15811 ;
  assign n37031 = n27669 ^ n16073 ^ n4352 ;
  assign n37032 = ~n874 & n1665 ;
  assign n37033 = n1065 | n37032 ;
  assign n37034 = n4215 & ~n37033 ;
  assign n37035 = n16874 ^ n6961 ^ n4869 ;
  assign n37036 = n37035 ^ n34928 ^ n24252 ;
  assign n37037 = n15271 ^ n13702 ^ n2819 ;
  assign n37038 = n37037 ^ n3530 ^ n2455 ;
  assign n37039 = n738 | n4847 ;
  assign n37040 = n19730 ^ n7763 ^ n1987 ;
  assign n37042 = n11099 ^ n4261 ^ n2437 ;
  assign n37043 = x85 & ~n30065 ;
  assign n37044 = ~n37042 & n37043 ;
  assign n37041 = n14246 | n20992 ;
  assign n37045 = n37044 ^ n37041 ^ n33686 ;
  assign n37046 = n6206 & n19950 ;
  assign n37047 = ( ~n793 & n9349 ) | ( ~n793 & n15126 ) | ( n9349 & n15126 ) ;
  assign n37049 = ( ~n5549 & n9109 ) | ( ~n5549 & n12456 ) | ( n9109 & n12456 ) ;
  assign n37048 = ( n5993 & n10363 ) | ( n5993 & n16869 ) | ( n10363 & n16869 ) ;
  assign n37050 = n37049 ^ n37048 ^ 1'b0 ;
  assign n37051 = n10002 ^ n7559 ^ n1745 ;
  assign n37052 = n37051 ^ n33488 ^ n33317 ;
  assign n37053 = n25333 ^ n7997 ^ n4168 ;
  assign n37054 = ( n11390 & ~n15746 ) | ( n11390 & n28333 ) | ( ~n15746 & n28333 ) ;
  assign n37055 = n4658 & n9218 ;
  assign n37056 = ~n6690 & n37055 ;
  assign n37057 = ( n3162 & n9817 ) | ( n3162 & n37056 ) | ( n9817 & n37056 ) ;
  assign n37058 = n16784 ^ n16260 ^ n8240 ;
  assign n37059 = ( ~n3408 & n14752 ) | ( ~n3408 & n37058 ) | ( n14752 & n37058 ) ;
  assign n37060 = n37059 ^ n6234 ^ n3804 ;
  assign n37061 = n4775 & ~n31120 ;
  assign n37062 = n37061 ^ n28103 ^ n24882 ;
  assign n37063 = n2479 ^ n942 ^ 1'b0 ;
  assign n37064 = ( n11695 & n36093 ) | ( n11695 & ~n37063 ) | ( n36093 & ~n37063 ) ;
  assign n37065 = n30963 & ~n32288 ;
  assign n37066 = n37065 ^ n25106 ^ n8621 ;
  assign n37067 = ( ~n17882 & n18347 ) | ( ~n17882 & n20163 ) | ( n18347 & n20163 ) ;
  assign n37068 = ( n1465 & n29872 ) | ( n1465 & n37067 ) | ( n29872 & n37067 ) ;
  assign n37069 = ( n24420 & n36962 ) | ( n24420 & n37068 ) | ( n36962 & n37068 ) ;
  assign n37070 = ( n5286 & n5543 ) | ( n5286 & ~n7708 ) | ( n5543 & ~n7708 ) ;
  assign n37074 = ~n5623 & n32397 ;
  assign n37075 = n37074 ^ n10007 ^ 1'b0 ;
  assign n37071 = n15909 ^ n12814 ^ n5376 ;
  assign n37072 = n26101 | n37071 ;
  assign n37073 = n26923 & ~n37072 ;
  assign n37076 = n37075 ^ n37073 ^ 1'b0 ;
  assign n37080 = ( n7365 & n8593 ) | ( n7365 & ~n9333 ) | ( n8593 & ~n9333 ) ;
  assign n37081 = ( n4817 & n31161 ) | ( n4817 & n37080 ) | ( n31161 & n37080 ) ;
  assign n37077 = n5075 ^ n4921 ^ n4833 ;
  assign n37078 = n37077 ^ n18921 ^ 1'b0 ;
  assign n37079 = ~n23604 & n37078 ;
  assign n37082 = n37081 ^ n37079 ^ n8429 ;
  assign n37083 = ( n3779 & ~n5345 ) | ( n3779 & n7416 ) | ( ~n5345 & n7416 ) ;
  assign n37084 = n37083 ^ n857 ^ 1'b0 ;
  assign n37085 = n2756 | n37084 ;
  assign n37086 = ( n6763 & ~n14354 ) | ( n6763 & n22431 ) | ( ~n14354 & n22431 ) ;
  assign n37087 = ( ~n13999 & n22672 ) | ( ~n13999 & n37086 ) | ( n22672 & n37086 ) ;
  assign n37088 = n37087 ^ n33470 ^ n14638 ;
  assign n37089 = ( ~n4692 & n37085 ) | ( ~n4692 & n37088 ) | ( n37085 & n37088 ) ;
  assign n37090 = n21405 ^ n14321 ^ 1'b0 ;
  assign n37091 = n18548 & n37090 ;
  assign n37092 = n27282 & ~n36267 ;
  assign n37093 = ( ~n1739 & n9107 ) | ( ~n1739 & n29595 ) | ( n9107 & n29595 ) ;
  assign n37094 = n37093 ^ n25001 ^ n19742 ;
  assign n37095 = n3954 ^ n3062 ^ n2014 ;
  assign n37096 = ( n4761 & n7696 ) | ( n4761 & n37095 ) | ( n7696 & n37095 ) ;
  assign n37102 = ( ~n21690 & n23807 ) | ( ~n21690 & n32481 ) | ( n23807 & n32481 ) ;
  assign n37097 = n29295 ^ n6213 ^ n4090 ;
  assign n37098 = ( n6628 & n13365 ) | ( n6628 & ~n37097 ) | ( n13365 & ~n37097 ) ;
  assign n37099 = n37098 ^ n15378 ^ n9441 ;
  assign n37100 = n37099 ^ n2500 ^ 1'b0 ;
  assign n37101 = n8860 & ~n37100 ;
  assign n37103 = n37102 ^ n37101 ^ n28991 ;
  assign n37104 = ( n3224 & n12138 ) | ( n3224 & n35105 ) | ( n12138 & n35105 ) ;
  assign n37105 = ( n25607 & n31861 ) | ( n25607 & ~n37104 ) | ( n31861 & ~n37104 ) ;
  assign n37106 = n30547 ^ n26682 ^ n19989 ;
  assign n37107 = n22844 ^ n20863 ^ n6250 ;
  assign n37108 = n37107 ^ n6219 ^ n1347 ;
  assign n37109 = ( n30655 & n37106 ) | ( n30655 & ~n37108 ) | ( n37106 & ~n37108 ) ;
  assign n37110 = n36433 ^ n1003 ^ 1'b0 ;
  assign n37111 = n19598 ^ n13322 ^ n4410 ;
  assign n37112 = ( ~n12784 & n37110 ) | ( ~n12784 & n37111 ) | ( n37110 & n37111 ) ;
  assign n37113 = ( n4852 & n5123 ) | ( n4852 & n15866 ) | ( n5123 & n15866 ) ;
  assign n37114 = n15505 ^ n6766 ^ 1'b0 ;
  assign n37115 = n5297 & n37114 ;
  assign n37116 = n37115 ^ n27311 ^ n3575 ;
  assign n37117 = n26230 ^ n6871 ^ n734 ;
  assign n37118 = n25273 ^ n13445 ^ n3911 ;
  assign n37119 = ( n2089 & ~n9574 ) | ( n2089 & n18514 ) | ( ~n9574 & n18514 ) ;
  assign n37120 = ( ~x167 & n10171 ) | ( ~x167 & n17867 ) | ( n10171 & n17867 ) ;
  assign n37121 = n37120 ^ n16748 ^ n1841 ;
  assign n37122 = n959 & n37121 ;
  assign n37123 = ~n33738 & n37122 ;
  assign n37124 = ( ~n1620 & n4555 ) | ( ~n1620 & n18016 ) | ( n4555 & n18016 ) ;
  assign n37125 = ( n37119 & ~n37123 ) | ( n37119 & n37124 ) | ( ~n37123 & n37124 ) ;
  assign n37126 = ( n2237 & n9942 ) | ( n2237 & n21535 ) | ( n9942 & n21535 ) ;
  assign n37127 = n37126 ^ n10919 ^ n6497 ;
  assign n37128 = ( n6489 & n16968 ) | ( n6489 & ~n18610 ) | ( n16968 & ~n18610 ) ;
  assign n37129 = n37128 ^ n5844 ^ 1'b0 ;
  assign n37130 = n17836 | n37129 ;
  assign n37131 = n34015 ^ n2765 ^ x27 ;
  assign n37132 = n5186 & ~n7350 ;
  assign n37133 = n37132 ^ n12411 ^ n3798 ;
  assign n37134 = n30529 ^ n19488 ^ n1458 ;
  assign n37135 = n27398 ^ n11549 ^ n6608 ;
  assign n37136 = n31933 ^ n8417 ^ n1779 ;
  assign n37137 = n37136 ^ n25322 ^ n15737 ;
  assign n37138 = ( n37134 & ~n37135 ) | ( n37134 & n37137 ) | ( ~n37135 & n37137 ) ;
  assign n37139 = ( n18240 & ~n30364 ) | ( n18240 & n37138 ) | ( ~n30364 & n37138 ) ;
  assign n37140 = n1961 & ~n4977 ;
  assign n37141 = n4717 & ~n20982 ;
  assign n37142 = n37141 ^ n22633 ^ n324 ;
  assign n37143 = n10472 | n28720 ;
  assign n37144 = ( n37140 & n37142 ) | ( n37140 & ~n37143 ) | ( n37142 & ~n37143 ) ;
  assign n37145 = n28695 ^ n14895 ^ n1747 ;
  assign n37146 = ( n7075 & ~n18005 ) | ( n7075 & n33906 ) | ( ~n18005 & n33906 ) ;
  assign n37147 = ( n5042 & n12401 ) | ( n5042 & n37146 ) | ( n12401 & n37146 ) ;
  assign n37148 = ( ~n13973 & n29732 ) | ( ~n13973 & n33083 ) | ( n29732 & n33083 ) ;
  assign n37149 = n31458 ^ n2252 ^ n837 ;
  assign n37150 = ( n10323 & n35109 ) | ( n10323 & ~n37149 ) | ( n35109 & ~n37149 ) ;
  assign n37151 = n21559 ^ n16875 ^ n9584 ;
  assign n37152 = n37151 ^ n29193 ^ n15407 ;
  assign n37153 = ( n7844 & n19329 ) | ( n7844 & ~n23752 ) | ( n19329 & ~n23752 ) ;
  assign n37154 = n37153 ^ n13939 ^ n5580 ;
  assign n37155 = ( n9421 & n22254 ) | ( n9421 & ~n34826 ) | ( n22254 & ~n34826 ) ;
  assign n37156 = n15243 ^ n5871 ^ n2760 ;
  assign n37157 = ( n6959 & n14161 ) | ( n6959 & ~n32920 ) | ( n14161 & ~n32920 ) ;
  assign n37158 = ( n1709 & n7642 ) | ( n1709 & n8849 ) | ( n7642 & n8849 ) ;
  assign n37159 = n22406 ^ n16161 ^ n13012 ;
  assign n37160 = ( n27413 & ~n37158 ) | ( n27413 & n37159 ) | ( ~n37158 & n37159 ) ;
  assign n37161 = n37160 ^ n7190 ^ n3962 ;
  assign n37162 = ( n2228 & ~n27485 ) | ( n2228 & n37161 ) | ( ~n27485 & n37161 ) ;
  assign n37163 = ( n3816 & ~n20419 ) | ( n3816 & n33933 ) | ( ~n20419 & n33933 ) ;
  assign n37164 = ( n1262 & n2828 ) | ( n1262 & ~n37163 ) | ( n2828 & ~n37163 ) ;
  assign n37165 = n17668 ^ n13087 ^ n970 ;
  assign n37170 = n36331 ^ n34509 ^ n16016 ;
  assign n37166 = n12396 ^ n988 ^ n676 ;
  assign n37167 = n37166 ^ n30439 ^ n14065 ;
  assign n37168 = ( n10209 & ~n33711 ) | ( n10209 & n37167 ) | ( ~n33711 & n37167 ) ;
  assign n37169 = n37168 ^ n22724 ^ x55 ;
  assign n37171 = n37170 ^ n37169 ^ 1'b0 ;
  assign n37172 = ~n37165 & n37171 ;
  assign n37176 = ( n5871 & ~n21293 ) | ( n5871 & n27365 ) | ( ~n21293 & n27365 ) ;
  assign n37173 = n36425 ^ n7606 ^ n6536 ;
  assign n37174 = ( ~n3347 & n26861 ) | ( ~n3347 & n37173 ) | ( n26861 & n37173 ) ;
  assign n37175 = n37174 ^ n3980 ^ 1'b0 ;
  assign n37177 = n37176 ^ n37175 ^ 1'b0 ;
  assign n37178 = ( ~n17451 & n27363 ) | ( ~n17451 & n31590 ) | ( n27363 & n31590 ) ;
  assign n37179 = ( n16264 & n21223 ) | ( n16264 & ~n25669 ) | ( n21223 & ~n25669 ) ;
  assign n37180 = ( n23294 & n26432 ) | ( n23294 & n37179 ) | ( n26432 & n37179 ) ;
  assign n37181 = ( n407 & n8703 ) | ( n407 & n37180 ) | ( n8703 & n37180 ) ;
  assign n37182 = n14884 | n19332 ;
  assign n37183 = n37182 ^ n33055 ^ n22104 ;
  assign n37184 = n16417 ^ n13069 ^ 1'b0 ;
  assign n37185 = n11093 | n26677 ;
  assign n37186 = n30059 ^ n25558 ^ n6178 ;
  assign n37187 = n16205 | n37186 ;
  assign n37188 = n20240 & ~n37187 ;
  assign n37189 = ( n9767 & n24728 ) | ( n9767 & n26214 ) | ( n24728 & n26214 ) ;
  assign n37190 = n27460 & ~n37189 ;
  assign n37191 = n33633 ^ n4533 ^ n2995 ;
  assign n37192 = n37191 ^ n34497 ^ n26560 ;
  assign n37193 = ( n8074 & n8522 ) | ( n8074 & ~n12001 ) | ( n8522 & ~n12001 ) ;
  assign n37194 = n2933 & n33313 ;
  assign n37195 = n37193 & n37194 ;
  assign n37196 = n14001 ^ n4315 ^ 1'b0 ;
  assign n37197 = ( n7227 & ~n14278 ) | ( n7227 & n37196 ) | ( ~n14278 & n37196 ) ;
  assign n37198 = n8618 ^ n7135 ^ n681 ;
  assign n37199 = n26846 ^ n24006 ^ n19914 ;
  assign n37200 = ( n17763 & n37198 ) | ( n17763 & ~n37199 ) | ( n37198 & ~n37199 ) ;
  assign n37201 = ( n7526 & n26414 ) | ( n7526 & ~n29782 ) | ( n26414 & ~n29782 ) ;
  assign n37202 = n10661 ^ n7140 ^ 1'b0 ;
  assign n37203 = n37202 ^ n28791 ^ n9879 ;
  assign n37204 = ( n9460 & ~n24009 ) | ( n9460 & n29367 ) | ( ~n24009 & n29367 ) ;
  assign n37205 = ( ~n16020 & n36720 ) | ( ~n16020 & n37204 ) | ( n36720 & n37204 ) ;
  assign n37207 = n33785 ^ n29122 ^ n9573 ;
  assign n37206 = n30371 ^ n11852 ^ n6811 ;
  assign n37208 = n37207 ^ n37206 ^ n6406 ;
  assign n37209 = ~n24806 & n35503 ;
  assign n37210 = n37209 ^ x0 ^ 1'b0 ;
  assign n37215 = ( n2237 & n2968 ) | ( n2237 & ~n7958 ) | ( n2968 & ~n7958 ) ;
  assign n37214 = n17597 ^ n16349 ^ n3619 ;
  assign n37211 = n3742 & n27466 ;
  assign n37212 = n37211 ^ n20560 ^ 1'b0 ;
  assign n37213 = ( ~n11230 & n12695 ) | ( ~n11230 & n37212 ) | ( n12695 & n37212 ) ;
  assign n37216 = n37215 ^ n37214 ^ n37213 ;
  assign n37217 = ( ~n4964 & n9924 ) | ( ~n4964 & n31849 ) | ( n9924 & n31849 ) ;
  assign n37218 = n37217 ^ n15230 ^ n13582 ;
  assign n37219 = ( n8208 & n12389 ) | ( n8208 & ~n37218 ) | ( n12389 & ~n37218 ) ;
  assign n37220 = n37219 ^ n21012 ^ 1'b0 ;
  assign n37222 = n16938 ^ n14611 ^ n12611 ;
  assign n37221 = n16414 ^ n12183 ^ 1'b0 ;
  assign n37223 = n37222 ^ n37221 ^ 1'b0 ;
  assign n37224 = n30615 ^ n28897 ^ n1132 ;
  assign n37225 = ( n12381 & n23042 ) | ( n12381 & n37224 ) | ( n23042 & n37224 ) ;
  assign n37226 = ~n29309 & n37225 ;
  assign n37227 = n12659 ^ n8030 ^ 1'b0 ;
  assign n37228 = ~n14428 & n37227 ;
  assign n37229 = n19295 ^ n3713 ^ n2108 ;
  assign n37230 = ( n11869 & n33836 ) | ( n11869 & n37229 ) | ( n33836 & n37229 ) ;
  assign n37231 = n27810 ^ n10277 ^ n5480 ;
  assign n37232 = n37231 ^ n30706 ^ n10622 ;
  assign n37233 = ~n13774 & n17723 ;
  assign n37234 = ~n37232 & n37233 ;
  assign n37235 = ( n18237 & n19629 ) | ( n18237 & ~n20315 ) | ( n19629 & ~n20315 ) ;
  assign n37237 = n15841 ^ n8995 ^ n1049 ;
  assign n37236 = n24383 ^ n18764 ^ n7064 ;
  assign n37238 = n37237 ^ n37236 ^ 1'b0 ;
  assign n37239 = n31836 ^ n30281 ^ n17370 ;
  assign n37240 = n36937 ^ n11890 ^ 1'b0 ;
  assign n37241 = x175 & n37240 ;
  assign n37242 = n2945 & n37241 ;
  assign n37243 = n9688 ^ n3693 ^ n3126 ;
  assign n37244 = n37243 ^ n31038 ^ n23793 ;
  assign n37245 = n11893 ^ n1572 ^ n1519 ;
  assign n37246 = n37245 ^ n20254 ^ n11334 ;
  assign n37247 = n37246 ^ n9948 ^ 1'b0 ;
  assign n37248 = n3349 & n37247 ;
  assign n37249 = n27999 ^ n22310 ^ n1927 ;
  assign n37250 = n37249 ^ n20439 ^ n14547 ;
  assign n37251 = n37250 ^ n30808 ^ n13553 ;
  assign n37252 = ( n10304 & n18980 ) | ( n10304 & ~n26601 ) | ( n18980 & ~n26601 ) ;
  assign n37253 = n13084 ^ n10582 ^ 1'b0 ;
  assign n37254 = n37253 ^ n9613 ^ n4083 ;
  assign n37255 = n14891 ^ n5881 ^ 1'b0 ;
  assign n37256 = n15860 & ~n37255 ;
  assign n37257 = ( n9741 & ~n15169 ) | ( n9741 & n37256 ) | ( ~n15169 & n37256 ) ;
  assign n37258 = n17844 ^ n16022 ^ n9449 ;
  assign n37259 = ( n7178 & ~n10657 ) | ( n7178 & n14717 ) | ( ~n10657 & n14717 ) ;
  assign n37262 = n28346 ^ n5814 ^ n1911 ;
  assign n37261 = n36175 ^ n15687 ^ n3532 ;
  assign n37263 = n37262 ^ n37261 ^ n2659 ;
  assign n37260 = ( n2733 & n16893 ) | ( n2733 & n22701 ) | ( n16893 & n22701 ) ;
  assign n37264 = n37263 ^ n37260 ^ n7384 ;
  assign n37265 = ( n4871 & n19479 ) | ( n4871 & ~n37264 ) | ( n19479 & ~n37264 ) ;
  assign n37266 = n37265 ^ n4462 ^ x33 ;
  assign n37267 = n26673 ^ n25883 ^ n12331 ;
  assign n37268 = n10418 ^ n1449 ^ 1'b0 ;
  assign n37269 = n26619 | n37268 ;
  assign n37270 = ( ~n11448 & n27086 ) | ( ~n11448 & n37269 ) | ( n27086 & n37269 ) ;
  assign n37271 = n31896 ^ n21625 ^ n2174 ;
  assign n37272 = n37271 ^ n6906 ^ 1'b0 ;
  assign n37273 = n24030 ^ n9538 ^ n9047 ;
  assign n37274 = n3004 & ~n21694 ;
  assign n37275 = ~n20054 & n37274 ;
  assign n37276 = n22219 ^ n11248 ^ n3694 ;
  assign n37277 = n7142 ^ n4943 ^ n1395 ;
  assign n37278 = ( n13533 & ~n37276 ) | ( n13533 & n37277 ) | ( ~n37276 & n37277 ) ;
  assign n37279 = ( n6317 & ~n20518 ) | ( n6317 & n28080 ) | ( ~n20518 & n28080 ) ;
  assign n37281 = ( n2204 & n7735 ) | ( n2204 & n12335 ) | ( n7735 & n12335 ) ;
  assign n37282 = n37281 ^ n22516 ^ n9619 ;
  assign n37280 = n20483 ^ n18282 ^ n5796 ;
  assign n37283 = n37282 ^ n37280 ^ n35039 ;
  assign n37285 = n15927 | n26104 ;
  assign n37284 = n25893 ^ n10304 ^ n5970 ;
  assign n37286 = n37285 ^ n37284 ^ n22706 ;
  assign n37287 = ( n3740 & n26595 ) | ( n3740 & n37286 ) | ( n26595 & n37286 ) ;
  assign n37288 = ( n12240 & ~n15872 ) | ( n12240 & n19468 ) | ( ~n15872 & n19468 ) ;
  assign n37289 = n37288 ^ n21033 ^ n15201 ;
  assign n37290 = ( n1662 & n4285 ) | ( n1662 & ~n33518 ) | ( n4285 & ~n33518 ) ;
  assign n37293 = n11172 ^ n8054 ^ n6861 ;
  assign n37294 = n37293 ^ n20982 ^ n4164 ;
  assign n37291 = ( n21478 & n26160 ) | ( n21478 & ~n30081 ) | ( n26160 & ~n30081 ) ;
  assign n37292 = n23832 | n37291 ;
  assign n37295 = n37294 ^ n37292 ^ n21450 ;
  assign n37296 = ( n1339 & ~n2811 ) | ( n1339 & n27347 ) | ( ~n2811 & n27347 ) ;
  assign n37297 = n6733 | n12028 ;
  assign n37298 = n20427 ^ n11156 ^ n2968 ;
  assign n37299 = n9289 & n19111 ;
  assign n37300 = n37299 ^ x124 ^ 1'b0 ;
  assign n37301 = n6561 & ~n37300 ;
  assign n37302 = ~n37298 & n37301 ;
  assign n37303 = n8550 ^ n2451 ^ 1'b0 ;
  assign n37304 = ~n8426 & n37303 ;
  assign n37305 = ~x216 & n2529 ;
  assign n37306 = ( n3947 & ~n5725 ) | ( n3947 & n11499 ) | ( ~n5725 & n11499 ) ;
  assign n37307 = n37306 ^ n27853 ^ n4405 ;
  assign n37308 = ( n7783 & n19383 ) | ( n7783 & ~n37307 ) | ( n19383 & ~n37307 ) ;
  assign n37309 = ( n32525 & ~n37305 ) | ( n32525 & n37308 ) | ( ~n37305 & n37308 ) ;
  assign n37314 = ( ~n12172 & n19519 ) | ( ~n12172 & n21091 ) | ( n19519 & n21091 ) ;
  assign n37315 = n37314 ^ n34810 ^ n19261 ;
  assign n37311 = n17636 ^ n1943 ^ x150 ;
  assign n37310 = n35006 ^ n14891 ^ n6231 ;
  assign n37312 = n37311 ^ n37310 ^ n22609 ;
  assign n37313 = ( ~n8425 & n17318 ) | ( ~n8425 & n37312 ) | ( n17318 & n37312 ) ;
  assign n37316 = n37315 ^ n37313 ^ n6681 ;
  assign n37317 = ( n10694 & n17884 ) | ( n10694 & n19052 ) | ( n17884 & n19052 ) ;
  assign n37318 = n37317 ^ n11358 ^ n8543 ;
  assign n37319 = n37318 ^ n31303 ^ n15190 ;
  assign n37320 = n27191 ^ n5964 ^ n1633 ;
  assign n37321 = ( n14753 & ~n29897 ) | ( n14753 & n37320 ) | ( ~n29897 & n37320 ) ;
  assign n37322 = n30414 ^ n20433 ^ n15440 ;
  assign n37323 = n18038 ^ n13469 ^ n7641 ;
  assign n37324 = n37323 ^ n27403 ^ n11625 ;
  assign n37325 = n23663 ^ n11651 ^ n7486 ;
  assign n37326 = n19255 ^ n15014 ^ x215 ;
  assign n37327 = n35066 ^ n13139 ^ n11553 ;
  assign n37328 = ( n18456 & n37326 ) | ( n18456 & n37327 ) | ( n37326 & n37327 ) ;
  assign n37329 = n37328 ^ n21696 ^ n15927 ;
  assign n37330 = ( n10726 & ~n34308 ) | ( n10726 & n37329 ) | ( ~n34308 & n37329 ) ;
  assign n37331 = ( n23518 & n37325 ) | ( n23518 & ~n37330 ) | ( n37325 & ~n37330 ) ;
  assign n37332 = n29827 ^ n15850 ^ n13671 ;
  assign n37333 = n29514 ^ n26407 ^ n22788 ;
  assign n37334 = ( n6013 & n37332 ) | ( n6013 & n37333 ) | ( n37332 & n37333 ) ;
  assign n37335 = n37334 ^ n26754 ^ n12404 ;
  assign n37336 = n31589 ^ n26675 ^ n16135 ;
  assign n37337 = ( n12588 & n28983 ) | ( n12588 & n32738 ) | ( n28983 & n32738 ) ;
  assign n37338 = n23785 ^ n23414 ^ n12839 ;
  assign n37339 = ( n27441 & n34971 ) | ( n27441 & ~n37338 ) | ( n34971 & ~n37338 ) ;
  assign n37341 = ( n1783 & n12824 ) | ( n1783 & ~n34407 ) | ( n12824 & ~n34407 ) ;
  assign n37340 = ( ~n773 & n24624 ) | ( ~n773 & n34589 ) | ( n24624 & n34589 ) ;
  assign n37342 = n37341 ^ n37340 ^ n12783 ;
  assign n37343 = ( n11652 & ~n25586 ) | ( n11652 & n37342 ) | ( ~n25586 & n37342 ) ;
  assign n37344 = n36092 ^ n16806 ^ n8026 ;
  assign n37345 = n33566 ^ n20307 ^ 1'b0 ;
  assign n37346 = ( ~n17946 & n19802 ) | ( ~n17946 & n34768 ) | ( n19802 & n34768 ) ;
  assign n37347 = ( n16692 & n23118 ) | ( n16692 & ~n37346 ) | ( n23118 & ~n37346 ) ;
  assign n37348 = ~n505 & n37347 ;
  assign n37349 = n37348 ^ n14001 ^ 1'b0 ;
  assign n37350 = ( ~n1370 & n6351 ) | ( ~n1370 & n22030 ) | ( n6351 & n22030 ) ;
  assign n37351 = ( n3974 & n24160 ) | ( n3974 & ~n33430 ) | ( n24160 & ~n33430 ) ;
  assign n37352 = ( n17547 & n31264 ) | ( n17547 & n37351 ) | ( n31264 & n37351 ) ;
  assign n37355 = n9132 ^ n8552 ^ n4826 ;
  assign n37353 = n1081 & ~n4703 ;
  assign n37354 = ~n8513 & n37353 ;
  assign n37356 = n37355 ^ n37354 ^ n27520 ;
  assign n37359 = ( n681 & ~n9667 ) | ( n681 & n10940 ) | ( ~n9667 & n10940 ) ;
  assign n37357 = ( n6342 & n7253 ) | ( n6342 & n10043 ) | ( n7253 & n10043 ) ;
  assign n37358 = ( n2494 & n6932 ) | ( n2494 & ~n37357 ) | ( n6932 & ~n37357 ) ;
  assign n37360 = n37359 ^ n37358 ^ n25037 ;
  assign n37361 = n15311 ^ n3816 ^ 1'b0 ;
  assign n37362 = n16417 & ~n37361 ;
  assign n37363 = ( n9319 & ~n17652 ) | ( n9319 & n20150 ) | ( ~n17652 & n20150 ) ;
  assign n37364 = ( n3762 & n31389 ) | ( n3762 & n37363 ) | ( n31389 & n37363 ) ;
  assign n37365 = n14790 & ~n37364 ;
  assign n37366 = n17047 ^ n1734 ^ n1030 ;
  assign n37367 = ( ~n2311 & n17047 ) | ( ~n2311 & n37366 ) | ( n17047 & n37366 ) ;
  assign n37368 = ~n15557 & n22078 ;
  assign n37373 = ~n8430 & n17123 ;
  assign n37374 = n1634 & n37373 ;
  assign n37369 = n10884 ^ n7251 ^ 1'b0 ;
  assign n37370 = n36429 | n37369 ;
  assign n37371 = n13579 | n37370 ;
  assign n37372 = n15142 | n37371 ;
  assign n37375 = n37374 ^ n37372 ^ n5264 ;
  assign n37376 = n18170 & ~n37375 ;
  assign n37377 = ( n4294 & ~n7267 ) | ( n4294 & n35799 ) | ( ~n7267 & n35799 ) ;
  assign n37378 = ~n13898 & n28139 ;
  assign n37379 = n8893 & n37378 ;
  assign n37380 = n3675 ^ x139 ^ x9 ;
  assign n37381 = n13693 ^ n7179 ^ n936 ;
  assign n37382 = ( n21488 & n37380 ) | ( n21488 & n37381 ) | ( n37380 & n37381 ) ;
  assign n37383 = n21407 ^ n10608 ^ n2412 ;
  assign n37384 = ( n8191 & n14246 ) | ( n8191 & n37383 ) | ( n14246 & n37383 ) ;
  assign n37385 = ( ~n5220 & n6531 ) | ( ~n5220 & n37384 ) | ( n6531 & n37384 ) ;
  assign n37386 = ( n10169 & n37382 ) | ( n10169 & ~n37385 ) | ( n37382 & ~n37385 ) ;
  assign n37387 = ( n4134 & ~n7012 ) | ( n4134 & n9178 ) | ( ~n7012 & n9178 ) ;
  assign n37388 = n37387 ^ n25804 ^ n14042 ;
  assign n37389 = n19134 ^ n7045 ^ n5321 ;
  assign n37390 = n37389 ^ n2012 ^ n563 ;
  assign n37391 = n37390 ^ n35963 ^ n33765 ;
  assign n37392 = ~n716 & n2673 ;
  assign n37393 = n37392 ^ n32098 ^ 1'b0 ;
  assign n37394 = n21893 ^ n20697 ^ n6406 ;
  assign n37395 = n6492 & n37394 ;
  assign n37396 = ( n1346 & n10808 ) | ( n1346 & ~n19126 ) | ( n10808 & ~n19126 ) ;
  assign n37397 = n21382 ^ n5323 ^ n4462 ;
  assign n37398 = n11458 ^ n4798 ^ n2237 ;
  assign n37399 = n11855 ^ n2468 ^ 1'b0 ;
  assign n37400 = n37399 ^ n3300 ^ n2146 ;
  assign n37401 = ( ~n3211 & n17065 ) | ( ~n3211 & n17554 ) | ( n17065 & n17554 ) ;
  assign n37402 = n14317 & n37401 ;
  assign n37403 = n37402 ^ n24457 ^ n12587 ;
  assign n37404 = ( n5154 & ~n16791 ) | ( n5154 & n22197 ) | ( ~n16791 & n22197 ) ;
  assign n37405 = n37404 ^ n3022 ^ 1'b0 ;
  assign n37406 = n7451 | n37405 ;
  assign n37407 = n37406 ^ n8673 ^ 1'b0 ;
  assign n37408 = n24462 & n37407 ;
  assign n37409 = ( ~n8586 & n13537 ) | ( ~n8586 & n17475 ) | ( n13537 & n17475 ) ;
  assign n37410 = n10722 ^ x108 ^ 1'b0 ;
  assign n37411 = n35620 ^ n27058 ^ n4801 ;
  assign n37412 = n24189 ^ n23682 ^ n1822 ;
  assign n37413 = n37412 ^ n18002 ^ n17767 ;
  assign n37414 = ( n12827 & n23340 ) | ( n12827 & n37413 ) | ( n23340 & n37413 ) ;
  assign n37416 = ( n10694 & n12426 ) | ( n10694 & ~n18093 ) | ( n12426 & ~n18093 ) ;
  assign n37415 = n18263 ^ n17040 ^ 1'b0 ;
  assign n37417 = n37416 ^ n37415 ^ n2088 ;
  assign n37418 = n32028 ^ n25367 ^ n1189 ;
  assign n37419 = n15315 ^ n14077 ^ n6176 ;
  assign n37420 = n37418 | n37419 ;
  assign n37421 = ~n8384 & n31802 ;
  assign n37422 = n14687 & n37421 ;
  assign n37423 = n37422 ^ x65 ^ 1'b0 ;
  assign n37424 = ( ~n787 & n1670 ) | ( ~n787 & n37423 ) | ( n1670 & n37423 ) ;
  assign n37426 = ( n2990 & ~n19041 ) | ( n2990 & n35518 ) | ( ~n19041 & n35518 ) ;
  assign n37425 = ( ~n12566 & n19336 ) | ( ~n12566 & n34956 ) | ( n19336 & n34956 ) ;
  assign n37427 = n37426 ^ n37425 ^ n898 ;
  assign n37428 = ( n16589 & n25016 ) | ( n16589 & n37427 ) | ( n25016 & n37427 ) ;
  assign n37429 = ( n6085 & ~n7944 ) | ( n6085 & n19026 ) | ( ~n7944 & n19026 ) ;
  assign n37430 = n37429 ^ n25235 ^ n19625 ;
  assign n37431 = ( ~n6477 & n11827 ) | ( ~n6477 & n25167 ) | ( n11827 & n25167 ) ;
  assign n37432 = n8082 & n29569 ;
  assign n37433 = ~n7255 & n37432 ;
  assign n37434 = ( n23875 & ~n37431 ) | ( n23875 & n37433 ) | ( ~n37431 & n37433 ) ;
  assign n37436 = ( n1636 & ~n3732 ) | ( n1636 & n6223 ) | ( ~n3732 & n6223 ) ;
  assign n37435 = n2001 & n33894 ;
  assign n37437 = n37436 ^ n37435 ^ n28657 ;
  assign n37438 = n20071 ^ n17948 ^ n7096 ;
  assign n37439 = n37438 ^ n15429 ^ n14467 ;
  assign n37440 = n355 & ~n37439 ;
  assign n37441 = ( n12198 & ~n25378 ) | ( n12198 & n29176 ) | ( ~n25378 & n29176 ) ;
  assign n37442 = n16459 ^ n5940 ^ x220 ;
  assign n37443 = ( ~n22147 & n23656 ) | ( ~n22147 & n37442 ) | ( n23656 & n37442 ) ;
  assign n37444 = n33056 ^ n28339 ^ n11770 ;
  assign n37445 = ( n5693 & ~n18958 ) | ( n5693 & n24346 ) | ( ~n18958 & n24346 ) ;
  assign n37446 = ( n37443 & n37444 ) | ( n37443 & n37445 ) | ( n37444 & n37445 ) ;
  assign n37447 = n23032 ^ n21679 ^ n10358 ;
  assign n37448 = n37447 ^ n34510 ^ 1'b0 ;
  assign n37449 = n22468 | n25666 ;
  assign n37450 = n37449 ^ n6050 ^ 1'b0 ;
  assign n37451 = n37450 ^ n32953 ^ n4774 ;
  assign n37452 = ( n1081 & n25222 ) | ( n1081 & n25273 ) | ( n25222 & n25273 ) ;
  assign n37453 = ( n12470 & n26577 ) | ( n12470 & ~n37452 ) | ( n26577 & ~n37452 ) ;
  assign n37459 = ( n2493 & n8271 ) | ( n2493 & ~n13222 ) | ( n8271 & ~n13222 ) ;
  assign n37454 = n9746 ^ n7944 ^ n1088 ;
  assign n37455 = ( n12463 & n21842 ) | ( n12463 & ~n37454 ) | ( n21842 & ~n37454 ) ;
  assign n37456 = ( n3617 & n8731 ) | ( n3617 & n16989 ) | ( n8731 & n16989 ) ;
  assign n37457 = n37456 ^ n18494 ^ 1'b0 ;
  assign n37458 = ~n37455 & n37457 ;
  assign n37460 = n37459 ^ n37458 ^ n2368 ;
  assign n37461 = ( n4852 & n9865 ) | ( n4852 & n37460 ) | ( n9865 & n37460 ) ;
  assign n37462 = n36824 ^ n26935 ^ n23143 ;
  assign n37463 = n10057 ^ n4609 ^ 1'b0 ;
  assign n37464 = ~n37462 & n37463 ;
  assign n37465 = n24685 ^ n4027 ^ 1'b0 ;
  assign n37466 = n3207 | n37465 ;
  assign n37467 = ( n5709 & ~n17741 ) | ( n5709 & n23026 ) | ( ~n17741 & n23026 ) ;
  assign n37468 = ( n865 & n3381 ) | ( n865 & ~n8142 ) | ( n3381 & ~n8142 ) ;
  assign n37469 = ( ~n4418 & n31977 ) | ( ~n4418 & n37468 ) | ( n31977 & n37468 ) ;
  assign n37470 = n12233 ^ n1430 ^ 1'b0 ;
  assign n37471 = n16223 & n37470 ;
  assign n37472 = n37471 ^ n34960 ^ n21668 ;
  assign n37473 = n27915 ^ n19324 ^ n16414 ;
  assign n37474 = ( n953 & n22533 ) | ( n953 & ~n37059 ) | ( n22533 & ~n37059 ) ;
  assign n37475 = ( n2901 & n33477 ) | ( n2901 & n37474 ) | ( n33477 & n37474 ) ;
  assign n37476 = ( n18117 & ~n29893 ) | ( n18117 & n37475 ) | ( ~n29893 & n37475 ) ;
  assign n37477 = n22773 ^ n16471 ^ n4625 ;
  assign n37478 = ( n37473 & n37476 ) | ( n37473 & n37477 ) | ( n37476 & n37477 ) ;
  assign n37479 = n37478 ^ n31048 ^ n2168 ;
  assign n37480 = ( ~x247 & n7833 ) | ( ~x247 & n15373 ) | ( n7833 & n15373 ) ;
  assign n37481 = ( n7506 & n22033 ) | ( n7506 & n32329 ) | ( n22033 & n32329 ) ;
  assign n37482 = n36127 ^ n3107 ^ 1'b0 ;
  assign n37483 = ~n12507 & n37482 ;
  assign n37484 = n3131 & ~n8924 ;
  assign n37485 = n4318 & n11113 ;
  assign n37486 = n1593 & n37485 ;
  assign n37487 = n2259 & ~n37486 ;
  assign n37488 = n37487 ^ n4415 ^ 1'b0 ;
  assign n37489 = n37488 ^ n10865 ^ n4077 ;
  assign n37490 = ( n11736 & n16023 ) | ( n11736 & n37489 ) | ( n16023 & n37489 ) ;
  assign n37491 = n37490 ^ n27544 ^ n12373 ;
  assign n37492 = ~n5368 & n31338 ;
  assign n37493 = n37492 ^ n23295 ^ n8152 ;
  assign n37494 = ( n6561 & n10010 ) | ( n6561 & n34691 ) | ( n10010 & n34691 ) ;
  assign n37495 = n32178 ^ n13940 ^ n10063 ;
  assign n37496 = n37495 ^ n4835 ^ n3859 ;
  assign n37497 = ( ~n22205 & n37494 ) | ( ~n22205 & n37496 ) | ( n37494 & n37496 ) ;
  assign n37498 = n37497 ^ n15594 ^ n6481 ;
  assign n37499 = n28732 ^ n26845 ^ n8228 ;
  assign n37500 = x95 & n18871 ;
  assign n37501 = ( n22840 & n37499 ) | ( n22840 & ~n37500 ) | ( n37499 & ~n37500 ) ;
  assign n37502 = ( n9279 & n11879 ) | ( n9279 & ~n12825 ) | ( n11879 & ~n12825 ) ;
  assign n37503 = n37502 ^ n11265 ^ n2757 ;
  assign n37504 = ( n1621 & ~n2613 ) | ( n1621 & n37503 ) | ( ~n2613 & n37503 ) ;
  assign n37505 = n22538 ^ n18480 ^ 1'b0 ;
  assign n37506 = n32606 & n37505 ;
  assign n37507 = n37506 ^ n24427 ^ n14012 ;
  assign n37508 = n33187 ^ n29429 ^ n17489 ;
  assign n37509 = ( ~n8424 & n27231 ) | ( ~n8424 & n37508 ) | ( n27231 & n37508 ) ;
  assign n37510 = n2407 ^ n2284 ^ 1'b0 ;
  assign n37511 = ~n22955 & n37510 ;
  assign n37512 = ~n2335 & n37511 ;
  assign n37513 = n37512 ^ n4203 ^ 1'b0 ;
  assign n37514 = n27437 | n37513 ;
  assign n37515 = n26097 ^ n1936 ^ n990 ;
  assign n37516 = n37515 ^ n30595 ^ n3962 ;
  assign n37517 = n9285 ^ n3637 ^ 1'b0 ;
  assign n37518 = n15144 & ~n37517 ;
  assign n37519 = n25372 ^ n10167 ^ n5607 ;
  assign n37520 = n37519 ^ n23646 ^ 1'b0 ;
  assign n37521 = n11563 & n37520 ;
  assign n37522 = ( n23855 & ~n37518 ) | ( n23855 & n37521 ) | ( ~n37518 & n37521 ) ;
  assign n37523 = ( ~n4155 & n11759 ) | ( ~n4155 & n11975 ) | ( n11759 & n11975 ) ;
  assign n37524 = ( x139 & n16322 ) | ( x139 & ~n37523 ) | ( n16322 & ~n37523 ) ;
  assign n37525 = n23273 ^ n2011 ^ n1150 ;
  assign n37526 = n37525 ^ n27955 ^ n25856 ;
  assign n37527 = ( n20557 & n37524 ) | ( n20557 & ~n37526 ) | ( n37524 & ~n37526 ) ;
  assign n37528 = n10230 ^ n5161 ^ x190 ;
  assign n37529 = n37528 ^ n30859 ^ n11358 ;
  assign n37530 = n37529 ^ n21315 ^ n12938 ;
  assign n37532 = ( n5475 & ~n8603 ) | ( n5475 & n8629 ) | ( ~n8603 & n8629 ) ;
  assign n37531 = n3257 & n33713 ;
  assign n37533 = n37532 ^ n37531 ^ 1'b0 ;
  assign n37534 = n37533 ^ n34673 ^ n19520 ;
  assign n37535 = ( n12955 & n29661 ) | ( n12955 & n37534 ) | ( n29661 & n37534 ) ;
  assign n37537 = n11076 ^ n7122 ^ n1120 ;
  assign n37538 = ( n16015 & ~n29716 ) | ( n16015 & n37537 ) | ( ~n29716 & n37537 ) ;
  assign n37536 = n15754 & n23874 ;
  assign n37539 = n37538 ^ n37536 ^ 1'b0 ;
  assign n37540 = n13999 ^ n7772 ^ n1356 ;
  assign n37541 = n37540 ^ n33249 ^ n13867 ;
  assign n37542 = n24827 ^ n19851 ^ n6694 ;
  assign n37543 = ( n27318 & n32771 ) | ( n27318 & n33226 ) | ( n32771 & n33226 ) ;
  assign n37544 = n4351 & n20728 ;
  assign n37545 = ( n12906 & n13884 ) | ( n12906 & n19974 ) | ( n13884 & n19974 ) ;
  assign n37549 = n18547 & n28704 ;
  assign n37548 = ( n22029 & n25605 ) | ( n22029 & n33099 ) | ( n25605 & n33099 ) ;
  assign n37546 = n11582 & n26107 ;
  assign n37547 = ~n32188 & n37546 ;
  assign n37550 = n37549 ^ n37548 ^ n37547 ;
  assign n37551 = ( n3271 & ~n15775 ) | ( n3271 & n32485 ) | ( ~n15775 & n32485 ) ;
  assign n37552 = ~n31153 & n37551 ;
  assign n37553 = ~n9913 & n37552 ;
  assign n37554 = n37553 ^ n30479 ^ n30379 ;
  assign n37555 = n31476 ^ n20697 ^ n4242 ;
  assign n37556 = n29555 & ~n37555 ;
  assign n37557 = n37556 ^ n1651 ^ 1'b0 ;
  assign n37558 = n23936 ^ n16722 ^ 1'b0 ;
  assign n37559 = ( n1050 & n6836 ) | ( n1050 & n32249 ) | ( n6836 & n32249 ) ;
  assign n37560 = n37559 ^ n18816 ^ n4171 ;
  assign n37561 = ( n9892 & n34401 ) | ( n9892 & n37560 ) | ( n34401 & n37560 ) ;
  assign n37563 = n17787 ^ n17434 ^ 1'b0 ;
  assign n37564 = n7384 & ~n37563 ;
  assign n37562 = ( n17165 & ~n19370 ) | ( n17165 & n25235 ) | ( ~n19370 & n25235 ) ;
  assign n37565 = n37564 ^ n37562 ^ n36182 ;
  assign n37566 = n6858 ^ n6668 ^ 1'b0 ;
  assign n37567 = ( n5033 & ~n24272 ) | ( n5033 & n37566 ) | ( ~n24272 & n37566 ) ;
  assign n37568 = n21901 ^ n6490 ^ n3291 ;
  assign n37569 = n10285 & ~n11341 ;
  assign n37570 = n5958 & n37569 ;
  assign n37571 = n17947 ^ n3498 ^ n2723 ;
  assign n37572 = ( ~n18215 & n21222 ) | ( ~n18215 & n37571 ) | ( n21222 & n37571 ) ;
  assign n37573 = ( n12897 & n17959 ) | ( n12897 & ~n36944 ) | ( n17959 & ~n36944 ) ;
  assign n37574 = n14939 | n24423 ;
  assign n37575 = n37574 ^ x189 ^ 1'b0 ;
  assign n37576 = n37575 ^ n24495 ^ n17164 ;
  assign n37577 = ( n6790 & n21408 ) | ( n6790 & n37576 ) | ( n21408 & n37576 ) ;
  assign n37578 = ( x110 & n12831 ) | ( x110 & n14664 ) | ( n12831 & n14664 ) ;
  assign n37579 = n37578 ^ n24776 ^ n16974 ;
  assign n37580 = n25552 ^ n25129 ^ n16161 ;
  assign n37585 = n6106 ^ n5745 ^ n964 ;
  assign n37582 = n7880 & n12384 ;
  assign n37583 = n37582 ^ n11386 ^ 1'b0 ;
  assign n37584 = ( ~n6923 & n15530 ) | ( ~n6923 & n37583 ) | ( n15530 & n37583 ) ;
  assign n37581 = ( n5346 & n25311 ) | ( n5346 & n27166 ) | ( n25311 & n27166 ) ;
  assign n37586 = n37585 ^ n37584 ^ n37581 ;
  assign n37587 = ( ~n1537 & n16916 ) | ( ~n1537 & n21949 ) | ( n16916 & n21949 ) ;
  assign n37588 = n24541 ^ n3920 ^ n3327 ;
  assign n37589 = n37587 & ~n37588 ;
  assign n37590 = n22696 & n33892 ;
  assign n37591 = n12283 & n37590 ;
  assign n37592 = ( n8011 & ~n17517 ) | ( n8011 & n37140 ) | ( ~n17517 & n37140 ) ;
  assign n37593 = ( n34444 & n37591 ) | ( n34444 & ~n37592 ) | ( n37591 & ~n37592 ) ;
  assign n37594 = n37170 ^ n14611 ^ x2 ;
  assign n37595 = ( n993 & ~n5655 ) | ( n993 & n6093 ) | ( ~n5655 & n6093 ) ;
  assign n37596 = ( n4469 & ~n5752 ) | ( n4469 & n37595 ) | ( ~n5752 & n37595 ) ;
  assign n37597 = n37596 ^ n36723 ^ n5581 ;
  assign n37598 = n25893 ^ n3071 ^ n593 ;
  assign n37599 = n31786 ^ n24753 ^ n16434 ;
  assign n37600 = ( n3607 & n11720 ) | ( n3607 & ~n37599 ) | ( n11720 & ~n37599 ) ;
  assign n37601 = n13401 ^ n4663 ^ 1'b0 ;
  assign n37602 = n37601 ^ n33537 ^ n15013 ;
  assign n37603 = n31764 ^ n19290 ^ n5356 ;
  assign n37609 = ( n4310 & n5225 ) | ( n4310 & n22895 ) | ( n5225 & n22895 ) ;
  assign n37610 = n37609 ^ n17395 ^ n14022 ;
  assign n37611 = n37610 ^ n35199 ^ n1631 ;
  assign n37604 = n34562 ^ n22348 ^ n18717 ;
  assign n37605 = n37604 ^ n22467 ^ n14344 ;
  assign n37606 = n37605 ^ n26037 ^ n21490 ;
  assign n37607 = n16208 & n17203 ;
  assign n37608 = ( n11012 & n37606 ) | ( n11012 & ~n37607 ) | ( n37606 & ~n37607 ) ;
  assign n37612 = n37611 ^ n37608 ^ n27045 ;
  assign n37613 = ( x201 & n3793 ) | ( x201 & ~n5010 ) | ( n3793 & ~n5010 ) ;
  assign n37617 = ( n1201 & ~n6994 ) | ( n1201 & n31406 ) | ( ~n6994 & n31406 ) ;
  assign n37618 = n37617 ^ n17788 ^ n12089 ;
  assign n37614 = n32567 ^ n6173 ^ 1'b0 ;
  assign n37615 = n37614 ^ n37575 ^ n10567 ;
  assign n37616 = n37615 ^ n27912 ^ n15967 ;
  assign n37619 = n37618 ^ n37616 ^ 1'b0 ;
  assign n37620 = n37613 & n37619 ;
  assign n37621 = ( ~n7949 & n22490 ) | ( ~n7949 & n28858 ) | ( n22490 & n28858 ) ;
  assign n37622 = n13436 ^ n13434 ^ n2865 ;
  assign n37623 = n37622 ^ n19026 ^ n3465 ;
  assign n37624 = n37623 ^ n10167 ^ n7293 ;
  assign n37625 = ( n18576 & ~n31603 ) | ( n18576 & n37624 ) | ( ~n31603 & n37624 ) ;
  assign n37626 = n37625 ^ n28592 ^ n11231 ;
  assign n37627 = ( n12362 & n33985 ) | ( n12362 & n37161 ) | ( n33985 & n37161 ) ;
  assign n37628 = n9778 & n37627 ;
  assign n37632 = n13034 ^ n5368 ^ n3132 ;
  assign n37631 = ( n5800 & ~n9128 ) | ( n5800 & n29631 ) | ( ~n9128 & n29631 ) ;
  assign n37629 = n14389 ^ n10178 ^ n1302 ;
  assign n37630 = ( n1434 & n22722 ) | ( n1434 & ~n37629 ) | ( n22722 & ~n37629 ) ;
  assign n37633 = n37632 ^ n37631 ^ n37630 ;
  assign n37634 = n27347 ^ n16491 ^ n6617 ;
  assign n37635 = ( n20156 & n27867 ) | ( n20156 & ~n37634 ) | ( n27867 & ~n37634 ) ;
  assign n37636 = n2674 | n7708 ;
  assign n37637 = n37636 ^ n36779 ^ 1'b0 ;
  assign n37638 = n37637 ^ n17255 ^ n12978 ;
  assign n37639 = ( n7902 & n12454 ) | ( n7902 & n14886 ) | ( n12454 & n14886 ) ;
  assign n37640 = n16275 & ~n37639 ;
  assign n37641 = n36382 ^ n12536 ^ n11125 ;
  assign n37642 = n12294 ^ n10810 ^ 1'b0 ;
  assign n37643 = n25294 & n37642 ;
  assign n37644 = ( n11022 & n37641 ) | ( n11022 & n37643 ) | ( n37641 & n37643 ) ;
  assign n37645 = n8604 ^ n319 ^ 1'b0 ;
  assign n37646 = ( n11924 & ~n12560 ) | ( n11924 & n14654 ) | ( ~n12560 & n14654 ) ;
  assign n37647 = n6365 | n23858 ;
  assign n37648 = n37646 | n37647 ;
  assign n37649 = ( ~n1967 & n37645 ) | ( ~n1967 & n37648 ) | ( n37645 & n37648 ) ;
  assign n37650 = n33444 ^ n32613 ^ n29221 ;
  assign n37651 = n37650 ^ n28192 ^ n793 ;
  assign n37653 = n21547 ^ n14171 ^ 1'b0 ;
  assign n37654 = ( n865 & n2432 ) | ( n865 & n37653 ) | ( n2432 & n37653 ) ;
  assign n37652 = n23238 ^ n6381 ^ 1'b0 ;
  assign n37655 = n37654 ^ n37652 ^ n22900 ;
  assign n37660 = n25526 ^ n3543 ^ n399 ;
  assign n37656 = n14249 ^ n980 ^ 1'b0 ;
  assign n37657 = n3251 | n37656 ;
  assign n37658 = n13677 & n16742 ;
  assign n37659 = n37657 & n37658 ;
  assign n37661 = n37660 ^ n37659 ^ n25586 ;
  assign n37662 = ( ~n7738 & n12901 ) | ( ~n7738 & n19089 ) | ( n12901 & n19089 ) ;
  assign n37663 = ~n28345 & n37662 ;
  assign n37664 = n37663 ^ n27164 ^ 1'b0 ;
  assign n37665 = n37664 ^ n11556 ^ 1'b0 ;
  assign n37666 = ( n3198 & n11073 ) | ( n3198 & ~n16927 ) | ( n11073 & ~n16927 ) ;
  assign n37667 = n12637 & n37666 ;
  assign n37668 = n17964 & n37667 ;
  assign n37669 = n19671 & n22076 ;
  assign n37670 = ~n2883 & n37669 ;
  assign n37671 = ( n1869 & n9270 ) | ( n1869 & n36713 ) | ( n9270 & n36713 ) ;
  assign n37672 = n16812 | n37671 ;
  assign n37673 = n37672 ^ n7292 ^ n1985 ;
  assign n37674 = n9638 | n37673 ;
  assign n37675 = n30987 ^ n21687 ^ 1'b0 ;
  assign n37678 = n7172 & ~n22633 ;
  assign n37679 = n5572 & n37678 ;
  assign n37676 = n16096 ^ n14838 ^ n2011 ;
  assign n37677 = n30459 & ~n37676 ;
  assign n37680 = n37679 ^ n37677 ^ 1'b0 ;
  assign n37681 = n37680 ^ n21119 ^ n18116 ;
  assign n37682 = ( x247 & n2491 ) | ( x247 & n7338 ) | ( n2491 & n7338 ) ;
  assign n37683 = ( n1687 & n22128 ) | ( n1687 & n37682 ) | ( n22128 & n37682 ) ;
  assign n37684 = n13248 & ~n37683 ;
  assign n37685 = ~n35642 & n37684 ;
  assign n37686 = n5642 | n18096 ;
  assign n37687 = ( ~n22170 & n37685 ) | ( ~n22170 & n37686 ) | ( n37685 & n37686 ) ;
  assign n37688 = n26608 ^ n4527 ^ n3683 ;
  assign n37689 = ( n3677 & n9441 ) | ( n3677 & ~n37688 ) | ( n9441 & ~n37688 ) ;
  assign n37690 = n37689 ^ n32875 ^ n1835 ;
  assign n37691 = n11329 & n37690 ;
  assign n37692 = ~n26041 & n37691 ;
  assign n37693 = ( ~n12262 & n12612 ) | ( ~n12262 & n13185 ) | ( n12612 & n13185 ) ;
  assign n37694 = ( n11604 & ~n12332 ) | ( n11604 & n17816 ) | ( ~n12332 & n17816 ) ;
  assign n37695 = n28370 ^ n17572 ^ n4969 ;
  assign n37699 = ~n12947 & n15757 ;
  assign n37700 = n37699 ^ n8846 ^ 1'b0 ;
  assign n37696 = ( n10800 & n11652 ) | ( n10800 & ~n13006 ) | ( n11652 & ~n13006 ) ;
  assign n37697 = n7652 & ~n33591 ;
  assign n37698 = n37696 & ~n37697 ;
  assign n37701 = n37700 ^ n37698 ^ n35269 ;
  assign n37702 = n32831 ^ n19602 ^ n12901 ;
  assign n37703 = n23427 ^ n5481 ^ n5401 ;
  assign n37704 = n35443 ^ n33793 ^ x3 ;
  assign n37705 = ( n15328 & ~n37703 ) | ( n15328 & n37704 ) | ( ~n37703 & n37704 ) ;
  assign n37706 = n31272 ^ n2124 ^ n1532 ;
  assign n37707 = ( ~n5470 & n20510 ) | ( ~n5470 & n21898 ) | ( n20510 & n21898 ) ;
  assign n37708 = n16082 ^ n10877 ^ n6748 ;
  assign n37711 = n13898 ^ n11053 ^ n617 ;
  assign n37710 = ( n8338 & n9924 ) | ( n8338 & ~n19354 ) | ( n9924 & ~n19354 ) ;
  assign n37709 = n14673 ^ n8068 ^ n1265 ;
  assign n37712 = n37711 ^ n37710 ^ n37709 ;
  assign n37713 = ( n12326 & ~n13498 ) | ( n12326 & n14587 ) | ( ~n13498 & n14587 ) ;
  assign n37717 = n17957 ^ n16295 ^ n6025 ;
  assign n37718 = n37717 ^ n3347 ^ n2096 ;
  assign n37714 = n13534 ^ n5968 ^ n805 ;
  assign n37715 = ( n3137 & n7173 ) | ( n3137 & n37714 ) | ( n7173 & n37714 ) ;
  assign n37716 = n37603 & ~n37715 ;
  assign n37719 = n37718 ^ n37716 ^ 1'b0 ;
  assign n37720 = n336 | n17286 ;
  assign n37721 = n37720 ^ n11383 ^ 1'b0 ;
  assign n37722 = n34114 & n37721 ;
  assign n37723 = n19512 & n37722 ;
  assign n37724 = n31387 ^ n27362 ^ n11089 ;
  assign n37725 = n17822 ^ n11067 ^ n4824 ;
  assign n37726 = ( n3656 & n34315 ) | ( n3656 & n35691 ) | ( n34315 & n35691 ) ;
  assign n37727 = ( n5339 & n27819 ) | ( n5339 & ~n37726 ) | ( n27819 & ~n37726 ) ;
  assign n37728 = ( ~n13927 & n15108 ) | ( ~n13927 & n15808 ) | ( n15108 & n15808 ) ;
  assign n37729 = ( n524 & n11317 ) | ( n524 & n30127 ) | ( n11317 & n30127 ) ;
  assign n37730 = n15546 ^ n2012 ^ 1'b0 ;
  assign n37731 = n4742 | n37730 ;
  assign n37732 = ( n3572 & n37729 ) | ( n3572 & n37731 ) | ( n37729 & n37731 ) ;
  assign n37733 = ( n11834 & n14427 ) | ( n11834 & ~n37732 ) | ( n14427 & ~n37732 ) ;
  assign n37734 = ( n7883 & n23377 ) | ( n7883 & n31190 ) | ( n23377 & n31190 ) ;
  assign n37735 = ( n11130 & n37733 ) | ( n11130 & n37734 ) | ( n37733 & n37734 ) ;
  assign n37736 = ( n11768 & n18506 ) | ( n11768 & n26337 ) | ( n18506 & n26337 ) ;
  assign n37737 = n37736 ^ n19538 ^ 1'b0 ;
  assign n37738 = ( ~n14269 & n16302 ) | ( ~n14269 & n31741 ) | ( n16302 & n31741 ) ;
  assign n37739 = n37738 ^ n25482 ^ n9502 ;
  assign n37740 = n20813 ^ n13387 ^ n7905 ;
  assign n37741 = ( n8585 & n37739 ) | ( n8585 & ~n37740 ) | ( n37739 & ~n37740 ) ;
  assign n37742 = x180 & ~n37741 ;
  assign n37743 = n37737 & n37742 ;
  assign n37744 = ( x222 & ~n31177 ) | ( x222 & n31420 ) | ( ~n31177 & n31420 ) ;
  assign n37745 = n37744 ^ n7610 ^ n6553 ;
  assign n37746 = n26698 ^ n17317 ^ n7785 ;
  assign n37747 = n37746 ^ n8885 ^ n2425 ;
  assign n37748 = n18474 ^ n18351 ^ 1'b0 ;
  assign n37749 = n3981 | n37748 ;
  assign n37754 = n9105 ^ n2687 ^ n781 ;
  assign n37752 = n15178 ^ n9876 ^ n2914 ;
  assign n37751 = ( n1994 & n3653 ) | ( n1994 & n30160 ) | ( n3653 & n30160 ) ;
  assign n37753 = n37752 ^ n37751 ^ n14258 ;
  assign n37750 = ( n2587 & n13152 ) | ( n2587 & ~n29394 ) | ( n13152 & ~n29394 ) ;
  assign n37755 = n37754 ^ n37753 ^ n37750 ;
  assign n37756 = ( n727 & ~n3090 ) | ( n727 & n23704 ) | ( ~n3090 & n23704 ) ;
  assign n37757 = ( n5442 & n15222 ) | ( n5442 & ~n15238 ) | ( n15222 & ~n15238 ) ;
  assign n37758 = ( n13184 & n13783 ) | ( n13184 & ~n37757 ) | ( n13783 & ~n37757 ) ;
  assign n37759 = ( n13541 & ~n30258 ) | ( n13541 & n37758 ) | ( ~n30258 & n37758 ) ;
  assign n37760 = n33595 ^ n8595 ^ n2852 ;
  assign n37761 = ( ~n12733 & n29026 ) | ( ~n12733 & n37760 ) | ( n29026 & n37760 ) ;
  assign n37762 = ( ~x192 & n1571 ) | ( ~x192 & n13187 ) | ( n1571 & n13187 ) ;
  assign n37763 = n33036 ^ n13766 ^ n6011 ;
  assign n37764 = ~n1965 & n19477 ;
  assign n37765 = n37764 ^ n31630 ^ 1'b0 ;
  assign n37766 = ( n6248 & ~n8240 ) | ( n6248 & n27594 ) | ( ~n8240 & n27594 ) ;
  assign n37767 = ~n5534 & n37766 ;
  assign n37768 = n12619 & ~n17234 ;
  assign n37769 = ~n33726 & n37768 ;
  assign n37770 = n37769 ^ n4241 ^ 1'b0 ;
  assign n37771 = ( n5782 & n8932 ) | ( n5782 & n37770 ) | ( n8932 & n37770 ) ;
  assign n37772 = n20605 ^ n7941 ^ n4379 ;
  assign n37773 = n20985 ^ n7335 ^ 1'b0 ;
  assign n37774 = ( n33672 & n37772 ) | ( n33672 & n37773 ) | ( n37772 & n37773 ) ;
  assign n37775 = n33194 ^ n31744 ^ n28186 ;
  assign n37778 = ( n1213 & ~n8951 ) | ( n1213 & n11162 ) | ( ~n8951 & n11162 ) ;
  assign n37776 = ( n17951 & n19448 ) | ( n17951 & ~n23642 ) | ( n19448 & ~n23642 ) ;
  assign n37777 = n37776 ^ n32105 ^ n28407 ;
  assign n37779 = n37778 ^ n37777 ^ n36280 ;
  assign n37780 = ( n9287 & n15350 ) | ( n9287 & ~n30578 ) | ( n15350 & ~n30578 ) ;
  assign n37781 = ( n5296 & n18812 ) | ( n5296 & ~n33162 ) | ( n18812 & ~n33162 ) ;
  assign n37782 = n37780 | n37781 ;
  assign n37783 = n26568 | n37782 ;
  assign n37784 = ( n5403 & n8106 ) | ( n5403 & ~n13874 ) | ( n8106 & ~n13874 ) ;
  assign n37785 = ( ~n840 & n12160 ) | ( ~n840 & n16335 ) | ( n12160 & n16335 ) ;
  assign n37786 = ( n3346 & ~n37784 ) | ( n3346 & n37785 ) | ( ~n37784 & n37785 ) ;
  assign n37787 = ( n17741 & n28490 ) | ( n17741 & n37786 ) | ( n28490 & n37786 ) ;
  assign n37788 = ( n27358 & n30515 ) | ( n27358 & n31936 ) | ( n30515 & n31936 ) ;
  assign n37789 = ~n24318 & n25861 ;
  assign n37790 = ~n19188 & n20048 ;
  assign n37791 = n37790 ^ n32917 ^ 1'b0 ;
  assign n37792 = n37791 ^ n28801 ^ n3098 ;
  assign n37793 = ~n37789 & n37792 ;
  assign n37794 = ( n11406 & n23412 ) | ( n11406 & ~n24517 ) | ( n23412 & ~n24517 ) ;
  assign n37796 = n20592 ^ n13831 ^ n341 ;
  assign n37795 = n33694 ^ n27595 ^ n4187 ;
  assign n37797 = n37796 ^ n37795 ^ n31475 ;
  assign n37798 = n37797 ^ n18675 ^ n18380 ;
  assign n37799 = n35793 ^ n25319 ^ n8808 ;
  assign n37800 = n5203 ^ n2277 ^ n365 ;
  assign n37801 = n35337 ^ n33640 ^ n819 ;
  assign n37802 = n22037 ^ n20050 ^ n11194 ;
  assign n37803 = n37802 ^ n28773 ^ n21027 ;
  assign n37804 = n15425 ^ n3710 ^ n2061 ;
  assign n37805 = n37804 ^ n12922 ^ n4234 ;
  assign n37806 = n37805 ^ n16111 ^ n14046 ;
  assign n37807 = n37806 ^ n12521 ^ n3667 ;
  assign n37808 = ( n4783 & n17294 ) | ( n4783 & ~n23494 ) | ( n17294 & ~n23494 ) ;
  assign n37809 = n12345 & ~n37808 ;
  assign n37810 = n37807 & n37809 ;
  assign n37811 = n34912 ^ n25986 ^ n14300 ;
  assign n37812 = ( n4403 & ~n20447 ) | ( n4403 & n37811 ) | ( ~n20447 & n37811 ) ;
  assign n37813 = n6574 & ~n28287 ;
  assign n37814 = ~n37812 & n37813 ;
  assign n37816 = n21759 ^ n4441 ^ n3462 ;
  assign n37817 = ( x115 & n5030 ) | ( x115 & n10515 ) | ( n5030 & n10515 ) ;
  assign n37818 = ( n4688 & n18662 ) | ( n4688 & n37817 ) | ( n18662 & n37817 ) ;
  assign n37819 = ( n10804 & n37816 ) | ( n10804 & ~n37818 ) | ( n37816 & ~n37818 ) ;
  assign n37815 = ( n857 & n21557 ) | ( n857 & ~n33187 ) | ( n21557 & ~n33187 ) ;
  assign n37820 = n37819 ^ n37815 ^ n8693 ;
  assign n37821 = n34726 ^ n21434 ^ n16658 ;
  assign n37822 = ( n1514 & n6228 ) | ( n1514 & ~n19070 ) | ( n6228 & ~n19070 ) ;
  assign n37823 = ( x122 & n5540 ) | ( x122 & n37822 ) | ( n5540 & n37822 ) ;
  assign n37824 = n24631 ^ n8660 ^ n3443 ;
  assign n37826 = n28580 ^ n14652 ^ n12310 ;
  assign n37825 = n16811 ^ n13984 ^ n12664 ;
  assign n37827 = n37826 ^ n37825 ^ n7479 ;
  assign n37828 = ( ~n320 & n2138 ) | ( ~n320 & n25050 ) | ( n2138 & n25050 ) ;
  assign n37829 = n30462 ^ n17159 ^ n11043 ;
  assign n37830 = n36594 ^ n28013 ^ n8464 ;
  assign n37831 = n28951 ^ n9050 ^ n3796 ;
  assign n37833 = ( n20728 & n21044 ) | ( n20728 & ~n25626 ) | ( n21044 & ~n25626 ) ;
  assign n37832 = n12601 ^ n480 ^ 1'b0 ;
  assign n37834 = n37833 ^ n37832 ^ n17424 ;
  assign n37841 = n6744 ^ n5716 ^ 1'b0 ;
  assign n37842 = ~n272 & n37841 ;
  assign n37838 = n7229 ^ n2475 ^ 1'b0 ;
  assign n37839 = n4218 & n37838 ;
  assign n37835 = n8007 | n18157 ;
  assign n37836 = n37835 ^ n19256 ^ 1'b0 ;
  assign n37837 = ( n4488 & n5699 ) | ( n4488 & n37836 ) | ( n5699 & n37836 ) ;
  assign n37840 = n37839 ^ n37837 ^ n10797 ;
  assign n37843 = n37842 ^ n37840 ^ n665 ;
  assign n37844 = n25962 ^ n17699 ^ n5044 ;
  assign n37845 = n37844 ^ n30170 ^ n7880 ;
  assign n37846 = n37845 ^ n27172 ^ n24105 ;
  assign n37847 = n16906 ^ n8957 ^ n8307 ;
  assign n37848 = ~n6046 & n37847 ;
  assign n37849 = n37848 ^ n34578 ^ n31587 ;
  assign n37851 = n5889 & n11847 ;
  assign n37852 = n37851 ^ n15421 ^ n15241 ;
  assign n37850 = n27827 ^ n3648 ^ n1069 ;
  assign n37853 = n37852 ^ n37850 ^ n13322 ;
  assign n37854 = n18330 & ~n36832 ;
  assign n37855 = n35861 ^ n33098 ^ n7523 ;
  assign n37857 = ( n657 & n693 ) | ( n657 & ~n25359 ) | ( n693 & ~n25359 ) ;
  assign n37856 = n14213 ^ n11564 ^ n7535 ;
  assign n37858 = n37857 ^ n37856 ^ n2722 ;
  assign n37859 = n37858 ^ n16473 ^ n9985 ;
  assign n37860 = ( n4408 & n27014 ) | ( n4408 & n34315 ) | ( n27014 & n34315 ) ;
  assign n37861 = n3092 & n9165 ;
  assign n37862 = ( ~n21009 & n37860 ) | ( ~n21009 & n37861 ) | ( n37860 & n37861 ) ;
  assign n37863 = n35637 ^ n26273 ^ n2703 ;
  assign n37864 = ( ~n21568 & n25689 ) | ( ~n21568 & n37863 ) | ( n25689 & n37863 ) ;
  assign n37865 = n31522 ^ n27052 ^ n25592 ;
  assign n37866 = n8056 & n23200 ;
  assign n37867 = n37866 ^ n10494 ^ n5642 ;
  assign n37868 = ( ~n9424 & n9872 ) | ( ~n9424 & n37867 ) | ( n9872 & n37867 ) ;
  assign n37869 = n26184 ^ n20384 ^ 1'b0 ;
  assign n37870 = n15345 & ~n37869 ;
  assign n37871 = ( n9831 & n16481 ) | ( n9831 & ~n37870 ) | ( n16481 & ~n37870 ) ;
  assign n37872 = n37871 ^ n19968 ^ n942 ;
  assign n37873 = ( ~n23651 & n37868 ) | ( ~n23651 & n37872 ) | ( n37868 & n37872 ) ;
  assign n37874 = n31015 ^ n20627 ^ n5470 ;
  assign n37875 = n6170 ^ n297 ^ 1'b0 ;
  assign n37876 = n37874 | n37875 ;
  assign n37877 = ( n9299 & n25832 ) | ( n9299 & n37876 ) | ( n25832 & n37876 ) ;
  assign n37878 = ( ~n8336 & n31675 ) | ( ~n8336 & n35595 ) | ( n31675 & n35595 ) ;
  assign n37879 = ( ~n5296 & n23538 ) | ( ~n5296 & n29101 ) | ( n23538 & n29101 ) ;
  assign n37880 = n19741 | n34288 ;
  assign n37881 = ( ~n8151 & n13261 ) | ( ~n8151 & n24531 ) | ( n13261 & n24531 ) ;
  assign n37887 = n22600 ^ n13164 ^ n2580 ;
  assign n37882 = ( n1606 & n2845 ) | ( n1606 & n22627 ) | ( n2845 & n22627 ) ;
  assign n37883 = n37882 ^ n13602 ^ n11577 ;
  assign n37884 = n37883 ^ n37128 ^ n3159 ;
  assign n37885 = ( ~n14455 & n17211 ) | ( ~n14455 & n37884 ) | ( n17211 & n37884 ) ;
  assign n37886 = ( n3565 & n24554 ) | ( n3565 & n37885 ) | ( n24554 & n37885 ) ;
  assign n37888 = n37887 ^ n37886 ^ n24663 ;
  assign n37889 = ( n20461 & ~n37881 ) | ( n20461 & n37888 ) | ( ~n37881 & n37888 ) ;
  assign n37890 = ( n2016 & ~n6840 ) | ( n2016 & n10940 ) | ( ~n6840 & n10940 ) ;
  assign n37891 = n21623 ^ n15968 ^ n8248 ;
  assign n37892 = n31422 ^ n10131 ^ n342 ;
  assign n37893 = n37892 ^ n31815 ^ 1'b0 ;
  assign n37894 = n32053 ^ n15235 ^ 1'b0 ;
  assign n37895 = n37894 ^ n10418 ^ n4698 ;
  assign n37896 = ( n30556 & n35946 ) | ( n30556 & n37895 ) | ( n35946 & n37895 ) ;
  assign n37897 = ( n3669 & n29856 ) | ( n3669 & ~n37896 ) | ( n29856 & ~n37896 ) ;
  assign n37898 = ~n12091 & n15090 ;
  assign n37899 = ~n2821 & n37898 ;
  assign n37900 = n37899 ^ n26839 ^ n7022 ;
  assign n37901 = n30866 ^ n8820 ^ 1'b0 ;
  assign n37902 = n34703 & ~n37901 ;
  assign n37903 = n29825 ^ n29315 ^ 1'b0 ;
  assign n37904 = n19424 | n37903 ;
  assign n37905 = ~n8912 & n13064 ;
  assign n37906 = n37905 ^ n627 ^ 1'b0 ;
  assign n37907 = n34267 ^ n17231 ^ n12280 ;
  assign n37908 = ~n7195 & n14187 ;
  assign n37909 = n1092 & n37908 ;
  assign n37910 = ( ~n5360 & n20665 ) | ( ~n5360 & n29153 ) | ( n20665 & n29153 ) ;
  assign n37911 = ~n4424 & n8695 ;
  assign n37912 = ( n37909 & n37910 ) | ( n37909 & n37911 ) | ( n37910 & n37911 ) ;
  assign n37913 = ( n37906 & ~n37907 ) | ( n37906 & n37912 ) | ( ~n37907 & n37912 ) ;
  assign n37916 = n20847 ^ n7968 ^ n1159 ;
  assign n37914 = n6488 ^ n3863 ^ 1'b0 ;
  assign n37915 = n37914 ^ n20214 ^ n4811 ;
  assign n37917 = n37916 ^ n37915 ^ n6555 ;
  assign n37921 = n27363 ^ n9066 ^ 1'b0 ;
  assign n37920 = ( n20276 & ~n24407 ) | ( n20276 & n24679 ) | ( ~n24407 & n24679 ) ;
  assign n37918 = n22727 ^ n14790 ^ n8818 ;
  assign n37919 = ( n4384 & ~n16270 ) | ( n4384 & n37918 ) | ( ~n16270 & n37918 ) ;
  assign n37922 = n37921 ^ n37920 ^ n37919 ;
  assign n37923 = n18773 ^ n13992 ^ n6778 ;
  assign n37924 = ( n2817 & n11736 ) | ( n2817 & n19068 ) | ( n11736 & n19068 ) ;
  assign n37925 = ( ~n1615 & n18016 ) | ( ~n1615 & n23707 ) | ( n18016 & n23707 ) ;
  assign n37926 = n21298 & n37925 ;
  assign n37927 = n37926 ^ n32239 ^ n8337 ;
  assign n37928 = ( n3234 & n37924 ) | ( n3234 & n37927 ) | ( n37924 & n37927 ) ;
  assign n37929 = ( ~n14410 & n24633 ) | ( ~n14410 & n37928 ) | ( n24633 & n37928 ) ;
  assign n37930 = n37929 ^ n26133 ^ n7814 ;
  assign n37931 = ~n3511 & n22281 ;
  assign n37932 = n37931 ^ n26673 ^ 1'b0 ;
  assign n37933 = ( n21130 & n21778 ) | ( n21130 & ~n22112 ) | ( n21778 & ~n22112 ) ;
  assign n37934 = ( ~n689 & n10652 ) | ( ~n689 & n37549 ) | ( n10652 & n37549 ) ;
  assign n37935 = ( n7312 & n17848 ) | ( n7312 & ~n37934 ) | ( n17848 & ~n37934 ) ;
  assign n37936 = ( ~n5248 & n6334 ) | ( ~n5248 & n11720 ) | ( n6334 & n11720 ) ;
  assign n37937 = ( ~n4944 & n23926 ) | ( ~n4944 & n37936 ) | ( n23926 & n37936 ) ;
  assign n37938 = ( n17877 & n19989 ) | ( n17877 & n34707 ) | ( n19989 & n34707 ) ;
  assign n37939 = ~n6848 & n33836 ;
  assign n37940 = n10144 & n37939 ;
  assign n37942 = n32232 ^ n29972 ^ n13637 ;
  assign n37941 = n16175 | n25014 ;
  assign n37943 = n37942 ^ n37941 ^ 1'b0 ;
  assign n37944 = n37943 ^ n28679 ^ n16576 ;
  assign n37945 = ( n2954 & n9004 ) | ( n2954 & ~n18780 ) | ( n9004 & ~n18780 ) ;
  assign n37946 = ( ~n11183 & n17776 ) | ( ~n11183 & n37945 ) | ( n17776 & n37945 ) ;
  assign n37947 = ( ~n730 & n36617 ) | ( ~n730 & n37946 ) | ( n36617 & n37946 ) ;
  assign n37948 = ( n4611 & n17415 ) | ( n4611 & n37947 ) | ( n17415 & n37947 ) ;
  assign n37949 = ~n3239 & n5014 ;
  assign n37950 = ~n33353 & n37949 ;
  assign n37951 = n19618 & ~n37950 ;
  assign n37952 = n37951 ^ n18423 ^ 1'b0 ;
  assign n37953 = ( n8802 & ~n14344 ) | ( n8802 & n37952 ) | ( ~n14344 & n37952 ) ;
  assign n37955 = n4071 | n10948 ;
  assign n37956 = n9402 & ~n37955 ;
  assign n37954 = ( ~n4133 & n28805 ) | ( ~n4133 & n35420 ) | ( n28805 & n35420 ) ;
  assign n37957 = n37956 ^ n37954 ^ n12125 ;
  assign n37958 = n20662 ^ n19440 ^ x14 ;
  assign n37959 = ( n10647 & n10769 ) | ( n10647 & n37958 ) | ( n10769 & n37958 ) ;
  assign n37960 = ~n20698 & n37959 ;
  assign n37961 = n33578 ^ n15714 ^ n1261 ;
  assign n37962 = n13578 ^ n11135 ^ n10938 ;
  assign n37963 = ( x203 & n16920 ) | ( x203 & ~n37962 ) | ( n16920 & ~n37962 ) ;
  assign n37964 = n37963 ^ n35562 ^ n11214 ;
  assign n37965 = n37964 ^ n32632 ^ n29593 ;
  assign n37966 = n18552 | n26901 ;
  assign n37967 = n9719 & ~n37966 ;
  assign n37968 = n37967 ^ n32244 ^ n24185 ;
  assign n37969 = ( ~n2612 & n4314 ) | ( ~n2612 & n17479 ) | ( n4314 & n17479 ) ;
  assign n37970 = n37969 ^ n36833 ^ n15483 ;
  assign n37971 = n37970 ^ n9338 ^ n8881 ;
  assign n37972 = ( n20111 & ~n22400 ) | ( n20111 & n37971 ) | ( ~n22400 & n37971 ) ;
  assign n37973 = n25104 ^ n12545 ^ 1'b0 ;
  assign n37974 = ~n12283 & n37973 ;
  assign n37975 = n37974 ^ n21396 ^ n14224 ;
  assign n37976 = ( n7590 & ~n8724 ) | ( n7590 & n34948 ) | ( ~n8724 & n34948 ) ;
  assign n37977 = ( n11786 & n37717 ) | ( n11786 & n37976 ) | ( n37717 & n37976 ) ;
  assign n37978 = n13375 & ~n24384 ;
  assign n37979 = n37978 ^ n6585 ^ 1'b0 ;
  assign n37980 = ( n7809 & n31115 ) | ( n7809 & n37909 ) | ( n31115 & n37909 ) ;
  assign n37981 = n33760 ^ n14902 ^ n14129 ;
  assign n37982 = ( ~n12993 & n24182 ) | ( ~n12993 & n30169 ) | ( n24182 & n30169 ) ;
  assign n37983 = n3368 ^ n2000 ^ n635 ;
  assign n37984 = n37983 ^ n13354 ^ n11557 ;
  assign n37985 = n37984 ^ n16737 ^ n2224 ;
  assign n37986 = ( ~n7549 & n26944 ) | ( ~n7549 & n36395 ) | ( n26944 & n36395 ) ;
  assign n37987 = n37986 ^ n22924 ^ n13077 ;
  assign n37988 = ( ~n21481 & n37985 ) | ( ~n21481 & n37987 ) | ( n37985 & n37987 ) ;
  assign n37989 = n33848 ^ n17623 ^ n3886 ;
  assign n37990 = ( n21748 & n24371 ) | ( n21748 & n35838 ) | ( n24371 & n35838 ) ;
  assign n37991 = n37990 ^ n13437 ^ n2759 ;
  assign n37992 = n2708 | n37991 ;
  assign n37993 = n37992 ^ n23437 ^ 1'b0 ;
  assign n37994 = n37993 ^ n28880 ^ n19840 ;
  assign n37995 = ( n19448 & n37989 ) | ( n19448 & n37994 ) | ( n37989 & n37994 ) ;
  assign n37996 = n1499 & n10784 ;
  assign n37997 = n16514 ^ n10516 ^ 1'b0 ;
  assign n37998 = n13896 & n17394 ;
  assign n37999 = n37997 & n37998 ;
  assign n38000 = n37999 ^ n18948 ^ 1'b0 ;
  assign n38001 = n14469 | n38000 ;
  assign n38002 = n19160 ^ n18717 ^ n11493 ;
  assign n38003 = ( n16767 & n38001 ) | ( n16767 & n38002 ) | ( n38001 & n38002 ) ;
  assign n38007 = n23168 ^ n17220 ^ x153 ;
  assign n38005 = n14202 ^ n8448 ^ x115 ;
  assign n38006 = ( n12226 & n15798 ) | ( n12226 & n38005 ) | ( n15798 & n38005 ) ;
  assign n38004 = n32315 ^ n22278 ^ n2235 ;
  assign n38008 = n38007 ^ n38006 ^ n38004 ;
  assign n38009 = n38008 ^ n32650 ^ n18093 ;
  assign n38010 = n11535 & ~n34578 ;
  assign n38011 = ( n12729 & ~n21498 ) | ( n12729 & n36579 ) | ( ~n21498 & n36579 ) ;
  assign n38012 = n31404 | n38011 ;
  assign n38013 = n38012 ^ n24739 ^ n17088 ;
  assign n38014 = ( ~n7392 & n7574 ) | ( ~n7392 & n27481 ) | ( n7574 & n27481 ) ;
  assign n38015 = ( ~n4039 & n27414 ) | ( ~n4039 & n34907 ) | ( n27414 & n34907 ) ;
  assign n38016 = n38015 ^ n31114 ^ n22977 ;
  assign n38020 = ( n1986 & n22985 ) | ( n1986 & n29462 ) | ( n22985 & n29462 ) ;
  assign n38019 = n12499 ^ n10880 ^ n10253 ;
  assign n38021 = n38020 ^ n38019 ^ n11698 ;
  assign n38017 = ( n4098 & n19139 ) | ( n4098 & n21449 ) | ( n19139 & n21449 ) ;
  assign n38018 = ( ~n7488 & n18199 ) | ( ~n7488 & n38017 ) | ( n18199 & n38017 ) ;
  assign n38022 = n38021 ^ n38018 ^ n8964 ;
  assign n38023 = ( ~n15864 & n31084 ) | ( ~n15864 & n38022 ) | ( n31084 & n38022 ) ;
  assign n38024 = ( n5570 & ~n7819 ) | ( n5570 & n15877 ) | ( ~n7819 & n15877 ) ;
  assign n38025 = ( n1380 & n13655 ) | ( n1380 & ~n38024 ) | ( n13655 & ~n38024 ) ;
  assign n38026 = ( n1430 & n23469 ) | ( n1430 & n38025 ) | ( n23469 & n38025 ) ;
  assign n38027 = n6964 & n22977 ;
  assign n38028 = n38027 ^ n19263 ^ 1'b0 ;
  assign n38029 = n38028 ^ n16335 ^ n6776 ;
  assign n38030 = n38029 ^ n24017 ^ 1'b0 ;
  assign n38031 = n38026 | n38030 ;
  assign n38033 = n9651 & n16135 ;
  assign n38032 = ( ~n4116 & n11118 ) | ( ~n4116 & n22288 ) | ( n11118 & n22288 ) ;
  assign n38034 = n38033 ^ n38032 ^ n28550 ;
  assign n38039 = ( n1980 & n11580 ) | ( n1980 & ~n28301 ) | ( n11580 & ~n28301 ) ;
  assign n38035 = ( n7582 & n8802 ) | ( n7582 & n10098 ) | ( n8802 & n10098 ) ;
  assign n38036 = ( n2954 & ~n3137 ) | ( n2954 & n16544 ) | ( ~n3137 & n16544 ) ;
  assign n38037 = n38035 & n38036 ;
  assign n38038 = n38037 ^ n3920 ^ 1'b0 ;
  assign n38040 = n38039 ^ n38038 ^ n6841 ;
  assign n38043 = ( n3874 & n5278 ) | ( n3874 & n9217 ) | ( n5278 & n9217 ) ;
  assign n38044 = n11871 & n38043 ;
  assign n38045 = ~n26156 & n38044 ;
  assign n38041 = ( n13435 & n27672 ) | ( n13435 & ~n32717 ) | ( n27672 & ~n32717 ) ;
  assign n38042 = n30156 & n38041 ;
  assign n38046 = n38045 ^ n38042 ^ 1'b0 ;
  assign n38047 = ( n4401 & ~n10102 ) | ( n4401 & n30839 ) | ( ~n10102 & n30839 ) ;
  assign n38048 = ( ~n10935 & n19502 ) | ( ~n10935 & n38047 ) | ( n19502 & n38047 ) ;
  assign n38049 = n38048 ^ n17402 ^ 1'b0 ;
  assign n38054 = n29357 ^ n23206 ^ n3281 ;
  assign n38052 = ( x184 & n5452 ) | ( x184 & ~n11724 ) | ( n5452 & ~n11724 ) ;
  assign n38050 = n17947 ^ n7467 ^ n4627 ;
  assign n38051 = ( n6028 & ~n12341 ) | ( n6028 & n38050 ) | ( ~n12341 & n38050 ) ;
  assign n38053 = n38052 ^ n38051 ^ 1'b0 ;
  assign n38055 = n38054 ^ n38053 ^ n4612 ;
  assign n38056 = x169 & ~n9610 ;
  assign n38057 = n38056 ^ n13272 ^ n13069 ;
  assign n38058 = ( ~n9293 & n26461 ) | ( ~n9293 & n32239 ) | ( n26461 & n32239 ) ;
  assign n38059 = ( n31709 & ~n35316 ) | ( n31709 & n38058 ) | ( ~n35316 & n38058 ) ;
  assign n38060 = ~n19905 & n38059 ;
  assign n38061 = n38060 ^ n34696 ^ 1'b0 ;
  assign n38062 = ( n12713 & n14234 ) | ( n12713 & n28779 ) | ( n14234 & n28779 ) ;
  assign n38063 = ~n12503 & n38062 ;
  assign n38064 = n12912 & n38063 ;
  assign n38065 = ~n23250 & n38064 ;
  assign n38066 = n8623 ^ n1014 ^ 1'b0 ;
  assign n38067 = ( n10605 & n11233 ) | ( n10605 & n26360 ) | ( n11233 & n26360 ) ;
  assign n38070 = n6096 ^ n2384 ^ 1'b0 ;
  assign n38068 = ( n1122 & n6497 ) | ( n1122 & n13669 ) | ( n6497 & n13669 ) ;
  assign n38069 = ( n1891 & n28360 ) | ( n1891 & ~n38068 ) | ( n28360 & ~n38068 ) ;
  assign n38071 = n38070 ^ n38069 ^ n3739 ;
  assign n38072 = ( ~n4508 & n38067 ) | ( ~n4508 & n38071 ) | ( n38067 & n38071 ) ;
  assign n38073 = ( n23093 & n35451 ) | ( n23093 & n36833 ) | ( n35451 & n36833 ) ;
  assign n38074 = n34222 ^ n8205 ^ n4617 ;
  assign n38075 = ( n6789 & ~n11968 ) | ( n6789 & n38074 ) | ( ~n11968 & n38074 ) ;
  assign n38076 = n17130 & n38075 ;
  assign n38077 = n2443 | n23365 ;
  assign n38078 = n7163 & ~n38077 ;
  assign n38079 = n38078 ^ n11678 ^ 1'b0 ;
  assign n38080 = n11152 ^ n9463 ^ 1'b0 ;
  assign n38081 = n5588 & n14137 ;
  assign n38082 = n3673 | n34850 ;
  assign n38083 = n25219 ^ n14587 ^ n1793 ;
  assign n38084 = n38083 ^ n7702 ^ 1'b0 ;
  assign n38085 = n11331 ^ n6604 ^ n3123 ;
  assign n38086 = ( n7861 & n21258 ) | ( n7861 & n36240 ) | ( n21258 & n36240 ) ;
  assign n38087 = ( n5562 & n38085 ) | ( n5562 & ~n38086 ) | ( n38085 & ~n38086 ) ;
  assign n38088 = n10491 ^ n6176 ^ n2165 ;
  assign n38089 = ~n758 & n18659 ;
  assign n38090 = n38089 ^ n24101 ^ 1'b0 ;
  assign n38091 = n38090 ^ n13835 ^ n12764 ;
  assign n38092 = ( n4391 & ~n38088 ) | ( n4391 & n38091 ) | ( ~n38088 & n38091 ) ;
  assign n38093 = n34151 ^ n5777 ^ n2431 ;
  assign n38094 = n36402 ^ n16826 ^ n5065 ;
  assign n38095 = ( ~n9111 & n30511 ) | ( ~n9111 & n37119 ) | ( n30511 & n37119 ) ;
  assign n38096 = ( ~n15478 & n31134 ) | ( ~n15478 & n38095 ) | ( n31134 & n38095 ) ;
  assign n38097 = n10689 & ~n31625 ;
  assign n38098 = n4217 | n19793 ;
  assign n38099 = n38097 & ~n38098 ;
  assign n38100 = n38099 ^ n15339 ^ 1'b0 ;
  assign n38101 = ~n38096 & n38100 ;
  assign n38102 = n38101 ^ n34422 ^ n30001 ;
  assign n38103 = ( n25965 & ~n31324 ) | ( n25965 & n38102 ) | ( ~n31324 & n38102 ) ;
  assign n38104 = ( n31214 & n38094 ) | ( n31214 & ~n38103 ) | ( n38094 & ~n38103 ) ;
  assign n38105 = n30837 ^ n30624 ^ n27506 ;
  assign n38106 = n18245 ^ n6575 ^ n6231 ;
  assign n38107 = ( ~n4831 & n26698 ) | ( ~n4831 & n38106 ) | ( n26698 & n38106 ) ;
  assign n38108 = n35527 & n38107 ;
  assign n38114 = ( ~n2797 & n4696 ) | ( ~n2797 & n5781 ) | ( n4696 & n5781 ) ;
  assign n38112 = ( n3888 & n25906 ) | ( n3888 & n35079 ) | ( n25906 & n35079 ) ;
  assign n38111 = ( n15404 & n26750 ) | ( n15404 & ~n34617 ) | ( n26750 & ~n34617 ) ;
  assign n38109 = n21818 ^ n21572 ^ 1'b0 ;
  assign n38110 = ~n6201 & n38109 ;
  assign n38113 = n38112 ^ n38111 ^ n38110 ;
  assign n38115 = n38114 ^ n38113 ^ n22835 ;
  assign n38116 = ( ~n610 & n6878 ) | ( ~n610 & n10724 ) | ( n6878 & n10724 ) ;
  assign n38117 = ( n1354 & ~n7728 ) | ( n1354 & n17565 ) | ( ~n7728 & n17565 ) ;
  assign n38118 = n38117 ^ n8473 ^ n2968 ;
  assign n38119 = n38118 ^ n27668 ^ n2303 ;
  assign n38120 = n38119 ^ n28658 ^ n16538 ;
  assign n38121 = ( n33502 & n38116 ) | ( n33502 & n38120 ) | ( n38116 & n38120 ) ;
  assign n38123 = n21182 ^ n12819 ^ n8524 ;
  assign n38122 = n28704 ^ n25347 ^ n11919 ;
  assign n38124 = n38123 ^ n38122 ^ n32075 ;
  assign n38125 = n38124 ^ n15867 ^ n5656 ;
  assign n38126 = n13174 ^ n5406 ^ 1'b0 ;
  assign n38127 = n17554 & ~n38126 ;
  assign n38128 = ~n1603 & n38127 ;
  assign n38129 = n38128 ^ n28773 ^ 1'b0 ;
  assign n38130 = n33135 ^ n7775 ^ 1'b0 ;
  assign n38131 = ~n18681 & n38130 ;
  assign n38132 = ~n21130 & n24363 ;
  assign n38133 = n1382 & n31703 ;
  assign n38134 = ~n3724 & n38133 ;
  assign n38135 = n38134 ^ n17291 ^ n4994 ;
  assign n38136 = n8319 & n17907 ;
  assign n38137 = ~n21650 & n38136 ;
  assign n38138 = ( n29680 & ~n30631 ) | ( n29680 & n38137 ) | ( ~n30631 & n38137 ) ;
  assign n38139 = ( n5134 & n28115 ) | ( n5134 & ~n38020 ) | ( n28115 & ~n38020 ) ;
  assign n38140 = n10173 ^ n1900 ^ 1'b0 ;
  assign n38141 = n3828 & ~n38140 ;
  assign n38142 = ( ~n27912 & n31350 ) | ( ~n27912 & n38141 ) | ( n31350 & n38141 ) ;
  assign n38143 = n31153 ^ n21833 ^ 1'b0 ;
  assign n38144 = ~n5685 & n38143 ;
  assign n38145 = ( ~n2949 & n17389 ) | ( ~n2949 & n38144 ) | ( n17389 & n38144 ) ;
  assign n38146 = n38145 ^ n14771 ^ n3508 ;
  assign n38148 = ( ~n3706 & n3755 ) | ( ~n3706 & n16568 ) | ( n3755 & n16568 ) ;
  assign n38147 = n24139 ^ n18696 ^ n11651 ;
  assign n38149 = n38148 ^ n38147 ^ n21883 ;
  assign n38150 = ( n4477 & n5990 ) | ( n4477 & n17593 ) | ( n5990 & n17593 ) ;
  assign n38151 = ( n2949 & n22174 ) | ( n2949 & n38150 ) | ( n22174 & n38150 ) ;
  assign n38152 = ( n12553 & n33531 ) | ( n12553 & n38151 ) | ( n33531 & n38151 ) ;
  assign n38153 = n38152 ^ n32575 ^ n1583 ;
  assign n38154 = ( n16473 & n35577 ) | ( n16473 & n38153 ) | ( n35577 & n38153 ) ;
  assign n38155 = n9006 ^ n7930 ^ 1'b0 ;
  assign n38156 = n38155 ^ n23840 ^ n7688 ;
  assign n38157 = n38156 ^ n16510 ^ n4022 ;
  assign n38162 = n24384 ^ n15925 ^ n14410 ;
  assign n38163 = ( n4494 & ~n5237 ) | ( n4494 & n38162 ) | ( ~n5237 & n38162 ) ;
  assign n38160 = ( ~n2284 & n8578 ) | ( ~n2284 & n13600 ) | ( n8578 & n13600 ) ;
  assign n38158 = ( n3199 & n8818 ) | ( n3199 & ~n16632 ) | ( n8818 & ~n16632 ) ;
  assign n38159 = ( n14647 & n21883 ) | ( n14647 & n38158 ) | ( n21883 & n38158 ) ;
  assign n38161 = n38160 ^ n38159 ^ n22473 ;
  assign n38164 = n38163 ^ n38161 ^ 1'b0 ;
  assign n38165 = n29313 ^ n27616 ^ n9808 ;
  assign n38166 = ( ~x157 & n13843 ) | ( ~x157 & n19621 ) | ( n13843 & n19621 ) ;
  assign n38167 = n18045 ^ n11557 ^ 1'b0 ;
  assign n38168 = n24910 ^ n897 ^ 1'b0 ;
  assign n38169 = n1541 & ~n38168 ;
  assign n38170 = n11265 | n31362 ;
  assign n38174 = ( ~n1074 & n12947 ) | ( ~n1074 & n14521 ) | ( n12947 & n14521 ) ;
  assign n38175 = ( n6224 & ~n8573 ) | ( n6224 & n38174 ) | ( ~n8573 & n38174 ) ;
  assign n38171 = n19403 ^ n17197 ^ n9996 ;
  assign n38172 = n20646 & n38171 ;
  assign n38173 = n38172 ^ n13127 ^ 1'b0 ;
  assign n38176 = n38175 ^ n38173 ^ n10043 ;
  assign n38177 = n38176 ^ n17150 ^ n15698 ;
  assign n38178 = ( ~n10136 & n11343 ) | ( ~n10136 & n14717 ) | ( n11343 & n14717 ) ;
  assign n38179 = ( ~n1866 & n20503 ) | ( ~n1866 & n38178 ) | ( n20503 & n38178 ) ;
  assign n38180 = ( n17026 & ~n26610 ) | ( n17026 & n37106 ) | ( ~n26610 & n37106 ) ;
  assign n38181 = ( n6706 & n16608 ) | ( n6706 & n28750 ) | ( n16608 & n28750 ) ;
  assign n38182 = ( n21747 & n32087 ) | ( n21747 & n38181 ) | ( n32087 & n38181 ) ;
  assign n38183 = n38182 ^ n6485 ^ n3713 ;
  assign n38184 = n17387 ^ n13043 ^ n9464 ;
  assign n38185 = ( n13736 & n13966 ) | ( n13736 & ~n38184 ) | ( n13966 & ~n38184 ) ;
  assign n38186 = n18358 ^ n3249 ^ n3043 ;
  assign n38187 = ( ~n18822 & n33760 ) | ( ~n18822 & n38186 ) | ( n33760 & n38186 ) ;
  assign n38189 = n1960 & n32798 ;
  assign n38188 = n26694 ^ n25028 ^ 1'b0 ;
  assign n38190 = n38189 ^ n38188 ^ 1'b0 ;
  assign n38191 = n31057 ^ n19858 ^ n11389 ;
  assign n38192 = n25893 ^ n11710 ^ n2535 ;
  assign n38193 = ( n4306 & ~n11487 ) | ( n4306 & n18983 ) | ( ~n11487 & n18983 ) ;
  assign n38194 = ~n11334 & n38193 ;
  assign n38195 = ~n20323 & n25681 ;
  assign n38196 = ( n993 & n2750 ) | ( n993 & n20859 ) | ( n2750 & n20859 ) ;
  assign n38197 = n33016 ^ n23909 ^ 1'b0 ;
  assign n38198 = n1423 | n38197 ;
  assign n38199 = ( n7959 & n16438 ) | ( n7959 & ~n38198 ) | ( n16438 & ~n38198 ) ;
  assign n38200 = ( n3449 & n38196 ) | ( n3449 & n38199 ) | ( n38196 & n38199 ) ;
  assign n38201 = ( n19720 & ~n30114 ) | ( n19720 & n38200 ) | ( ~n30114 & n38200 ) ;
  assign n38202 = n38201 ^ n13751 ^ 1'b0 ;
  assign n38203 = n26265 ^ n10903 ^ n10582 ;
  assign n38204 = n28732 | n38054 ;
  assign n38205 = n38204 ^ n11807 ^ 1'b0 ;
  assign n38209 = ( n7732 & ~n15453 ) | ( n7732 & n23643 ) | ( ~n15453 & n23643 ) ;
  assign n38206 = n1906 & n17307 ;
  assign n38207 = n4387 & n38206 ;
  assign n38208 = n38207 ^ n35437 ^ n2004 ;
  assign n38210 = n38209 ^ n38208 ^ n21091 ;
  assign n38213 = ( ~n5495 & n17732 ) | ( ~n5495 & n33896 ) | ( n17732 & n33896 ) ;
  assign n38211 = ~n3176 & n12943 ;
  assign n38212 = ( n3908 & n10299 ) | ( n3908 & n38211 ) | ( n10299 & n38211 ) ;
  assign n38214 = n38213 ^ n38212 ^ n12772 ;
  assign n38215 = ( n2010 & ~n18654 ) | ( n2010 & n25484 ) | ( ~n18654 & n25484 ) ;
  assign n38216 = n38215 ^ n17425 ^ 1'b0 ;
  assign n38217 = ~n6520 & n6929 ;
  assign n38218 = ( n38214 & n38216 ) | ( n38214 & n38217 ) | ( n38216 & n38217 ) ;
  assign n38219 = ( ~n38205 & n38210 ) | ( ~n38205 & n38218 ) | ( n38210 & n38218 ) ;
  assign n38220 = n21231 ^ n1764 ^ n388 ;
  assign n38221 = ( n685 & n2320 ) | ( n685 & n3414 ) | ( n2320 & n3414 ) ;
  assign n38222 = n38221 ^ n4708 ^ 1'b0 ;
  assign n38223 = ~n6068 & n38222 ;
  assign n38224 = ( n872 & ~n5990 ) | ( n872 & n38223 ) | ( ~n5990 & n38223 ) ;
  assign n38225 = ( n788 & n38220 ) | ( n788 & n38224 ) | ( n38220 & n38224 ) ;
  assign n38226 = n38225 ^ n25513 ^ n22087 ;
  assign n38227 = n16670 ^ n7727 ^ n4216 ;
  assign n38228 = n38227 ^ n35792 ^ n14428 ;
  assign n38229 = n38228 ^ n23940 ^ n13324 ;
  assign n38230 = ( n21408 & n29099 ) | ( n21408 & n38229 ) | ( n29099 & n38229 ) ;
  assign n38231 = n32774 ^ n9876 ^ n9464 ;
  assign n38232 = ( n4118 & ~n29233 ) | ( n4118 & n38231 ) | ( ~n29233 & n38231 ) ;
  assign n38233 = n30016 ^ n22281 ^ n9209 ;
  assign n38234 = n37717 & ~n38233 ;
  assign n38235 = n10476 ^ n9854 ^ n9509 ;
  assign n38236 = n38234 & ~n38235 ;
  assign n38237 = ~n14623 & n16258 ;
  assign n38238 = ~n9999 & n38237 ;
  assign n38239 = ( ~n9812 & n11395 ) | ( ~n9812 & n27271 ) | ( n11395 & n27271 ) ;
  assign n38240 = n33433 ^ n26604 ^ n19144 ;
  assign n38241 = n20233 & n38240 ;
  assign n38243 = n20182 ^ n363 ^ 1'b0 ;
  assign n38244 = n8201 & ~n38243 ;
  assign n38242 = ( n3283 & n7063 ) | ( n3283 & n10582 ) | ( n7063 & n10582 ) ;
  assign n38245 = n38244 ^ n38242 ^ n28583 ;
  assign n38246 = ( n3281 & ~n24352 ) | ( n3281 & n30594 ) | ( ~n24352 & n30594 ) ;
  assign n38247 = ( n980 & ~n14954 ) | ( n980 & n23197 ) | ( ~n14954 & n23197 ) ;
  assign n38248 = ( n773 & ~n7833 ) | ( n773 & n32107 ) | ( ~n7833 & n32107 ) ;
  assign n38249 = ~n1979 & n24060 ;
  assign n38250 = n29335 ^ n8855 ^ n409 ;
  assign n38251 = ( n36303 & ~n38249 ) | ( n36303 & n38250 ) | ( ~n38249 & n38250 ) ;
  assign n38252 = n15171 ^ n13651 ^ n5946 ;
  assign n38253 = n36770 & ~n38252 ;
  assign n38254 = n38253 ^ n4241 ^ 1'b0 ;
  assign n38255 = n11048 ^ n6332 ^ 1'b0 ;
  assign n38256 = n8116 | n38255 ;
  assign n38257 = ~n3832 & n32038 ;
  assign n38258 = n3003 & n38257 ;
  assign n38260 = n9094 ^ n8236 ^ 1'b0 ;
  assign n38261 = n9778 & ~n38260 ;
  assign n38259 = n511 & n626 ;
  assign n38262 = n38261 ^ n38259 ^ n28077 ;
  assign n38263 = ( n38256 & ~n38258 ) | ( n38256 & n38262 ) | ( ~n38258 & n38262 ) ;
  assign n38264 = n38263 ^ n17789 ^ n7833 ;
  assign n38265 = n32361 ^ n14926 ^ n8230 ;
  assign n38266 = ( ~n1670 & n9844 ) | ( ~n1670 & n38265 ) | ( n9844 & n38265 ) ;
  assign n38267 = ( ~n5136 & n7591 ) | ( ~n5136 & n10973 ) | ( n7591 & n10973 ) ;
  assign n38268 = n38267 ^ n30797 ^ n3711 ;
  assign n38269 = n38268 ^ n35682 ^ n4878 ;
  assign n38270 = n1344 & n16751 ;
  assign n38271 = ( ~n18541 & n20886 ) | ( ~n18541 & n38270 ) | ( n20886 & n38270 ) ;
  assign n38272 = ( n23081 & n34625 ) | ( n23081 & n38271 ) | ( n34625 & n38271 ) ;
  assign n38273 = n28451 ^ n18634 ^ n4608 ;
  assign n38274 = n38273 ^ n24080 ^ n10248 ;
  assign n38275 = ( ~n8095 & n13296 ) | ( ~n8095 & n25722 ) | ( n13296 & n25722 ) ;
  assign n38276 = ( n5326 & n23958 ) | ( n5326 & n38275 ) | ( n23958 & n38275 ) ;
  assign n38277 = ( ~n13232 & n22000 ) | ( ~n13232 & n38276 ) | ( n22000 & n38276 ) ;
  assign n38278 = ( ~x159 & n5547 ) | ( ~x159 & n15901 ) | ( n5547 & n15901 ) ;
  assign n38279 = ( n11855 & n36459 ) | ( n11855 & ~n38278 ) | ( n36459 & ~n38278 ) ;
  assign n38280 = n38279 ^ n22246 ^ n7790 ;
  assign n38281 = n3820 | n11535 ;
  assign n38282 = n38281 ^ n33403 ^ 1'b0 ;
  assign n38283 = n38282 ^ n9633 ^ 1'b0 ;
  assign n38284 = ( ~n6824 & n14330 ) | ( ~n6824 & n22864 ) | ( n14330 & n22864 ) ;
  assign n38285 = n33667 | n38284 ;
  assign n38286 = n20160 ^ n13743 ^ n1751 ;
  assign n38287 = ( n27599 & n36921 ) | ( n27599 & ~n38286 ) | ( n36921 & ~n38286 ) ;
  assign n38288 = n28061 ^ n10010 ^ n8498 ;
  assign n38290 = n18739 ^ n18222 ^ n2210 ;
  assign n38289 = ( n2196 & n17517 ) | ( n2196 & n18605 ) | ( n17517 & n18605 ) ;
  assign n38291 = n38290 ^ n38289 ^ n28641 ;
  assign n38292 = n14030 & n33836 ;
  assign n38293 = n38292 ^ n8966 ^ 1'b0 ;
  assign n38294 = ( n7728 & n38291 ) | ( n7728 & ~n38293 ) | ( n38291 & ~n38293 ) ;
  assign n38295 = ( x246 & n4616 ) | ( x246 & ~n18624 ) | ( n4616 & ~n18624 ) ;
  assign n38296 = n38295 ^ n31779 ^ n23844 ;
  assign n38300 = n24726 ^ n20953 ^ n15677 ;
  assign n38298 = ( ~n2118 & n7712 ) | ( ~n2118 & n12781 ) | ( n7712 & n12781 ) ;
  assign n38299 = n38298 ^ n10938 ^ n450 ;
  assign n38301 = n38300 ^ n38299 ^ n3469 ;
  assign n38297 = n36335 ^ n33590 ^ n33011 ;
  assign n38302 = n38301 ^ n38297 ^ n16035 ;
  assign n38303 = ~n21251 & n31177 ;
  assign n38304 = ( ~n552 & n1774 ) | ( ~n552 & n24117 ) | ( n1774 & n24117 ) ;
  assign n38305 = n17901 ^ n16085 ^ n11546 ;
  assign n38306 = n38305 ^ n25255 ^ n16084 ;
  assign n38307 = n3143 | n33497 ;
  assign n38308 = n38307 ^ n11614 ^ 1'b0 ;
  assign n38309 = n16705 & ~n38308 ;
  assign n38310 = n38309 ^ n18334 ^ n7371 ;
  assign n38311 = ( n6465 & n38306 ) | ( n6465 & ~n38310 ) | ( n38306 & ~n38310 ) ;
  assign n38312 = n1805 & n13973 ;
  assign n38313 = ~n14545 & n38312 ;
  assign n38314 = ( n11676 & ~n14168 ) | ( n11676 & n34745 ) | ( ~n14168 & n34745 ) ;
  assign n38315 = ( n7776 & ~n10308 ) | ( n7776 & n38314 ) | ( ~n10308 & n38314 ) ;
  assign n38316 = n38315 ^ n26568 ^ n24221 ;
  assign n38317 = ( ~n10835 & n23333 ) | ( ~n10835 & n31985 ) | ( n23333 & n31985 ) ;
  assign n38318 = ( n6139 & n10103 ) | ( n6139 & n38317 ) | ( n10103 & n38317 ) ;
  assign n38319 = n38318 ^ n36468 ^ n32420 ;
  assign n38320 = n38319 ^ n10225 ^ 1'b0 ;
  assign n38321 = n23367 ^ n9588 ^ n7941 ;
  assign n38322 = n38321 ^ n11575 ^ n6702 ;
  assign n38323 = ( n18692 & ~n20844 ) | ( n18692 & n35112 ) | ( ~n20844 & n35112 ) ;
  assign n38324 = ( n804 & n18139 ) | ( n804 & n38323 ) | ( n18139 & n38323 ) ;
  assign n38325 = n38324 ^ n10999 ^ n10595 ;
  assign n38326 = ( ~n14356 & n22812 ) | ( ~n14356 & n25602 ) | ( n22812 & n25602 ) ;
  assign n38327 = n38326 ^ n17594 ^ n16570 ;
  assign n38328 = ( n1979 & ~n10248 ) | ( n1979 & n28687 ) | ( ~n10248 & n28687 ) ;
  assign n38329 = ( n5360 & n7994 ) | ( n5360 & ~n34279 ) | ( n7994 & ~n34279 ) ;
  assign n38330 = ( n4058 & n11826 ) | ( n4058 & ~n38329 ) | ( n11826 & ~n38329 ) ;
  assign n38331 = ( n3199 & ~n31618 ) | ( n3199 & n38330 ) | ( ~n31618 & n38330 ) ;
  assign n38332 = n9033 & ~n32576 ;
  assign n38333 = n38332 ^ n34682 ^ n32571 ;
  assign n38334 = n3155 & n24200 ;
  assign n38335 = n14191 & n38334 ;
  assign n38338 = n15909 ^ n6635 ^ n1588 ;
  assign n38336 = n28936 ^ n1709 ^ n559 ;
  assign n38337 = ( n15468 & n16696 ) | ( n15468 & n38336 ) | ( n16696 & n38336 ) ;
  assign n38339 = n38338 ^ n38337 ^ 1'b0 ;
  assign n38340 = n9148 & ~n38339 ;
  assign n38341 = n38340 ^ n31407 ^ n21936 ;
  assign n38342 = n37587 ^ n6810 ^ 1'b0 ;
  assign n38343 = n38341 & n38342 ;
  assign n38344 = ~n3019 & n20733 ;
  assign n38345 = n12732 | n38344 ;
  assign n38346 = ~n4685 & n32756 ;
  assign n38347 = n38346 ^ n27342 ^ 1'b0 ;
  assign n38348 = ( n15934 & n27208 ) | ( n15934 & ~n38347 ) | ( n27208 & ~n38347 ) ;
  assign n38349 = n6865 ^ n3984 ^ n3552 ;
  assign n38350 = ( n4216 & ~n7544 ) | ( n4216 & n28867 ) | ( ~n7544 & n28867 ) ;
  assign n38351 = n38350 ^ n20593 ^ n513 ;
  assign n38352 = n38351 ^ n19018 ^ n1749 ;
  assign n38353 = n22915 ^ n18538 ^ n15034 ;
  assign n38354 = n9379 & n18513 ;
  assign n38355 = n11768 & n38354 ;
  assign n38356 = ( n6939 & n10144 ) | ( n6939 & ~n15610 ) | ( n10144 & ~n15610 ) ;
  assign n38357 = n13803 ^ n4924 ^ n3624 ;
  assign n38358 = n19440 ^ n18632 ^ n6792 ;
  assign n38359 = ( n32851 & n38357 ) | ( n32851 & n38358 ) | ( n38357 & n38358 ) ;
  assign n38360 = ( n4502 & n38356 ) | ( n4502 & n38359 ) | ( n38356 & n38359 ) ;
  assign n38361 = ( n2280 & ~n8078 ) | ( n2280 & n30190 ) | ( ~n8078 & n30190 ) ;
  assign n38362 = n22104 & n35264 ;
  assign n38363 = n38362 ^ n23030 ^ 1'b0 ;
  assign n38364 = n38361 & ~n38363 ;
  assign n38365 = n38364 ^ n31547 ^ 1'b0 ;
  assign n38366 = n27390 ^ n24981 ^ 1'b0 ;
  assign n38367 = n38366 ^ n28097 ^ n1915 ;
  assign n38368 = ( n1746 & ~n31969 ) | ( n1746 & n38367 ) | ( ~n31969 & n38367 ) ;
  assign n38369 = ( n3303 & n9538 ) | ( n3303 & ~n22454 ) | ( n9538 & ~n22454 ) ;
  assign n38376 = ( n2820 & ~n4271 ) | ( n2820 & n11051 ) | ( ~n4271 & n11051 ) ;
  assign n38375 = n860 | n28887 ;
  assign n38377 = n38376 ^ n38375 ^ 1'b0 ;
  assign n38372 = x89 & n22247 ;
  assign n38373 = n11508 & n38372 ;
  assign n38374 = n38373 ^ n11035 ^ 1'b0 ;
  assign n38370 = ( n8129 & ~n13843 ) | ( n8129 & n17496 ) | ( ~n13843 & n17496 ) ;
  assign n38371 = ( n9386 & ~n31868 ) | ( n9386 & n38370 ) | ( ~n31868 & n38370 ) ;
  assign n38378 = n38377 ^ n38374 ^ n38371 ;
  assign n38379 = ~n6729 & n35154 ;
  assign n38380 = n38379 ^ n6890 ^ 1'b0 ;
  assign n38381 = ( n14620 & n20398 ) | ( n14620 & ~n32753 ) | ( n20398 & ~n32753 ) ;
  assign n38382 = n38381 ^ n18732 ^ n17948 ;
  assign n38383 = ~n7501 & n28117 ;
  assign n38384 = n1889 & n6829 ;
  assign n38385 = n38384 ^ n32913 ^ 1'b0 ;
  assign n38386 = n38385 ^ n35929 ^ n27565 ;
  assign n38387 = ( n33404 & n36952 ) | ( n33404 & ~n38386 ) | ( n36952 & ~n38386 ) ;
  assign n38390 = ( n1440 & n21728 ) | ( n1440 & ~n27302 ) | ( n21728 & ~n27302 ) ;
  assign n38388 = n4072 ^ n2141 ^ n1034 ;
  assign n38389 = ( n19069 & n37204 ) | ( n19069 & n38388 ) | ( n37204 & n38388 ) ;
  assign n38391 = n38390 ^ n38389 ^ n23854 ;
  assign n38392 = n4305 & ~n8524 ;
  assign n38393 = n38392 ^ n13530 ^ 1'b0 ;
  assign n38394 = ( n23082 & ~n23280 ) | ( n23082 & n26528 ) | ( ~n23280 & n26528 ) ;
  assign n38400 = n13291 | n24586 ;
  assign n38401 = ( n3540 & n19583 ) | ( n3540 & ~n38400 ) | ( n19583 & ~n38400 ) ;
  assign n38395 = ( n2866 & ~n5818 ) | ( n2866 & n25360 ) | ( ~n5818 & n25360 ) ;
  assign n38396 = ( ~n12143 & n16304 ) | ( ~n12143 & n31024 ) | ( n16304 & n31024 ) ;
  assign n38397 = ~n23879 & n38396 ;
  assign n38398 = ~n7231 & n38397 ;
  assign n38399 = ( n17599 & n38395 ) | ( n17599 & ~n38398 ) | ( n38395 & ~n38398 ) ;
  assign n38402 = n38401 ^ n38399 ^ n13363 ;
  assign n38403 = ( n13864 & ~n32257 ) | ( n13864 & n37496 ) | ( ~n32257 & n37496 ) ;
  assign n38404 = n38403 ^ n25638 ^ n9897 ;
  assign n38405 = n38404 ^ n34412 ^ n4082 ;
  assign n38406 = n37499 ^ n36382 ^ n12200 ;
  assign n38407 = n15263 ^ n2761 ^ 1'b0 ;
  assign n38408 = ~n21651 & n38407 ;
  assign n38409 = n38408 ^ n10205 ^ n7409 ;
  assign n38413 = ~n736 & n10689 ;
  assign n38414 = n38413 ^ n6633 ^ 1'b0 ;
  assign n38410 = ~n13822 & n20063 ;
  assign n38411 = ~n17555 & n38410 ;
  assign n38412 = ( n8737 & n20952 ) | ( n8737 & ~n38411 ) | ( n20952 & ~n38411 ) ;
  assign n38415 = n38414 ^ n38412 ^ 1'b0 ;
  assign n38416 = ( n6584 & ~n38409 ) | ( n6584 & n38415 ) | ( ~n38409 & n38415 ) ;
  assign n38417 = n13999 ^ n13592 ^ n3327 ;
  assign n38418 = ( n1560 & ~n29858 ) | ( n1560 & n38417 ) | ( ~n29858 & n38417 ) ;
  assign n38419 = n33093 ^ n9192 ^ 1'b0 ;
  assign n38420 = n14076 | n38419 ;
  assign n38421 = n12555 ^ n8277 ^ 1'b0 ;
  assign n38422 = ( n377 & n25488 ) | ( n377 & n38421 ) | ( n25488 & n38421 ) ;
  assign n38423 = ( n10152 & n33621 ) | ( n10152 & n38422 ) | ( n33621 & n38422 ) ;
  assign n38426 = ( n467 & n12951 ) | ( n467 & n24276 ) | ( n12951 & n24276 ) ;
  assign n38427 = ( n19773 & n37341 ) | ( n19773 & n38426 ) | ( n37341 & n38426 ) ;
  assign n38428 = ( n6866 & n21837 ) | ( n6866 & n38427 ) | ( n21837 & n38427 ) ;
  assign n38424 = n4534 & n25828 ;
  assign n38425 = ( ~n5894 & n32530 ) | ( ~n5894 & n38424 ) | ( n32530 & n38424 ) ;
  assign n38429 = n38428 ^ n38425 ^ n5598 ;
  assign n38430 = ( n6656 & ~n12636 ) | ( n6656 & n14570 ) | ( ~n12636 & n14570 ) ;
  assign n38431 = ( n5495 & n12465 ) | ( n5495 & n38430 ) | ( n12465 & n38430 ) ;
  assign n38432 = n38431 ^ n36406 ^ n12630 ;
  assign n38433 = n38432 ^ n35060 ^ n433 ;
  assign n38434 = n38433 ^ n29339 ^ n9650 ;
  assign n38435 = n27913 ^ n20417 ^ n11022 ;
  assign n38436 = ( ~n18980 & n19819 ) | ( ~n18980 & n29666 ) | ( n19819 & n29666 ) ;
  assign n38437 = ( n1578 & n8081 ) | ( n1578 & n38436 ) | ( n8081 & n38436 ) ;
  assign n38438 = n2203 ^ n1993 ^ 1'b0 ;
  assign n38440 = n21651 ^ n16501 ^ n4412 ;
  assign n38439 = ( ~n19364 & n19737 ) | ( ~n19364 & n29381 ) | ( n19737 & n29381 ) ;
  assign n38441 = n38440 ^ n38439 ^ n31440 ;
  assign n38442 = ( n2644 & ~n38438 ) | ( n2644 & n38441 ) | ( ~n38438 & n38441 ) ;
  assign n38443 = ( n3501 & n3734 ) | ( n3501 & ~n8142 ) | ( n3734 & ~n8142 ) ;
  assign n38444 = ( n7754 & n27733 ) | ( n7754 & ~n34636 ) | ( n27733 & ~n34636 ) ;
  assign n38445 = n2059 | n11653 ;
  assign n38446 = ( n11536 & n30076 ) | ( n11536 & ~n38445 ) | ( n30076 & ~n38445 ) ;
  assign n38447 = ( x224 & n12884 ) | ( x224 & ~n38446 ) | ( n12884 & ~n38446 ) ;
  assign n38448 = ( ~n38443 & n38444 ) | ( ~n38443 & n38447 ) | ( n38444 & n38447 ) ;
  assign n38449 = ( n27364 & ~n30455 ) | ( n27364 & n34728 ) | ( ~n30455 & n34728 ) ;
  assign n38450 = ( n2491 & n35751 ) | ( n2491 & n38449 ) | ( n35751 & n38449 ) ;
  assign n38451 = n38450 ^ n34572 ^ n23406 ;
  assign n38452 = n38451 ^ n20202 ^ n11932 ;
  assign n38453 = n8989 ^ n265 ^ 1'b0 ;
  assign n38454 = n38453 ^ n35957 ^ n7717 ;
  assign n38457 = n25399 ^ n22481 ^ n22048 ;
  assign n38455 = ( n2047 & ~n12849 ) | ( n2047 & n17801 ) | ( ~n12849 & n17801 ) ;
  assign n38456 = n38455 ^ n22613 ^ n19176 ;
  assign n38458 = n38457 ^ n38456 ^ n11388 ;
  assign n38459 = n985 & ~n15690 ;
  assign n38460 = n38459 ^ n8892 ^ n7595 ;
  assign n38461 = ( n631 & ~n2059 ) | ( n631 & n38460 ) | ( ~n2059 & n38460 ) ;
  assign n38462 = n31596 ^ n24647 ^ n18929 ;
  assign n38463 = n20511 ^ n17030 ^ n15513 ;
  assign n38464 = ( ~n34377 & n34631 ) | ( ~n34377 & n38463 ) | ( n34631 & n38463 ) ;
  assign n38465 = n20234 ^ n6078 ^ n426 ;
  assign n38466 = n38465 ^ n6833 ^ n3904 ;
  assign n38467 = n2320 | n38466 ;
  assign n38468 = ( n24076 & n34253 ) | ( n24076 & ~n38467 ) | ( n34253 & ~n38467 ) ;
  assign n38469 = n18394 ^ n4519 ^ 1'b0 ;
  assign n38470 = n8824 & n38469 ;
  assign n38471 = ( n2875 & ~n3829 ) | ( n2875 & n6679 ) | ( ~n3829 & n6679 ) ;
  assign n38472 = n38471 ^ n17373 ^ n4298 ;
  assign n38473 = ( n8429 & n19846 ) | ( n8429 & n20697 ) | ( n19846 & n20697 ) ;
  assign n38474 = ( n15197 & n16090 ) | ( n15197 & n27751 ) | ( n16090 & n27751 ) ;
  assign n38475 = ( ~n23378 & n38473 ) | ( ~n23378 & n38474 ) | ( n38473 & n38474 ) ;
  assign n38476 = n11420 ^ n10207 ^ n331 ;
  assign n38477 = n38476 ^ n31278 ^ n12203 ;
  assign n38478 = ( n8003 & n9056 ) | ( n8003 & ~n38477 ) | ( n9056 & ~n38477 ) ;
  assign n38479 = ( n6660 & n20746 ) | ( n6660 & n37955 ) | ( n20746 & n37955 ) ;
  assign n38480 = ( ~n9197 & n13104 ) | ( ~n9197 & n22588 ) | ( n13104 & n22588 ) ;
  assign n38481 = ( n1451 & n15917 ) | ( n1451 & n38480 ) | ( n15917 & n38480 ) ;
  assign n38484 = ( n21764 & ~n28537 ) | ( n21764 & n33753 ) | ( ~n28537 & n33753 ) ;
  assign n38482 = n21446 ^ n18938 ^ n581 ;
  assign n38483 = n20348 | n38482 ;
  assign n38485 = n38484 ^ n38483 ^ 1'b0 ;
  assign n38486 = ( n6834 & ~n17593 ) | ( n6834 & n19582 ) | ( ~n17593 & n19582 ) ;
  assign n38487 = n9298 & ~n21046 ;
  assign n38488 = ~n17871 & n38487 ;
  assign n38489 = ~n38486 & n38488 ;
  assign n38490 = ( n5110 & n6355 ) | ( n5110 & ~n29758 ) | ( n6355 & ~n29758 ) ;
  assign n38491 = n16386 ^ n4678 ^ 1'b0 ;
  assign n38492 = ( ~n23399 & n38490 ) | ( ~n23399 & n38491 ) | ( n38490 & n38491 ) ;
  assign n38493 = n24803 ^ n12712 ^ n10736 ;
  assign n38494 = ( ~n6536 & n14389 ) | ( ~n6536 & n23747 ) | ( n14389 & n23747 ) ;
  assign n38495 = n38494 ^ n7889 ^ n4896 ;
  assign n38496 = ( n37174 & n38493 ) | ( n37174 & ~n38495 ) | ( n38493 & ~n38495 ) ;
  assign n38497 = ( ~n6162 & n7972 ) | ( ~n6162 & n10833 ) | ( n7972 & n10833 ) ;
  assign n38498 = ( n17901 & n30289 ) | ( n17901 & n38497 ) | ( n30289 & n38497 ) ;
  assign n38499 = x152 & ~n8174 ;
  assign n38500 = n38499 ^ n8970 ^ 1'b0 ;
  assign n38501 = ( n16239 & ~n20443 ) | ( n16239 & n38062 ) | ( ~n20443 & n38062 ) ;
  assign n38502 = n38501 ^ n5874 ^ 1'b0 ;
  assign n38503 = n38502 ^ n21713 ^ n20007 ;
  assign n38504 = n10507 & n14945 ;
  assign n38505 = ~n38503 & n38504 ;
  assign n38507 = n1879 & ~n5573 ;
  assign n38508 = n17259 & n38507 ;
  assign n38509 = n38508 ^ n33099 ^ n6099 ;
  assign n38510 = n7248 & n38509 ;
  assign n38506 = ( n15273 & n26102 ) | ( n15273 & ~n36670 ) | ( n26102 & ~n36670 ) ;
  assign n38511 = n38510 ^ n38506 ^ n13632 ;
  assign n38512 = ( n3905 & ~n13932 ) | ( n3905 & n38511 ) | ( ~n13932 & n38511 ) ;
  assign n38513 = n10220 ^ n6037 ^ 1'b0 ;
  assign n38514 = ( n12807 & ~n14227 ) | ( n12807 & n38513 ) | ( ~n14227 & n38513 ) ;
  assign n38515 = ( n1488 & n6488 ) | ( n1488 & ~n9364 ) | ( n6488 & ~n9364 ) ;
  assign n38516 = n38515 ^ n6470 ^ n536 ;
  assign n38517 = n22160 ^ x0 ^ 1'b0 ;
  assign n38518 = n38516 & n38517 ;
  assign n38519 = ( n326 & ~n15515 ) | ( n326 & n38518 ) | ( ~n15515 & n38518 ) ;
  assign n38520 = ( n9188 & n10951 ) | ( n9188 & n14396 ) | ( n10951 & n14396 ) ;
  assign n38521 = ( n29792 & n38519 ) | ( n29792 & n38520 ) | ( n38519 & n38520 ) ;
  assign n38522 = ( ~n16587 & n26655 ) | ( ~n16587 & n38521 ) | ( n26655 & n38521 ) ;
  assign n38523 = ( n9739 & ~n18672 ) | ( n9739 & n20346 ) | ( ~n18672 & n20346 ) ;
  assign n38524 = n28361 ^ n23054 ^ n19448 ;
  assign n38525 = n30950 ^ n30414 ^ n21599 ;
  assign n38526 = n15173 ^ n11153 ^ n6836 ;
  assign n38527 = ( ~n4094 & n7047 ) | ( ~n4094 & n38526 ) | ( n7047 & n38526 ) ;
  assign n38528 = ( ~n17303 & n25379 ) | ( ~n17303 & n38527 ) | ( n25379 & n38527 ) ;
  assign n38529 = n38528 ^ n37140 ^ n35312 ;
  assign n38530 = n38529 ^ n22255 ^ n3702 ;
  assign n38531 = n38530 ^ n24110 ^ n21088 ;
  assign n38532 = ( n4187 & n11113 ) | ( n4187 & ~n13687 ) | ( n11113 & ~n13687 ) ;
  assign n38534 = n28532 ^ n9215 ^ n7883 ;
  assign n38533 = ( n7188 & n23734 ) | ( n7188 & n27172 ) | ( n23734 & n27172 ) ;
  assign n38535 = n38534 ^ n38533 ^ n27240 ;
  assign n38536 = ( n825 & n6828 ) | ( n825 & ~n9628 ) | ( n6828 & ~n9628 ) ;
  assign n38537 = n38536 ^ n16993 ^ n14652 ;
  assign n38538 = n38537 ^ n32833 ^ n29745 ;
  assign n38539 = n38538 ^ n25910 ^ n13132 ;
  assign n38540 = n13973 ^ n4274 ^ 1'b0 ;
  assign n38541 = ~n19156 & n38540 ;
  assign n38542 = ~n13324 & n20626 ;
  assign n38543 = ~n38541 & n38542 ;
  assign n38544 = n38543 ^ n22688 ^ n22568 ;
  assign n38545 = ( n38535 & ~n38539 ) | ( n38535 & n38544 ) | ( ~n38539 & n38544 ) ;
  assign n38546 = ( n14892 & n21881 ) | ( n14892 & ~n29370 ) | ( n21881 & ~n29370 ) ;
  assign n38547 = n38546 ^ n17340 ^ n15046 ;
  assign n38548 = n26800 ^ n17860 ^ n11120 ;
  assign n38549 = n26691 & n38548 ;
  assign n38550 = ~n10249 & n38549 ;
  assign n38551 = ( ~n8129 & n22794 ) | ( ~n8129 & n38244 ) | ( n22794 & n38244 ) ;
  assign n38552 = n7892 & ~n12552 ;
  assign n38553 = n9964 & ~n27709 ;
  assign n38554 = n38553 ^ n13998 ^ 1'b0 ;
  assign n38555 = ( ~n6090 & n9248 ) | ( ~n6090 & n12672 ) | ( n9248 & n12672 ) ;
  assign n38556 = ( n18149 & n22461 ) | ( n18149 & ~n38555 ) | ( n22461 & ~n38555 ) ;
  assign n38557 = n38556 ^ n23986 ^ n18860 ;
  assign n38558 = ( n32760 & n32891 ) | ( n32760 & ~n38557 ) | ( n32891 & ~n38557 ) ;
  assign n38559 = ( n30725 & ~n38554 ) | ( n30725 & n38558 ) | ( ~n38554 & n38558 ) ;
  assign n38560 = ( n9790 & n38552 ) | ( n9790 & n38559 ) | ( n38552 & n38559 ) ;
  assign n38561 = n24488 ^ n14240 ^ n3336 ;
  assign n38562 = n37870 ^ n462 ^ 1'b0 ;
  assign n38563 = ( n15232 & n20521 ) | ( n15232 & n26838 ) | ( n20521 & n26838 ) ;
  assign n38564 = n38563 ^ n36436 ^ n27701 ;
  assign n38565 = ( n29126 & n38562 ) | ( n29126 & n38564 ) | ( n38562 & n38564 ) ;
  assign n38566 = ( ~n2590 & n3074 ) | ( ~n2590 & n23270 ) | ( n3074 & n23270 ) ;
  assign n38567 = n38566 ^ n37277 ^ n3334 ;
  assign n38568 = ( n38561 & n38565 ) | ( n38561 & n38567 ) | ( n38565 & n38567 ) ;
  assign n38569 = n1662 & n7771 ;
  assign n38570 = ( n4493 & ~n10146 ) | ( n4493 & n38569 ) | ( ~n10146 & n38569 ) ;
  assign n38571 = ( n5794 & n16629 ) | ( n5794 & ~n21554 ) | ( n16629 & ~n21554 ) ;
  assign n38572 = n38571 ^ n25316 ^ n9633 ;
  assign n38573 = n17740 ^ n17218 ^ n11897 ;
  assign n38575 = ( ~n7388 & n7588 ) | ( ~n7388 & n14740 ) | ( n7588 & n14740 ) ;
  assign n38576 = n7702 & n38575 ;
  assign n38577 = n38576 ^ n11940 ^ 1'b0 ;
  assign n38578 = n5656 ^ n5265 ^ n340 ;
  assign n38579 = ( n7145 & ~n16006 ) | ( n7145 & n33444 ) | ( ~n16006 & n33444 ) ;
  assign n38580 = ( ~n18090 & n38578 ) | ( ~n18090 & n38579 ) | ( n38578 & n38579 ) ;
  assign n38581 = ~n13931 & n38580 ;
  assign n38582 = n38577 & n38581 ;
  assign n38574 = n25878 & ~n35781 ;
  assign n38583 = n38582 ^ n38574 ^ n4488 ;
  assign n38584 = n22190 ^ n11600 ^ 1'b0 ;
  assign n38585 = ~n7332 & n38584 ;
  assign n38586 = ( n15940 & ~n29644 ) | ( n15940 & n38585 ) | ( ~n29644 & n38585 ) ;
  assign n38587 = ( n20688 & ~n24924 ) | ( n20688 & n38586 ) | ( ~n24924 & n38586 ) ;
  assign n38588 = ( n406 & n2183 ) | ( n406 & n31254 ) | ( n2183 & n31254 ) ;
  assign n38589 = n38588 ^ n16722 ^ n4795 ;
  assign n38590 = ( n7048 & n9704 ) | ( n7048 & n38589 ) | ( n9704 & n38589 ) ;
  assign n38591 = n23480 ^ n19487 ^ n16742 ;
  assign n38592 = n38591 ^ n25146 ^ n16822 ;
  assign n38593 = n1722 & ~n32971 ;
  assign n38594 = n38593 ^ n14565 ^ 1'b0 ;
  assign n38595 = n38594 ^ n14920 ^ n10420 ;
  assign n38596 = ~n36730 & n38595 ;
  assign n38597 = ~n11827 & n18116 ;
  assign n38598 = n38597 ^ n13521 ^ 1'b0 ;
  assign n38599 = ( n1990 & n15344 ) | ( n1990 & n38598 ) | ( n15344 & n38598 ) ;
  assign n38600 = ( ~n22163 & n35669 ) | ( ~n22163 & n36771 ) | ( n35669 & n36771 ) ;
  assign n38601 = ( ~n6128 & n38599 ) | ( ~n6128 & n38600 ) | ( n38599 & n38600 ) ;
  assign n38602 = n8357 ^ n1575 ^ 1'b0 ;
  assign n38603 = ~n22207 & n38602 ;
  assign n38604 = n2370 | n4653 ;
  assign n38605 = n38604 ^ n20478 ^ 1'b0 ;
  assign n38606 = n6527 & ~n34296 ;
  assign n38607 = n38606 ^ n1502 ^ 1'b0 ;
  assign n38608 = n32069 ^ n17640 ^ n13647 ;
  assign n38609 = n38608 ^ n28981 ^ n26750 ;
  assign n38610 = n17534 ^ n7415 ^ 1'b0 ;
  assign n38611 = n38610 ^ n19189 ^ n17411 ;
  assign n38612 = n13647 ^ n6756 ^ 1'b0 ;
  assign n38613 = n1983 & n38612 ;
  assign n38614 = ( n31803 & n38611 ) | ( n31803 & ~n38613 ) | ( n38611 & ~n38613 ) ;
  assign n38615 = n30333 ^ n25045 ^ n8653 ;
  assign n38616 = n20815 ^ n11566 ^ n7790 ;
  assign n38617 = n36093 ^ n32774 ^ 1'b0 ;
  assign n38618 = n38616 & n38617 ;
  assign n38619 = n6849 & n16520 ;
  assign n38620 = n38619 ^ n13411 ^ n5271 ;
  assign n38621 = n38620 ^ n2046 ^ x205 ;
  assign n38622 = n32381 ^ n28251 ^ n7930 ;
  assign n38623 = n12037 ^ n8156 ^ 1'b0 ;
  assign n38624 = ( n4058 & n8064 ) | ( n4058 & n11487 ) | ( n8064 & n11487 ) ;
  assign n38625 = ( ~n769 & n5584 ) | ( ~n769 & n9565 ) | ( n5584 & n9565 ) ;
  assign n38626 = ( n3816 & n38624 ) | ( n3816 & ~n38625 ) | ( n38624 & ~n38625 ) ;
  assign n38627 = ~n445 & n38626 ;
  assign n38628 = n18293 ^ n17422 ^ 1'b0 ;
  assign n38629 = n31145 ^ n17110 ^ n9575 ;
  assign n38632 = n3250 & n25607 ;
  assign n38633 = n38632 ^ n18270 ^ 1'b0 ;
  assign n38630 = n30353 ^ n5120 ^ 1'b0 ;
  assign n38631 = n30170 & ~n38630 ;
  assign n38634 = n38633 ^ n38631 ^ n2775 ;
  assign n38635 = ( n38628 & ~n38629 ) | ( n38628 & n38634 ) | ( ~n38629 & n38634 ) ;
  assign n38637 = ( n7045 & n20439 ) | ( n7045 & ~n31487 ) | ( n20439 & ~n31487 ) ;
  assign n38636 = n6594 ^ n4830 ^ 1'b0 ;
  assign n38638 = n38637 ^ n38636 ^ 1'b0 ;
  assign n38639 = n36617 & n38638 ;
  assign n38640 = ( n9196 & ~n28890 ) | ( n9196 & n31222 ) | ( ~n28890 & n31222 ) ;
  assign n38641 = ( n7612 & ~n21837 ) | ( n7612 & n22454 ) | ( ~n21837 & n22454 ) ;
  assign n38642 = n25358 ^ n24849 ^ n6972 ;
  assign n38643 = n20640 ^ n20248 ^ n1075 ;
  assign n38644 = ( n14216 & n38642 ) | ( n14216 & n38643 ) | ( n38642 & n38643 ) ;
  assign n38645 = ( ~n7248 & n7584 ) | ( ~n7248 & n20241 ) | ( n7584 & n20241 ) ;
  assign n38646 = n2310 & ~n35642 ;
  assign n38647 = ( n4071 & n8277 ) | ( n4071 & ~n38646 ) | ( n8277 & ~n38646 ) ;
  assign n38648 = n38647 ^ n26340 ^ 1'b0 ;
  assign n38649 = n35933 | n38648 ;
  assign n38650 = ( n11854 & n26908 ) | ( n11854 & ~n35541 ) | ( n26908 & ~n35541 ) ;
  assign n38651 = n38650 ^ n1759 ^ 1'b0 ;
  assign n38652 = n15503 | n24242 ;
  assign n38653 = n38652 ^ n24285 ^ 1'b0 ;
  assign n38654 = n38653 ^ n37575 ^ n33950 ;
  assign n38655 = ( ~n10732 & n14129 ) | ( ~n10732 & n14921 ) | ( n14129 & n14921 ) ;
  assign n38656 = ( n18808 & n36942 ) | ( n18808 & n38655 ) | ( n36942 & n38655 ) ;
  assign n38657 = n38656 ^ n23004 ^ n1956 ;
  assign n38659 = n31915 ^ n23669 ^ 1'b0 ;
  assign n38660 = n38659 ^ n22011 ^ n1744 ;
  assign n38661 = ( n4638 & ~n12580 ) | ( n4638 & n38660 ) | ( ~n12580 & n38660 ) ;
  assign n38658 = n34400 ^ n28033 ^ n2857 ;
  assign n38662 = n38661 ^ n38658 ^ 1'b0 ;
  assign n38663 = n38662 ^ n16984 ^ n14077 ;
  assign n38664 = n21824 & ~n33592 ;
  assign n38665 = n38664 ^ n3696 ^ 1'b0 ;
  assign n38670 = ~n15926 & n18187 ;
  assign n38666 = ( n3048 & n8183 ) | ( n3048 & n15275 ) | ( n8183 & n15275 ) ;
  assign n38667 = n36284 ^ n11248 ^ n7242 ;
  assign n38668 = ~n35898 & n38667 ;
  assign n38669 = n38666 & n38668 ;
  assign n38671 = n38670 ^ n38669 ^ n6656 ;
  assign n38672 = n38671 ^ n16322 ^ n6635 ;
  assign n38673 = n16528 ^ n8630 ^ n311 ;
  assign n38674 = ( n20679 & n27999 ) | ( n20679 & n31734 ) | ( n27999 & n31734 ) ;
  assign n38675 = n38674 ^ n27283 ^ n12627 ;
  assign n38676 = ( ~n18636 & n38673 ) | ( ~n18636 & n38675 ) | ( n38673 & n38675 ) ;
  assign n38677 = ( n38665 & n38672 ) | ( n38665 & ~n38676 ) | ( n38672 & ~n38676 ) ;
  assign n38678 = ~n3024 & n8012 ;
  assign n38679 = n38678 ^ n16016 ^ n9618 ;
  assign n38680 = ( n2695 & ~n3479 ) | ( n2695 & n4094 ) | ( ~n3479 & n4094 ) ;
  assign n38689 = n3121 & n33881 ;
  assign n38690 = n11617 & n38689 ;
  assign n38684 = n22416 ^ n15764 ^ n12455 ;
  assign n38685 = n38684 ^ n31664 ^ n16086 ;
  assign n38682 = n34499 ^ n27807 ^ n6578 ;
  assign n38683 = n38682 ^ n25205 ^ n22953 ;
  assign n38686 = n38685 ^ n38683 ^ n25937 ;
  assign n38687 = ( n9073 & ~n35668 ) | ( n9073 & n38686 ) | ( ~n35668 & n38686 ) ;
  assign n38688 = n38687 ^ n29853 ^ n23342 ;
  assign n38681 = n22509 ^ n17424 ^ n15159 ;
  assign n38691 = n38690 ^ n38688 ^ n38681 ;
  assign n38692 = n34296 ^ n25920 ^ n19076 ;
  assign n38693 = ( n24184 & n30638 ) | ( n24184 & ~n38692 ) | ( n30638 & ~n38692 ) ;
  assign n38694 = n38693 ^ n17530 ^ n9380 ;
  assign n38695 = n28103 ^ n26411 ^ n17493 ;
  assign n38696 = n38695 ^ n29334 ^ n14150 ;
  assign n38697 = ( n685 & n4082 ) | ( n685 & n11013 ) | ( n4082 & n11013 ) ;
  assign n38698 = n30627 ^ n28180 ^ n11130 ;
  assign n38699 = ( ~n13065 & n38697 ) | ( ~n13065 & n38698 ) | ( n38697 & n38698 ) ;
  assign n38700 = ( ~n9758 & n11479 ) | ( ~n9758 & n14008 ) | ( n11479 & n14008 ) ;
  assign n38701 = n31248 ^ n28955 ^ n13986 ;
  assign n38702 = n21526 ^ n9813 ^ 1'b0 ;
  assign n38703 = ( n38700 & n38701 ) | ( n38700 & n38702 ) | ( n38701 & n38702 ) ;
  assign n38704 = n20093 | n25236 ;
  assign n38705 = n38704 ^ n15125 ^ 1'b0 ;
  assign n38706 = n9472 ^ n2982 ^ n2819 ;
  assign n38707 = n25823 ^ n13894 ^ n13557 ;
  assign n38708 = n11919 ^ n8567 ^ n6403 ;
  assign n38709 = ( n14778 & ~n18546 ) | ( n14778 & n38708 ) | ( ~n18546 & n38708 ) ;
  assign n38710 = n38709 ^ n14700 ^ n273 ;
  assign n38711 = n27704 | n38710 ;
  assign n38712 = ( ~n6345 & n22680 ) | ( ~n6345 & n34939 ) | ( n22680 & n34939 ) ;
  assign n38713 = ( ~n1054 & n6183 ) | ( ~n1054 & n21698 ) | ( n6183 & n21698 ) ;
  assign n38714 = ( ~n5703 & n25381 ) | ( ~n5703 & n38713 ) | ( n25381 & n38713 ) ;
  assign n38715 = n6689 & n38714 ;
  assign n38716 = n38715 ^ n11384 ^ 1'b0 ;
  assign n38717 = n19054 ^ n16704 ^ x190 ;
  assign n38718 = n2756 | n38717 ;
  assign n38719 = n8239 & ~n38718 ;
  assign n38720 = ~n1000 & n9758 ;
  assign n38721 = n38720 ^ n27506 ^ n8223 ;
  assign n38722 = ( n6985 & n9185 ) | ( n6985 & ~n36942 ) | ( n9185 & ~n36942 ) ;
  assign n38723 = ( ~n8024 & n23807 ) | ( ~n8024 & n38722 ) | ( n23807 & n38722 ) ;
  assign n38724 = n38723 ^ n36367 ^ n32637 ;
  assign n38725 = ( n10185 & n22630 ) | ( n10185 & n35315 ) | ( n22630 & n35315 ) ;
  assign n38726 = n38725 ^ n16814 ^ n4922 ;
  assign n38727 = n12245 ^ n7021 ^ n5255 ;
  assign n38728 = n22865 ^ n18609 ^ 1'b0 ;
  assign n38729 = n3194 | n38728 ;
  assign n38730 = ( ~n12150 & n23767 ) | ( ~n12150 & n38729 ) | ( n23767 & n38729 ) ;
  assign n38731 = n9934 ^ n7363 ^ n6144 ;
  assign n38733 = n15819 ^ n13276 ^ n9107 ;
  assign n38732 = ( n8291 & ~n14895 ) | ( n8291 & n31918 ) | ( ~n14895 & n31918 ) ;
  assign n38734 = n38733 ^ n38732 ^ n6958 ;
  assign n38735 = ( n4102 & ~n12921 ) | ( n4102 & n17128 ) | ( ~n12921 & n17128 ) ;
  assign n38736 = n32808 ^ n7615 ^ n1491 ;
  assign n38737 = ( ~n31053 & n38735 ) | ( ~n31053 & n38736 ) | ( n38735 & n38736 ) ;
  assign n38738 = ( n859 & ~n24746 ) | ( n859 & n38737 ) | ( ~n24746 & n38737 ) ;
  assign n38740 = n37857 ^ n19916 ^ n17299 ;
  assign n38741 = ~n8972 & n38740 ;
  assign n38742 = n38741 ^ n4208 ^ 1'b0 ;
  assign n38743 = n38742 ^ n34712 ^ n14515 ;
  assign n38739 = ( n462 & ~n13843 ) | ( n462 & n22186 ) | ( ~n13843 & n22186 ) ;
  assign n38744 = n38743 ^ n38739 ^ n6309 ;
  assign n38745 = n3032 & n5827 ;
  assign n38746 = n38745 ^ n36579 ^ 1'b0 ;
  assign n38747 = n6398 ^ x135 ^ 1'b0 ;
  assign n38748 = n2838 | n38747 ;
  assign n38749 = ~n1367 & n3898 ;
  assign n38750 = n38749 ^ n16291 ^ 1'b0 ;
  assign n38751 = ( n31434 & n38748 ) | ( n31434 & n38750 ) | ( n38748 & n38750 ) ;
  assign n38752 = ( n12736 & ~n38746 ) | ( n12736 & n38751 ) | ( ~n38746 & n38751 ) ;
  assign n38754 = n1341 & n19365 ;
  assign n38753 = ( n9682 & ~n9845 ) | ( n9682 & n22831 ) | ( ~n9845 & n22831 ) ;
  assign n38755 = n38754 ^ n38753 ^ n3957 ;
  assign n38756 = ( n10979 & n14817 ) | ( n10979 & n27915 ) | ( n14817 & n27915 ) ;
  assign n38757 = n17532 ^ n15133 ^ 1'b0 ;
  assign n38758 = n38756 | n38757 ;
  assign n38759 = n38758 ^ n33682 ^ n521 ;
  assign n38760 = ( n3595 & ~n4835 ) | ( n3595 & n31840 ) | ( ~n4835 & n31840 ) ;
  assign n38761 = ( n5876 & n30895 ) | ( n5876 & n38760 ) | ( n30895 & n38760 ) ;
  assign n38764 = n9316 ^ n4495 ^ n294 ;
  assign n38765 = ( n26382 & ~n33955 ) | ( n26382 & n38764 ) | ( ~n33955 & n38764 ) ;
  assign n38762 = ( ~n7094 & n10168 ) | ( ~n7094 & n15357 ) | ( n10168 & n15357 ) ;
  assign n38763 = n38762 ^ n2685 ^ 1'b0 ;
  assign n38766 = n38765 ^ n38763 ^ 1'b0 ;
  assign n38771 = n9092 | n19119 ;
  assign n38770 = n24035 ^ n18326 ^ n11726 ;
  assign n38767 = n5060 ^ n627 ^ 1'b0 ;
  assign n38768 = n38767 ^ n27196 ^ n4435 ;
  assign n38769 = ~n19691 & n38768 ;
  assign n38772 = n38771 ^ n38770 ^ n38769 ;
  assign n38773 = ~n6902 & n28978 ;
  assign n38774 = n38773 ^ n4602 ^ 1'b0 ;
  assign n38779 = n21674 ^ n8298 ^ 1'b0 ;
  assign n38780 = n12290 | n38779 ;
  assign n38778 = n30892 ^ n7907 ^ n5303 ;
  assign n38775 = n20023 & ~n37650 ;
  assign n38776 = n38775 ^ n32475 ^ 1'b0 ;
  assign n38777 = ( n7459 & ~n12179 ) | ( n7459 & n38776 ) | ( ~n12179 & n38776 ) ;
  assign n38781 = n38780 ^ n38778 ^ n38777 ;
  assign n38782 = n9713 ^ n6318 ^ 1'b0 ;
  assign n38783 = n6654 & ~n38782 ;
  assign n38784 = n38783 ^ n29595 ^ n10900 ;
  assign n38785 = ( n21214 & n38750 ) | ( n21214 & n38784 ) | ( n38750 & n38784 ) ;
  assign n38786 = n36296 ^ n4344 ^ 1'b0 ;
  assign n38787 = n18066 & n38786 ;
  assign n38788 = ( ~n19858 & n33360 ) | ( ~n19858 & n38787 ) | ( n33360 & n38787 ) ;
  assign n38789 = ( n10491 & n12682 ) | ( n10491 & ~n38788 ) | ( n12682 & ~n38788 ) ;
  assign n38790 = n38789 ^ n13395 ^ n9848 ;
  assign n38791 = n15864 ^ n9704 ^ n5422 ;
  assign n38792 = ( n14979 & ~n31923 ) | ( n14979 & n31965 ) | ( ~n31923 & n31965 ) ;
  assign n38793 = n2062 & n3898 ;
  assign n38794 = n18090 & n38793 ;
  assign n38795 = n13292 ^ n6517 ^ n2995 ;
  assign n38796 = n38795 ^ n26160 ^ n7239 ;
  assign n38797 = ( ~n9425 & n34151 ) | ( ~n9425 & n38796 ) | ( n34151 & n38796 ) ;
  assign n38798 = n17415 ^ n16164 ^ n9888 ;
  assign n38799 = ( n389 & ~n2274 ) | ( n389 & n5599 ) | ( ~n2274 & n5599 ) ;
  assign n38800 = ( n15510 & n38563 ) | ( n15510 & ~n38799 ) | ( n38563 & ~n38799 ) ;
  assign n38801 = ( n13067 & ~n38798 ) | ( n13067 & n38800 ) | ( ~n38798 & n38800 ) ;
  assign n38802 = n30076 ^ n8268 ^ n471 ;
  assign n38803 = n36835 ^ n28584 ^ n12251 ;
  assign n38805 = n11389 ^ n5215 ^ n1514 ;
  assign n38806 = ( ~n5501 & n22548 ) | ( ~n5501 & n38805 ) | ( n22548 & n38805 ) ;
  assign n38807 = n38806 ^ n13328 ^ n5109 ;
  assign n38804 = n19722 ^ n7969 ^ n7273 ;
  assign n38808 = n38807 ^ n38804 ^ n17150 ;
  assign n38809 = n32741 ^ n25006 ^ n19786 ;
  assign n38810 = ( n6685 & n9044 ) | ( n6685 & ~n38809 ) | ( n9044 & ~n38809 ) ;
  assign n38811 = ( n26669 & n33694 ) | ( n26669 & ~n38810 ) | ( n33694 & ~n38810 ) ;
  assign n38812 = ( n22010 & n38808 ) | ( n22010 & ~n38811 ) | ( n38808 & ~n38811 ) ;
  assign n38813 = n24117 ^ n5909 ^ 1'b0 ;
  assign n38814 = n3291 & ~n12122 ;
  assign n38815 = n38814 ^ n29011 ^ 1'b0 ;
  assign n38816 = ( n1518 & n3272 ) | ( n1518 & ~n7464 ) | ( n3272 & ~n7464 ) ;
  assign n38817 = ( n9609 & n12591 ) | ( n9609 & ~n38816 ) | ( n12591 & ~n38816 ) ;
  assign n38821 = n3685 & n5948 ;
  assign n38822 = n38821 ^ n3259 ^ 1'b0 ;
  assign n38818 = n15728 ^ n1513 ^ 1'b0 ;
  assign n38819 = n18306 | n38818 ;
  assign n38820 = n5452 | n38819 ;
  assign n38823 = n38822 ^ n38820 ^ 1'b0 ;
  assign n38824 = ( n10690 & ~n38817 ) | ( n10690 & n38823 ) | ( ~n38817 & n38823 ) ;
  assign n38825 = ( ~n27347 & n29561 ) | ( ~n27347 & n38824 ) | ( n29561 & n38824 ) ;
  assign n38826 = ( n2686 & n10173 ) | ( n2686 & ~n12318 ) | ( n10173 & ~n12318 ) ;
  assign n38827 = n21007 & ~n38826 ;
  assign n38828 = n38827 ^ n27466 ^ n433 ;
  assign n38829 = n36480 ^ n14001 ^ n5778 ;
  assign n38830 = ( ~n10999 & n28363 ) | ( ~n10999 & n38829 ) | ( n28363 & n38829 ) ;
  assign n38839 = ( ~n3502 & n19084 ) | ( ~n3502 & n36334 ) | ( n19084 & n36334 ) ;
  assign n38832 = n6250 & n16876 ;
  assign n38833 = n38832 ^ n5014 ^ 1'b0 ;
  assign n38834 = ~n7316 & n12098 ;
  assign n38835 = n38833 & n38834 ;
  assign n38831 = n23924 ^ n1498 ^ n829 ;
  assign n38836 = n38835 ^ n38831 ^ n13053 ;
  assign n38837 = n38148 ^ n31728 ^ n31020 ;
  assign n38838 = n38836 & ~n38837 ;
  assign n38840 = n38839 ^ n38838 ^ n14828 ;
  assign n38841 = ~n14245 & n15310 ;
  assign n38842 = ( x159 & ~n22413 ) | ( x159 & n38841 ) | ( ~n22413 & n38841 ) ;
  assign n38843 = ~n11512 & n38842 ;
  assign n38844 = ( n11282 & n17334 ) | ( n11282 & ~n24904 ) | ( n17334 & ~n24904 ) ;
  assign n38845 = ( ~n10513 & n10661 ) | ( ~n10513 & n38844 ) | ( n10661 & n38844 ) ;
  assign n38846 = ( ~n6641 & n14726 ) | ( ~n6641 & n26288 ) | ( n14726 & n26288 ) ;
  assign n38847 = ( ~n13119 & n20894 ) | ( ~n13119 & n38846 ) | ( n20894 & n38846 ) ;
  assign n38848 = n38847 ^ n13298 ^ n6536 ;
  assign n38849 = n31664 ^ n25192 ^ n23547 ;
  assign n38850 = n28367 ^ n22555 ^ x81 ;
  assign n38851 = n19540 ^ n12161 ^ n5414 ;
  assign n38852 = n25202 ^ n13220 ^ n3718 ;
  assign n38853 = n38852 ^ n3448 ^ n1996 ;
  assign n38854 = n10116 & ~n38853 ;
  assign n38855 = ( n18822 & ~n19358 ) | ( n18822 & n38854 ) | ( ~n19358 & n38854 ) ;
  assign n38856 = ~n7152 & n35221 ;
  assign n38857 = n38856 ^ n19729 ^ 1'b0 ;
  assign n38858 = n29213 ^ n26961 ^ n1607 ;
  assign n38859 = n38858 ^ n11456 ^ n7110 ;
  assign n38860 = ( n6154 & n8119 ) | ( n6154 & ~n38859 ) | ( n8119 & ~n38859 ) ;
  assign n38862 = n21313 ^ n20040 ^ n11936 ;
  assign n38861 = ( n5665 & ~n10002 ) | ( n5665 & n13983 ) | ( ~n10002 & n13983 ) ;
  assign n38863 = n38862 ^ n38861 ^ n22074 ;
  assign n38864 = n38863 ^ n3833 ^ 1'b0 ;
  assign n38865 = n38860 | n38864 ;
  assign n38866 = ( ~n19610 & n32070 ) | ( ~n19610 & n38047 ) | ( n32070 & n38047 ) ;
  assign n38867 = ( ~n12597 & n28083 ) | ( ~n12597 & n29568 ) | ( n28083 & n29568 ) ;
  assign n38868 = n22564 ^ n19504 ^ n13239 ;
  assign n38869 = ( n2732 & n9397 ) | ( n2732 & n20640 ) | ( n9397 & n20640 ) ;
  assign n38870 = n38869 ^ n15092 ^ 1'b0 ;
  assign n38871 = n11657 & n38870 ;
  assign n38872 = n38871 ^ n18774 ^ n6255 ;
  assign n38873 = n38872 ^ n27358 ^ n6414 ;
  assign n38874 = n38868 & ~n38873 ;
  assign n38875 = n38874 ^ n26709 ^ 1'b0 ;
  assign n38876 = n18460 ^ n5097 ^ 1'b0 ;
  assign n38877 = ( n6799 & n22512 ) | ( n6799 & ~n38876 ) | ( n22512 & ~n38876 ) ;
  assign n38878 = n28409 ^ n28367 ^ n5844 ;
  assign n38879 = n4100 | n25301 ;
  assign n38881 = ( n956 & ~n7071 ) | ( n956 & n35958 ) | ( ~n7071 & n35958 ) ;
  assign n38880 = n12365 | n34157 ;
  assign n38882 = n38881 ^ n38880 ^ 1'b0 ;
  assign n38883 = n38882 ^ n29858 ^ n19593 ;
  assign n38884 = ( n2421 & ~n13884 ) | ( n2421 & n15058 ) | ( ~n13884 & n15058 ) ;
  assign n38885 = ( n1948 & n32170 ) | ( n1948 & ~n35778 ) | ( n32170 & ~n35778 ) ;
  assign n38886 = n38885 ^ n38196 ^ n6744 ;
  assign n38887 = n15145 ^ n14137 ^ n6972 ;
  assign n38888 = ( n11264 & n14051 ) | ( n11264 & ~n38887 ) | ( n14051 & ~n38887 ) ;
  assign n38889 = n7288 | n9008 ;
  assign n38890 = n6428 | n38889 ;
  assign n38892 = ~n26952 & n30015 ;
  assign n38891 = ( n2459 & ~n11721 ) | ( n2459 & n21978 ) | ( ~n11721 & n21978 ) ;
  assign n38893 = n38892 ^ n38891 ^ n21585 ;
  assign n38894 = n10697 ^ n2886 ^ n657 ;
  assign n38895 = ( n4504 & n33663 ) | ( n4504 & n38894 ) | ( n33663 & n38894 ) ;
  assign n38896 = n20288 ^ n12929 ^ n11817 ;
  assign n38898 = ( n5344 & ~n8951 ) | ( n5344 & n9741 ) | ( ~n8951 & n9741 ) ;
  assign n38897 = ( ~n10783 & n23604 ) | ( ~n10783 & n27093 ) | ( n23604 & n27093 ) ;
  assign n38899 = n38898 ^ n38897 ^ n15308 ;
  assign n38900 = ( ~n3809 & n9098 ) | ( ~n3809 & n15201 ) | ( n9098 & n15201 ) ;
  assign n38901 = n38900 ^ n30400 ^ 1'b0 ;
  assign n38902 = n8619 ^ n5519 ^ n2029 ;
  assign n38903 = n38902 ^ n3184 ^ 1'b0 ;
  assign n38904 = n38903 ^ n24751 ^ 1'b0 ;
  assign n38905 = n20075 & n38904 ;
  assign n38906 = ( ~n5759 & n9865 ) | ( ~n5759 & n13055 ) | ( n9865 & n13055 ) ;
  assign n38907 = ( n7338 & n33892 ) | ( n7338 & n38906 ) | ( n33892 & n38906 ) ;
  assign n38908 = n36331 ^ n24830 ^ n20059 ;
  assign n38909 = ( n11716 & n17644 ) | ( n11716 & n30013 ) | ( n17644 & n30013 ) ;
  assign n38910 = ( n5906 & n8926 ) | ( n5906 & ~n10861 ) | ( n8926 & ~n10861 ) ;
  assign n38911 = n38910 ^ n37416 ^ n583 ;
  assign n38912 = ( n21501 & n38909 ) | ( n21501 & ~n38911 ) | ( n38909 & ~n38911 ) ;
  assign n38913 = ( ~n31658 & n38908 ) | ( ~n31658 & n38912 ) | ( n38908 & n38912 ) ;
  assign n38918 = ( ~n4287 & n6546 ) | ( ~n4287 & n19375 ) | ( n6546 & n19375 ) ;
  assign n38919 = ~n37585 & n38918 ;
  assign n38920 = ~n10885 & n38919 ;
  assign n38916 = n8105 & n11144 ;
  assign n38917 = ( ~n918 & n31481 ) | ( ~n918 & n38916 ) | ( n31481 & n38916 ) ;
  assign n38914 = ~n3686 & n18909 ;
  assign n38915 = n38914 ^ n32678 ^ 1'b0 ;
  assign n38921 = n38920 ^ n38917 ^ n38915 ;
  assign n38923 = n23080 ^ n7087 ^ n2470 ;
  assign n38922 = n12951 & n14813 ;
  assign n38924 = n38923 ^ n38922 ^ n3560 ;
  assign n38925 = ( n3998 & n21474 ) | ( n3998 & n38329 ) | ( n21474 & n38329 ) ;
  assign n38926 = n13253 ^ n7312 ^ n2259 ;
  assign n38927 = n34536 | n35775 ;
  assign n38928 = ( n38925 & n38926 ) | ( n38925 & ~n38927 ) | ( n38926 & ~n38927 ) ;
  assign n38929 = n8553 & n35356 ;
  assign n38930 = n38929 ^ n13856 ^ n5564 ;
  assign n38931 = ( n2784 & ~n9267 ) | ( n2784 & n38930 ) | ( ~n9267 & n38930 ) ;
  assign n38932 = ( ~n14859 & n16066 ) | ( ~n14859 & n24958 ) | ( n16066 & n24958 ) ;
  assign n38933 = n38932 ^ n26767 ^ n3277 ;
  assign n38934 = ( n26270 & n34858 ) | ( n26270 & ~n38417 ) | ( n34858 & ~n38417 ) ;
  assign n38935 = ( ~n5576 & n7674 ) | ( ~n5576 & n38934 ) | ( n7674 & n38934 ) ;
  assign n38936 = n38933 | n38935 ;
  assign n38937 = n6168 | n38936 ;
  assign n38938 = ( n10892 & n16876 ) | ( n10892 & ~n17734 ) | ( n16876 & ~n17734 ) ;
  assign n38939 = n23243 ^ n19284 ^ n15243 ;
  assign n38940 = n38939 ^ n27263 ^ n26602 ;
  assign n38941 = n22431 ^ n9176 ^ n3066 ;
  assign n38942 = ( n343 & n10657 ) | ( n343 & n38941 ) | ( n10657 & n38941 ) ;
  assign n38943 = ( n1624 & n10988 ) | ( n1624 & n38942 ) | ( n10988 & n38942 ) ;
  assign n38944 = n38735 ^ n34191 ^ 1'b0 ;
  assign n38945 = n10218 | n38944 ;
  assign n38946 = ~n2113 & n38945 ;
  assign n38947 = n29414 ^ n27183 ^ n20810 ;
  assign n38948 = ( n17233 & n38946 ) | ( n17233 & ~n38947 ) | ( n38946 & ~n38947 ) ;
  assign n38949 = ( n21653 & n38943 ) | ( n21653 & ~n38948 ) | ( n38943 & ~n38948 ) ;
  assign n38950 = n38949 ^ n27914 ^ n762 ;
  assign n38951 = n38950 ^ n16037 ^ n1982 ;
  assign n38952 = ( n7631 & n10933 ) | ( n7631 & n22394 ) | ( n10933 & n22394 ) ;
  assign n38953 = ( n13863 & ~n25670 ) | ( n13863 & n38952 ) | ( ~n25670 & n38952 ) ;
  assign n38954 = ( ~n5019 & n5683 ) | ( ~n5019 & n11017 ) | ( n5683 & n11017 ) ;
  assign n38955 = n26118 ^ n25517 ^ 1'b0 ;
  assign n38956 = ~n21575 & n38955 ;
  assign n38957 = n38956 ^ n24280 ^ n11119 ;
  assign n38958 = ( n3689 & ~n7275 ) | ( n3689 & n33777 ) | ( ~n7275 & n33777 ) ;
  assign n38959 = ( n1082 & n8732 ) | ( n1082 & ~n38958 ) | ( n8732 & ~n38958 ) ;
  assign n38961 = ( n12296 & ~n21790 ) | ( n12296 & n31149 ) | ( ~n21790 & n31149 ) ;
  assign n38960 = n13063 | n14300 ;
  assign n38962 = n38961 ^ n38960 ^ 1'b0 ;
  assign n38963 = n38962 ^ n32093 ^ n25839 ;
  assign n38964 = n12839 & n37945 ;
  assign n38965 = n7257 & ~n20849 ;
  assign n38966 = n38965 ^ n34200 ^ 1'b0 ;
  assign n38967 = ( n17147 & ~n25630 ) | ( n17147 & n26247 ) | ( ~n25630 & n26247 ) ;
  assign n38968 = n10521 ^ n3915 ^ n2570 ;
  assign n38969 = n38968 ^ n37300 ^ n1521 ;
  assign n38970 = ( n3632 & n24814 ) | ( n3632 & ~n38969 ) | ( n24814 & ~n38969 ) ;
  assign n38971 = ( n37462 & n38967 ) | ( n37462 & n38970 ) | ( n38967 & n38970 ) ;
  assign n38972 = n25360 ^ n25173 ^ n14590 ;
  assign n38973 = n38972 ^ n21740 ^ n17471 ;
  assign n38974 = ( x85 & n2114 ) | ( x85 & n5209 ) | ( n2114 & n5209 ) ;
  assign n38975 = ( ~n4303 & n8857 ) | ( ~n4303 & n38974 ) | ( n8857 & n38974 ) ;
  assign n38976 = ( n4324 & n8558 ) | ( n4324 & ~n38975 ) | ( n8558 & ~n38975 ) ;
  assign n38977 = n17113 ^ n1117 ^ 1'b0 ;
  assign n38978 = n38976 & ~n38977 ;
  assign n38979 = ( ~n17402 & n18645 ) | ( ~n17402 & n38978 ) | ( n18645 & n38978 ) ;
  assign n38980 = n10121 | n22125 ;
  assign n38981 = n38980 ^ n37894 ^ 1'b0 ;
  assign n38982 = n38981 ^ n23249 ^ n13563 ;
  assign n38983 = n24565 | n31312 ;
  assign n38984 = n10649 | n38983 ;
  assign n38985 = n38984 ^ n14566 ^ 1'b0 ;
  assign n38986 = ( n894 & n2217 ) | ( n894 & n8186 ) | ( n2217 & n8186 ) ;
  assign n38987 = ( n2036 & n14065 ) | ( n2036 & n17486 ) | ( n14065 & n17486 ) ;
  assign n38988 = n38987 ^ n28251 ^ n10277 ;
  assign n38989 = n21608 ^ n12922 ^ n9339 ;
  assign n38990 = n12549 & ~n38989 ;
  assign n38991 = n38990 ^ n7546 ^ 1'b0 ;
  assign n38992 = ( n38986 & n38988 ) | ( n38986 & ~n38991 ) | ( n38988 & ~n38991 ) ;
  assign n38993 = n10490 ^ n1850 ^ 1'b0 ;
  assign n38994 = n14274 | n38993 ;
  assign n38995 = ( ~n416 & n9841 ) | ( ~n416 & n38994 ) | ( n9841 & n38994 ) ;
  assign n38996 = ( n5045 & n16436 ) | ( n5045 & ~n17247 ) | ( n16436 & ~n17247 ) ;
  assign n38997 = n38996 ^ n30730 ^ n29449 ;
  assign n38998 = ( ~n8259 & n38262 ) | ( ~n8259 & n38997 ) | ( n38262 & n38997 ) ;
  assign n38999 = n26345 ^ n26106 ^ 1'b0 ;
  assign n39000 = n25063 | n35330 ;
  assign n39001 = n18904 ^ n13900 ^ n9617 ;
  assign n39002 = ~n7875 & n9197 ;
  assign n39003 = n39002 ^ n24791 ^ 1'b0 ;
  assign n39011 = n11159 & n22847 ;
  assign n39012 = ~n19991 & n39011 ;
  assign n39004 = n24145 ^ n23283 ^ n9829 ;
  assign n39005 = n39004 ^ n20257 ^ n3401 ;
  assign n39006 = ( ~n13770 & n15927 ) | ( ~n13770 & n23805 ) | ( n15927 & n23805 ) ;
  assign n39007 = n39006 ^ n33930 ^ n31176 ;
  assign n39008 = ( n23132 & n39005 ) | ( n23132 & n39007 ) | ( n39005 & n39007 ) ;
  assign n39009 = n26366 ^ n2538 ^ 1'b0 ;
  assign n39010 = n39008 | n39009 ;
  assign n39013 = n39012 ^ n39010 ^ n23254 ;
  assign n39014 = ( n39001 & ~n39003 ) | ( n39001 & n39013 ) | ( ~n39003 & n39013 ) ;
  assign n39015 = ~n364 & n675 ;
  assign n39016 = ( n7225 & ~n35474 ) | ( n7225 & n39015 ) | ( ~n35474 & n39015 ) ;
  assign n39017 = ( ~n14788 & n16991 ) | ( ~n14788 & n39016 ) | ( n16991 & n39016 ) ;
  assign n39018 = ( ~n20988 & n31856 ) | ( ~n20988 & n34330 ) | ( n31856 & n34330 ) ;
  assign n39019 = n14423 ^ n4752 ^ n3928 ;
  assign n39020 = ( n21470 & n26857 ) | ( n21470 & ~n39019 ) | ( n26857 & ~n39019 ) ;
  assign n39021 = n16019 ^ n496 ^ 1'b0 ;
  assign n39022 = n39021 ^ n13752 ^ n1863 ;
  assign n39023 = n39022 ^ n7149 ^ 1'b0 ;
  assign n39024 = n37732 ^ n22302 ^ 1'b0 ;
  assign n39025 = ( ~n1217 & n5891 ) | ( ~n1217 & n25638 ) | ( n5891 & n25638 ) ;
  assign n39026 = n34135 ^ n22985 ^ n17454 ;
  assign n39027 = ( n3910 & n7207 ) | ( n3910 & n32093 ) | ( n7207 & n32093 ) ;
  assign n39028 = n24006 ^ n9116 ^ n5803 ;
  assign n39029 = n26862 ^ n8418 ^ 1'b0 ;
  assign n39030 = n2897 & ~n39029 ;
  assign n39031 = ~n28755 & n39030 ;
  assign n39032 = n13287 & n39031 ;
  assign n39034 = n23855 ^ n10304 ^ n5301 ;
  assign n39033 = ( n9440 & ~n12176 ) | ( n9440 & n12525 ) | ( ~n12176 & n12525 ) ;
  assign n39035 = n39034 ^ n39033 ^ 1'b0 ;
  assign n39036 = n16830 & ~n33704 ;
  assign n39037 = ~n39035 & n39036 ;
  assign n39038 = n23080 | n38196 ;
  assign n39039 = ( n4355 & ~n39037 ) | ( n4355 & n39038 ) | ( ~n39037 & n39038 ) ;
  assign n39040 = ( n14251 & ~n21632 ) | ( n14251 & n35725 ) | ( ~n21632 & n35725 ) ;
  assign n39041 = n1937 & ~n10952 ;
  assign n39042 = ( ~n18879 & n39040 ) | ( ~n18879 & n39041 ) | ( n39040 & n39041 ) ;
  assign n39043 = n14891 ^ n10766 ^ n3860 ;
  assign n39044 = n8099 | n18196 ;
  assign n39045 = n39044 ^ n35814 ^ n10907 ;
  assign n39046 = n1008 & ~n21018 ;
  assign n39047 = ( n2492 & n21852 ) | ( n2492 & ~n39046 ) | ( n21852 & ~n39046 ) ;
  assign n39048 = n26840 ^ n14112 ^ n8804 ;
  assign n39049 = n665 & ~n39048 ;
  assign n39050 = n39049 ^ n26018 ^ n13424 ;
  assign n39051 = n25703 ^ n18271 ^ 1'b0 ;
  assign n39052 = n39051 ^ n29704 ^ n6270 ;
  assign n39053 = ( n15469 & n24804 ) | ( n15469 & n32265 ) | ( n24804 & n32265 ) ;
  assign n39056 = x121 & n21846 ;
  assign n39057 = n39056 ^ n1255 ^ 1'b0 ;
  assign n39058 = n39057 ^ n27165 ^ n3628 ;
  assign n39054 = n23121 ^ n3074 ^ n2336 ;
  assign n39055 = n39054 ^ n24415 ^ n21805 ;
  assign n39059 = n39058 ^ n39055 ^ n19140 ;
  assign n39060 = n19857 ^ n9531 ^ 1'b0 ;
  assign n39062 = n37165 ^ n19399 ^ n10946 ;
  assign n39063 = ( n16788 & ~n28882 ) | ( n16788 & n39062 ) | ( ~n28882 & n39062 ) ;
  assign n39061 = n13402 & ~n17316 ;
  assign n39064 = n39063 ^ n39061 ^ 1'b0 ;
  assign n39067 = n20737 ^ n19938 ^ x74 ;
  assign n39065 = ( n2790 & ~n15738 ) | ( n2790 & n25484 ) | ( ~n15738 & n25484 ) ;
  assign n39066 = n39065 ^ n18582 ^ n4238 ;
  assign n39068 = n39067 ^ n39066 ^ n11303 ;
  assign n39069 = n21219 ^ n15845 ^ n8047 ;
  assign n39070 = n39069 ^ n18245 ^ n8869 ;
  assign n39071 = n5995 ^ n2983 ^ n1808 ;
  assign n39072 = n39071 ^ n5066 ^ 1'b0 ;
  assign n39073 = n39072 ^ n18296 ^ n16805 ;
  assign n39074 = ( n33324 & n39070 ) | ( n33324 & ~n39073 ) | ( n39070 & ~n39073 ) ;
  assign n39075 = n37657 ^ n3245 ^ n1810 ;
  assign n39076 = n39075 ^ n32837 ^ n2473 ;
  assign n39077 = n39076 ^ n30316 ^ n22433 ;
  assign n39078 = n39077 ^ n21436 ^ n1541 ;
  assign n39083 = n13337 ^ n10878 ^ 1'b0 ;
  assign n39084 = ~n38767 & n39083 ;
  assign n39080 = n9018 | n34390 ;
  assign n39081 = n39080 ^ n25446 ^ 1'b0 ;
  assign n39082 = n39081 ^ n28832 ^ n14579 ;
  assign n39079 = ( n4076 & n14400 ) | ( n4076 & ~n38678 ) | ( n14400 & ~n38678 ) ;
  assign n39085 = n39084 ^ n39082 ^ n39079 ;
  assign n39086 = ( n2093 & ~n14189 ) | ( n2093 & n20217 ) | ( ~n14189 & n20217 ) ;
  assign n39087 = n39086 ^ n11323 ^ 1'b0 ;
  assign n39088 = n29838 ^ n16261 ^ n14452 ;
  assign n39089 = n39088 ^ n16696 ^ n7844 ;
  assign n39094 = n8141 ^ n5364 ^ 1'b0 ;
  assign n39095 = n13583 & n39094 ;
  assign n39096 = ~n10389 & n39095 ;
  assign n39090 = n4476 ^ n3514 ^ n1567 ;
  assign n39091 = n14450 & n39090 ;
  assign n39092 = n39091 ^ n37786 ^ 1'b0 ;
  assign n39093 = ( ~n22688 & n27612 ) | ( ~n22688 & n39092 ) | ( n27612 & n39092 ) ;
  assign n39097 = n39096 ^ n39093 ^ n38396 ;
  assign n39098 = n37298 ^ n34400 ^ n21973 ;
  assign n39099 = n39098 ^ n35343 ^ n29168 ;
  assign n39100 = n8288 ^ n5405 ^ n3836 ;
  assign n39101 = n12881 ^ n5765 ^ n3509 ;
  assign n39102 = n39096 ^ n23100 ^ n934 ;
  assign n39103 = ( n39100 & ~n39101 ) | ( n39100 & n39102 ) | ( ~n39101 & n39102 ) ;
  assign n39106 = n28176 ^ n27414 ^ n15262 ;
  assign n39104 = ( n2122 & n7314 ) | ( n2122 & ~n16105 ) | ( n7314 & ~n16105 ) ;
  assign n39105 = ( n3649 & n18974 ) | ( n3649 & ~n39104 ) | ( n18974 & ~n39104 ) ;
  assign n39107 = n39106 ^ n39105 ^ n7148 ;
  assign n39110 = n28367 ^ n10286 ^ 1'b0 ;
  assign n39111 = n8412 & n39110 ;
  assign n39108 = ( n17554 & n19519 ) | ( n17554 & ~n31101 ) | ( n19519 & ~n31101 ) ;
  assign n39109 = ( n10964 & n33849 ) | ( n10964 & ~n39108 ) | ( n33849 & ~n39108 ) ;
  assign n39112 = n39111 ^ n39109 ^ n29877 ;
  assign n39113 = n39112 ^ n32301 ^ n14659 ;
  assign n39116 = n25114 ^ n17736 ^ 1'b0 ;
  assign n39117 = n17889 | n39116 ;
  assign n39114 = n24506 ^ n16946 ^ n6926 ;
  assign n39115 = n5406 | n39114 ;
  assign n39118 = n39117 ^ n39115 ^ 1'b0 ;
  assign n39119 = ( ~n12384 & n16458 ) | ( ~n12384 & n23109 ) | ( n16458 & n23109 ) ;
  assign n39120 = n33368 ^ n4091 ^ n2731 ;
  assign n39121 = ( n1300 & n10080 ) | ( n1300 & n16050 ) | ( n10080 & n16050 ) ;
  assign n39122 = n39121 ^ n20598 ^ n18802 ;
  assign n39123 = n33146 ^ n6424 ^ n1496 ;
  assign n39124 = n2744 | n35751 ;
  assign n39125 = n39124 ^ n31357 ^ 1'b0 ;
  assign n39126 = ~n39123 & n39125 ;
  assign n39127 = ( n22426 & ~n25273 ) | ( n22426 & n39126 ) | ( ~n25273 & n39126 ) ;
  assign n39128 = ( n12117 & ~n35792 ) | ( n12117 & n39127 ) | ( ~n35792 & n39127 ) ;
  assign n39129 = ( x184 & n39122 ) | ( x184 & n39128 ) | ( n39122 & n39128 ) ;
  assign n39130 = ( n6484 & n22637 ) | ( n6484 & ~n26160 ) | ( n22637 & ~n26160 ) ;
  assign n39131 = ( ~n3832 & n26934 ) | ( ~n3832 & n39130 ) | ( n26934 & n39130 ) ;
  assign n39132 = ( n5264 & n7855 ) | ( n5264 & ~n39131 ) | ( n7855 & ~n39131 ) ;
  assign n39133 = n3553 | n13449 ;
  assign n39134 = n39133 ^ n28999 ^ n2055 ;
  assign n39135 = n38527 ^ n22238 ^ n4553 ;
  assign n39136 = ( n12049 & n32390 ) | ( n12049 & ~n34064 ) | ( n32390 & ~n34064 ) ;
  assign n39137 = ( ~n5115 & n14296 ) | ( ~n5115 & n24629 ) | ( n14296 & n24629 ) ;
  assign n39138 = n31163 ^ n6139 ^ n3838 ;
  assign n39139 = ( n23527 & n39137 ) | ( n23527 & ~n39138 ) | ( n39137 & ~n39138 ) ;
  assign n39140 = ( n5957 & ~n9630 ) | ( n5957 & n11600 ) | ( ~n9630 & n11600 ) ;
  assign n39141 = n34359 ^ n17267 ^ n1706 ;
  assign n39142 = n39141 ^ n32301 ^ n8728 ;
  assign n39143 = n26429 | n39142 ;
  assign n39144 = n22777 & ~n39143 ;
  assign n39145 = ( n19504 & n23219 ) | ( n19504 & ~n25477 ) | ( n23219 & ~n25477 ) ;
  assign n39146 = n29839 ^ n28910 ^ n21748 ;
  assign n39147 = ( ~n18501 & n20498 ) | ( ~n18501 & n39146 ) | ( n20498 & n39146 ) ;
  assign n39151 = ( ~n7127 & n13807 ) | ( ~n7127 & n36951 ) | ( n13807 & n36951 ) ;
  assign n39152 = n39151 ^ n26538 ^ n19231 ;
  assign n39153 = ( n1987 & n24178 ) | ( n1987 & n39152 ) | ( n24178 & n39152 ) ;
  assign n39154 = n39153 ^ n13670 ^ n9165 ;
  assign n39148 = n28558 ^ n15058 ^ n673 ;
  assign n39149 = n17973 ^ n1495 ^ 1'b0 ;
  assign n39150 = n39148 | n39149 ;
  assign n39155 = n39154 ^ n39150 ^ n13595 ;
  assign n39156 = n13016 ^ n11709 ^ n2976 ;
  assign n39157 = n2552 | n35163 ;
  assign n39158 = n6508 | n39157 ;
  assign n39159 = ( n1900 & n3252 ) | ( n1900 & n39158 ) | ( n3252 & n39158 ) ;
  assign n39160 = ( n5954 & n39156 ) | ( n5954 & n39159 ) | ( n39156 & n39159 ) ;
  assign n39161 = n22374 ^ n5845 ^ 1'b0 ;
  assign n39162 = ~n10285 & n39161 ;
  assign n39163 = n31716 ^ n16548 ^ n8210 ;
  assign n39164 = ( n10006 & ~n26741 ) | ( n10006 & n30297 ) | ( ~n26741 & n30297 ) ;
  assign n39165 = ( ~n10174 & n21030 ) | ( ~n10174 & n39164 ) | ( n21030 & n39164 ) ;
  assign n39166 = n39165 ^ n27355 ^ 1'b0 ;
  assign n39167 = n39163 & n39166 ;
  assign n39170 = n6269 | n13914 ;
  assign n39168 = n14599 ^ n14558 ^ n1496 ;
  assign n39169 = ( n6528 & n34778 ) | ( n6528 & n39168 ) | ( n34778 & n39168 ) ;
  assign n39171 = n39170 ^ n39169 ^ n22244 ;
  assign n39172 = n31145 ^ n25238 ^ n18983 ;
  assign n39173 = n26394 ^ n19965 ^ n4845 ;
  assign n39174 = ( n7735 & ~n21984 ) | ( n7735 & n39173 ) | ( ~n21984 & n39173 ) ;
  assign n39175 = n31145 ^ n6423 ^ n1294 ;
  assign n39176 = n39175 ^ n16919 ^ n6905 ;
  assign n39177 = n4888 & n20410 ;
  assign n39178 = n32494 & n39177 ;
  assign n39179 = n30725 ^ n26155 ^ n4178 ;
  assign n39180 = n18831 ^ n6067 ^ n2927 ;
  assign n39181 = n39180 ^ n17381 ^ n8243 ;
  assign n39182 = ( n39178 & ~n39179 ) | ( n39178 & n39181 ) | ( ~n39179 & n39181 ) ;
  assign n39183 = ( n15868 & n26917 ) | ( n15868 & ~n39182 ) | ( n26917 & ~n39182 ) ;
  assign n39184 = n2589 & n14913 ;
  assign n39185 = ~n768 & n19960 ;
  assign n39186 = ~n39184 & n39185 ;
  assign n39187 = n39186 ^ n13005 ^ n11987 ;
  assign n39190 = n23824 ^ n1644 ^ x171 ;
  assign n39191 = ( ~n3393 & n24904 ) | ( ~n3393 & n39190 ) | ( n24904 & n39190 ) ;
  assign n39188 = ~n2528 & n3702 ;
  assign n39189 = ( n24177 & n38722 ) | ( n24177 & n39188 ) | ( n38722 & n39188 ) ;
  assign n39192 = n39191 ^ n39189 ^ n6960 ;
  assign n39193 = ( n12676 & ~n18487 ) | ( n12676 & n24508 ) | ( ~n18487 & n24508 ) ;
  assign n39194 = n15349 ^ n9679 ^ n5468 ;
  assign n39195 = n5215 & ~n39194 ;
  assign n39196 = ( ~n12840 & n19415 ) | ( ~n12840 & n39195 ) | ( n19415 & n39195 ) ;
  assign n39197 = ( n35477 & ~n39193 ) | ( n35477 & n39196 ) | ( ~n39193 & n39196 ) ;
  assign n39198 = n39197 ^ n9565 ^ n2745 ;
  assign n39201 = ( n1135 & n7542 ) | ( n1135 & n26788 ) | ( n7542 & n26788 ) ;
  assign n39199 = n24467 ^ n21641 ^ n20728 ;
  assign n39200 = n39199 ^ n5347 ^ n4961 ;
  assign n39202 = n39201 ^ n39200 ^ 1'b0 ;
  assign n39203 = n1875 & n39202 ;
  assign n39204 = ( n26181 & n34930 ) | ( n26181 & n39203 ) | ( n34930 & n39203 ) ;
  assign n39205 = n2383 | n8679 ;
  assign n39206 = n5798 & ~n39205 ;
  assign n39207 = n39206 ^ n8589 ^ 1'b0 ;
  assign n39208 = n6261 & n39207 ;
  assign n39209 = ( n5908 & n39204 ) | ( n5908 & n39208 ) | ( n39204 & n39208 ) ;
  assign n39210 = n17888 ^ n15089 ^ 1'b0 ;
  assign n39211 = ( n14463 & n20166 ) | ( n14463 & ~n39210 ) | ( n20166 & ~n39210 ) ;
  assign n39212 = n35803 ^ n32782 ^ 1'b0 ;
  assign n39213 = ~n37032 & n39212 ;
  assign n39214 = n13242 ^ n1834 ^ n536 ;
  assign n39215 = ( n1578 & n2424 ) | ( n1578 & ~n5572 ) | ( n2424 & ~n5572 ) ;
  assign n39216 = ( n3408 & ~n14140 ) | ( n3408 & n39215 ) | ( ~n14140 & n39215 ) ;
  assign n39217 = ( n15678 & ~n39214 ) | ( n15678 & n39216 ) | ( ~n39214 & n39216 ) ;
  assign n39218 = n25583 ^ n7273 ^ 1'b0 ;
  assign n39219 = ~n39217 & n39218 ;
  assign n39223 = n6195 & ~n12369 ;
  assign n39224 = n39223 ^ n11258 ^ 1'b0 ;
  assign n39221 = n14859 ^ n8941 ^ n6917 ;
  assign n39222 = n39221 ^ n32860 ^ 1'b0 ;
  assign n39220 = ( n10534 & n11039 ) | ( n10534 & n36790 ) | ( n11039 & n36790 ) ;
  assign n39225 = n39224 ^ n39222 ^ n39220 ;
  assign n39226 = n35771 ^ n12364 ^ n2488 ;
  assign n39227 = ( n4173 & n23651 ) | ( n4173 & n39226 ) | ( n23651 & n39226 ) ;
  assign n39228 = n36758 ^ n10528 ^ n3244 ;
  assign n39229 = ( n15857 & n27188 ) | ( n15857 & ~n31951 ) | ( n27188 & ~n31951 ) ;
  assign n39230 = n39229 ^ n12826 ^ n6800 ;
  assign n39234 = n10340 ^ n9697 ^ n8790 ;
  assign n39231 = ~n3367 & n5437 ;
  assign n39232 = n16609 & ~n19005 ;
  assign n39233 = ( n8504 & n39231 ) | ( n8504 & ~n39232 ) | ( n39231 & ~n39232 ) ;
  assign n39235 = n39234 ^ n39233 ^ 1'b0 ;
  assign n39241 = n15065 ^ n13437 ^ n10444 ;
  assign n39242 = ( n5987 & n21162 ) | ( n5987 & n39241 ) | ( n21162 & n39241 ) ;
  assign n39239 = n33560 ^ n24405 ^ n7256 ;
  assign n39240 = ( ~n21502 & n27774 ) | ( ~n21502 & n39239 ) | ( n27774 & n39239 ) ;
  assign n39237 = n15515 ^ n14887 ^ 1'b0 ;
  assign n39236 = ( ~n1599 & n21243 ) | ( ~n1599 & n36740 ) | ( n21243 & n36740 ) ;
  assign n39238 = n39237 ^ n39236 ^ 1'b0 ;
  assign n39243 = n39242 ^ n39240 ^ n39238 ;
  assign n39244 = ( n2823 & ~n39235 ) | ( n2823 & n39243 ) | ( ~n39235 & n39243 ) ;
  assign n39245 = n11120 ^ n7954 ^ n1428 ;
  assign n39246 = n39245 ^ n2055 ^ 1'b0 ;
  assign n39247 = n10174 & ~n39246 ;
  assign n39248 = n21826 ^ n16880 ^ 1'b0 ;
  assign n39249 = n11624 & n39248 ;
  assign n39250 = n33781 ^ n6774 ^ 1'b0 ;
  assign n39251 = n18142 ^ n12765 ^ n8334 ;
  assign n39252 = ( n17262 & n17916 ) | ( n17262 & ~n39251 ) | ( n17916 & ~n39251 ) ;
  assign n39253 = ( n7559 & n21792 ) | ( n7559 & ~n38932 ) | ( n21792 & ~n38932 ) ;
  assign n39254 = n39253 ^ n24557 ^ 1'b0 ;
  assign n39255 = n36392 ^ n34280 ^ n24915 ;
  assign n39256 = ( ~n4306 & n27842 ) | ( ~n4306 & n30379 ) | ( n27842 & n30379 ) ;
  assign n39257 = ( n687 & n6584 ) | ( n687 & n7299 ) | ( n6584 & n7299 ) ;
  assign n39258 = n39257 ^ n16160 ^ 1'b0 ;
  assign n39259 = n30264 ^ n17662 ^ n1929 ;
  assign n39260 = ( ~n17016 & n39258 ) | ( ~n17016 & n39259 ) | ( n39258 & n39259 ) ;
  assign n39261 = n36085 ^ n24475 ^ n23452 ;
  assign n39262 = ( n3666 & n9466 ) | ( n3666 & ~n39261 ) | ( n9466 & ~n39261 ) ;
  assign n39263 = n17197 ^ n6896 ^ 1'b0 ;
  assign n39264 = ~n5008 & n39263 ;
  assign n39265 = n39264 ^ n21408 ^ n19336 ;
  assign n39266 = ( n25022 & ~n26117 ) | ( n25022 & n36329 ) | ( ~n26117 & n36329 ) ;
  assign n39267 = ( ~n9040 & n24031 ) | ( ~n9040 & n39266 ) | ( n24031 & n39266 ) ;
  assign n39268 = n15116 & n16344 ;
  assign n39269 = n39268 ^ n10523 ^ n6743 ;
  assign n39270 = n24850 ^ n23173 ^ n3452 ;
  assign n39271 = ( n19351 & n33335 ) | ( n19351 & ~n39270 ) | ( n33335 & ~n39270 ) ;
  assign n39272 = ( ~n1100 & n28115 ) | ( ~n1100 & n32884 ) | ( n28115 & n32884 ) ;
  assign n39273 = n39272 ^ n6377 ^ 1'b0 ;
  assign n39274 = n39271 & ~n39273 ;
  assign n39275 = n39274 ^ n38344 ^ n36566 ;
  assign n39276 = ( ~n21592 & n39269 ) | ( ~n21592 & n39275 ) | ( n39269 & n39275 ) ;
  assign n39277 = ( n2427 & n3498 ) | ( n2427 & n25753 ) | ( n3498 & n25753 ) ;
  assign n39278 = ( n16574 & n16626 ) | ( n16574 & ~n32984 ) | ( n16626 & ~n32984 ) ;
  assign n39281 = ( n9372 & n18483 ) | ( n9372 & ~n20448 ) | ( n18483 & ~n20448 ) ;
  assign n39279 = ~n6921 & n29259 ;
  assign n39280 = n3419 & n39279 ;
  assign n39282 = n39281 ^ n39280 ^ 1'b0 ;
  assign n39283 = n39282 ^ n5680 ^ n1779 ;
  assign n39286 = n30755 ^ n14518 ^ n2122 ;
  assign n39284 = n38665 ^ n18488 ^ n3847 ;
  assign n39285 = n39284 ^ n22081 ^ n4611 ;
  assign n39287 = n39286 ^ n39285 ^ n14365 ;
  assign n39288 = n20167 ^ n4071 ^ 1'b0 ;
  assign n39289 = n651 & n39288 ;
  assign n39293 = n19281 ^ n17197 ^ n13391 ;
  assign n39294 = n39293 ^ n16989 ^ n2793 ;
  assign n39295 = ~n2645 & n39294 ;
  assign n39296 = n39295 ^ n11954 ^ 1'b0 ;
  assign n39292 = n26524 ^ n24248 ^ n9635 ;
  assign n39290 = ( ~n5063 & n15341 ) | ( ~n5063 & n23291 ) | ( n15341 & n23291 ) ;
  assign n39291 = ( n13538 & n25811 ) | ( n13538 & ~n39290 ) | ( n25811 & ~n39290 ) ;
  assign n39297 = n39296 ^ n39292 ^ n39291 ;
  assign n39298 = n39289 & n39297 ;
  assign n39299 = n39298 ^ n2053 ^ 1'b0 ;
  assign n39300 = n16496 ^ n11452 ^ n9033 ;
  assign n39301 = ( n9119 & n13842 ) | ( n9119 & n39300 ) | ( n13842 & n39300 ) ;
  assign n39302 = ( n4356 & ~n10626 ) | ( n4356 & n31427 ) | ( ~n10626 & n31427 ) ;
  assign n39303 = n9335 | n33398 ;
  assign n39304 = ( n35044 & ~n39302 ) | ( n35044 & n39303 ) | ( ~n39302 & n39303 ) ;
  assign n39307 = ( n8387 & n11103 ) | ( n8387 & ~n35212 ) | ( n11103 & ~n35212 ) ;
  assign n39305 = n16669 ^ n1172 ^ n831 ;
  assign n39306 = ( n13741 & n38932 ) | ( n13741 & ~n39305 ) | ( n38932 & ~n39305 ) ;
  assign n39308 = n39307 ^ n39306 ^ n35797 ;
  assign n39309 = ~n6901 & n31510 ;
  assign n39310 = n8406 & n39309 ;
  assign n39311 = n12153 ^ n8743 ^ 1'b0 ;
  assign n39312 = n2641 & n25863 ;
  assign n39313 = n39312 ^ n17717 ^ 1'b0 ;
  assign n39314 = n23465 ^ n3375 ^ 1'b0 ;
  assign n39315 = n39314 ^ n30028 ^ 1'b0 ;
  assign n39316 = ( n10006 & ~n22452 ) | ( n10006 & n36445 ) | ( ~n22452 & n36445 ) ;
  assign n39317 = n11464 ^ n4865 ^ n2249 ;
  assign n39318 = n39317 ^ n12755 ^ 1'b0 ;
  assign n39319 = ( n5682 & ~n16086 ) | ( n5682 & n26080 ) | ( ~n16086 & n26080 ) ;
  assign n39320 = n19553 ^ n15190 ^ n9503 ;
  assign n39321 = ( n4802 & n39319 ) | ( n4802 & n39320 ) | ( n39319 & n39320 ) ;
  assign n39322 = ( n18408 & ~n22279 ) | ( n18408 & n39321 ) | ( ~n22279 & n39321 ) ;
  assign n39323 = ( ~n916 & n6397 ) | ( ~n916 & n32951 ) | ( n6397 & n32951 ) ;
  assign n39324 = n35245 ^ n11245 ^ n6648 ;
  assign n39328 = n25480 ^ n18117 ^ n8003 ;
  assign n39327 = ( ~n3498 & n9943 ) | ( ~n3498 & n32026 ) | ( n9943 & n32026 ) ;
  assign n39325 = n34024 ^ n33688 ^ n6240 ;
  assign n39326 = ( n14286 & n15118 ) | ( n14286 & n39325 ) | ( n15118 & n39325 ) ;
  assign n39329 = n39328 ^ n39327 ^ n39326 ;
  assign n39330 = n9005 & ~n12012 ;
  assign n39331 = n16318 & n39330 ;
  assign n39332 = n4349 & ~n32314 ;
  assign n39333 = n23228 & n39332 ;
  assign n39334 = n39333 ^ n7573 ^ 1'b0 ;
  assign n39335 = n33892 ^ n23780 ^ n12027 ;
  assign n39336 = n39335 ^ n32063 ^ n19282 ;
  assign n39338 = n34041 ^ n28782 ^ n4243 ;
  assign n39337 = n28017 ^ n25386 ^ n23467 ;
  assign n39339 = n39338 ^ n39337 ^ n8585 ;
  assign n39340 = ( n5734 & ~n6526 ) | ( n5734 & n16227 ) | ( ~n6526 & n16227 ) ;
  assign n39341 = ( n28597 & ~n37591 ) | ( n28597 & n39340 ) | ( ~n37591 & n39340 ) ;
  assign n39342 = n17403 | n22163 ;
  assign n39343 = ( n8857 & ~n20282 ) | ( n8857 & n39342 ) | ( ~n20282 & n39342 ) ;
  assign n39344 = ( n37048 & ~n39341 ) | ( n37048 & n39343 ) | ( ~n39341 & n39343 ) ;
  assign n39345 = n20714 ^ n6000 ^ n5540 ;
  assign n39346 = ( n23778 & n30089 ) | ( n23778 & n39345 ) | ( n30089 & n39345 ) ;
  assign n39347 = n39346 ^ n5558 ^ n3739 ;
  assign n39348 = n5719 | n14122 ;
  assign n39349 = n9079 | n39348 ;
  assign n39350 = n39349 ^ n24688 ^ n24199 ;
  assign n39351 = ( ~n4018 & n4135 ) | ( ~n4018 & n6575 ) | ( n4135 & n6575 ) ;
  assign n39352 = n33384 & n39351 ;
  assign n39353 = ( n9939 & ~n22449 ) | ( n9939 & n23713 ) | ( ~n22449 & n23713 ) ;
  assign n39354 = n39353 ^ n21760 ^ n15087 ;
  assign n39355 = n32822 & n38340 ;
  assign n39356 = ( ~n9895 & n11727 ) | ( ~n9895 & n24123 ) | ( n11727 & n24123 ) ;
  assign n39357 = n25490 ^ n8354 ^ 1'b0 ;
  assign n39358 = n38119 & n39357 ;
  assign n39359 = n39358 ^ n21227 ^ n707 ;
  assign n39360 = n19757 & n19938 ;
  assign n39361 = ~n34158 & n39360 ;
  assign n39362 = n39361 ^ n22197 ^ n16738 ;
  assign n39363 = n39362 ^ n6753 ^ 1'b0 ;
  assign n39364 = ( n2599 & n16681 ) | ( n2599 & ~n27288 ) | ( n16681 & ~n27288 ) ;
  assign n39365 = n39364 ^ n36782 ^ n21970 ;
  assign n39366 = ( ~n9238 & n22773 ) | ( ~n9238 & n25367 ) | ( n22773 & n25367 ) ;
  assign n39367 = n29281 ^ n23180 ^ n23143 ;
  assign n39368 = n39367 ^ n38853 ^ n4676 ;
  assign n39369 = n39368 ^ n22950 ^ n11970 ;
  assign n39370 = ( n11174 & ~n39366 ) | ( n11174 & n39369 ) | ( ~n39366 & n39369 ) ;
  assign n39371 = ( ~n464 & n12858 ) | ( ~n464 & n39370 ) | ( n12858 & n39370 ) ;
  assign n39372 = ( ~n766 & n13799 ) | ( ~n766 & n27939 ) | ( n13799 & n27939 ) ;
  assign n39374 = ( x116 & n6663 ) | ( x116 & n22713 ) | ( n6663 & n22713 ) ;
  assign n39373 = ( ~n2102 & n6591 ) | ( ~n2102 & n14386 ) | ( n6591 & n14386 ) ;
  assign n39375 = n39374 ^ n39373 ^ n3975 ;
  assign n39376 = n39375 ^ n7941 ^ n1133 ;
  assign n39377 = ( n12612 & n18738 ) | ( n12612 & n31576 ) | ( n18738 & n31576 ) ;
  assign n39378 = ( n15271 & ~n19305 ) | ( n15271 & n39377 ) | ( ~n19305 & n39377 ) ;
  assign n39379 = ( n4210 & n7045 ) | ( n4210 & n9948 ) | ( n7045 & n9948 ) ;
  assign n39380 = n39379 ^ n23946 ^ 1'b0 ;
  assign n39381 = ~n34223 & n39380 ;
  assign n39382 = n8157 ^ n3761 ^ 1'b0 ;
  assign n39387 = n12443 ^ n4390 ^ n2967 ;
  assign n39388 = ( ~x93 & n11718 ) | ( ~x93 & n39387 ) | ( n11718 & n39387 ) ;
  assign n39386 = ( ~n933 & n4717 ) | ( ~n933 & n11448 ) | ( n4717 & n11448 ) ;
  assign n39383 = ( ~n19654 & n24104 ) | ( ~n19654 & n38961 ) | ( n24104 & n38961 ) ;
  assign n39384 = n28048 ^ n7696 ^ n6258 ;
  assign n39385 = ( n34792 & ~n39383 ) | ( n34792 & n39384 ) | ( ~n39383 & n39384 ) ;
  assign n39389 = n39388 ^ n39386 ^ n39385 ;
  assign n39390 = n35896 ^ n21066 ^ n13012 ;
  assign n39391 = n28074 ^ n19553 ^ n13116 ;
  assign n39395 = n18455 ^ n14356 ^ n3009 ;
  assign n39392 = ( ~n11577 & n17564 ) | ( ~n11577 & n33374 ) | ( n17564 & n33374 ) ;
  assign n39393 = n39392 ^ n30691 ^ n23049 ;
  assign n39394 = n39393 ^ n20812 ^ n11661 ;
  assign n39396 = n39395 ^ n39394 ^ n11812 ;
  assign n39397 = n30095 ^ n4723 ^ 1'b0 ;
  assign n39398 = n36495 | n39397 ;
  assign n39399 = ( n6459 & n8986 ) | ( n6459 & n18529 ) | ( n8986 & n18529 ) ;
  assign n39400 = n39399 ^ n28680 ^ 1'b0 ;
  assign n39401 = n25915 & n39400 ;
  assign n39402 = ( n10197 & n14012 ) | ( n10197 & ~n24723 ) | ( n14012 & ~n24723 ) ;
  assign n39403 = ~n23253 & n31422 ;
  assign n39404 = n39403 ^ n10671 ^ 1'b0 ;
  assign n39405 = ( n8799 & n18882 ) | ( n8799 & ~n39404 ) | ( n18882 & ~n39404 ) ;
  assign n39406 = n8670 ^ n5264 ^ n3770 ;
  assign n39407 = n39406 ^ n38332 ^ n17606 ;
  assign n39409 = n23463 ^ n7898 ^ n4958 ;
  assign n39408 = n25146 ^ n21602 ^ n16015 ;
  assign n39410 = n39409 ^ n39408 ^ n16956 ;
  assign n39411 = n21415 ^ n18768 ^ n7825 ;
  assign n39412 = n39411 ^ n30023 ^ n15484 ;
  assign n39413 = ( n17194 & ~n21083 ) | ( n17194 & n21829 ) | ( ~n21083 & n21829 ) ;
  assign n39414 = ( n11194 & n13545 ) | ( n11194 & ~n19796 ) | ( n13545 & ~n19796 ) ;
  assign n39415 = n39414 ^ n5853 ^ n1236 ;
  assign n39416 = n6370 & n33329 ;
  assign n39417 = ~n3854 & n39416 ;
  assign n39418 = n4992 ^ n4862 ^ n4260 ;
  assign n39419 = n39418 ^ n32130 ^ x24 ;
  assign n39420 = n24493 ^ n5483 ^ 1'b0 ;
  assign n39422 = n38817 ^ n10702 ^ n5783 ;
  assign n39421 = ( ~n3217 & n22039 ) | ( ~n3217 & n35568 ) | ( n22039 & n35568 ) ;
  assign n39423 = n39422 ^ n39421 ^ n4314 ;
  assign n39424 = ( n39419 & n39420 ) | ( n39419 & ~n39423 ) | ( n39420 & ~n39423 ) ;
  assign n39432 = ( n1638 & n8525 ) | ( n1638 & ~n18821 ) | ( n8525 & ~n18821 ) ;
  assign n39431 = n26894 ^ n12156 ^ n5286 ;
  assign n39426 = n17917 ^ n8404 ^ n1290 ;
  assign n39425 = n18466 & n24725 ;
  assign n39427 = n39426 ^ n39425 ^ n13590 ;
  assign n39428 = ( n4361 & ~n10814 ) | ( n4361 & n39427 ) | ( ~n10814 & n39427 ) ;
  assign n39429 = ( n5367 & ~n5653 ) | ( n5367 & n19702 ) | ( ~n5653 & n19702 ) ;
  assign n39430 = ( n16275 & n39428 ) | ( n16275 & n39429 ) | ( n39428 & n39429 ) ;
  assign n39433 = n39432 ^ n39431 ^ n39430 ;
  assign n39434 = ( x32 & ~n5027 ) | ( x32 & n19984 ) | ( ~n5027 & n19984 ) ;
  assign n39435 = n16616 ^ n5050 ^ n430 ;
  assign n39436 = n39435 ^ n10669 ^ n7811 ;
  assign n39437 = n648 & n30368 ;
  assign n39438 = n28497 ^ n10253 ^ n5733 ;
  assign n39439 = n14888 ^ n9673 ^ 1'b0 ;
  assign n39440 = n8934 & ~n39439 ;
  assign n39441 = ( n1050 & ~n39438 ) | ( n1050 & n39440 ) | ( ~n39438 & n39440 ) ;
  assign n39442 = n17620 & ~n39441 ;
  assign n39443 = n35085 ^ n13585 ^ n5364 ;
  assign n39444 = n13914 & ~n39443 ;
  assign n39445 = ~n24212 & n39444 ;
  assign n39446 = ~n4926 & n26455 ;
  assign n39447 = ( n21115 & n31839 ) | ( n21115 & n39446 ) | ( n31839 & n39446 ) ;
  assign n39448 = ( x253 & ~n9174 ) | ( x253 & n20894 ) | ( ~n9174 & n20894 ) ;
  assign n39449 = n16878 & n39448 ;
  assign n39450 = n5091 & n39449 ;
  assign n39451 = n39450 ^ n34979 ^ 1'b0 ;
  assign n39452 = ~n39447 & n39451 ;
  assign n39453 = ( n1243 & ~n16511 ) | ( n1243 & n36982 ) | ( ~n16511 & n36982 ) ;
  assign n39454 = ( n21718 & n24424 ) | ( n21718 & n39453 ) | ( n24424 & n39453 ) ;
  assign n39455 = n39454 ^ n33522 ^ n25426 ;
  assign n39456 = n22394 ^ n16035 ^ n13848 ;
  assign n39463 = ( n4877 & n18259 ) | ( n4877 & n22262 ) | ( n18259 & n22262 ) ;
  assign n39461 = n6304 & n21279 ;
  assign n39462 = n7919 & n39461 ;
  assign n39457 = ( ~n8865 & n19005 ) | ( ~n8865 & n32837 ) | ( n19005 & n32837 ) ;
  assign n39458 = ( n3307 & n5347 ) | ( n3307 & ~n14914 ) | ( n5347 & ~n14914 ) ;
  assign n39459 = ( ~n8181 & n23972 ) | ( ~n8181 & n39458 ) | ( n23972 & n39458 ) ;
  assign n39460 = n39457 | n39459 ;
  assign n39464 = n39463 ^ n39462 ^ n39460 ;
  assign n39465 = ( n9895 & n15209 ) | ( n9895 & n19907 ) | ( n15209 & n19907 ) ;
  assign n39471 = n6350 ^ n3562 ^ n971 ;
  assign n39467 = x171 ^ x42 ^ 1'b0 ;
  assign n39468 = ~n6254 & n39467 ;
  assign n39469 = ~n16211 & n39468 ;
  assign n39470 = n23030 & n39469 ;
  assign n39466 = ( n10809 & ~n24849 ) | ( n10809 & n33288 ) | ( ~n24849 & n33288 ) ;
  assign n39472 = n39471 ^ n39470 ^ n39466 ;
  assign n39473 = n39472 ^ n17053 ^ n14804 ;
  assign n39474 = ( n19546 & n20923 ) | ( n19546 & n39473 ) | ( n20923 & n39473 ) ;
  assign n39475 = ( n33363 & n38873 ) | ( n33363 & ~n39178 ) | ( n38873 & ~n39178 ) ;
  assign n39476 = n27614 ^ n268 ^ 1'b0 ;
  assign n39477 = n3308 | n39476 ;
  assign n39481 = n5336 ^ n2518 ^ x146 ;
  assign n39482 = ( n14931 & n15496 ) | ( n14931 & ~n39481 ) | ( n15496 & ~n39481 ) ;
  assign n39483 = n39482 ^ n19858 ^ n15171 ;
  assign n39480 = n14931 & n32130 ;
  assign n39478 = n18713 ^ n7270 ^ n4694 ;
  assign n39479 = n39478 ^ n37502 ^ n15177 ;
  assign n39484 = n39483 ^ n39480 ^ n39479 ;
  assign n39485 = ( n17652 & n20578 ) | ( n17652 & n39484 ) | ( n20578 & n39484 ) ;
  assign n39486 = n10438 ^ n7264 ^ n3242 ;
  assign n39487 = ( n6536 & ~n9151 ) | ( n6536 & n36943 ) | ( ~n9151 & n36943 ) ;
  assign n39488 = ( n1339 & ~n37914 ) | ( n1339 & n39487 ) | ( ~n37914 & n39487 ) ;
  assign n39489 = ( n6557 & ~n8590 ) | ( n6557 & n9576 ) | ( ~n8590 & n9576 ) ;
  assign n39490 = ( ~n2537 & n14101 ) | ( ~n2537 & n39489 ) | ( n14101 & n39489 ) ;
  assign n39491 = ( ~n2853 & n14424 ) | ( ~n2853 & n17743 ) | ( n14424 & n17743 ) ;
  assign n39492 = ~n1278 & n39491 ;
  assign n39494 = n22950 ^ n707 ^ 1'b0 ;
  assign n39495 = x54 & ~n39494 ;
  assign n39496 = ( n16043 & ~n26966 ) | ( n16043 & n39495 ) | ( ~n26966 & n39495 ) ;
  assign n39493 = ( n2761 & ~n8170 ) | ( n2761 & n10148 ) | ( ~n8170 & n10148 ) ;
  assign n39497 = n39496 ^ n39493 ^ n2069 ;
  assign n39498 = n2098 ^ n733 ^ 1'b0 ;
  assign n39499 = ( n8937 & n12755 ) | ( n8937 & ~n39498 ) | ( n12755 & ~n39498 ) ;
  assign n39500 = n31149 ^ n18081 ^ n7290 ;
  assign n39501 = n23473 | n39500 ;
  assign n39502 = n39501 ^ n13478 ^ 1'b0 ;
  assign n39504 = ( ~n6374 & n8356 ) | ( ~n6374 & n29801 ) | ( n8356 & n29801 ) ;
  assign n39503 = n32438 ^ n21432 ^ n17133 ;
  assign n39505 = n39504 ^ n39503 ^ n30962 ;
  assign n39506 = n39505 ^ n27500 ^ n13285 ;
  assign n39507 = n23514 ^ n17973 ^ n2101 ;
  assign n39508 = ( n34529 & ~n39450 ) | ( n34529 & n39507 ) | ( ~n39450 & n39507 ) ;
  assign n39509 = n17683 ^ n15096 ^ 1'b0 ;
  assign n39510 = ~n13357 & n39509 ;
  assign n39511 = ( n13067 & n29582 ) | ( n13067 & n39510 ) | ( n29582 & n39510 ) ;
  assign n39512 = n39511 ^ n34131 ^ n30154 ;
  assign n39518 = n33263 ^ n27531 ^ n25969 ;
  assign n39519 = n39518 ^ n38918 ^ n14817 ;
  assign n39515 = n37587 ^ n5067 ^ 1'b0 ;
  assign n39516 = n2143 & ~n39515 ;
  assign n39517 = n39516 ^ n27125 ^ 1'b0 ;
  assign n39513 = n8573 ^ n8143 ^ n3807 ;
  assign n39514 = n20608 & ~n39513 ;
  assign n39520 = n39519 ^ n39517 ^ n39514 ;
  assign n39521 = n39520 ^ n22673 ^ n6077 ;
  assign n39522 = ( ~n3948 & n7824 ) | ( ~n3948 & n23634 ) | ( n7824 & n23634 ) ;
  assign n39523 = n5914 & ~n7304 ;
  assign n39524 = n39523 ^ n10843 ^ 1'b0 ;
  assign n39525 = n39524 ^ n11112 ^ n9550 ;
  assign n39526 = n4279 & n39525 ;
  assign n39527 = n22308 & n39526 ;
  assign n39528 = n4437 & n11319 ;
  assign n39529 = n16545 & n39528 ;
  assign n39530 = n8103 ^ n6488 ^ n755 ;
  assign n39531 = n39530 ^ n19069 ^ 1'b0 ;
  assign n39532 = n9828 & n25318 ;
  assign n39533 = ( n1846 & ~n22451 ) | ( n1846 & n39532 ) | ( ~n22451 & n39532 ) ;
  assign n39534 = n39533 ^ n16161 ^ n15174 ;
  assign n39535 = n39534 ^ n12308 ^ n2582 ;
  assign n39536 = ~n9941 & n31476 ;
  assign n39537 = ~n29906 & n39536 ;
  assign n39538 = ~n12824 & n14190 ;
  assign n39539 = n39537 & n39538 ;
  assign n39540 = n39539 ^ n31648 ^ n13511 ;
  assign n39541 = ( n5918 & n6425 ) | ( n5918 & ~n22047 ) | ( n6425 & ~n22047 ) ;
  assign n39542 = ~n2516 & n12184 ;
  assign n39543 = n39541 & n39542 ;
  assign n39544 = n39543 ^ n29347 ^ n14892 ;
  assign n39545 = n39544 ^ n36339 ^ n22582 ;
  assign n39546 = ( n11340 & ~n20733 ) | ( n11340 & n39545 ) | ( ~n20733 & n39545 ) ;
  assign n39548 = n19467 ^ n5285 ^ n1696 ;
  assign n39549 = n39548 ^ n8377 ^ n828 ;
  assign n39550 = n39549 ^ n22137 ^ n15264 ;
  assign n39551 = n39550 ^ n13105 ^ n10729 ;
  assign n39547 = ( n4210 & n4859 ) | ( n4210 & ~n22996 ) | ( n4859 & ~n22996 ) ;
  assign n39552 = n39551 ^ n39547 ^ n520 ;
  assign n39553 = ( n4005 & n6776 ) | ( n4005 & n31938 ) | ( n6776 & n31938 ) ;
  assign n39554 = ( n10502 & n25094 ) | ( n10502 & ~n32196 ) | ( n25094 & ~n32196 ) ;
  assign n39555 = n39554 ^ n23140 ^ 1'b0 ;
  assign n39556 = n39555 ^ n12974 ^ 1'b0 ;
  assign n39557 = ~n9355 & n39556 ;
  assign n39558 = ( n9204 & n21899 ) | ( n9204 & n39557 ) | ( n21899 & n39557 ) ;
  assign n39559 = n27817 ^ n11720 ^ n3278 ;
  assign n39560 = ( ~n6252 & n19243 ) | ( ~n6252 & n39559 ) | ( n19243 & n39559 ) ;
  assign n39561 = ( n4583 & n11958 ) | ( n4583 & ~n39560 ) | ( n11958 & ~n39560 ) ;
  assign n39562 = n39561 ^ n28616 ^ n6469 ;
  assign n39563 = ~n3650 & n18037 ;
  assign n39564 = ~n14842 & n39563 ;
  assign n39565 = n37130 | n39564 ;
  assign n39566 = n39562 & ~n39565 ;
  assign n39567 = ( n4926 & n11788 ) | ( n4926 & ~n19875 ) | ( n11788 & ~n19875 ) ;
  assign n39568 = n39567 ^ n17676 ^ n4890 ;
  assign n39569 = n21359 ^ n14067 ^ n5270 ;
  assign n39570 = ( n1106 & n35313 ) | ( n1106 & n37473 ) | ( n35313 & n37473 ) ;
  assign n39571 = n39570 ^ n18177 ^ n12228 ;
  assign n39572 = ( n3213 & n16440 ) | ( n3213 & n28212 ) | ( n16440 & n28212 ) ;
  assign n39573 = n20073 ^ n8815 ^ x66 ;
  assign n39574 = ( n1511 & ~n2310 ) | ( n1511 & n2552 ) | ( ~n2310 & n2552 ) ;
  assign n39575 = n39574 ^ n39207 ^ n37160 ;
  assign n39576 = ( n11883 & n32463 ) | ( n11883 & n39575 ) | ( n32463 & n39575 ) ;
  assign n39577 = n39576 ^ n31213 ^ n10169 ;
  assign n39578 = n30515 ^ n17524 ^ n3573 ;
  assign n39579 = n750 & ~n5609 ;
  assign n39580 = ( n21002 & ~n24751 ) | ( n21002 & n39579 ) | ( ~n24751 & n39579 ) ;
  assign n39581 = n3891 | n25360 ;
  assign n39582 = n14421 | n38987 ;
  assign n39583 = n39582 ^ n9873 ^ 1'b0 ;
  assign n39585 = ( n2225 & n11748 ) | ( n2225 & n36790 ) | ( n11748 & n36790 ) ;
  assign n39584 = ( n294 & n18782 ) | ( n294 & ~n26228 ) | ( n18782 & ~n26228 ) ;
  assign n39586 = n39585 ^ n39584 ^ n13848 ;
  assign n39587 = n37697 ^ n29494 ^ n27757 ;
  assign n39588 = n39587 ^ n12007 ^ n1805 ;
  assign n39589 = ( n10704 & n14085 ) | ( n10704 & ~n39588 ) | ( n14085 & ~n39588 ) ;
  assign n39590 = n19198 ^ n16269 ^ n8878 ;
  assign n39591 = ( ~n26310 & n32131 ) | ( ~n26310 & n39590 ) | ( n32131 & n39590 ) ;
  assign n39592 = n39591 ^ n37928 ^ n26199 ;
  assign n39593 = n11463 ^ n10293 ^ n10278 ;
  assign n39594 = ( n1129 & n29788 ) | ( n1129 & n39593 ) | ( n29788 & n39593 ) ;
  assign n39595 = ( n14184 & n31979 ) | ( n14184 & ~n36224 ) | ( n31979 & ~n36224 ) ;
  assign n39596 = n22352 & ~n39595 ;
  assign n39597 = n36378 ^ n6453 ^ n2333 ;
  assign n39598 = n24196 ^ n8846 ^ n1346 ;
  assign n39600 = n37653 ^ n21363 ^ n3339 ;
  assign n39601 = n39600 ^ n26271 ^ n20235 ;
  assign n39602 = n39601 ^ n29860 ^ n8469 ;
  assign n39599 = n19499 ^ n14996 ^ n7884 ;
  assign n39603 = n39602 ^ n39599 ^ 1'b0 ;
  assign n39604 = n26410 | n39603 ;
  assign n39605 = n33907 ^ n25714 ^ 1'b0 ;
  assign n39607 = n11678 ^ n10407 ^ n4739 ;
  assign n39608 = n39607 ^ n2860 ^ n1760 ;
  assign n39609 = n39608 ^ n4990 ^ n4051 ;
  assign n39606 = n22473 ^ n13171 ^ n7202 ;
  assign n39610 = n39609 ^ n39606 ^ n34483 ;
  assign n39611 = ( n6068 & ~n39605 ) | ( n6068 & n39610 ) | ( ~n39605 & n39610 ) ;
  assign n39612 = ( n9462 & n12152 ) | ( n9462 & ~n21210 ) | ( n12152 & ~n21210 ) ;
  assign n39613 = n39612 ^ n19943 ^ 1'b0 ;
  assign n39614 = n39611 | n39613 ;
  assign n39615 = n16522 ^ n9921 ^ 1'b0 ;
  assign n39616 = n34168 ^ n19023 ^ n2371 ;
  assign n39617 = ( n28170 & n30761 ) | ( n28170 & n39616 ) | ( n30761 & n39616 ) ;
  assign n39618 = ( n21011 & n39615 ) | ( n21011 & n39617 ) | ( n39615 & n39617 ) ;
  assign n39623 = n35052 ^ n15341 ^ n4170 ;
  assign n39624 = n11224 & ~n39623 ;
  assign n39625 = n39624 ^ n17565 ^ 1'b0 ;
  assign n39626 = n35655 & ~n39625 ;
  assign n39627 = ( ~n14039 & n17976 ) | ( ~n14039 & n39626 ) | ( n17976 & n39626 ) ;
  assign n39619 = n37887 ^ n20787 ^ n8996 ;
  assign n39620 = ( n9155 & n29169 ) | ( n9155 & n39619 ) | ( n29169 & n39619 ) ;
  assign n39621 = n30503 & n39620 ;
  assign n39622 = ( n8716 & n39620 ) | ( n8716 & ~n39621 ) | ( n39620 & ~n39621 ) ;
  assign n39628 = n39627 ^ n39622 ^ n3830 ;
  assign n39630 = n17874 ^ n12455 ^ n11286 ;
  assign n39631 = n33825 ^ n16305 ^ n3895 ;
  assign n39632 = n39631 ^ n34948 ^ n6173 ;
  assign n39633 = ( n6087 & ~n39630 ) | ( n6087 & n39632 ) | ( ~n39630 & n39632 ) ;
  assign n39629 = ( ~n3565 & n26891 ) | ( ~n3565 & n28004 ) | ( n26891 & n28004 ) ;
  assign n39634 = n39633 ^ n39629 ^ 1'b0 ;
  assign n39635 = n35389 ^ n8305 ^ n1283 ;
  assign n39636 = n25333 ^ n24694 ^ n17922 ;
  assign n39637 = ( n12984 & ~n20737 ) | ( n12984 & n39636 ) | ( ~n20737 & n39636 ) ;
  assign n39638 = ( n9584 & n34135 ) | ( n9584 & ~n39637 ) | ( n34135 & ~n39637 ) ;
  assign n39639 = ( n38200 & n39635 ) | ( n38200 & ~n39638 ) | ( n39635 & ~n39638 ) ;
  assign n39640 = n17881 ^ n8463 ^ n3305 ;
  assign n39641 = ( n2524 & n18489 ) | ( n2524 & n35568 ) | ( n18489 & n35568 ) ;
  assign n39642 = ( n17513 & n39640 ) | ( n17513 & ~n39641 ) | ( n39640 & ~n39641 ) ;
  assign n39643 = ( ~n3329 & n15769 ) | ( ~n3329 & n39642 ) | ( n15769 & n39642 ) ;
  assign n39644 = n18018 ^ n16947 ^ n7514 ;
  assign n39645 = n7768 & ~n17933 ;
  assign n39646 = ~n39644 & n39645 ;
  assign n39647 = n23073 ^ n5764 ^ x204 ;
  assign n39648 = ( n342 & n17218 ) | ( n342 & n23243 ) | ( n17218 & n23243 ) ;
  assign n39649 = ( n13272 & n39647 ) | ( n13272 & n39648 ) | ( n39647 & n39648 ) ;
  assign n39650 = n11157 & n34267 ;
  assign n39651 = n39650 ^ n23915 ^ n704 ;
  assign n39652 = n12814 | n36016 ;
  assign n39653 = ( n14904 & ~n23813 ) | ( n14904 & n39652 ) | ( ~n23813 & n39652 ) ;
  assign n39654 = n39653 ^ n4171 ^ 1'b0 ;
  assign n39655 = ( n4941 & n18910 ) | ( n4941 & n31034 ) | ( n18910 & n31034 ) ;
  assign n39656 = ( n2951 & n3664 ) | ( n2951 & n9617 ) | ( n3664 & n9617 ) ;
  assign n39657 = n39656 ^ n9029 ^ 1'b0 ;
  assign n39658 = n16427 ^ n2441 ^ 1'b0 ;
  assign n39659 = n36883 & n39658 ;
  assign n39660 = n23263 ^ n20162 ^ n13663 ;
  assign n39661 = ( ~n28631 & n35381 ) | ( ~n28631 & n39660 ) | ( n35381 & n39660 ) ;
  assign n39662 = ( ~n7927 & n30353 ) | ( ~n7927 & n39661 ) | ( n30353 & n39661 ) ;
  assign n39663 = n38188 ^ n32664 ^ 1'b0 ;
  assign n39664 = n12036 | n39663 ;
  assign n39665 = n37311 | n39664 ;
  assign n39666 = n39665 ^ n23579 ^ n2743 ;
  assign n39667 = n22802 | n22996 ;
  assign n39668 = n39667 ^ n10200 ^ 1'b0 ;
  assign n39669 = ( n3019 & ~n8773 ) | ( n3019 & n39668 ) | ( ~n8773 & n39668 ) ;
  assign n39670 = n10889 ^ n404 ^ 1'b0 ;
  assign n39671 = ~n3619 & n39670 ;
  assign n39672 = ( n804 & ~n1368 ) | ( n804 & n39671 ) | ( ~n1368 & n39671 ) ;
  assign n39673 = ( ~n767 & n23212 ) | ( ~n767 & n35114 ) | ( n23212 & n35114 ) ;
  assign n39674 = n33657 ^ n20493 ^ n6141 ;
  assign n39675 = ( ~n12341 & n33211 ) | ( ~n12341 & n35028 ) | ( n33211 & n35028 ) ;
  assign n39676 = ( n649 & n9256 ) | ( n649 & ~n31147 ) | ( n9256 & ~n31147 ) ;
  assign n39677 = ( n12558 & ~n18723 ) | ( n12558 & n39676 ) | ( ~n18723 & n39676 ) ;
  assign n39678 = ( ~n7441 & n19574 ) | ( ~n7441 & n39677 ) | ( n19574 & n39677 ) ;
  assign n39679 = ( n2511 & n13009 ) | ( n2511 & ~n16565 ) | ( n13009 & ~n16565 ) ;
  assign n39680 = n39679 ^ n20698 ^ n20375 ;
  assign n39681 = ~n2792 & n39680 ;
  assign n39685 = ( ~n11241 & n14527 ) | ( ~n11241 & n33118 ) | ( n14527 & n33118 ) ;
  assign n39682 = n17415 ^ n15863 ^ n10222 ;
  assign n39683 = n14045 & n39682 ;
  assign n39684 = n7963 & n39683 ;
  assign n39686 = n39685 ^ n39684 ^ n3079 ;
  assign n39687 = ( n6609 & n8145 ) | ( n6609 & ~n18113 ) | ( n8145 & ~n18113 ) ;
  assign n39688 = ( n18809 & n24135 ) | ( n18809 & ~n39687 ) | ( n24135 & ~n39687 ) ;
  assign n39689 = n39688 ^ n23307 ^ n9996 ;
  assign n39690 = ( ~n9095 & n9971 ) | ( ~n9095 & n11007 ) | ( n9971 & n11007 ) ;
  assign n39691 = ( n2275 & n4366 ) | ( n2275 & n39690 ) | ( n4366 & n39690 ) ;
  assign n39692 = n4508 ^ n1145 ^ n605 ;
  assign n39693 = n17428 ^ n7093 ^ n4321 ;
  assign n39694 = ( n27966 & n39692 ) | ( n27966 & ~n39693 ) | ( n39692 & ~n39693 ) ;
  assign n39695 = n23919 ^ n20076 ^ n7040 ;
  assign n39696 = n24920 ^ n3586 ^ n335 ;
  assign n39697 = ( n18593 & ~n34422 ) | ( n18593 & n39696 ) | ( ~n34422 & n39696 ) ;
  assign n39698 = n38476 ^ n18337 ^ 1'b0 ;
  assign n39699 = ( n2184 & n9060 ) | ( n2184 & ~n39698 ) | ( n9060 & ~n39698 ) ;
  assign n39700 = ( n31625 & n39697 ) | ( n31625 & ~n39699 ) | ( n39697 & ~n39699 ) ;
  assign n39701 = n36155 ^ n11894 ^ 1'b0 ;
  assign n39702 = ~n15169 & n39701 ;
  assign n39703 = n30642 ^ n4448 ^ n2589 ;
  assign n39704 = n828 & n39703 ;
  assign n39705 = ~n39702 & n39704 ;
  assign n39706 = ( n7977 & n10411 ) | ( n7977 & n14811 ) | ( n10411 & n14811 ) ;
  assign n39707 = n39706 ^ n26157 ^ n22368 ;
  assign n39708 = n39707 ^ n33568 ^ n8761 ;
  assign n39709 = n39708 ^ n9854 ^ 1'b0 ;
  assign n39710 = n38778 & n39709 ;
  assign n39711 = ( n2958 & n7397 ) | ( n2958 & ~n36206 ) | ( n7397 & ~n36206 ) ;
  assign n39712 = n39711 ^ n25195 ^ 1'b0 ;
  assign n39713 = ( ~n10121 & n22870 ) | ( ~n10121 & n39712 ) | ( n22870 & n39712 ) ;
  assign n39715 = n23874 ^ x175 ^ 1'b0 ;
  assign n39716 = n13874 & n39715 ;
  assign n39717 = ( n7261 & n31472 ) | ( n7261 & ~n39716 ) | ( n31472 & ~n39716 ) ;
  assign n39714 = ( n19664 & ~n28434 ) | ( n19664 & n36962 ) | ( ~n28434 & n36962 ) ;
  assign n39718 = n39717 ^ n39714 ^ n20325 ;
  assign n39719 = ( n1817 & n4176 ) | ( n1817 & n35325 ) | ( n4176 & n35325 ) ;
  assign n39720 = n21497 ^ n15108 ^ n258 ;
  assign n39721 = ( n7724 & n25640 ) | ( n7724 & n35938 ) | ( n25640 & n35938 ) ;
  assign n39722 = n39721 ^ n39539 ^ n32114 ;
  assign n39723 = ( n3185 & ~n3382 ) | ( n3185 & n25736 ) | ( ~n3382 & n25736 ) ;
  assign n39726 = n22689 ^ n5865 ^ n1382 ;
  assign n39724 = n4407 & n5541 ;
  assign n39725 = n39724 ^ n7908 ^ 1'b0 ;
  assign n39727 = n39726 ^ n39725 ^ n12712 ;
  assign n39728 = ( n3546 & ~n17781 ) | ( n3546 & n23276 ) | ( ~n17781 & n23276 ) ;
  assign n39729 = n7303 ^ n1645 ^ 1'b0 ;
  assign n39730 = n39729 ^ n16290 ^ 1'b0 ;
  assign n39731 = ~n39728 & n39730 ;
  assign n39732 = n31770 ^ n27369 ^ 1'b0 ;
  assign n39733 = ( ~n4254 & n29619 ) | ( ~n4254 & n39732 ) | ( n29619 & n39732 ) ;
  assign n39734 = ( n13615 & n27957 ) | ( n13615 & n39733 ) | ( n27957 & n39733 ) ;
  assign n39735 = ( n3139 & ~n11452 ) | ( n3139 & n19280 ) | ( ~n11452 & n19280 ) ;
  assign n39736 = ( n901 & n5956 ) | ( n901 & n10531 ) | ( n5956 & n10531 ) ;
  assign n39737 = ( n5340 & n10457 ) | ( n5340 & ~n21574 ) | ( n10457 & ~n21574 ) ;
  assign n39738 = ( n31127 & n39736 ) | ( n31127 & ~n39737 ) | ( n39736 & ~n39737 ) ;
  assign n39739 = ( n647 & ~n3242 ) | ( n647 & n4760 ) | ( ~n3242 & n4760 ) ;
  assign n39740 = n955 | n22299 ;
  assign n39741 = n12976 | n39740 ;
  assign n39742 = n39741 ^ n20542 ^ n1775 ;
  assign n39743 = n6766 | n13459 ;
  assign n39744 = n25740 & ~n39743 ;
  assign n39745 = ( n10381 & n11147 ) | ( n10381 & n39744 ) | ( n11147 & n39744 ) ;
  assign n39746 = ( ~n11653 & n32525 ) | ( ~n11653 & n39745 ) | ( n32525 & n39745 ) ;
  assign n39747 = n4355 | n38376 ;
  assign n39748 = n37258 ^ n9635 ^ 1'b0 ;
  assign n39749 = n39747 & ~n39748 ;
  assign n39751 = n15430 ^ n13493 ^ n3657 ;
  assign n39752 = n39751 ^ n16990 ^ n9201 ;
  assign n39753 = ( n402 & ~n14673 ) | ( n402 & n39752 ) | ( ~n14673 & n39752 ) ;
  assign n39750 = n5737 & n30733 ;
  assign n39754 = n39753 ^ n39750 ^ 1'b0 ;
  assign n39759 = n10077 ^ n8980 ^ n3613 ;
  assign n39755 = ( ~n3318 & n9368 ) | ( ~n3318 & n15834 ) | ( n9368 & n15834 ) ;
  assign n39756 = n39755 ^ n5563 ^ n636 ;
  assign n39757 = n18108 | n18481 ;
  assign n39758 = n39756 & ~n39757 ;
  assign n39760 = n39759 ^ n39758 ^ n3483 ;
  assign n39761 = n18154 ^ n14485 ^ n2918 ;
  assign n39762 = ( n2591 & n8472 ) | ( n2591 & n39761 ) | ( n8472 & n39761 ) ;
  assign n39763 = n9847 ^ n2593 ^ 1'b0 ;
  assign n39764 = n39763 ^ n21553 ^ n17143 ;
  assign n39767 = ( ~n9643 & n12481 ) | ( ~n9643 & n30443 ) | ( n12481 & n30443 ) ;
  assign n39765 = ( n14510 & n24611 ) | ( n14510 & ~n33362 ) | ( n24611 & ~n33362 ) ;
  assign n39766 = n39765 ^ n38561 ^ n5935 ;
  assign n39768 = n39767 ^ n39766 ^ n8742 ;
  assign n39769 = ( n10626 & n19621 ) | ( n10626 & n21689 ) | ( n19621 & n21689 ) ;
  assign n39770 = n39769 ^ n32967 ^ n26523 ;
  assign n39771 = n29251 | n39136 ;
  assign n39772 = n28141 | n39771 ;
  assign n39773 = n26568 ^ n20748 ^ n15892 ;
  assign n39775 = ( n6405 & n14861 ) | ( n6405 & ~n16754 ) | ( n14861 & ~n16754 ) ;
  assign n39774 = n5834 ^ n5748 ^ 1'b0 ;
  assign n39776 = n39775 ^ n39774 ^ n16808 ;
  assign n39777 = n29754 ^ n29122 ^ n6551 ;
  assign n39778 = n25321 | n29651 ;
  assign n39779 = n35828 ^ n30168 ^ n16282 ;
  assign n39780 = ( n13776 & n24276 ) | ( n13776 & ~n39779 ) | ( n24276 & ~n39779 ) ;
  assign n39781 = n39780 ^ n36938 ^ n24390 ;
  assign n39782 = ( ~n8323 & n10579 ) | ( ~n8323 & n33968 ) | ( n10579 & n33968 ) ;
  assign n39783 = ( n5199 & n18110 ) | ( n5199 & ~n39782 ) | ( n18110 & ~n39782 ) ;
  assign n39784 = ( n26649 & ~n27593 ) | ( n26649 & n38503 ) | ( ~n27593 & n38503 ) ;
  assign n39792 = n9598 | n10741 ;
  assign n39793 = n23977 | n39792 ;
  assign n39789 = n12651 & n13441 ;
  assign n39790 = n19196 & n39789 ;
  assign n39788 = ( n1336 & ~n8404 ) | ( n1336 & n10377 ) | ( ~n8404 & n10377 ) ;
  assign n39791 = n39790 ^ n39788 ^ n31606 ;
  assign n39785 = ( ~n14243 & n24434 ) | ( ~n14243 & n32315 ) | ( n24434 & n32315 ) ;
  assign n39786 = ( n8854 & n19312 ) | ( n8854 & n39785 ) | ( n19312 & n39785 ) ;
  assign n39787 = n39786 ^ n38300 ^ n10311 ;
  assign n39794 = n39793 ^ n39791 ^ n39787 ;
  assign n39798 = ( ~n1548 & n28444 ) | ( ~n1548 & n34722 ) | ( n28444 & n34722 ) ;
  assign n39795 = n16565 ^ n1613 ^ 1'b0 ;
  assign n39796 = n3533 & ~n39795 ;
  assign n39797 = ( n3601 & n37962 ) | ( n3601 & n39796 ) | ( n37962 & n39796 ) ;
  assign n39799 = n39798 ^ n39797 ^ 1'b0 ;
  assign n39800 = ( ~n22609 & n26991 ) | ( ~n22609 & n36544 ) | ( n26991 & n36544 ) ;
  assign n39801 = n39800 ^ n910 ^ 1'b0 ;
  assign n39802 = n35261 ^ n10973 ^ 1'b0 ;
  assign n39803 = n39377 ^ n6588 ^ 1'b0 ;
  assign n39804 = n2379 | n39803 ;
  assign n39805 = n27984 ^ n11104 ^ x189 ;
  assign n39806 = n39805 ^ n12716 ^ n5607 ;
  assign n39807 = n19709 ^ n1113 ^ x6 ;
  assign n39808 = n26739 ^ n17912 ^ n4862 ;
  assign n39809 = ( ~n5169 & n8450 ) | ( ~n5169 & n39808 ) | ( n8450 & n39808 ) ;
  assign n39810 = n21796 ^ n8215 ^ n6728 ;
  assign n39811 = n30761 ^ n8734 ^ n1756 ;
  assign n39812 = ( ~n26530 & n39810 ) | ( ~n26530 & n39811 ) | ( n39810 & n39811 ) ;
  assign n39813 = n34923 ^ n8720 ^ 1'b0 ;
  assign n39815 = n14371 ^ n11020 ^ 1'b0 ;
  assign n39816 = n39815 ^ n17905 ^ n10005 ;
  assign n39814 = ( ~n7654 & n14748 ) | ( ~n7654 & n31964 ) | ( n14748 & n31964 ) ;
  assign n39817 = n39816 ^ n39814 ^ n11122 ;
  assign n39818 = n39817 ^ n31638 ^ 1'b0 ;
  assign n39819 = n27206 ^ n10793 ^ n4385 ;
  assign n39820 = n39819 ^ n21636 ^ n19850 ;
  assign n39821 = n39820 ^ n28264 ^ n2642 ;
  assign n39822 = ~n25043 & n33390 ;
  assign n39823 = n39822 ^ n9585 ^ 1'b0 ;
  assign n39824 = ~n6009 & n13780 ;
  assign n39825 = n39824 ^ n26959 ^ 1'b0 ;
  assign n39826 = ( n13293 & n15151 ) | ( n13293 & ~n36594 ) | ( n15151 & ~n36594 ) ;
  assign n39827 = n39826 ^ n30913 ^ n28090 ;
  assign n39830 = n11043 ^ n9763 ^ n7518 ;
  assign n39831 = n39830 ^ n12690 ^ n9852 ;
  assign n39828 = ( n10820 & n19736 ) | ( n10820 & ~n23182 ) | ( n19736 & ~n23182 ) ;
  assign n39829 = n39828 ^ n11891 ^ n8663 ;
  assign n39832 = n39831 ^ n39829 ^ n25554 ;
  assign n39833 = n34175 ^ n20455 ^ n6705 ;
  assign n39834 = n36883 ^ n36376 ^ n9525 ;
  assign n39835 = n39834 ^ n23778 ^ n18084 ;
  assign n39836 = n5996 ^ x235 ^ 1'b0 ;
  assign n39837 = n39836 ^ n28762 ^ n5791 ;
  assign n39838 = ( n551 & ~n27065 ) | ( n551 & n33463 ) | ( ~n27065 & n33463 ) ;
  assign n39839 = ( ~n26265 & n39837 ) | ( ~n26265 & n39838 ) | ( n39837 & n39838 ) ;
  assign n39840 = ( n24241 & n38881 ) | ( n24241 & n39839 ) | ( n38881 & n39839 ) ;
  assign n39842 = ~n26374 & n37622 ;
  assign n39841 = n15555 ^ n12442 ^ n11408 ;
  assign n39843 = n39842 ^ n39841 ^ n11100 ;
  assign n39844 = ( n4110 & n6028 ) | ( n4110 & ~n6923 ) | ( n6028 & ~n6923 ) ;
  assign n39845 = n39844 ^ n19101 ^ n8042 ;
  assign n39846 = n3732 | n17278 ;
  assign n39847 = n39846 ^ n24845 ^ n1265 ;
  assign n39848 = n16389 ^ n13835 ^ n9737 ;
  assign n39849 = ~n27240 & n39848 ;
  assign n39850 = n39849 ^ n15077 ^ 1'b0 ;
  assign n39851 = n39847 | n39850 ;
  assign n39852 = n33021 ^ n25352 ^ n15879 ;
  assign n39853 = n6731 ^ n5871 ^ 1'b0 ;
  assign n39854 = ( ~n13442 & n39775 ) | ( ~n13442 & n39853 ) | ( n39775 & n39853 ) ;
  assign n39855 = n9624 & n32040 ;
  assign n39856 = n15260 & n18596 ;
  assign n39857 = n39856 ^ n2686 ^ 1'b0 ;
  assign n39858 = n28840 ^ n27330 ^ n17238 ;
  assign n39859 = ~n30365 & n39858 ;
  assign n39860 = n39859 ^ n36068 ^ 1'b0 ;
  assign n39861 = ( ~n10642 & n39857 ) | ( ~n10642 & n39860 ) | ( n39857 & n39860 ) ;
  assign n39862 = ( ~n31812 & n39855 ) | ( ~n31812 & n39861 ) | ( n39855 & n39861 ) ;
  assign n39864 = n25079 ^ n7242 ^ n4487 ;
  assign n39865 = n39864 ^ n24090 ^ n2462 ;
  assign n39863 = n37035 ^ n27636 ^ n22125 ;
  assign n39866 = n39865 ^ n39863 ^ n25886 ;
  assign n39867 = n15469 ^ n1945 ^ 1'b0 ;
  assign n39868 = ( n14919 & ~n27862 ) | ( n14919 & n31475 ) | ( ~n27862 & n31475 ) ;
  assign n39869 = ( n4010 & n16790 ) | ( n4010 & n39868 ) | ( n16790 & n39868 ) ;
  assign n39870 = ( n13892 & ~n27963 ) | ( n13892 & n39869 ) | ( ~n27963 & n39869 ) ;
  assign n39871 = ( ~n1181 & n4120 ) | ( ~n1181 & n29100 ) | ( n4120 & n29100 ) ;
  assign n39872 = n39871 ^ n38636 ^ x193 ;
  assign n39879 = n28236 ^ n25988 ^ n1831 ;
  assign n39880 = ( x51 & n28117 ) | ( x51 & n39879 ) | ( n28117 & n39879 ) ;
  assign n39877 = n30973 ^ n25650 ^ n15264 ;
  assign n39875 = ( n13992 & n15674 ) | ( n13992 & n23073 ) | ( n15674 & n23073 ) ;
  assign n39874 = ( ~n4985 & n5882 ) | ( ~n4985 & n19593 ) | ( n5882 & n19593 ) ;
  assign n39876 = n39875 ^ n39874 ^ n1341 ;
  assign n39878 = n39877 ^ n39876 ^ n38398 ;
  assign n39873 = ( n17359 & n35736 ) | ( n17359 & ~n39725 ) | ( n35736 & ~n39725 ) ;
  assign n39881 = n39880 ^ n39878 ^ n39873 ;
  assign n39882 = ( ~n11689 & n21089 ) | ( ~n11689 & n38991 ) | ( n21089 & n38991 ) ;
  assign n39883 = n1098 | n31839 ;
  assign n39884 = n1332 | n39883 ;
  assign n39885 = n39884 ^ n7343 ^ n4599 ;
  assign n39886 = n39885 ^ n4374 ^ 1'b0 ;
  assign n39887 = n33278 ^ n23534 ^ n19929 ;
  assign n39888 = n39887 ^ n11897 ^ n9939 ;
  assign n39889 = n39888 ^ n34503 ^ n8844 ;
  assign n39890 = ( n23587 & n26388 ) | ( n23587 & n39889 ) | ( n26388 & n39889 ) ;
  assign n39891 = n16443 & ~n39890 ;
  assign n39892 = n15369 ^ n10261 ^ n6211 ;
  assign n39893 = ( n13731 & ~n13893 ) | ( n13731 & n39892 ) | ( ~n13893 & n39892 ) ;
  assign n39894 = n39893 ^ n15799 ^ 1'b0 ;
  assign n39895 = n39891 & ~n39894 ;
  assign n39896 = ( n5064 & n9807 ) | ( n5064 & n39385 ) | ( n9807 & n39385 ) ;
  assign n39897 = n7690 & n29556 ;
  assign n39898 = n39897 ^ n16168 ^ n326 ;
  assign n39899 = ( n4909 & n17181 ) | ( n4909 & ~n39898 ) | ( n17181 & ~n39898 ) ;
  assign n39900 = ( n9509 & n20107 ) | ( n9509 & n20968 ) | ( n20107 & n20968 ) ;
  assign n39901 = ~n5916 & n39900 ;
  assign n39902 = ~n20907 & n39901 ;
  assign n39903 = n30931 | n39902 ;
  assign n39904 = ~n2730 & n12827 ;
  assign n39905 = n39904 ^ n11567 ^ n7407 ;
  assign n39906 = ( ~n6653 & n12521 ) | ( ~n6653 & n38768 ) | ( n12521 & n38768 ) ;
  assign n39907 = ( n6392 & ~n7757 ) | ( n6392 & n16160 ) | ( ~n7757 & n16160 ) ;
  assign n39908 = ( ~n2196 & n15710 ) | ( ~n2196 & n39907 ) | ( n15710 & n39907 ) ;
  assign n39909 = n25611 & ~n39908 ;
  assign n39910 = ( n4052 & ~n39906 ) | ( n4052 & n39909 ) | ( ~n39906 & n39909 ) ;
  assign n39911 = ( n2785 & n31522 ) | ( n2785 & ~n39392 ) | ( n31522 & ~n39392 ) ;
  assign n39912 = n39911 ^ n16248 ^ n14462 ;
  assign n39913 = n30660 ^ n11566 ^ n5224 ;
  assign n39914 = ( n6744 & n7535 ) | ( n6744 & ~n39913 ) | ( n7535 & ~n39913 ) ;
  assign n39915 = n2463 & n17415 ;
  assign n39916 = n28574 & n39915 ;
  assign n39917 = ( n3467 & ~n5636 ) | ( n3467 & n30152 ) | ( ~n5636 & n30152 ) ;
  assign n39918 = ( n5944 & ~n17174 ) | ( n5944 & n39917 ) | ( ~n17174 & n39917 ) ;
  assign n39919 = n11286 & n28815 ;
  assign n39920 = ~n28426 & n39919 ;
  assign n39921 = n39920 ^ n28978 ^ n10024 ;
  assign n39925 = n26702 ^ n10218 ^ 1'b0 ;
  assign n39922 = ~n2167 & n18584 ;
  assign n39923 = n39922 ^ n859 ^ 1'b0 ;
  assign n39924 = n39923 ^ n29153 ^ 1'b0 ;
  assign n39926 = n39925 ^ n39924 ^ n3828 ;
  assign n39927 = n20821 ^ n10534 ^ 1'b0 ;
  assign n39928 = n32990 ^ n10565 ^ 1'b0 ;
  assign n39929 = n18483 ^ n9813 ^ n6468 ;
  assign n39930 = ( n11425 & ~n14946 ) | ( n11425 & n39929 ) | ( ~n14946 & n39929 ) ;
  assign n39931 = n28866 ^ n23692 ^ n14950 ;
  assign n39932 = n37660 ^ n32672 ^ n17653 ;
  assign n39933 = n25713 ^ n24226 ^ n22263 ;
  assign n39934 = n39933 ^ n18663 ^ 1'b0 ;
  assign n39935 = ( n24378 & ~n39932 ) | ( n24378 & n39934 ) | ( ~n39932 & n39934 ) ;
  assign n39938 = n21382 ^ n6117 ^ n2451 ;
  assign n39937 = n28373 ^ n20859 ^ n7238 ;
  assign n39936 = n29196 ^ n26846 ^ n25745 ;
  assign n39939 = n39938 ^ n39937 ^ n39936 ;
  assign n39940 = n8488 ^ n5297 ^ 1'b0 ;
  assign n39941 = n7483 & ~n12836 ;
  assign n39942 = ( n11657 & ~n12913 ) | ( n11657 & n22494 ) | ( ~n12913 & n22494 ) ;
  assign n39943 = n32984 & n39942 ;
  assign n39944 = ~n36338 & n39943 ;
  assign n39945 = n11616 ^ n10334 ^ n2129 ;
  assign n39946 = n39945 ^ n30370 ^ n14692 ;
  assign n39947 = n17145 ^ n14867 ^ n1406 ;
  assign n39948 = ( ~n13253 & n16245 ) | ( ~n13253 & n21640 ) | ( n16245 & n21640 ) ;
  assign n39949 = n13783 & ~n39948 ;
  assign n39950 = ( n6025 & n39947 ) | ( n6025 & n39949 ) | ( n39947 & n39949 ) ;
  assign n39951 = ( n2871 & ~n17770 ) | ( n2871 & n39844 ) | ( ~n17770 & n39844 ) ;
  assign n39952 = n12938 ^ n9128 ^ 1'b0 ;
  assign n39953 = n39952 ^ n17504 ^ n4608 ;
  assign n39954 = ( n10156 & ~n10745 ) | ( n10156 & n18871 ) | ( ~n10745 & n18871 ) ;
  assign n39955 = ( n935 & n14767 ) | ( n935 & n26150 ) | ( n14767 & n26150 ) ;
  assign n39956 = ( n2127 & n39954 ) | ( n2127 & n39955 ) | ( n39954 & n39955 ) ;
  assign n39957 = n9679 & n11796 ;
  assign n39958 = ( n7862 & n15503 ) | ( n7862 & ~n17742 ) | ( n15503 & ~n17742 ) ;
  assign n39959 = ( n28466 & n39957 ) | ( n28466 & ~n39958 ) | ( n39957 & ~n39958 ) ;
  assign n39960 = n21592 ^ n10290 ^ n403 ;
  assign n39961 = n39960 ^ n36331 ^ n8290 ;
  assign n39962 = n8014 ^ n7483 ^ 1'b0 ;
  assign n39963 = ( ~n21897 & n30160 ) | ( ~n21897 & n39962 ) | ( n30160 & n39962 ) ;
  assign n39967 = n24994 ^ n16939 ^ n14441 ;
  assign n39964 = n4423 | n20236 ;
  assign n39965 = n39964 ^ n28218 ^ 1'b0 ;
  assign n39966 = ( ~n2198 & n4347 ) | ( ~n2198 & n39965 ) | ( n4347 & n39965 ) ;
  assign n39968 = n39967 ^ n39966 ^ n3986 ;
  assign n39969 = ( ~n12781 & n14779 ) | ( ~n12781 & n18181 ) | ( n14779 & n18181 ) ;
  assign n39970 = n26970 ^ n18304 ^ 1'b0 ;
  assign n39971 = ( n5949 & n39969 ) | ( n5949 & ~n39970 ) | ( n39969 & ~n39970 ) ;
  assign n39972 = ( n10411 & n19200 ) | ( n10411 & ~n32335 ) | ( n19200 & ~n32335 ) ;
  assign n39973 = ( n2586 & ~n27161 ) | ( n2586 & n39972 ) | ( ~n27161 & n39972 ) ;
  assign n39974 = n7294 ^ n6921 ^ n5840 ;
  assign n39975 = ( n24060 & n35727 ) | ( n24060 & n39974 ) | ( n35727 & n39974 ) ;
  assign n39978 = ( ~n2714 & n7876 ) | ( ~n2714 & n14239 ) | ( n7876 & n14239 ) ;
  assign n39979 = ( n17355 & n20534 ) | ( n17355 & ~n39978 ) | ( n20534 & ~n39978 ) ;
  assign n39976 = n13694 ^ n8765 ^ n5743 ;
  assign n39977 = ( n23767 & n34301 ) | ( n23767 & ~n39976 ) | ( n34301 & ~n39976 ) ;
  assign n39980 = n39979 ^ n39977 ^ n30217 ;
  assign n39981 = ( n22909 & n31440 ) | ( n22909 & n34997 ) | ( n31440 & n34997 ) ;
  assign n39982 = n35431 ^ n26351 ^ n13068 ;
  assign n39983 = n21824 ^ n6921 ^ n4909 ;
  assign n39984 = ~n11096 & n39983 ;
  assign n39985 = ~n7312 & n39984 ;
  assign n39986 = ( n2373 & n10674 ) | ( n2373 & ~n10934 ) | ( n10674 & ~n10934 ) ;
  assign n39987 = n39986 ^ n38910 ^ n27827 ;
  assign n39988 = ( n3755 & ~n6347 ) | ( n3755 & n39987 ) | ( ~n6347 & n39987 ) ;
  assign n39989 = ( n2932 & n13987 ) | ( n2932 & ~n20843 ) | ( n13987 & ~n20843 ) ;
  assign n39990 = ( n17659 & n24640 ) | ( n17659 & ~n39989 ) | ( n24640 & ~n39989 ) ;
  assign n39991 = ( n4917 & n13779 ) | ( n4917 & n34287 ) | ( n13779 & n34287 ) ;
  assign n39992 = ( ~n6911 & n34183 ) | ( ~n6911 & n39991 ) | ( n34183 & n39991 ) ;
  assign n39993 = n28537 ^ n12325 ^ n7989 ;
  assign n39994 = n24839 ^ n22678 ^ n21166 ;
  assign n39995 = n39994 ^ n20907 ^ 1'b0 ;
  assign n39996 = n39995 ^ n10855 ^ 1'b0 ;
  assign n39997 = n26217 | n39996 ;
  assign n39998 = ( n2351 & n8655 ) | ( n2351 & ~n39997 ) | ( n8655 & ~n39997 ) ;
  assign n40001 = n17307 ^ n10544 ^ n4324 ;
  assign n40002 = ( ~n1597 & n23805 ) | ( ~n1597 & n40001 ) | ( n23805 & n40001 ) ;
  assign n40003 = n40002 ^ n30603 ^ n15648 ;
  assign n39999 = ( n2913 & ~n7132 ) | ( n2913 & n22503 ) | ( ~n7132 & n22503 ) ;
  assign n40000 = n39999 ^ n23258 ^ 1'b0 ;
  assign n40004 = n40003 ^ n40000 ^ n15794 ;
  assign n40005 = n40004 ^ n39127 ^ n24803 ;
  assign n40006 = n40005 ^ n30169 ^ n6703 ;
  assign n40007 = n21619 ^ n7911 ^ 1'b0 ;
  assign n40008 = n40007 ^ n13182 ^ n11233 ;
  assign n40009 = ( n2609 & n25885 ) | ( n2609 & ~n40008 ) | ( n25885 & ~n40008 ) ;
  assign n40010 = ( n24885 & n35372 ) | ( n24885 & n40009 ) | ( n35372 & n40009 ) ;
  assign n40011 = n1881 ^ n1779 ^ x56 ;
  assign n40012 = n14195 & ~n40011 ;
  assign n40013 = n40012 ^ n2388 ^ 1'b0 ;
  assign n40014 = n40013 ^ n15785 ^ 1'b0 ;
  assign n40015 = ~n16330 & n40014 ;
  assign n40016 = n32258 ^ n30863 ^ n865 ;
  assign n40018 = ~n1284 & n25888 ;
  assign n40019 = n13788 & n40018 ;
  assign n40017 = n10884 ^ n1333 ^ x71 ;
  assign n40020 = n40019 ^ n40017 ^ n17850 ;
  assign n40021 = ( n18931 & ~n30547 ) | ( n18931 & n40020 ) | ( ~n30547 & n40020 ) ;
  assign n40022 = ( n19834 & n26327 ) | ( n19834 & n38449 ) | ( n26327 & n38449 ) ;
  assign n40023 = n39693 ^ n23089 ^ n6969 ;
  assign n40024 = ( ~n7267 & n40022 ) | ( ~n7267 & n40023 ) | ( n40022 & n40023 ) ;
  assign n40025 = n40024 ^ n26767 ^ n10767 ;
  assign n40026 = n34617 ^ n18674 ^ n471 ;
  assign n40027 = n27238 ^ n2074 ^ 1'b0 ;
  assign n40028 = ( ~n26051 & n40026 ) | ( ~n26051 & n40027 ) | ( n40026 & n40027 ) ;
  assign n40029 = n40028 ^ n14209 ^ n1473 ;
  assign n40030 = n39815 ^ n9697 ^ n969 ;
  assign n40031 = n40030 ^ n17121 ^ n6097 ;
  assign n40032 = ~n7921 & n16831 ;
  assign n40033 = n40032 ^ n19047 ^ 1'b0 ;
  assign n40034 = ( n4373 & ~n20524 ) | ( n4373 & n39150 ) | ( ~n20524 & n39150 ) ;
  assign n40035 = n36245 ^ n24317 ^ n3118 ;
  assign n40036 = ( ~n7281 & n12771 ) | ( ~n7281 & n40035 ) | ( n12771 & n40035 ) ;
  assign n40037 = ( n1473 & n22953 ) | ( n1473 & n24979 ) | ( n22953 & n24979 ) ;
  assign n40038 = n40037 ^ n33604 ^ n8827 ;
  assign n40039 = ( n15296 & ~n28338 ) | ( n15296 & n40038 ) | ( ~n28338 & n40038 ) ;
  assign n40045 = n36315 ^ n707 ^ 1'b0 ;
  assign n40043 = ( n7404 & ~n12969 ) | ( n7404 & n14196 ) | ( ~n12969 & n14196 ) ;
  assign n40044 = n3090 & ~n40043 ;
  assign n40040 = n1634 | n33356 ;
  assign n40041 = n37261 | n40040 ;
  assign n40042 = ( ~n10485 & n34330 ) | ( ~n10485 & n40041 ) | ( n34330 & n40041 ) ;
  assign n40046 = n40045 ^ n40044 ^ n40042 ;
  assign n40047 = ( n1893 & ~n8299 ) | ( n1893 & n13713 ) | ( ~n8299 & n13713 ) ;
  assign n40048 = ( ~n8671 & n9200 ) | ( ~n8671 & n40047 ) | ( n9200 & n40047 ) ;
  assign n40049 = n37690 ^ n22671 ^ n7188 ;
  assign n40050 = n40049 ^ n24426 ^ n14271 ;
  assign n40051 = n40050 ^ n8254 ^ 1'b0 ;
  assign n40052 = n7064 ^ n4242 ^ n473 ;
  assign n40053 = n40052 ^ n39152 ^ n13820 ;
  assign n40054 = ( n14452 & ~n19194 ) | ( n14452 & n25082 ) | ( ~n19194 & n25082 ) ;
  assign n40055 = n33605 ^ n14628 ^ 1'b0 ;
  assign n40056 = n13702 & ~n40055 ;
  assign n40057 = n40056 ^ n31935 ^ 1'b0 ;
  assign n40061 = n37634 ^ n9601 ^ 1'b0 ;
  assign n40059 = n33329 | n33759 ;
  assign n40060 = n40059 ^ n13400 ^ n7957 ;
  assign n40058 = ( ~n6055 & n8413 ) | ( ~n6055 & n16821 ) | ( n8413 & n16821 ) ;
  assign n40062 = n40061 ^ n40060 ^ n40058 ;
  assign n40063 = ( ~n1374 & n1500 ) | ( ~n1374 & n37717 ) | ( n1500 & n37717 ) ;
  assign n40066 = n25839 ^ n1563 ^ 1'b0 ;
  assign n40067 = n40066 ^ n27568 ^ n16048 ;
  assign n40065 = x33 & n6922 ;
  assign n40068 = n40067 ^ n40065 ^ 1'b0 ;
  assign n40069 = n1459 | n40068 ;
  assign n40064 = ~x189 & n23874 ;
  assign n40070 = n40069 ^ n40064 ^ n781 ;
  assign n40072 = n16008 ^ n13122 ^ n12337 ;
  assign n40071 = n30875 ^ n15350 ^ n10150 ;
  assign n40073 = n40072 ^ n40071 ^ n9888 ;
  assign n40074 = n25309 ^ n9736 ^ n1939 ;
  assign n40075 = ( n20080 & ~n25109 ) | ( n20080 & n40074 ) | ( ~n25109 & n40074 ) ;
  assign n40077 = n20928 ^ n19753 ^ n6169 ;
  assign n40076 = ( x205 & n15346 ) | ( x205 & ~n19975 ) | ( n15346 & ~n19975 ) ;
  assign n40078 = n40077 ^ n40076 ^ n28619 ;
  assign n40079 = n37051 ^ n20177 ^ n10341 ;
  assign n40080 = n37486 ^ n13290 ^ 1'b0 ;
  assign n40081 = n2892 & n40080 ;
  assign n40082 = ( n21288 & n33404 ) | ( n21288 & n40081 ) | ( n33404 & n40081 ) ;
  assign n40083 = n39986 ^ n33518 ^ 1'b0 ;
  assign n40084 = ( n1033 & n8903 ) | ( n1033 & ~n17510 ) | ( n8903 & ~n17510 ) ;
  assign n40085 = ~n17916 & n39711 ;
  assign n40086 = ~n40084 & n40085 ;
  assign n40087 = ( ~n29109 & n40083 ) | ( ~n29109 & n40086 ) | ( n40083 & n40086 ) ;
  assign n40088 = n24435 ^ n12305 ^ n12085 ;
  assign n40089 = n40088 ^ n30627 ^ n30265 ;
  assign n40090 = n21595 ^ n16885 ^ n3461 ;
  assign n40091 = n20684 ^ n9786 ^ n4091 ;
  assign n40092 = ( ~n10168 & n12029 ) | ( ~n10168 & n24675 ) | ( n12029 & n24675 ) ;
  assign n40093 = ( n14114 & ~n21066 ) | ( n14114 & n40092 ) | ( ~n21066 & n40092 ) ;
  assign n40094 = n40093 ^ n37459 ^ n3785 ;
  assign n40095 = n40094 ^ n34807 ^ n27860 ;
  assign n40099 = n17519 ^ n12648 ^ n6348 ;
  assign n40100 = n7956 & ~n40099 ;
  assign n40101 = ~n14584 & n40100 ;
  assign n40102 = ( x15 & n30102 ) | ( x15 & n35458 ) | ( n30102 & n35458 ) ;
  assign n40103 = ( n5601 & ~n7668 ) | ( n5601 & n40102 ) | ( ~n7668 & n40102 ) ;
  assign n40104 = ~n40101 & n40103 ;
  assign n40105 = n40104 ^ n6628 ^ 1'b0 ;
  assign n40106 = ( n25311 & n33061 ) | ( n25311 & ~n40105 ) | ( n33061 & ~n40105 ) ;
  assign n40096 = n36404 ^ n5886 ^ 1'b0 ;
  assign n40097 = n19643 | n40096 ;
  assign n40098 = ( n7814 & n19412 ) | ( n7814 & n40097 ) | ( n19412 & n40097 ) ;
  assign n40107 = n40106 ^ n40098 ^ n20026 ;
  assign n40110 = n21238 ^ n14070 ^ n9218 ;
  assign n40108 = n27912 ^ n19996 ^ n10896 ;
  assign n40109 = n32348 & ~n40108 ;
  assign n40111 = n40110 ^ n40109 ^ 1'b0 ;
  assign n40112 = n8618 & ~n27668 ;
  assign n40113 = n5087 ^ n4428 ^ n1712 ;
  assign n40114 = ( n6143 & n8918 ) | ( n6143 & ~n32741 ) | ( n8918 & ~n32741 ) ;
  assign n40115 = n22190 & ~n40114 ;
  assign n40116 = n40115 ^ n10853 ^ 1'b0 ;
  assign n40117 = n40116 ^ n20302 ^ n2652 ;
  assign n40118 = ~n40113 & n40117 ;
  assign n40119 = ( n386 & ~n8140 ) | ( n386 & n10670 ) | ( ~n8140 & n10670 ) ;
  assign n40120 = ( n2411 & n4740 ) | ( n2411 & n8876 ) | ( n4740 & n8876 ) ;
  assign n40121 = n40120 ^ n17296 ^ 1'b0 ;
  assign n40122 = n40119 | n40121 ;
  assign n40123 = ( ~n14664 & n17019 ) | ( ~n14664 & n40122 ) | ( n17019 & n40122 ) ;
  assign n40124 = ~n19372 & n24086 ;
  assign n40125 = n21415 & n32755 ;
  assign n40126 = n40125 ^ n25051 ^ 1'b0 ;
  assign n40127 = ( n11770 & n13270 ) | ( n11770 & ~n39779 ) | ( n13270 & ~n39779 ) ;
  assign n40128 = n40127 ^ n38674 ^ 1'b0 ;
  assign n40129 = n7902 & ~n40128 ;
  assign n40130 = n39190 & n40129 ;
  assign n40137 = ( n2016 & n2705 ) | ( n2016 & ~n27221 ) | ( n2705 & ~n27221 ) ;
  assign n40138 = ( n20022 & n38561 ) | ( n20022 & n40137 ) | ( n38561 & n40137 ) ;
  assign n40133 = ( n3263 & n16227 ) | ( n3263 & ~n30998 ) | ( n16227 & ~n30998 ) ;
  assign n40134 = ( n3770 & n14561 ) | ( n3770 & ~n40133 ) | ( n14561 & ~n40133 ) ;
  assign n40135 = n40134 ^ n12385 ^ n1937 ;
  assign n40131 = n21691 ^ n19534 ^ 1'b0 ;
  assign n40132 = n23435 | n40131 ;
  assign n40136 = n40135 ^ n40132 ^ 1'b0 ;
  assign n40139 = n40138 ^ n40136 ^ n4459 ;
  assign n40140 = n28000 ^ n25942 ^ n13077 ;
  assign n40143 = n37614 ^ n27403 ^ n26796 ;
  assign n40141 = n18961 ^ n13017 ^ n6754 ;
  assign n40142 = ( ~n13309 & n19532 ) | ( ~n13309 & n40141 ) | ( n19532 & n40141 ) ;
  assign n40144 = n40143 ^ n40142 ^ n18001 ;
  assign n40145 = ( n13996 & n20869 ) | ( n13996 & ~n40144 ) | ( n20869 & ~n40144 ) ;
  assign n40146 = ( n24273 & n40140 ) | ( n24273 & n40145 ) | ( n40140 & n40145 ) ;
  assign n40147 = n27292 ^ n22940 ^ n5232 ;
  assign n40148 = ( n26923 & ~n37752 ) | ( n26923 & n40147 ) | ( ~n37752 & n40147 ) ;
  assign n40149 = n40148 ^ n38262 ^ 1'b0 ;
  assign n40150 = n37355 & ~n40149 ;
  assign n40151 = ( n6921 & n27669 ) | ( n6921 & ~n29525 ) | ( n27669 & ~n29525 ) ;
  assign n40152 = ( n30917 & n39994 ) | ( n30917 & n40151 ) | ( n39994 & n40151 ) ;
  assign n40153 = n19608 ^ n13886 ^ 1'b0 ;
  assign n40154 = n3383 & ~n40153 ;
  assign n40155 = n16282 ^ n10530 ^ 1'b0 ;
  assign n40156 = n40154 & n40155 ;
  assign n40157 = n34094 ^ n24489 ^ n741 ;
  assign n40161 = ( n5427 & ~n5633 ) | ( n5427 & n7423 ) | ( ~n5633 & n7423 ) ;
  assign n40162 = n40161 ^ n17799 ^ n11736 ;
  assign n40163 = ( ~n18727 & n22975 ) | ( ~n18727 & n40162 ) | ( n22975 & n40162 ) ;
  assign n40160 = n7459 | n12539 ;
  assign n40164 = n40163 ^ n40160 ^ 1'b0 ;
  assign n40158 = ( n6711 & n18500 ) | ( n6711 & ~n25828 ) | ( n18500 & ~n25828 ) ;
  assign n40159 = ( n10579 & n18175 ) | ( n10579 & n40158 ) | ( n18175 & n40158 ) ;
  assign n40165 = n40164 ^ n40159 ^ n28841 ;
  assign n40166 = n38123 ^ n29123 ^ n23984 ;
  assign n40167 = ( n7352 & n10130 ) | ( n7352 & ~n24448 ) | ( n10130 & ~n24448 ) ;
  assign n40168 = n21535 ^ n4391 ^ 1'b0 ;
  assign n40169 = ~n9458 & n40168 ;
  assign n40170 = n40169 ^ n26113 ^ n13065 ;
  assign n40171 = ( ~n2744 & n24624 ) | ( ~n2744 & n40170 ) | ( n24624 & n40170 ) ;
  assign n40172 = ( ~n3687 & n7565 ) | ( ~n3687 & n8006 ) | ( n7565 & n8006 ) ;
  assign n40173 = ( ~n9930 & n19023 ) | ( ~n9930 & n40172 ) | ( n19023 & n40172 ) ;
  assign n40179 = n19063 ^ n16245 ^ n7027 ;
  assign n40175 = n24881 ^ n2689 ^ n2569 ;
  assign n40174 = ( n4529 & n9404 ) | ( n4529 & n16574 ) | ( n9404 & n16574 ) ;
  assign n40176 = n40175 ^ n40174 ^ n8669 ;
  assign n40177 = ( n7625 & n38869 ) | ( n7625 & n40176 ) | ( n38869 & n40176 ) ;
  assign n40178 = n40177 ^ n22073 ^ n1150 ;
  assign n40180 = n40179 ^ n40178 ^ 1'b0 ;
  assign n40185 = n16198 ^ n6218 ^ n5149 ;
  assign n40186 = ( n7672 & n30092 ) | ( n7672 & n40185 ) | ( n30092 & n40185 ) ;
  assign n40183 = n30604 ^ n14991 ^ 1'b0 ;
  assign n40184 = n35386 & ~n40183 ;
  assign n40187 = n40186 ^ n40184 ^ 1'b0 ;
  assign n40181 = n27731 ^ n15911 ^ n13532 ;
  assign n40182 = ~n3332 & n40181 ;
  assign n40188 = n40187 ^ n40182 ^ 1'b0 ;
  assign n40189 = n11528 ^ n8805 ^ n6676 ;
  assign n40190 = n1464 & n14760 ;
  assign n40191 = n40190 ^ n1047 ^ 1'b0 ;
  assign n40192 = ( n37253 & n40189 ) | ( n37253 & ~n40191 ) | ( n40189 & ~n40191 ) ;
  assign n40193 = n40120 ^ n12978 ^ n9762 ;
  assign n40195 = ( n16346 & n20656 ) | ( n16346 & ~n38869 ) | ( n20656 & ~n38869 ) ;
  assign n40196 = ( n1415 & ~n16333 ) | ( n1415 & n40195 ) | ( ~n16333 & n40195 ) ;
  assign n40194 = ~n4109 & n22085 ;
  assign n40197 = n40196 ^ n40194 ^ 1'b0 ;
  assign n40198 = n27073 ^ n9608 ^ n9078 ;
  assign n40199 = ( n12884 & ~n27452 ) | ( n12884 & n40198 ) | ( ~n27452 & n40198 ) ;
  assign n40200 = ( ~n10011 & n17128 ) | ( ~n10011 & n40199 ) | ( n17128 & n40199 ) ;
  assign n40201 = ( n11137 & ~n25595 ) | ( n11137 & n35289 ) | ( ~n25595 & n35289 ) ;
  assign n40203 = n11919 ^ n11801 ^ n7055 ;
  assign n40202 = n13382 & n13813 ;
  assign n40204 = n40203 ^ n40202 ^ 1'b0 ;
  assign n40205 = ( n6152 & ~n6302 ) | ( n6152 & n17443 ) | ( ~n6302 & n17443 ) ;
  assign n40206 = n22827 ^ n12369 ^ n5443 ;
  assign n40207 = n34889 ^ n14611 ^ 1'b0 ;
  assign n40208 = ( n25464 & n31318 ) | ( n25464 & n40207 ) | ( n31318 & n40207 ) ;
  assign n40209 = ( ~n1762 & n11831 ) | ( ~n1762 & n31830 ) | ( n11831 & n31830 ) ;
  assign n40210 = n40209 ^ n26724 ^ n6768 ;
  assign n40211 = ( ~n4905 & n28849 ) | ( ~n4905 & n37490 ) | ( n28849 & n37490 ) ;
  assign n40212 = ( n12941 & n20220 ) | ( n12941 & ~n20575 ) | ( n20220 & ~n20575 ) ;
  assign n40213 = ( n9061 & n20105 ) | ( n9061 & n40212 ) | ( n20105 & n40212 ) ;
  assign n40214 = n10891 ^ n8950 ^ n2921 ;
  assign n40215 = n40214 ^ n18479 ^ n10076 ;
  assign n40216 = ( n5914 & n18343 ) | ( n5914 & ~n40215 ) | ( n18343 & ~n40215 ) ;
  assign n40217 = ~n12080 & n14705 ;
  assign n40218 = n40217 ^ n1343 ^ 1'b0 ;
  assign n40219 = ( n11407 & n21062 ) | ( n11407 & ~n40218 ) | ( n21062 & ~n40218 ) ;
  assign n40220 = ( n7537 & n16134 ) | ( n7537 & n40219 ) | ( n16134 & n40219 ) ;
  assign n40221 = ~n30237 & n32925 ;
  assign n40222 = n40221 ^ n39631 ^ 1'b0 ;
  assign n40223 = ( n14885 & n21053 ) | ( n14885 & n38101 ) | ( n21053 & n38101 ) ;
  assign n40224 = n31719 ^ n28280 ^ 1'b0 ;
  assign n40225 = n8834 | n35860 ;
  assign n40226 = n40225 ^ n6810 ^ 1'b0 ;
  assign n40227 = n40226 ^ n12444 ^ n9234 ;
  assign n40228 = ( n1315 & n3941 ) | ( n1315 & ~n40227 ) | ( n3941 & ~n40227 ) ;
  assign n40229 = ( n3720 & n40224 ) | ( n3720 & n40228 ) | ( n40224 & n40228 ) ;
  assign n40230 = ( ~n343 & n6985 ) | ( ~n343 & n11498 ) | ( n6985 & n11498 ) ;
  assign n40231 = n40230 ^ n23112 ^ n21697 ;
  assign n40232 = ( n4801 & n34667 ) | ( n4801 & n40231 ) | ( n34667 & n40231 ) ;
  assign n40233 = ( n37529 & n39156 ) | ( n37529 & ~n40232 ) | ( n39156 & ~n40232 ) ;
  assign n40234 = n4638 ^ n3886 ^ n2034 ;
  assign n40235 = n40234 ^ n17853 ^ n1839 ;
  assign n40236 = ( n23874 & ~n26248 ) | ( n23874 & n40235 ) | ( ~n26248 & n40235 ) ;
  assign n40237 = n40236 ^ n31466 ^ n16975 ;
  assign n40238 = n32530 ^ n25699 ^ n10935 ;
  assign n40239 = ( ~n17899 & n20990 ) | ( ~n17899 & n40238 ) | ( n20990 & n40238 ) ;
  assign n40240 = n40239 ^ n17247 ^ n8480 ;
  assign n40241 = n38289 ^ n30844 ^ n23007 ;
  assign n40242 = n26210 ^ n24627 ^ n20094 ;
  assign n40243 = n40242 ^ n10294 ^ n9357 ;
  assign n40244 = n40243 ^ n34187 ^ n30911 ;
  assign n40245 = n7044 ^ n2849 ^ n2691 ;
  assign n40251 = n31264 ^ n23073 ^ n15862 ;
  assign n40248 = x52 & n11611 ;
  assign n40249 = ~n14492 & n40248 ;
  assign n40246 = n3024 | n32494 ;
  assign n40247 = n40246 ^ n24675 ^ 1'b0 ;
  assign n40250 = n40249 ^ n40247 ^ n25092 ;
  assign n40252 = n40251 ^ n40250 ^ n39122 ;
  assign n40253 = n38526 | n40252 ;
  assign n40254 = n40245 | n40253 ;
  assign n40255 = ( ~n674 & n1846 ) | ( ~n674 & n8734 ) | ( n1846 & n8734 ) ;
  assign n40256 = ~n7732 & n40255 ;
  assign n40257 = n11785 & n40256 ;
  assign n40258 = ( ~n685 & n14591 ) | ( ~n685 & n15792 ) | ( n14591 & n15792 ) ;
  assign n40259 = n7479 & ~n21432 ;
  assign n40260 = ( n8017 & n18097 ) | ( n8017 & ~n40259 ) | ( n18097 & ~n40259 ) ;
  assign n40261 = ( ~n13799 & n13919 ) | ( ~n13799 & n37851 ) | ( n13919 & n37851 ) ;
  assign n40262 = ( n6549 & n21033 ) | ( n6549 & n40261 ) | ( n21033 & n40261 ) ;
  assign n40263 = n7711 ^ n3169 ^ n482 ;
  assign n40264 = ( n5811 & n11580 ) | ( n5811 & n40263 ) | ( n11580 & n40263 ) ;
  assign n40265 = n8049 ^ n2256 ^ 1'b0 ;
  assign n40266 = n37518 & n40265 ;
  assign n40267 = ( ~n31596 & n40264 ) | ( ~n31596 & n40266 ) | ( n40264 & n40266 ) ;
  assign n40268 = n23626 ^ n18445 ^ n4390 ;
  assign n40269 = n32447 & n35417 ;
  assign n40270 = n40269 ^ n9864 ^ 1'b0 ;
  assign n40271 = ( ~n2249 & n8234 ) | ( ~n2249 & n40270 ) | ( n8234 & n40270 ) ;
  assign n40272 = n40271 ^ n9397 ^ n4751 ;
  assign n40273 = n9712 ^ n9000 ^ n1691 ;
  assign n40274 = n40273 ^ n28315 ^ n1577 ;
  assign n40275 = n40274 ^ n11308 ^ n6801 ;
  assign n40276 = n6080 ^ n5418 ^ n3724 ;
  assign n40277 = n40276 ^ n38122 ^ n4767 ;
  assign n40278 = n40277 ^ n18211 ^ n625 ;
  assign n40279 = ( n7653 & n35307 ) | ( n7653 & n40278 ) | ( n35307 & n40278 ) ;
  assign n40280 = ( n13035 & n14176 ) | ( n13035 & n20082 ) | ( n14176 & n20082 ) ;
  assign n40281 = n27672 ^ n17061 ^ n14019 ;
  assign n40282 = n14820 ^ n11137 ^ n3866 ;
  assign n40283 = ( ~n14025 & n17585 ) | ( ~n14025 & n40282 ) | ( n17585 & n40282 ) ;
  assign n40284 = n15631 ^ n4310 ^ n1279 ;
  assign n40285 = ( n3559 & n10499 ) | ( n3559 & ~n11591 ) | ( n10499 & ~n11591 ) ;
  assign n40286 = n40285 ^ n35052 ^ n12176 ;
  assign n40287 = ~n8403 & n40286 ;
  assign n40288 = n36378 & n40287 ;
  assign n40289 = ( n6240 & n28970 ) | ( n6240 & n37456 ) | ( n28970 & n37456 ) ;
  assign n40290 = n23932 ^ n15762 ^ n13493 ;
  assign n40291 = ( n21255 & ~n27788 ) | ( n21255 & n35228 ) | ( ~n27788 & n35228 ) ;
  assign n40292 = n40291 ^ n37474 ^ n9905 ;
  assign n40293 = ( n2647 & n40290 ) | ( n2647 & n40292 ) | ( n40290 & n40292 ) ;
  assign n40294 = n40293 ^ n18129 ^ n6864 ;
  assign n40295 = ( n8737 & n17000 ) | ( n8737 & n24640 ) | ( n17000 & n24640 ) ;
  assign n40296 = n40295 ^ n27639 ^ n24954 ;
  assign n40297 = ( n2122 & ~n2214 ) | ( n2122 & n40296 ) | ( ~n2214 & n40296 ) ;
  assign n40298 = ( ~n26792 & n31448 ) | ( ~n26792 & n33527 ) | ( n31448 & n33527 ) ;
  assign n40299 = ( ~n6847 & n23896 ) | ( ~n6847 & n30999 ) | ( n23896 & n30999 ) ;
  assign n40300 = ( n7293 & n21345 ) | ( n7293 & n25652 ) | ( n21345 & n25652 ) ;
  assign n40301 = n40300 ^ n30694 ^ n2036 ;
  assign n40302 = ~n29143 & n39183 ;
  assign n40303 = ~n3584 & n40302 ;
  assign n40304 = ( n2921 & n13424 ) | ( n2921 & n17373 ) | ( n13424 & n17373 ) ;
  assign n40305 = ( n4233 & n5539 ) | ( n4233 & ~n40304 ) | ( n5539 & ~n40304 ) ;
  assign n40306 = ( n9538 & n38508 ) | ( n9538 & ~n40305 ) | ( n38508 & ~n40305 ) ;
  assign n40307 = n18344 ^ n4475 ^ 1'b0 ;
  assign n40308 = ~n2013 & n40307 ;
  assign n40309 = n40308 ^ n20845 ^ n2236 ;
  assign n40310 = n40309 ^ n39443 ^ n18975 ;
  assign n40311 = ( ~n1814 & n14249 ) | ( ~n1814 & n21242 ) | ( n14249 & n21242 ) ;
  assign n40312 = ( ~n13466 & n21071 ) | ( ~n13466 & n26689 ) | ( n21071 & n26689 ) ;
  assign n40313 = n40311 | n40312 ;
  assign n40314 = n40310 | n40313 ;
  assign n40315 = ( n28239 & ~n40306 ) | ( n28239 & n40314 ) | ( ~n40306 & n40314 ) ;
  assign n40317 = n19473 | n27266 ;
  assign n40318 = n40317 ^ n33499 ^ 1'b0 ;
  assign n40316 = n20984 | n27615 ;
  assign n40319 = n40318 ^ n40316 ^ 1'b0 ;
  assign n40320 = ( ~n18597 & n38687 ) | ( ~n18597 & n40319 ) | ( n38687 & n40319 ) ;
  assign n40321 = n2286 & ~n38673 ;
  assign n40322 = n16310 & n40321 ;
  assign n40323 = n35709 ^ n32840 ^ n15313 ;
  assign n40324 = n29544 & n36093 ;
  assign n40325 = ( n8567 & n13096 ) | ( n8567 & ~n33926 ) | ( n13096 & ~n33926 ) ;
  assign n40326 = n40325 ^ n23651 ^ n10607 ;
  assign n40331 = n31037 ^ n20923 ^ 1'b0 ;
  assign n40332 = n8920 | n40331 ;
  assign n40333 = n2041 & ~n40332 ;
  assign n40330 = n32597 ^ n7408 ^ n4177 ;
  assign n40327 = n12102 ^ n7999 ^ n6548 ;
  assign n40328 = n22992 ^ n17672 ^ n9337 ;
  assign n40329 = ( ~n33908 & n40327 ) | ( ~n33908 & n40328 ) | ( n40327 & n40328 ) ;
  assign n40334 = n40333 ^ n40330 ^ n40329 ;
  assign n40335 = n9744 & n40334 ;
  assign n40336 = ( ~n16360 & n40326 ) | ( ~n16360 & n40335 ) | ( n40326 & n40335 ) ;
  assign n40337 = ( ~n355 & n3851 ) | ( ~n355 & n4718 ) | ( n3851 & n4718 ) ;
  assign n40338 = ( ~n1940 & n18988 ) | ( ~n1940 & n24091 ) | ( n18988 & n24091 ) ;
  assign n40339 = ( n31307 & n40337 ) | ( n31307 & ~n40338 ) | ( n40337 & ~n40338 ) ;
  assign n40340 = n12696 ^ n1094 ^ 1'b0 ;
  assign n40341 = ~n35054 & n40340 ;
  assign n40342 = ( ~n3168 & n36553 ) | ( ~n3168 & n40341 ) | ( n36553 & n40341 ) ;
  assign n40343 = ( ~n6718 & n11912 ) | ( ~n6718 & n12797 ) | ( n11912 & n12797 ) ;
  assign n40344 = n40343 ^ n24620 ^ n6767 ;
  assign n40345 = n8508 ^ n7544 ^ n4481 ;
  assign n40346 = n15738 ^ n4031 ^ n3384 ;
  assign n40347 = n38533 ^ n26830 ^ 1'b0 ;
  assign n40348 = n25796 | n40347 ;
  assign n40349 = n12761 & ~n40348 ;
  assign n40350 = ( n7721 & ~n16131 ) | ( n7721 & n40349 ) | ( ~n16131 & n40349 ) ;
  assign n40351 = ( ~n11853 & n14711 ) | ( ~n11853 & n19243 ) | ( n14711 & n19243 ) ;
  assign n40352 = n5925 & n40351 ;
  assign n40353 = ( n2468 & n4659 ) | ( n2468 & n10541 ) | ( n4659 & n10541 ) ;
  assign n40354 = ~n13404 & n40353 ;
  assign n40355 = ~n31681 & n40354 ;
  assign n40356 = ( n3322 & n16457 ) | ( n3322 & ~n21079 ) | ( n16457 & ~n21079 ) ;
  assign n40357 = ( n3408 & n5328 ) | ( n3408 & ~n40356 ) | ( n5328 & ~n40356 ) ;
  assign n40358 = n21040 ^ n9747 ^ n1805 ;
  assign n40359 = ( x109 & n18068 ) | ( x109 & n40358 ) | ( n18068 & n40358 ) ;
  assign n40360 = n37547 ^ n15753 ^ 1'b0 ;
  assign n40361 = n18029 ^ n11987 ^ n9399 ;
  assign n40362 = ~n17532 & n23731 ;
  assign n40363 = n31429 ^ n11368 ^ 1'b0 ;
  assign n40364 = n40363 ^ n34581 ^ n7567 ;
  assign n40365 = ( ~n6881 & n8068 ) | ( ~n6881 & n17918 ) | ( n8068 & n17918 ) ;
  assign n40366 = ~n275 & n40365 ;
  assign n40367 = ~n3387 & n28439 ;
  assign n40368 = n36999 & n40367 ;
  assign n40369 = n40368 ^ n11904 ^ 1'b0 ;
  assign n40370 = n27107 ^ n10893 ^ n1133 ;
  assign n40371 = n40370 ^ n34249 ^ n16842 ;
  assign n40372 = n36191 ^ n34843 ^ n11542 ;
  assign n40373 = n13078 & n35997 ;
  assign n40374 = n40373 ^ n33263 ^ 1'b0 ;
  assign n40375 = n40374 ^ n20924 ^ x173 ;
  assign n40376 = n40375 ^ n17795 ^ n3730 ;
  assign n40378 = n35145 ^ n7314 ^ 1'b0 ;
  assign n40379 = n40378 ^ n36275 ^ n999 ;
  assign n40380 = ( n25701 & ~n35273 ) | ( n25701 & n40379 ) | ( ~n35273 & n40379 ) ;
  assign n40381 = ( n1355 & n2410 ) | ( n1355 & n16091 ) | ( n2410 & n16091 ) ;
  assign n40382 = ( n2302 & n5417 ) | ( n2302 & ~n40381 ) | ( n5417 & ~n40381 ) ;
  assign n40383 = ( n18152 & n40380 ) | ( n18152 & n40382 ) | ( n40380 & n40382 ) ;
  assign n40377 = ( x66 & n15933 ) | ( x66 & ~n36352 ) | ( n15933 & ~n36352 ) ;
  assign n40384 = n40383 ^ n40377 ^ n23000 ;
  assign n40385 = ( ~n24454 & n40376 ) | ( ~n24454 & n40384 ) | ( n40376 & n40384 ) ;
  assign n40386 = n33157 ^ n17687 ^ n7093 ;
  assign n40387 = ( n3410 & n6017 ) | ( n3410 & n20606 ) | ( n6017 & n20606 ) ;
  assign n40388 = n27173 ^ n7657 ^ 1'b0 ;
  assign n40389 = ~n40387 & n40388 ;
  assign n40390 = ( ~n1012 & n6076 ) | ( ~n1012 & n40389 ) | ( n6076 & n40389 ) ;
  assign n40391 = ( x15 & n8996 ) | ( x15 & n30723 ) | ( n8996 & n30723 ) ;
  assign n40394 = n11546 ^ n11070 ^ n5709 ;
  assign n40392 = n11001 ^ n2355 ^ 1'b0 ;
  assign n40393 = n2982 & n40392 ;
  assign n40395 = n40394 ^ n40393 ^ n32226 ;
  assign n40396 = ( n11516 & ~n40391 ) | ( n11516 & n40395 ) | ( ~n40391 & n40395 ) ;
  assign n40397 = ( n17376 & n30565 ) | ( n17376 & n37384 ) | ( n30565 & n37384 ) ;
  assign n40398 = n3773 | n5170 ;
  assign n40399 = n40398 ^ n19127 ^ 1'b0 ;
  assign n40400 = n21653 ^ n16291 ^ n6913 ;
  assign n40401 = n40400 ^ n21022 ^ n8314 ;
  assign n40402 = n16556 & n31529 ;
  assign n40403 = n2405 ^ n2188 ^ x188 ;
  assign n40404 = n40403 ^ n38798 ^ n19291 ;
  assign n40405 = n35364 ^ n25823 ^ 1'b0 ;
  assign n40406 = ( n36439 & n40404 ) | ( n36439 & n40405 ) | ( n40404 & n40405 ) ;
  assign n40407 = ( n6203 & ~n10256 ) | ( n6203 & n11103 ) | ( ~n10256 & n11103 ) ;
  assign n40408 = ( ~n287 & n3472 ) | ( ~n287 & n30628 ) | ( n3472 & n30628 ) ;
  assign n40409 = n28473 ^ n4844 ^ 1'b0 ;
  assign n40410 = n40074 | n40409 ;
  assign n40411 = ( n656 & n1701 ) | ( n656 & ~n22888 ) | ( n1701 & ~n22888 ) ;
  assign n40412 = n14032 ^ n5388 ^ n4398 ;
  assign n40413 = ~n11114 & n40412 ;
  assign n40414 = n16199 | n39570 ;
  assign n40415 = n38961 ^ n7258 ^ n6340 ;
  assign n40416 = n40415 ^ n28597 ^ n26310 ;
  assign n40417 = n11895 ^ n2972 ^ n2347 ;
  assign n40418 = n40417 ^ n11091 ^ n6693 ;
  assign n40419 = n10822 & ~n19405 ;
  assign n40420 = ~n34562 & n40419 ;
  assign n40421 = n40420 ^ n28679 ^ n21783 ;
  assign n40422 = ~n7486 & n15026 ;
  assign n40423 = n40422 ^ n21524 ^ 1'b0 ;
  assign n40424 = n40423 ^ n11120 ^ n5367 ;
  assign n40425 = ( ~n11128 & n14294 ) | ( ~n11128 & n32310 ) | ( n14294 & n32310 ) ;
  assign n40426 = ~n14489 & n15952 ;
  assign n40427 = n36937 ^ n19322 ^ n13807 ;
  assign n40428 = n40427 ^ n21943 ^ 1'b0 ;
  assign n40429 = n40426 & n40428 ;
  assign n40430 = n9087 | n32244 ;
  assign n40431 = n40430 ^ n6137 ^ 1'b0 ;
  assign n40432 = ( ~n13293 & n13905 ) | ( ~n13293 & n33594 ) | ( n13905 & n33594 ) ;
  assign n40433 = n28481 ^ n21489 ^ n14521 ;
  assign n40436 = n17789 & ~n37399 ;
  assign n40435 = n33976 ^ n32523 ^ n14383 ;
  assign n40434 = ( n696 & n19614 ) | ( n696 & n38050 ) | ( n19614 & n38050 ) ;
  assign n40437 = n40436 ^ n40435 ^ n40434 ;
  assign n40438 = n39733 ^ n24408 ^ 1'b0 ;
  assign n40439 = ( ~n1645 & n17817 ) | ( ~n1645 & n27178 ) | ( n17817 & n27178 ) ;
  assign n40440 = ( n7289 & n36408 ) | ( n7289 & ~n40439 ) | ( n36408 & ~n40439 ) ;
  assign n40441 = ( n8421 & n9095 ) | ( n8421 & ~n34838 ) | ( n9095 & ~n34838 ) ;
  assign n40442 = n40441 ^ n10808 ^ n3247 ;
  assign n40443 = n19353 ^ n14094 ^ 1'b0 ;
  assign n40444 = ~n35241 & n40443 ;
  assign n40445 = ( n17743 & ~n28465 ) | ( n17743 & n40444 ) | ( ~n28465 & n40444 ) ;
  assign n40446 = n27008 | n38490 ;
  assign n40447 = n3874 | n40446 ;
  assign n40448 = ( n598 & ~n31127 ) | ( n598 & n40447 ) | ( ~n31127 & n40447 ) ;
  assign n40449 = ( n4048 & n4117 ) | ( n4048 & n13217 ) | ( n4117 & n13217 ) ;
  assign n40450 = ~n11742 & n40449 ;
  assign n40451 = ~n13632 & n40450 ;
  assign n40453 = ( n14344 & ~n15415 ) | ( n14344 & n15435 ) | ( ~n15415 & n15435 ) ;
  assign n40452 = n33408 ^ n30664 ^ n20608 ;
  assign n40454 = n40453 ^ n40452 ^ n13878 ;
  assign n40455 = n37587 ^ n15913 ^ n3097 ;
  assign n40456 = n36699 ^ n13887 ^ n519 ;
  assign n40457 = ( n35241 & n40455 ) | ( n35241 & n40456 ) | ( n40455 & n40456 ) ;
  assign n40458 = n3905 & ~n4782 ;
  assign n40459 = n40458 ^ n7403 ^ n6837 ;
  assign n40460 = n40457 & ~n40459 ;
  assign n40461 = n3371 & ~n27124 ;
  assign n40462 = ( n14334 & n14355 ) | ( n14334 & ~n40461 ) | ( n14355 & ~n40461 ) ;
  assign n40463 = ( n24636 & ~n33298 ) | ( n24636 & n40462 ) | ( ~n33298 & n40462 ) ;
  assign n40468 = ( ~x181 & n13481 ) | ( ~x181 & n27494 ) | ( n13481 & n27494 ) ;
  assign n40469 = n21489 ^ n17370 ^ n10105 ;
  assign n40470 = ( n11650 & n40468 ) | ( n11650 & n40469 ) | ( n40468 & n40469 ) ;
  assign n40464 = ( n5504 & n15973 ) | ( n5504 & n16708 ) | ( n15973 & n16708 ) ;
  assign n40465 = n20165 ^ n9604 ^ n9023 ;
  assign n40466 = ( ~n6004 & n7328 ) | ( ~n6004 & n40465 ) | ( n7328 & n40465 ) ;
  assign n40467 = ( n13775 & n40464 ) | ( n13775 & n40466 ) | ( n40464 & n40466 ) ;
  assign n40471 = n40470 ^ n40467 ^ 1'b0 ;
  assign n40473 = n10311 ^ n3414 ^ 1'b0 ;
  assign n40472 = ~n7752 & n19848 ;
  assign n40474 = n40473 ^ n40472 ^ 1'b0 ;
  assign n40475 = n40474 ^ n28139 ^ n28067 ;
  assign n40476 = n465 & ~n25401 ;
  assign n40477 = n40476 ^ n25231 ^ n13716 ;
  assign n40478 = ~n2577 & n18974 ;
  assign n40479 = n40478 ^ n3389 ^ 1'b0 ;
  assign n40480 = ( n26943 & ~n31127 ) | ( n26943 & n40479 ) | ( ~n31127 & n40479 ) ;
  assign n40481 = n40480 ^ n24743 ^ n9171 ;
  assign n40482 = n35824 ^ n6627 ^ 1'b0 ;
  assign n40483 = n27448 ^ n8634 ^ n5406 ;
  assign n40484 = n40483 ^ n14650 ^ x243 ;
  assign n40485 = n15218 ^ n15000 ^ n10957 ;
  assign n40486 = n40485 ^ n36310 ^ n22728 ;
  assign n40487 = n28740 ^ n5853 ^ 1'b0 ;
  assign n40488 = n2006 ^ x67 ^ 1'b0 ;
  assign n40489 = ( n6561 & n8073 ) | ( n6561 & ~n40488 ) | ( n8073 & ~n40488 ) ;
  assign n40490 = n40487 & n40489 ;
  assign n40491 = ( n13039 & n22714 ) | ( n13039 & ~n40490 ) | ( n22714 & ~n40490 ) ;
  assign n40492 = n9165 ^ n7519 ^ n5008 ;
  assign n40493 = ( n12312 & n14725 ) | ( n12312 & ~n40492 ) | ( n14725 & ~n40492 ) ;
  assign n40494 = ( ~n36578 & n40491 ) | ( ~n36578 & n40493 ) | ( n40491 & n40493 ) ;
  assign n40495 = n8828 & ~n19591 ;
  assign n40496 = ( n6980 & n12638 ) | ( n6980 & ~n19500 ) | ( n12638 & ~n19500 ) ;
  assign n40497 = n40013 ^ n7388 ^ n2327 ;
  assign n40498 = ( n24019 & n40496 ) | ( n24019 & n40497 ) | ( n40496 & n40497 ) ;
  assign n40499 = n40498 ^ n35814 ^ n14770 ;
  assign n40500 = ( ~n2754 & n19796 ) | ( ~n2754 & n23777 ) | ( n19796 & n23777 ) ;
  assign n40501 = ( n9256 & ~n15029 ) | ( n9256 & n40500 ) | ( ~n15029 & n40500 ) ;
  assign n40502 = ~n13457 & n23089 ;
  assign n40503 = n40502 ^ n7249 ^ 1'b0 ;
  assign n40504 = n6217 ^ n5977 ^ 1'b0 ;
  assign n40505 = ~n9613 & n40504 ;
  assign n40506 = n40505 ^ n21859 ^ n10379 ;
  assign n40507 = n40506 ^ n8903 ^ n7906 ;
  assign n40509 = n14921 ^ n1567 ^ 1'b0 ;
  assign n40508 = ( n17528 & n21016 ) | ( n17528 & n34076 ) | ( n21016 & n34076 ) ;
  assign n40510 = n40509 ^ n40508 ^ n17651 ;
  assign n40511 = ( n4029 & n15821 ) | ( n4029 & n40510 ) | ( n15821 & n40510 ) ;
  assign n40515 = n14386 ^ n4493 ^ 1'b0 ;
  assign n40512 = ( n3431 & n4126 ) | ( n3431 & ~n4517 ) | ( n4126 & ~n4517 ) ;
  assign n40513 = n20898 ^ n17146 ^ n3560 ;
  assign n40514 = ( ~n29735 & n40512 ) | ( ~n29735 & n40513 ) | ( n40512 & n40513 ) ;
  assign n40516 = n40515 ^ n40514 ^ n35883 ;
  assign n40517 = ( n9213 & n19838 ) | ( n9213 & n33358 ) | ( n19838 & n33358 ) ;
  assign n40518 = n40517 ^ n20425 ^ 1'b0 ;
  assign n40519 = n6269 & n40518 ;
  assign n40520 = ( n7689 & ~n28308 ) | ( n7689 & n33966 ) | ( ~n28308 & n33966 ) ;
  assign n40521 = n40520 ^ n34275 ^ n22024 ;
  assign n40522 = n30921 ^ n21731 ^ n1795 ;
  assign n40523 = ( n10346 & ~n17560 ) | ( n10346 & n40522 ) | ( ~n17560 & n40522 ) ;
  assign n40524 = n4826 ^ n3268 ^ n3084 ;
  assign n40525 = ( n3250 & ~n6859 ) | ( n3250 & n40524 ) | ( ~n6859 & n40524 ) ;
  assign n40526 = ( n13908 & n32580 ) | ( n13908 & ~n40525 ) | ( n32580 & ~n40525 ) ;
  assign n40527 = n22001 & n30912 ;
  assign n40528 = ( n18336 & n26370 ) | ( n18336 & ~n28604 ) | ( n26370 & ~n28604 ) ;
  assign n40529 = n7193 | n14535 ;
  assign n40530 = n40528 | n40529 ;
  assign n40531 = n21890 ^ n16743 ^ n1968 ;
  assign n40532 = n40531 ^ n34783 ^ n3851 ;
  assign n40533 = n19708 ^ n16023 ^ n4197 ;
  assign n40534 = ( n22204 & n31147 ) | ( n22204 & n40533 ) | ( n31147 & n40533 ) ;
  assign n40535 = n40534 ^ n21997 ^ 1'b0 ;
  assign n40536 = n10359 | n40535 ;
  assign n40537 = ( n3088 & ~n12999 ) | ( n3088 & n40536 ) | ( ~n12999 & n40536 ) ;
  assign n40538 = ( n4513 & n8299 ) | ( n4513 & ~n40537 ) | ( n8299 & ~n40537 ) ;
  assign n40539 = n9462 & n18868 ;
  assign n40540 = n35073 & n40539 ;
  assign n40541 = ( ~n8704 & n10232 ) | ( ~n8704 & n10524 ) | ( n10232 & n10524 ) ;
  assign n40542 = n40541 ^ n33092 ^ n13046 ;
  assign n40543 = ( ~n33330 & n40540 ) | ( ~n33330 & n40542 ) | ( n40540 & n40542 ) ;
  assign n40544 = x140 & n7922 ;
  assign n40545 = n2979 & n40544 ;
  assign n40546 = ( n11218 & n16129 ) | ( n11218 & n40545 ) | ( n16129 & n40545 ) ;
  assign n40547 = n19490 ^ n4122 ^ n3983 ;
  assign n40548 = ~n19955 & n40547 ;
  assign n40549 = ( n993 & n26854 ) | ( n993 & n34480 ) | ( n26854 & n34480 ) ;
  assign n40550 = n40549 ^ n1375 ^ 1'b0 ;
  assign n40551 = n19937 & n40550 ;
  assign n40552 = ( n19135 & n40548 ) | ( n19135 & n40551 ) | ( n40548 & n40551 ) ;
  assign n40553 = n35303 ^ n30410 ^ n29497 ;
  assign n40554 = n33400 ^ n6448 ^ n308 ;
  assign n40555 = n25049 ^ n23192 ^ n4682 ;
  assign n40556 = ( ~n10233 & n40554 ) | ( ~n10233 & n40555 ) | ( n40554 & n40555 ) ;
  assign n40557 = n40556 ^ n38619 ^ n614 ;
  assign n40561 = n4118 ^ n2353 ^ n1340 ;
  assign n40559 = n20143 ^ n8549 ^ 1'b0 ;
  assign n40560 = n23019 & ~n40559 ;
  assign n40558 = n27945 ^ n18594 ^ n11808 ;
  assign n40562 = n40561 ^ n40560 ^ n40558 ;
  assign n40563 = n39373 ^ n26666 ^ n6745 ;
  assign n40564 = ~n13114 & n35182 ;
  assign n40565 = n40564 ^ n33089 ^ n27815 ;
  assign n40566 = n33350 ^ n22923 ^ n10436 ;
  assign n40567 = n40566 ^ n14740 ^ 1'b0 ;
  assign n40568 = ( n9999 & n34151 ) | ( n9999 & ~n40567 ) | ( n34151 & ~n40567 ) ;
  assign n40569 = ~n18001 & n18808 ;
  assign n40570 = n6927 & n40569 ;
  assign n40571 = n19406 ^ n8082 ^ 1'b0 ;
  assign n40572 = n40570 | n40571 ;
  assign n40573 = n30408 & ~n34388 ;
  assign n40574 = n38559 ^ n26967 ^ n1019 ;
  assign n40575 = ( n2962 & n4852 ) | ( n2962 & n37338 ) | ( n4852 & n37338 ) ;
  assign n40577 = ( n1260 & ~n8869 ) | ( n1260 & n15612 ) | ( ~n8869 & n15612 ) ;
  assign n40578 = ( n9156 & n28905 ) | ( n9156 & n40577 ) | ( n28905 & n40577 ) ;
  assign n40576 = ~n3370 & n23496 ;
  assign n40579 = n40578 ^ n40576 ^ n29008 ;
  assign n40580 = ( ~n11980 & n15904 ) | ( ~n11980 & n40579 ) | ( n15904 & n40579 ) ;
  assign n40581 = n31153 ^ n9416 ^ n5310 ;
  assign n40582 = n24793 ^ n15698 ^ n9564 ;
  assign n40583 = n11976 | n40582 ;
  assign n40584 = n26927 | n40583 ;
  assign n40585 = n27452 | n40584 ;
  assign n40586 = ( n9082 & n23860 ) | ( n9082 & ~n29541 ) | ( n23860 & ~n29541 ) ;
  assign n40587 = n40586 ^ n27493 ^ n7475 ;
  assign n40588 = ( n7764 & n12595 ) | ( n7764 & ~n40587 ) | ( n12595 & ~n40587 ) ;
  assign n40589 = ( n10498 & n13275 ) | ( n10498 & ~n18110 ) | ( n13275 & ~n18110 ) ;
  assign n40590 = ( n9799 & ~n27501 ) | ( n9799 & n40589 ) | ( ~n27501 & n40589 ) ;
  assign n40591 = n29365 ^ n13438 ^ n6935 ;
  assign n40592 = n40591 ^ n13670 ^ n11929 ;
  assign n40593 = ( ~n6317 & n6552 ) | ( ~n6317 & n40592 ) | ( n6552 & n40592 ) ;
  assign n40594 = ( n14145 & n26245 ) | ( n14145 & ~n40593 ) | ( n26245 & ~n40593 ) ;
  assign n40595 = ( n6558 & n8418 ) | ( n6558 & ~n9382 ) | ( n8418 & ~n9382 ) ;
  assign n40596 = n20587 ^ n16268 ^ n2003 ;
  assign n40597 = ( n6064 & ~n36533 ) | ( n6064 & n40596 ) | ( ~n36533 & n40596 ) ;
  assign n40598 = n39702 ^ n30620 ^ n12724 ;
  assign n40599 = n25141 ^ n15090 ^ 1'b0 ;
  assign n40607 = n10134 & ~n26103 ;
  assign n40606 = ( n4333 & n12551 ) | ( n4333 & ~n13912 ) | ( n12551 & ~n13912 ) ;
  assign n40608 = n40607 ^ n40606 ^ 1'b0 ;
  assign n40605 = ( ~n16016 & n38459 ) | ( ~n16016 & n40013 ) | ( n38459 & n40013 ) ;
  assign n40609 = n40608 ^ n40605 ^ n19015 ;
  assign n40600 = ~n14843 & n25498 ;
  assign n40602 = n21714 ^ n8426 ^ n8053 ;
  assign n40601 = n12559 ^ n10187 ^ n8824 ;
  assign n40603 = n40602 ^ n40601 ^ n8437 ;
  assign n40604 = ( ~n31329 & n40600 ) | ( ~n31329 & n40603 ) | ( n40600 & n40603 ) ;
  assign n40610 = n40609 ^ n40604 ^ n23084 ;
  assign n40611 = n35672 ^ n33927 ^ n31412 ;
  assign n40612 = n3766 ^ n1393 ^ 1'b0 ;
  assign n40613 = n40612 ^ n34497 ^ n10568 ;
  assign n40614 = ( n10260 & ~n27351 ) | ( n10260 & n28781 ) | ( ~n27351 & n28781 ) ;
  assign n40615 = ( n22080 & ~n40613 ) | ( n22080 & n40614 ) | ( ~n40613 & n40614 ) ;
  assign n40616 = n40615 ^ n40381 ^ n29526 ;
  assign n40617 = ( n14548 & n40611 ) | ( n14548 & ~n40616 ) | ( n40611 & ~n40616 ) ;
  assign n40618 = n35472 ^ n10917 ^ n6373 ;
  assign n40619 = ( n2954 & n10210 ) | ( n2954 & ~n40618 ) | ( n10210 & ~n40618 ) ;
  assign n40620 = n40619 ^ n31601 ^ n30710 ;
  assign n40621 = ( ~n5758 & n16879 ) | ( ~n5758 & n18376 ) | ( n16879 & n18376 ) ;
  assign n40622 = n40621 ^ n13344 ^ n2575 ;
  assign n40628 = n39438 ^ n23381 ^ n1090 ;
  assign n40629 = n40628 ^ n16960 ^ n15620 ;
  assign n40623 = ( n2952 & ~n16868 ) | ( n2952 & n31127 ) | ( ~n16868 & n31127 ) ;
  assign n40624 = ~n12480 & n34182 ;
  assign n40625 = n40624 ^ n14886 ^ 1'b0 ;
  assign n40626 = ( n10410 & ~n40623 ) | ( n10410 & n40625 ) | ( ~n40623 & n40625 ) ;
  assign n40627 = ( n389 & n31862 ) | ( n389 & ~n40626 ) | ( n31862 & ~n40626 ) ;
  assign n40630 = n40629 ^ n40627 ^ n22801 ;
  assign n40631 = ( n27501 & n30065 ) | ( n27501 & ~n34736 ) | ( n30065 & ~n34736 ) ;
  assign n40632 = ( n1026 & n8281 ) | ( n1026 & ~n16028 ) | ( n8281 & ~n16028 ) ;
  assign n40633 = n40632 ^ n20236 ^ n2374 ;
  assign n40634 = n13755 & n17037 ;
  assign n40635 = n40634 ^ n26706 ^ 1'b0 ;
  assign n40636 = ( n23321 & ~n35250 ) | ( n23321 & n40635 ) | ( ~n35250 & n40635 ) ;
  assign n40637 = ( n9421 & ~n10730 ) | ( n9421 & n10767 ) | ( ~n10730 & n10767 ) ;
  assign n40638 = n20857 ^ n18244 ^ n2309 ;
  assign n40639 = ( n1293 & ~n11869 ) | ( n1293 & n24565 ) | ( ~n11869 & n24565 ) ;
  assign n40640 = n40639 ^ n5723 ^ 1'b0 ;
  assign n40641 = n40638 | n40640 ;
  assign n40642 = n40641 ^ n30510 ^ n27451 ;
  assign n40643 = n11926 ^ n11073 ^ 1'b0 ;
  assign n40644 = ( n3805 & ~n20535 ) | ( n3805 & n40643 ) | ( ~n20535 & n40643 ) ;
  assign n40645 = n40644 ^ n20985 ^ n7732 ;
  assign n40646 = n34997 ^ n14168 ^ n5359 ;
  assign n40647 = ( n2649 & ~n4300 ) | ( n2649 & n7837 ) | ( ~n4300 & n7837 ) ;
  assign n40648 = ( n8588 & n40646 ) | ( n8588 & ~n40647 ) | ( n40646 & ~n40647 ) ;
  assign n40649 = ( n6654 & n9584 ) | ( n6654 & ~n40648 ) | ( n9584 & ~n40648 ) ;
  assign n40650 = n23115 ^ n3959 ^ 1'b0 ;
  assign n40651 = n6103 & ~n40650 ;
  assign n40652 = n40651 ^ n14575 ^ n13898 ;
  assign n40653 = n37758 | n40652 ;
  assign n40654 = n40653 ^ n12907 ^ n8195 ;
  assign n40655 = n9198 ^ n5530 ^ n2911 ;
  assign n40656 = ( n607 & n4177 ) | ( n607 & n40655 ) | ( n4177 & n40655 ) ;
  assign n40657 = n35230 ^ n11688 ^ n8510 ;
  assign n40658 = ( n17128 & n36786 ) | ( n17128 & n40657 ) | ( n36786 & n40657 ) ;
  assign n40659 = ( ~n20162 & n40656 ) | ( ~n20162 & n40658 ) | ( n40656 & n40658 ) ;
  assign n40660 = n40659 ^ n36726 ^ 1'b0 ;
  assign n40661 = n40654 & n40660 ;
  assign n40662 = n13657 ^ n6691 ^ 1'b0 ;
  assign n40663 = n40662 ^ n19856 ^ n1502 ;
  assign n40664 = n11233 ^ n5786 ^ 1'b0 ;
  assign n40665 = n3981 | n6741 ;
  assign n40666 = n40665 ^ n19831 ^ n9422 ;
  assign n40667 = n40666 ^ n21545 ^ 1'b0 ;
  assign n40670 = n14974 | n19794 ;
  assign n40671 = n40670 ^ n38305 ^ 1'b0 ;
  assign n40672 = n40671 ^ n20556 ^ n13773 ;
  assign n40668 = n31001 ^ n23394 ^ n5288 ;
  assign n40669 = n1192 | n40668 ;
  assign n40673 = n40672 ^ n40669 ^ 1'b0 ;
  assign n40674 = ( ~n14925 & n20207 ) | ( ~n14925 & n40515 ) | ( n20207 & n40515 ) ;
  assign n40675 = ( n7169 & ~n28420 ) | ( n7169 & n40674 ) | ( ~n28420 & n40674 ) ;
  assign n40676 = n40675 ^ n35799 ^ n20038 ;
  assign n40677 = ( ~n10008 & n32124 ) | ( ~n10008 & n33326 ) | ( n32124 & n33326 ) ;
  assign n40678 = n40677 ^ n23559 ^ n7850 ;
  assign n40679 = n23682 ^ n17738 ^ n938 ;
  assign n40680 = n37744 ^ n37473 ^ n34805 ;
  assign n40681 = n7483 & n15868 ;
  assign n40682 = ~n28535 & n40681 ;
  assign n40683 = n3971 | n15574 ;
  assign n40684 = n32390 & ~n40683 ;
  assign n40685 = n40684 ^ n11661 ^ n2932 ;
  assign n40686 = n40685 ^ n28473 ^ n13398 ;
  assign n40687 = n33873 | n40686 ;
  assign n40688 = n40687 ^ n37680 ^ 1'b0 ;
  assign n40689 = n40688 ^ n39320 ^ n2620 ;
  assign n40690 = n40682 & n40689 ;
  assign n40691 = n38005 ^ n26991 ^ n19629 ;
  assign n40693 = ( n3498 & n7730 ) | ( n3498 & n26365 ) | ( n7730 & n26365 ) ;
  assign n40692 = ( n8894 & n25426 ) | ( n8894 & ~n31770 ) | ( n25426 & ~n31770 ) ;
  assign n40694 = n40693 ^ n40692 ^ n17138 ;
  assign n40695 = n40458 ^ n16005 ^ n9729 ;
  assign n40696 = n15264 ^ n14406 ^ n3114 ;
  assign n40697 = ( ~n2775 & n19625 ) | ( ~n2775 & n40696 ) | ( n19625 & n40696 ) ;
  assign n40698 = ( n13807 & n40695 ) | ( n13807 & n40697 ) | ( n40695 & n40697 ) ;
  assign n40699 = ( n2894 & n4099 ) | ( n2894 & ~n38088 ) | ( n4099 & ~n38088 ) ;
  assign n40700 = ( n5376 & ~n8981 ) | ( n5376 & n10010 ) | ( ~n8981 & n10010 ) ;
  assign n40701 = ( n24837 & n40699 ) | ( n24837 & ~n40700 ) | ( n40699 & ~n40700 ) ;
  assign n40702 = ( n1873 & ~n5540 ) | ( n1873 & n40701 ) | ( ~n5540 & n40701 ) ;
  assign n40703 = ( n1921 & n29521 ) | ( n1921 & ~n40389 ) | ( n29521 & ~n40389 ) ;
  assign n40704 = n40703 ^ n30194 ^ n4819 ;
  assign n40705 = ( n662 & n3384 ) | ( n662 & n25763 ) | ( n3384 & n25763 ) ;
  assign n40706 = n40705 ^ n11998 ^ 1'b0 ;
  assign n40707 = n2728 & n40706 ;
  assign n40708 = ( n7494 & n22043 ) | ( n7494 & n40707 ) | ( n22043 & n40707 ) ;
  assign n40709 = n13501 ^ n7524 ^ n5803 ;
  assign n40710 = ( ~n21734 & n32438 ) | ( ~n21734 & n40709 ) | ( n32438 & n40709 ) ;
  assign n40711 = ( n745 & ~n7130 ) | ( n745 & n38941 ) | ( ~n7130 & n38941 ) ;
  assign n40712 = n40711 ^ n26192 ^ n14249 ;
  assign n40713 = ( x82 & n31015 ) | ( x82 & ~n32477 ) | ( n31015 & ~n32477 ) ;
  assign n40714 = ( ~n5980 & n22087 ) | ( ~n5980 & n40713 ) | ( n22087 & n40713 ) ;
  assign n40715 = n19305 ^ n17711 ^ n13799 ;
  assign n40716 = n29071 ^ n26907 ^ n25201 ;
  assign n40717 = n26970 ^ n565 ^ 1'b0 ;
  assign n40718 = n710 & n1930 ;
  assign n40719 = n40718 ^ n6745 ^ 1'b0 ;
  assign n40720 = ( n40716 & ~n40717 ) | ( n40716 & n40719 ) | ( ~n40717 & n40719 ) ;
  assign n40721 = ( n18609 & ~n40715 ) | ( n18609 & n40720 ) | ( ~n40715 & n40720 ) ;
  assign n40722 = ( n12962 & n13342 ) | ( n12962 & ~n24834 ) | ( n13342 & ~n24834 ) ;
  assign n40723 = ( ~n38083 & n39156 ) | ( ~n38083 & n40722 ) | ( n39156 & n40722 ) ;
  assign n40724 = ( n3326 & n5964 ) | ( n3326 & n33267 ) | ( n5964 & n33267 ) ;
  assign n40725 = n40724 ^ n16330 ^ n15238 ;
  assign n40726 = ( n11693 & ~n34290 ) | ( n11693 & n40725 ) | ( ~n34290 & n40725 ) ;
  assign n40727 = n23313 ^ n4715 ^ 1'b0 ;
  assign n40728 = n19410 ^ n11539 ^ n5772 ;
  assign n40729 = n3885 & ~n22140 ;
  assign n40730 = n29941 ^ n17959 ^ n519 ;
  assign n40731 = ( n15612 & ~n40729 ) | ( n15612 & n40730 ) | ( ~n40729 & n40730 ) ;
  assign n40732 = ( n28206 & n40728 ) | ( n28206 & ~n40731 ) | ( n40728 & ~n40731 ) ;
  assign n40733 = ( ~x55 & n40727 ) | ( ~x55 & n40732 ) | ( n40727 & n40732 ) ;
  assign n40734 = n35400 ^ n25546 ^ n8713 ;
  assign n40735 = ( ~n20587 & n30820 ) | ( ~n20587 & n40734 ) | ( n30820 & n40734 ) ;
  assign n40736 = ( n10331 & ~n17771 ) | ( n10331 & n22714 ) | ( ~n17771 & n22714 ) ;
  assign n40737 = ( n19693 & n22803 ) | ( n19693 & n35962 ) | ( n22803 & n35962 ) ;
  assign n40738 = ( n12542 & ~n28894 ) | ( n12542 & n40737 ) | ( ~n28894 & n40737 ) ;
  assign n40739 = n40738 ^ n8372 ^ 1'b0 ;
  assign n40740 = n38395 | n40739 ;
  assign n40743 = ( n36011 & n37173 ) | ( n36011 & n40226 ) | ( n37173 & n40226 ) ;
  assign n40741 = ( n2160 & ~n8009 ) | ( n2160 & n25244 ) | ( ~n8009 & n25244 ) ;
  assign n40742 = n40741 ^ n25907 ^ n20726 ;
  assign n40744 = n40743 ^ n40742 ^ 1'b0 ;
  assign n40745 = n35168 ^ n628 ^ 1'b0 ;
  assign n40746 = n6506 & n40745 ;
  assign n40747 = n40746 ^ n21357 ^ 1'b0 ;
  assign n40748 = ( ~n8628 & n37711 ) | ( ~n8628 & n40747 ) | ( n37711 & n40747 ) ;
  assign n40749 = n17215 ^ n15541 ^ 1'b0 ;
  assign n40750 = n37575 ^ n20332 ^ n18033 ;
  assign n40751 = n40750 ^ n24533 ^ n24349 ;
  assign n40752 = n40751 ^ n25791 ^ n20969 ;
  assign n40753 = n40749 & ~n40752 ;
  assign n40754 = n36531 ^ n11651 ^ n10845 ;
  assign n40755 = ~n19677 & n30968 ;
  assign n40756 = n16008 & n40755 ;
  assign n40757 = ( ~n1760 & n15792 ) | ( ~n1760 & n20823 ) | ( n15792 & n20823 ) ;
  assign n40762 = n12343 ^ n12006 ^ n6129 ;
  assign n40763 = ( n11481 & n17043 ) | ( n11481 & ~n40762 ) | ( n17043 & ~n40762 ) ;
  assign n40758 = n36372 ^ n31661 ^ 1'b0 ;
  assign n40759 = n7995 ^ n5813 ^ n5097 ;
  assign n40760 = ~n8318 & n40759 ;
  assign n40761 = n40758 & n40760 ;
  assign n40764 = n40763 ^ n40761 ^ n5836 ;
  assign n40765 = n5863 & ~n17821 ;
  assign n40766 = n40765 ^ n34350 ^ 1'b0 ;
  assign n40767 = ( n9139 & n28858 ) | ( n9139 & n40766 ) | ( n28858 & n40766 ) ;
  assign n40768 = ( ~n3998 & n13384 ) | ( ~n3998 & n33604 ) | ( n13384 & n33604 ) ;
  assign n40769 = ( ~n23855 & n33600 ) | ( ~n23855 & n40768 ) | ( n33600 & n40768 ) ;
  assign n40770 = ( n2651 & ~n4597 ) | ( n2651 & n37772 ) | ( ~n4597 & n37772 ) ;
  assign n40771 = n40770 ^ n23588 ^ n13440 ;
  assign n40772 = ( ~n563 & n13609 ) | ( ~n563 & n24115 ) | ( n13609 & n24115 ) ;
  assign n40773 = ( n3013 & n40771 ) | ( n3013 & ~n40772 ) | ( n40771 & ~n40772 ) ;
  assign n40774 = n9620 | n25301 ;
  assign n40775 = n10165 & ~n40774 ;
  assign n40776 = ( ~n12302 & n13190 ) | ( ~n12302 & n14952 ) | ( n13190 & n14952 ) ;
  assign n40777 = ~n28023 & n40776 ;
  assign n40778 = n10181 ^ n5859 ^ n4518 ;
  assign n40779 = n40778 ^ n21548 ^ n6286 ;
  assign n40780 = ( ~n10193 & n11383 ) | ( ~n10193 & n18310 ) | ( n11383 & n18310 ) ;
  assign n40781 = n6623 | n40780 ;
  assign n40782 = ( n19753 & ~n24832 ) | ( n19753 & n40781 ) | ( ~n24832 & n40781 ) ;
  assign n40784 = n24130 ^ n19588 ^ n8415 ;
  assign n40785 = n40784 ^ n39435 ^ n20503 ;
  assign n40786 = ( ~n1492 & n10404 ) | ( ~n1492 & n40785 ) | ( n10404 & n40785 ) ;
  assign n40787 = ( n2489 & n37496 ) | ( n2489 & n40786 ) | ( n37496 & n40786 ) ;
  assign n40783 = n14846 & ~n39179 ;
  assign n40788 = n40787 ^ n40783 ^ n15378 ;
  assign n40789 = n38399 ^ n23237 ^ n3270 ;
  assign n40790 = ~n7706 & n24270 ;
  assign n40791 = n40790 ^ n11683 ^ 1'b0 ;
  assign n40792 = ( n14100 & n27497 ) | ( n14100 & n40452 ) | ( n27497 & n40452 ) ;
  assign n40793 = ( n2548 & ~n8550 ) | ( n2548 & n13904 ) | ( ~n8550 & n13904 ) ;
  assign n40794 = ( ~n1139 & n5761 ) | ( ~n1139 & n40793 ) | ( n5761 & n40793 ) ;
  assign n40795 = n40794 ^ n28756 ^ n19192 ;
  assign n40796 = n10956 & n40795 ;
  assign n40797 = n40796 ^ n7526 ^ 1'b0 ;
  assign n40798 = n40797 ^ n19608 ^ n13908 ;
  assign n40799 = ( n40791 & n40792 ) | ( n40791 & ~n40798 ) | ( n40792 & ~n40798 ) ;
  assign n40800 = n23620 ^ n6395 ^ n6324 ;
  assign n40801 = n26635 ^ n23197 ^ n15777 ;
  assign n40802 = ( ~n1683 & n36846 ) | ( ~n1683 & n40801 ) | ( n36846 & n40801 ) ;
  assign n40803 = n31626 ^ n14382 ^ n9361 ;
  assign n40804 = n40803 ^ n7967 ^ n5684 ;
  assign n40805 = ( n3110 & n39436 ) | ( n3110 & n40804 ) | ( n39436 & n40804 ) ;
  assign n40806 = n40805 ^ n14722 ^ n9365 ;
  assign n40807 = n40806 ^ n35991 ^ n20843 ;
  assign n40808 = n8071 | n40807 ;
  assign n40809 = n365 | n40808 ;
  assign n40810 = n30618 | n40809 ;
  assign n40811 = n40810 ^ n6016 ^ 1'b0 ;
  assign n40812 = n32046 ^ n25602 ^ 1'b0 ;
  assign n40813 = n22040 | n40812 ;
  assign n40814 = ( ~n10775 & n12012 ) | ( ~n10775 & n17090 ) | ( n12012 & n17090 ) ;
  assign n40815 = n40814 ^ n32041 ^ n30155 ;
  assign n40816 = ( ~n2237 & n28948 ) | ( ~n2237 & n40815 ) | ( n28948 & n40815 ) ;
  assign n40817 = n24699 ^ n18534 ^ n8879 ;
  assign n40818 = n40817 ^ n9347 ^ n8412 ;
  assign n40819 = ~n2510 & n25235 ;
  assign n40820 = n40819 ^ n2408 ^ 1'b0 ;
  assign n40821 = n6966 ^ n2108 ^ 1'b0 ;
  assign n40822 = ( n11704 & ~n40820 ) | ( n11704 & n40821 ) | ( ~n40820 & n40821 ) ;
  assign n40823 = n13816 & ~n40822 ;
  assign n40824 = n40818 & n40823 ;
  assign n40825 = ( n20656 & n35777 ) | ( n20656 & ~n40824 ) | ( n35777 & ~n40824 ) ;
  assign n40826 = ( n6608 & n14205 ) | ( n6608 & n19320 ) | ( n14205 & n19320 ) ;
  assign n40827 = n21943 ^ n15328 ^ n10441 ;
  assign n40828 = ( ~n11073 & n15694 ) | ( ~n11073 & n40827 ) | ( n15694 & n40827 ) ;
  assign n40829 = n40828 ^ n11362 ^ n3604 ;
  assign n40830 = ( ~n4093 & n18025 ) | ( ~n4093 & n21048 ) | ( n18025 & n21048 ) ;
  assign n40831 = n40309 ^ n27565 ^ 1'b0 ;
  assign n40832 = n8909 & n31754 ;
  assign n40833 = ~n40831 & n40832 ;
  assign n40834 = n27905 ^ n23803 ^ n17221 ;
  assign n40835 = ( n3180 & n20059 ) | ( n3180 & ~n33270 ) | ( n20059 & ~n33270 ) ;
  assign n40836 = ( n34785 & ~n40834 ) | ( n34785 & n40835 ) | ( ~n40834 & n40835 ) ;
  assign n40837 = n40836 ^ n29672 ^ n5768 ;
  assign n40838 = n31619 ^ n14897 ^ n14345 ;
  assign n40839 = ( n3092 & n19131 ) | ( n3092 & n40838 ) | ( n19131 & n40838 ) ;
  assign n40840 = n40839 ^ n19856 ^ 1'b0 ;
  assign n40841 = n40837 | n40840 ;
  assign n40842 = n24566 | n25869 ;
  assign n40843 = n40842 ^ n29843 ^ 1'b0 ;
  assign n40844 = n40843 ^ n34043 ^ n32575 ;
  assign n40845 = n40844 ^ n10096 ^ n2704 ;
  assign n40846 = n33263 ^ n7457 ^ n5734 ;
  assign n40847 = ( n15235 & n37087 ) | ( n15235 & ~n40846 ) | ( n37087 & ~n40846 ) ;
  assign n40850 = n17563 ^ n13519 ^ n10262 ;
  assign n40848 = n12991 & n28004 ;
  assign n40849 = ( ~n19658 & n23604 ) | ( ~n19658 & n40848 ) | ( n23604 & n40848 ) ;
  assign n40851 = n40850 ^ n40849 ^ n17022 ;
  assign n40852 = n20464 ^ n9956 ^ n3794 ;
  assign n40853 = ( n8625 & n15883 ) | ( n8625 & ~n29179 ) | ( n15883 & ~n29179 ) ;
  assign n40854 = ( ~n34095 & n40852 ) | ( ~n34095 & n40853 ) | ( n40852 & n40853 ) ;
  assign n40855 = n14594 & n18537 ;
  assign n40856 = ~n33859 & n40855 ;
  assign n40859 = n5983 ^ n1537 ^ n1325 ;
  assign n40858 = ( n1153 & ~n11493 ) | ( n1153 & n25570 ) | ( ~n11493 & n25570 ) ;
  assign n40860 = n40859 ^ n40858 ^ n14888 ;
  assign n40861 = ( n20796 & n26425 ) | ( n20796 & n40860 ) | ( n26425 & n40860 ) ;
  assign n40857 = n24300 ^ n21635 ^ n17545 ;
  assign n40862 = n40861 ^ n40857 ^ n40330 ;
  assign n40863 = ( n20837 & ~n23554 ) | ( n20837 & n38193 ) | ( ~n23554 & n38193 ) ;
  assign n40864 = n15708 ^ n8647 ^ n6467 ;
  assign n40865 = n6296 & ~n17289 ;
  assign n40866 = n2340 & n40865 ;
  assign n40867 = ( n2166 & n31204 ) | ( n2166 & ~n32523 ) | ( n31204 & ~n32523 ) ;
  assign n40868 = ( n7076 & n40866 ) | ( n7076 & ~n40867 ) | ( n40866 & ~n40867 ) ;
  assign n40869 = n30343 ^ n19429 ^ n16822 ;
  assign n40870 = n40869 ^ n18987 ^ n5147 ;
  assign n40871 = ( ~n7353 & n13966 ) | ( ~n7353 & n30052 ) | ( n13966 & n30052 ) ;
  assign n40872 = n28887 ^ n12188 ^ n9461 ;
  assign n40873 = n40872 ^ n6605 ^ n3023 ;
  assign n40874 = n40873 ^ n13491 ^ n13412 ;
  assign n40875 = n40874 ^ n17290 ^ n16300 ;
  assign n40876 = n40875 ^ n18234 ^ n9811 ;
  assign n40877 = ( ~n1086 & n19115 ) | ( ~n1086 & n25390 ) | ( n19115 & n25390 ) ;
  assign n40878 = ( n4709 & n14477 ) | ( n4709 & n40877 ) | ( n14477 & n40877 ) ;
  assign n40879 = n39063 ^ n11023 ^ n726 ;
  assign n40880 = n1716 & n36783 ;
  assign n40881 = n15346 ^ n14602 ^ n8860 ;
  assign n40882 = ( n6326 & n16504 ) | ( n6326 & n35167 ) | ( n16504 & n35167 ) ;
  assign n40883 = ( n39561 & n40881 ) | ( n39561 & ~n40882 ) | ( n40881 & ~n40882 ) ;
  assign n40886 = n33653 ^ n25738 ^ 1'b0 ;
  assign n40884 = n34836 ^ n33892 ^ n25629 ;
  assign n40885 = n40884 ^ n17732 ^ n7321 ;
  assign n40887 = n40886 ^ n40885 ^ n12268 ;
  assign n40888 = ( ~n5631 & n16501 ) | ( ~n5631 & n19091 ) | ( n16501 & n19091 ) ;
  assign n40889 = n6889 ^ n627 ^ 1'b0 ;
  assign n40890 = n6631 & n40889 ;
  assign n40891 = n40890 ^ n35933 ^ n9810 ;
  assign n40895 = ~n34676 & n39493 ;
  assign n40896 = n40895 ^ n13015 ^ 1'b0 ;
  assign n40892 = ( ~n1301 & n6426 ) | ( ~n1301 & n10869 ) | ( n6426 & n10869 ) ;
  assign n40893 = n40892 ^ n8042 ^ n4198 ;
  assign n40894 = ( n3601 & n19916 ) | ( n3601 & n40893 ) | ( n19916 & n40893 ) ;
  assign n40897 = n40896 ^ n40894 ^ n37618 ;
  assign n40898 = ( ~n11826 & n28585 ) | ( ~n11826 & n31037 ) | ( n28585 & n31037 ) ;
  assign n40899 = n3526 | n12857 ;
  assign n40900 = n40899 ^ n30186 ^ 1'b0 ;
  assign n40901 = ( n3080 & n6875 ) | ( n3080 & n18065 ) | ( n6875 & n18065 ) ;
  assign n40902 = n40901 ^ n32029 ^ n29669 ;
  assign n40903 = n25332 ^ n7009 ^ 1'b0 ;
  assign n40904 = ( n31318 & n36868 ) | ( n31318 & ~n40903 ) | ( n36868 & ~n40903 ) ;
  assign n40905 = n23862 ^ n13388 ^ 1'b0 ;
  assign n40906 = n40905 ^ n19907 ^ n6639 ;
  assign n40907 = ( n2626 & n18301 ) | ( n2626 & ~n40906 ) | ( n18301 & ~n40906 ) ;
  assign n40908 = n26302 ^ x47 ^ 1'b0 ;
  assign n40909 = n32827 & ~n40908 ;
  assign n40910 = n16662 & n18704 ;
  assign n40911 = ~n40909 & n40910 ;
  assign n40912 = n40911 ^ n19068 ^ n16687 ;
  assign n40913 = ( ~n23926 & n40907 ) | ( ~n23926 & n40912 ) | ( n40907 & n40912 ) ;
  assign n40914 = n40913 ^ n35232 ^ n14957 ;
  assign n40919 = ( n338 & n2638 ) | ( n338 & n21007 ) | ( n2638 & n21007 ) ;
  assign n40915 = n33139 ^ n16225 ^ 1'b0 ;
  assign n40916 = n5935 | n38145 ;
  assign n40917 = n40916 ^ n37497 ^ 1'b0 ;
  assign n40918 = ( ~n34423 & n40915 ) | ( ~n34423 & n40917 ) | ( n40915 & n40917 ) ;
  assign n40920 = n40919 ^ n40918 ^ n40119 ;
  assign n40921 = ( ~n7177 & n12798 ) | ( ~n7177 & n20361 ) | ( n12798 & n20361 ) ;
  assign n40922 = n15240 ^ n6109 ^ 1'b0 ;
  assign n40923 = n13887 ^ n10450 ^ n7162 ;
  assign n40924 = ( n32190 & ~n40922 ) | ( n32190 & n40923 ) | ( ~n40922 & n40923 ) ;
  assign n40925 = n6118 ^ n3717 ^ n2783 ;
  assign n40926 = n40925 ^ n33240 ^ n14195 ;
  assign n40927 = n40926 ^ n33437 ^ n18943 ;
  assign n40928 = ( n8945 & n10420 ) | ( n8945 & ~n14797 ) | ( n10420 & ~n14797 ) ;
  assign n40929 = ~n40927 & n40928 ;
  assign n40930 = ( ~n14014 & n20700 ) | ( ~n14014 & n40929 ) | ( n20700 & n40929 ) ;
  assign n40931 = ( n5085 & n20714 ) | ( n5085 & n28672 ) | ( n20714 & n28672 ) ;
  assign n40932 = ( n1067 & n13719 ) | ( n1067 & ~n21733 ) | ( n13719 & ~n21733 ) ;
  assign n40933 = n40932 ^ n20841 ^ n12188 ;
  assign n40934 = ( ~n16286 & n22466 ) | ( ~n16286 & n40933 ) | ( n22466 & n40933 ) ;
  assign n40935 = n1901 | n21265 ;
  assign n40936 = n13195 & ~n40935 ;
  assign n40937 = n2814 | n4322 ;
  assign n40938 = n7409 & ~n40937 ;
  assign n40939 = ( ~n5770 & n12707 ) | ( ~n5770 & n40938 ) | ( n12707 & n40938 ) ;
  assign n40940 = n40939 ^ n19170 ^ n9015 ;
  assign n40941 = ( n10777 & ~n12712 ) | ( n10777 & n40940 ) | ( ~n12712 & n40940 ) ;
  assign n40942 = n28739 ^ n16784 ^ n11965 ;
  assign n40943 = n40942 ^ n1477 ^ 1'b0 ;
  assign n40944 = n990 & n40943 ;
  assign n40945 = n40944 ^ n34749 ^ 1'b0 ;
  assign n40946 = x192 & ~n40945 ;
  assign n40947 = n18931 ^ n14354 ^ n3867 ;
  assign n40949 = ( n19739 & ~n22285 ) | ( n19739 & n23489 ) | ( ~n22285 & n23489 ) ;
  assign n40948 = n25728 ^ n9359 ^ n1700 ;
  assign n40950 = n40949 ^ n40948 ^ n20113 ;
  assign n40951 = n40950 ^ n20792 ^ n7972 ;
  assign n40952 = ( n16840 & n40947 ) | ( n16840 & n40951 ) | ( n40947 & n40951 ) ;
  assign n40953 = ( n15697 & n28782 ) | ( n15697 & n32961 ) | ( n28782 & n32961 ) ;
  assign n40954 = ( n40946 & n40952 ) | ( n40946 & n40953 ) | ( n40952 & n40953 ) ;
  assign n40955 = ( n19137 & n33346 ) | ( n19137 & n35409 ) | ( n33346 & n35409 ) ;
  assign n40956 = n30422 ^ n6977 ^ 1'b0 ;
  assign n40957 = ( n9878 & n17184 ) | ( n9878 & ~n29734 ) | ( n17184 & ~n29734 ) ;
  assign n40958 = ( n496 & n40956 ) | ( n496 & ~n40957 ) | ( n40956 & ~n40957 ) ;
  assign n40959 = ( n707 & n9262 ) | ( n707 & n15989 ) | ( n9262 & n15989 ) ;
  assign n40960 = n31361 ^ n19811 ^ n9104 ;
  assign n40961 = ( ~n13940 & n40959 ) | ( ~n13940 & n40960 ) | ( n40959 & n40960 ) ;
  assign n40962 = n31654 ^ n3613 ^ n428 ;
  assign n40963 = n40962 ^ n35688 ^ 1'b0 ;
  assign n40964 = n351 & n40963 ;
  assign n40965 = n4227 & n14819 ;
  assign n40966 = n40965 ^ n9357 ^ n9067 ;
  assign n40967 = n24263 ^ n17676 ^ n1893 ;
  assign n40968 = n26523 | n40967 ;
  assign n40969 = n8603 & ~n40968 ;
  assign n40970 = ( ~n5078 & n15069 ) | ( ~n5078 & n40969 ) | ( n15069 & n40969 ) ;
  assign n40971 = ( ~n6194 & n9449 ) | ( ~n6194 & n26199 ) | ( n9449 & n26199 ) ;
  assign n40972 = ( n16285 & ~n25279 ) | ( n16285 & n30961 ) | ( ~n25279 & n30961 ) ;
  assign n40973 = ( n8835 & ~n14718 ) | ( n8835 & n15709 ) | ( ~n14718 & n15709 ) ;
  assign n40974 = n40973 ^ n25102 ^ n5501 ;
  assign n40975 = ( ~n22524 & n40972 ) | ( ~n22524 & n40974 ) | ( n40972 & n40974 ) ;
  assign n40976 = ( n3725 & ~n26864 ) | ( n3725 & n30168 ) | ( ~n26864 & n30168 ) ;
  assign n40977 = ( ~n8501 & n19443 ) | ( ~n8501 & n31954 ) | ( n19443 & n31954 ) ;
  assign n40978 = ( ~n6471 & n8170 ) | ( ~n6471 & n40977 ) | ( n8170 & n40977 ) ;
  assign n40979 = n14581 | n19638 ;
  assign n40980 = n40979 ^ n5492 ^ 1'b0 ;
  assign n40981 = ( n2402 & n10536 ) | ( n2402 & n24098 ) | ( n10536 & n24098 ) ;
  assign n40982 = n26034 ^ n22218 ^ n12460 ;
  assign n40983 = ( n3138 & n10074 ) | ( n3138 & ~n40982 ) | ( n10074 & ~n40982 ) ;
  assign n40984 = n40983 ^ n17591 ^ n13551 ;
  assign n40985 = ( n16338 & n37852 ) | ( n16338 & ~n40984 ) | ( n37852 & ~n40984 ) ;
  assign n40986 = ( ~n7119 & n24194 ) | ( ~n7119 & n40985 ) | ( n24194 & n40985 ) ;
  assign n40987 = n2846 | n21368 ;
  assign n40988 = n12938 & ~n40987 ;
  assign n40989 = ( n826 & ~n16097 ) | ( n826 & n40988 ) | ( ~n16097 & n40988 ) ;
  assign n40990 = ( n1151 & n11406 ) | ( n1151 & n38493 ) | ( n11406 & n38493 ) ;
  assign n40991 = ( n6450 & ~n10519 ) | ( n6450 & n21860 ) | ( ~n10519 & n21860 ) ;
  assign n40992 = n36590 ^ n35898 ^ 1'b0 ;
  assign n40993 = ( n9685 & n40991 ) | ( n9685 & ~n40992 ) | ( n40991 & ~n40992 ) ;
  assign n40994 = n1917 & n10376 ;
  assign n40995 = n40994 ^ n2251 ^ 1'b0 ;
  assign n40996 = n15269 ^ n1193 ^ 1'b0 ;
  assign n40997 = n40996 ^ n7715 ^ n5421 ;
  assign n40998 = ( n26207 & n29146 ) | ( n26207 & n40997 ) | ( n29146 & n40997 ) ;
  assign n40999 = ( n1064 & n6040 ) | ( n1064 & ~n14651 ) | ( n6040 & ~n14651 ) ;
  assign n41000 = n10017 & ~n40999 ;
  assign n41001 = ( n19491 & n39828 ) | ( n19491 & n41000 ) | ( n39828 & n41000 ) ;
  assign n41002 = ( n7933 & n20858 ) | ( n7933 & ~n41001 ) | ( n20858 & ~n41001 ) ;
  assign n41003 = n41002 ^ n30595 ^ n25715 ;
  assign n41004 = ( n16226 & n35711 ) | ( n16226 & ~n41003 ) | ( n35711 & ~n41003 ) ;
  assign n41005 = n25829 ^ n5740 ^ x224 ;
  assign n41006 = ( n17487 & n39040 ) | ( n17487 & n41005 ) | ( n39040 & n41005 ) ;
  assign n41007 = ( n884 & ~n4795 ) | ( n884 & n8239 ) | ( ~n4795 & n8239 ) ;
  assign n41008 = n13069 ^ n6405 ^ 1'b0 ;
  assign n41009 = n588 & ~n41008 ;
  assign n41010 = ( n12004 & ~n30459 ) | ( n12004 & n41009 ) | ( ~n30459 & n41009 ) ;
  assign n41011 = ( ~n593 & n8698 ) | ( ~n593 & n41010 ) | ( n8698 & n41010 ) ;
  assign n41012 = ( n26574 & ~n41007 ) | ( n26574 & n41011 ) | ( ~n41007 & n41011 ) ;
  assign n41013 = n34453 ^ n24436 ^ n23337 ;
  assign n41014 = ( n665 & n21307 ) | ( n665 & ~n41013 ) | ( n21307 & ~n41013 ) ;
  assign n41015 = n33148 ^ n26770 ^ 1'b0 ;
  assign n41016 = n2333 | n41015 ;
  assign n41020 = ~n6755 & n12898 ;
  assign n41021 = n41020 ^ n28298 ^ 1'b0 ;
  assign n41017 = ( n6351 & ~n6763 ) | ( n6351 & n33520 ) | ( ~n6763 & n33520 ) ;
  assign n41018 = n41017 ^ n16315 ^ n2805 ;
  assign n41019 = n41018 ^ n24865 ^ n8000 ;
  assign n41022 = n41021 ^ n41019 ^ n14565 ;
  assign n41023 = n41022 ^ n34584 ^ n17717 ;
  assign n41024 = n5131 & ~n8859 ;
  assign n41025 = ~n36676 & n41024 ;
  assign n41026 = ( n1488 & n2138 ) | ( n1488 & n41025 ) | ( n2138 & n41025 ) ;
  assign n41027 = ( n3854 & n7597 ) | ( n3854 & n12332 ) | ( n7597 & n12332 ) ;
  assign n41028 = ( n26036 & n31509 ) | ( n26036 & n35330 ) | ( n31509 & n35330 ) ;
  assign n41029 = n41028 ^ n37851 ^ 1'b0 ;
  assign n41031 = ( x28 & ~n6444 ) | ( x28 & n22721 ) | ( ~n6444 & n22721 ) ;
  assign n41032 = ( ~n4411 & n11943 ) | ( ~n4411 & n41031 ) | ( n11943 & n41031 ) ;
  assign n41030 = n38910 ^ n27184 ^ n25092 ;
  assign n41033 = n41032 ^ n41030 ^ n2548 ;
  assign n41037 = n19970 ^ n6886 ^ n4482 ;
  assign n41035 = n24406 & n28327 ;
  assign n41036 = ~n19212 & n41035 ;
  assign n41034 = n25083 ^ x192 ^ 1'b0 ;
  assign n41038 = n41037 ^ n41036 ^ n41034 ;
  assign n41041 = n28687 ^ n13509 ^ n2588 ;
  assign n41039 = n26699 ^ n21129 ^ n20546 ;
  assign n41040 = n41039 ^ n18405 ^ n15640 ;
  assign n41042 = n41041 ^ n41040 ^ n39251 ;
  assign n41043 = ~n7554 & n38101 ;
  assign n41044 = n41042 & n41043 ;
  assign n41045 = n18874 ^ n1689 ^ 1'b0 ;
  assign n41046 = n41044 | n41045 ;
  assign n41047 = ( n15333 & ~n16698 ) | ( n15333 & n18700 ) | ( ~n16698 & n18700 ) ;
  assign n41048 = ( ~n17724 & n19272 ) | ( ~n17724 & n41047 ) | ( n19272 & n41047 ) ;
  assign n41049 = ( n12405 & n14532 ) | ( n12405 & n41048 ) | ( n14532 & n41048 ) ;
  assign n41050 = n41049 ^ n29770 ^ n16190 ;
  assign n41051 = n41050 ^ n35799 ^ 1'b0 ;
  assign n41052 = n18592 | n41051 ;
  assign n41053 = ( n4447 & n17526 ) | ( n4447 & n18981 ) | ( n17526 & n18981 ) ;
  assign n41054 = ( n9515 & n16081 ) | ( n9515 & n41053 ) | ( n16081 & n41053 ) ;
  assign n41055 = n6510 | n35605 ;
  assign n41056 = ( n24738 & ~n38805 ) | ( n24738 & n41055 ) | ( ~n38805 & n41055 ) ;
  assign n41057 = n23351 ^ n12888 ^ n8034 ;
  assign n41058 = n41057 ^ n31113 ^ n25859 ;
  assign n41059 = n8318 & n35264 ;
  assign n41060 = n41059 ^ n27885 ^ n22880 ;
  assign n41061 = ( n39133 & n40093 ) | ( n39133 & n41060 ) | ( n40093 & n41060 ) ;
  assign n41062 = ( n2864 & n6472 ) | ( n2864 & n15213 ) | ( n6472 & n15213 ) ;
  assign n41063 = ( ~n13750 & n28022 ) | ( ~n13750 & n41062 ) | ( n28022 & n41062 ) ;
  assign n41065 = n7816 ^ n7380 ^ n1825 ;
  assign n41064 = n14281 ^ n11051 ^ n572 ;
  assign n41066 = n41065 ^ n41064 ^ n26902 ;
  assign n41067 = n41066 ^ n13351 ^ n8460 ;
  assign n41068 = n41067 ^ n3527 ^ 1'b0 ;
  assign n41069 = n36396 ^ n15932 ^ n3714 ;
  assign n41070 = n11810 ^ n5265 ^ 1'b0 ;
  assign n41071 = n14245 & ~n41070 ;
  assign n41072 = n41071 ^ n12253 ^ 1'b0 ;
  assign n41073 = n40134 | n41072 ;
  assign n41074 = ~n1024 & n10543 ;
  assign n41075 = n41074 ^ n11257 ^ 1'b0 ;
  assign n41077 = n9347 ^ n7257 ^ n4946 ;
  assign n41076 = n27564 ^ n14233 ^ n12280 ;
  assign n41078 = n41077 ^ n41076 ^ n21016 ;
  assign n41079 = n41078 ^ n34991 ^ n5434 ;
  assign n41080 = ( n5549 & ~n9724 ) | ( n5549 & n19284 ) | ( ~n9724 & n19284 ) ;
  assign n41081 = n3419 ^ n878 ^ 1'b0 ;
  assign n41082 = n41080 & ~n41081 ;
  assign n41083 = n41082 ^ n29540 ^ n26149 ;
  assign n41084 = ~n3198 & n13360 ;
  assign n41085 = ~n21035 & n41084 ;
  assign n41086 = n41085 ^ n22235 ^ n944 ;
  assign n41087 = n7134 | n38685 ;
  assign n41088 = n22562 & ~n41087 ;
  assign n41089 = ( n10840 & n24596 ) | ( n10840 & ~n41088 ) | ( n24596 & ~n41088 ) ;
  assign n41090 = ( ~n2573 & n6824 ) | ( ~n2573 & n24624 ) | ( n6824 & n24624 ) ;
  assign n41091 = ( n439 & n14027 ) | ( n439 & n41090 ) | ( n14027 & n41090 ) ;
  assign n41092 = ( n1323 & n6021 ) | ( n1323 & n18485 ) | ( n6021 & n18485 ) ;
  assign n41093 = n41092 ^ n22214 ^ n16295 ;
  assign n41094 = ~n19252 & n23570 ;
  assign n41095 = ~n30570 & n41094 ;
  assign n41096 = ( n6737 & n9087 ) | ( n6737 & n17345 ) | ( n9087 & n17345 ) ;
  assign n41097 = ~n6800 & n41096 ;
  assign n41098 = n41097 ^ n26822 ^ 1'b0 ;
  assign n41099 = ~n1266 & n11225 ;
  assign n41100 = ( n3372 & n11726 ) | ( n3372 & ~n41099 ) | ( n11726 & ~n41099 ) ;
  assign n41107 = n12577 ^ n5850 ^ n1188 ;
  assign n41108 = n41107 ^ n18799 ^ n1522 ;
  assign n41109 = ( ~n4793 & n24826 ) | ( ~n4793 & n41108 ) | ( n24826 & n41108 ) ;
  assign n41101 = n11134 ^ n8359 ^ 1'b0 ;
  assign n41102 = n5022 & n41101 ;
  assign n41103 = ( n1668 & n13508 ) | ( n1668 & n41102 ) | ( n13508 & n41102 ) ;
  assign n41104 = n8703 & ~n17819 ;
  assign n41105 = n41104 ^ n34940 ^ 1'b0 ;
  assign n41106 = ~n41103 & n41105 ;
  assign n41110 = n41109 ^ n41106 ^ n26861 ;
  assign n41113 = n30199 ^ n22505 ^ n18577 ;
  assign n41114 = n41113 ^ n31437 ^ n25730 ;
  assign n41111 = ( n2494 & n15562 ) | ( n2494 & n16068 ) | ( n15562 & n16068 ) ;
  assign n41112 = ( n3420 & ~n8438 ) | ( n3420 & n41111 ) | ( ~n8438 & n41111 ) ;
  assign n41115 = n41114 ^ n41112 ^ n19631 ;
  assign n41116 = n24924 ^ n16038 ^ x68 ;
  assign n41117 = n41116 ^ n25717 ^ n17943 ;
  assign n41118 = n35502 ^ n15685 ^ n7287 ;
  assign n41119 = ( n18612 & ~n21187 ) | ( n18612 & n41118 ) | ( ~n21187 & n41118 ) ;
  assign n41120 = ( n3622 & n36253 ) | ( n3622 & n41119 ) | ( n36253 & n41119 ) ;
  assign n41121 = ~n22032 & n38693 ;
  assign n41122 = ( n4995 & ~n22323 ) | ( n4995 & n29736 ) | ( ~n22323 & n29736 ) ;
  assign n41123 = n41122 ^ n17668 ^ n1839 ;
  assign n41124 = n4621 & n14286 ;
  assign n41125 = ~n41123 & n41124 ;
  assign n41126 = ( n1967 & ~n41121 ) | ( n1967 & n41125 ) | ( ~n41121 & n41125 ) ;
  assign n41127 = n41126 ^ n24013 ^ n14440 ;
  assign n41128 = n16681 | n19179 ;
  assign n41129 = ( n10594 & n33444 ) | ( n10594 & n41128 ) | ( n33444 & n41128 ) ;
  assign n41133 = n36045 ^ n6269 ^ n3687 ;
  assign n41130 = ( ~n3244 & n4817 ) | ( ~n3244 & n5477 ) | ( n4817 & n5477 ) ;
  assign n41131 = n41130 ^ n17866 ^ n1289 ;
  assign n41132 = n5273 & ~n41131 ;
  assign n41134 = n41133 ^ n41132 ^ 1'b0 ;
  assign n41135 = n18690 ^ n3063 ^ 1'b0 ;
  assign n41136 = n41135 ^ n40827 ^ n22529 ;
  assign n41137 = n41136 ^ n29517 ^ n1268 ;
  assign n41138 = n13542 ^ n8201 ^ n556 ;
  assign n41139 = n41138 ^ n4965 ^ 1'b0 ;
  assign n41140 = ~n624 & n41139 ;
  assign n41141 = ~n15593 & n22360 ;
  assign n41142 = ( n33863 & ~n41140 ) | ( n33863 & n41141 ) | ( ~n41140 & n41141 ) ;
  assign n41143 = ~n16259 & n28476 ;
  assign n41144 = ~n16958 & n31014 ;
  assign n41145 = n41144 ^ n36905 ^ 1'b0 ;
  assign n41146 = ( n2543 & n31178 ) | ( n2543 & ~n32494 ) | ( n31178 & ~n32494 ) ;
  assign n41147 = n7923 | n17172 ;
  assign n41148 = ~n41146 & n41147 ;
  assign n41149 = n41148 ^ n13640 ^ 1'b0 ;
  assign n41150 = ( ~n23893 & n41145 ) | ( ~n23893 & n41149 ) | ( n41145 & n41149 ) ;
  assign n41151 = n9464 ^ n5544 ^ 1'b0 ;
  assign n41152 = n4003 & ~n41151 ;
  assign n41153 = ( n18637 & n29388 ) | ( n18637 & n41152 ) | ( n29388 & n41152 ) ;
  assign n41154 = n6809 ^ n6363 ^ n3105 ;
  assign n41155 = n7098 | n41154 ;
  assign n41156 = n1877 & ~n41155 ;
  assign n41157 = n41156 ^ n28866 ^ n19952 ;
  assign n41158 = ( n9534 & n35803 ) | ( n9534 & ~n41157 ) | ( n35803 & ~n41157 ) ;
  assign n41159 = ( n5855 & n15402 ) | ( n5855 & ~n23101 ) | ( n15402 & ~n23101 ) ;
  assign n41160 = n41159 ^ n5111 ^ n4283 ;
  assign n41161 = n9497 ^ n8001 ^ n6875 ;
  assign n41162 = ( n10310 & n16708 ) | ( n10310 & ~n37261 ) | ( n16708 & ~n37261 ) ;
  assign n41163 = ( n28175 & n41161 ) | ( n28175 & n41162 ) | ( n41161 & n41162 ) ;
  assign n41164 = ( x106 & n3706 ) | ( x106 & ~n41163 ) | ( n3706 & ~n41163 ) ;
  assign n41165 = ( n14581 & n30265 ) | ( n14581 & n41164 ) | ( n30265 & n41164 ) ;
  assign n41166 = n33950 ^ n32998 ^ n1763 ;
  assign n41167 = n16694 ^ n14048 ^ n739 ;
  assign n41168 = n41167 ^ n19753 ^ n18240 ;
  assign n41169 = ( n3573 & n10165 ) | ( n3573 & ~n41168 ) | ( n10165 & ~n41168 ) ;
  assign n41170 = ( n5291 & n35745 ) | ( n5291 & ~n41169 ) | ( n35745 & ~n41169 ) ;
  assign n41171 = ( n904 & n5910 ) | ( n904 & ~n35382 ) | ( n5910 & ~n35382 ) ;
  assign n41172 = ( n25947 & n33724 ) | ( n25947 & ~n35739 ) | ( n33724 & ~n35739 ) ;
  assign n41173 = n41172 ^ n25876 ^ n15687 ;
  assign n41174 = n41173 ^ n15050 ^ 1'b0 ;
  assign n41175 = n6671 & n41174 ;
  assign n41176 = n41175 ^ n27451 ^ n9750 ;
  assign n41177 = n25289 ^ n24435 ^ n21653 ;
  assign n41178 = n19996 ^ n11569 ^ 1'b0 ;
  assign n41179 = n41178 ^ n21968 ^ n3851 ;
  assign n41180 = n41179 ^ n40045 ^ n22997 ;
  assign n41181 = ( n3568 & n6783 ) | ( n3568 & ~n25230 ) | ( n6783 & ~n25230 ) ;
  assign n41182 = n28211 | n41181 ;
  assign n41183 = n4213 | n41182 ;
  assign n41185 = ( n3101 & ~n9114 ) | ( n3101 & n31062 ) | ( ~n9114 & n31062 ) ;
  assign n41184 = n11238 ^ n743 ^ 1'b0 ;
  assign n41186 = n41185 ^ n41184 ^ n4480 ;
  assign n41187 = ( n5851 & ~n12541 ) | ( n5851 & n41186 ) | ( ~n12541 & n41186 ) ;
  assign n41196 = n38039 ^ n16019 ^ n9565 ;
  assign n41190 = ( n293 & n3904 ) | ( n293 & ~n25410 ) | ( n3904 & ~n25410 ) ;
  assign n41191 = ( n11117 & n14780 ) | ( n11117 & ~n41190 ) | ( n14780 & ~n41190 ) ;
  assign n41192 = n41191 ^ n32918 ^ n18945 ;
  assign n41188 = n9681 ^ n9647 ^ n3524 ;
  assign n41189 = n41188 ^ n20915 ^ n12167 ;
  assign n41193 = n41192 ^ n41189 ^ n35828 ;
  assign n41194 = ( ~n9197 & n20680 ) | ( ~n9197 & n25436 ) | ( n20680 & n25436 ) ;
  assign n41195 = ( n8506 & ~n41193 ) | ( n8506 & n41194 ) | ( ~n41193 & n41194 ) ;
  assign n41197 = n41196 ^ n41195 ^ n9605 ;
  assign n41198 = n41197 ^ n756 ^ n658 ;
  assign n41199 = ( n14878 & n21143 ) | ( n14878 & n24192 ) | ( n21143 & n24192 ) ;
  assign n41200 = n4210 | n12288 ;
  assign n41201 = ( ~n11482 & n21939 ) | ( ~n11482 & n25581 ) | ( n21939 & n25581 ) ;
  assign n41202 = ( n5616 & ~n13141 ) | ( n5616 & n21019 ) | ( ~n13141 & n21019 ) ;
  assign n41203 = n41202 ^ n26133 ^ n293 ;
  assign n41204 = ( n35419 & n38527 ) | ( n35419 & n39408 ) | ( n38527 & n39408 ) ;
  assign n41205 = ( n3327 & n10072 ) | ( n3327 & ~n13577 ) | ( n10072 & ~n13577 ) ;
  assign n41206 = ( n8902 & ~n36193 ) | ( n8902 & n41205 ) | ( ~n36193 & n41205 ) ;
  assign n41207 = n15612 & n24261 ;
  assign n41208 = n41207 ^ n26654 ^ n530 ;
  assign n41209 = ( n3593 & ~n11815 ) | ( n3593 & n12782 ) | ( ~n11815 & n12782 ) ;
  assign n41210 = n12739 ^ n9108 ^ 1'b0 ;
  assign n41211 = n41209 | n41210 ;
  assign n41212 = ( n33919 & ~n35741 ) | ( n33919 & n41211 ) | ( ~n35741 & n41211 ) ;
  assign n41213 = ( n7202 & n14950 ) | ( n7202 & ~n41212 ) | ( n14950 & ~n41212 ) ;
  assign n41214 = ( n7543 & n41208 ) | ( n7543 & ~n41213 ) | ( n41208 & ~n41213 ) ;
  assign n41215 = n33479 ^ x187 ^ 1'b0 ;
  assign n41216 = n14729 ^ n9378 ^ n7324 ;
  assign n41217 = ( n808 & n36799 ) | ( n808 & n41216 ) | ( n36799 & n41216 ) ;
  assign n41218 = ( n3181 & n38758 ) | ( n3181 & n41217 ) | ( n38758 & n41217 ) ;
  assign n41219 = ( n2759 & n41215 ) | ( n2759 & ~n41218 ) | ( n41215 & ~n41218 ) ;
  assign n41220 = n23349 ^ n22696 ^ n3702 ;
  assign n41221 = n41220 ^ n2890 ^ n825 ;
  assign n41226 = n30199 ^ n15370 ^ n15276 ;
  assign n41222 = n10889 ^ n4617 ^ n1606 ;
  assign n41223 = ( n23934 & n26744 ) | ( n23934 & n26923 ) | ( n26744 & n26923 ) ;
  assign n41224 = n41223 ^ n28718 ^ n15055 ;
  assign n41225 = ( n21239 & n41222 ) | ( n21239 & ~n41224 ) | ( n41222 & ~n41224 ) ;
  assign n41227 = n41226 ^ n41225 ^ n14764 ;
  assign n41228 = ( n4871 & n10974 ) | ( n4871 & ~n19142 ) | ( n10974 & ~n19142 ) ;
  assign n41229 = ( ~n11955 & n25089 ) | ( ~n11955 & n37207 ) | ( n25089 & n37207 ) ;
  assign n41230 = n41229 ^ n15586 ^ n10289 ;
  assign n41231 = ( n31561 & n41228 ) | ( n31561 & n41230 ) | ( n41228 & n41230 ) ;
  assign n41232 = ( n351 & ~n15479 ) | ( n351 & n22262 ) | ( ~n15479 & n22262 ) ;
  assign n41233 = n41232 ^ n22255 ^ 1'b0 ;
  assign n41234 = n17196 & n25371 ;
  assign n41235 = n41234 ^ n10775 ^ 1'b0 ;
  assign n41236 = n37719 ^ n37406 ^ n989 ;
  assign n41237 = ( ~n9301 & n10555 ) | ( ~n9301 & n14205 ) | ( n10555 & n14205 ) ;
  assign n41238 = n38178 ^ n16658 ^ n891 ;
  assign n41239 = n32841 ^ n31164 ^ n28978 ;
  assign n41240 = ( ~n718 & n9866 ) | ( ~n718 & n17199 ) | ( n9866 & n17199 ) ;
  assign n41241 = n2216 & ~n4845 ;
  assign n41242 = n41240 & n41241 ;
  assign n41243 = n40516 ^ n25177 ^ 1'b0 ;
  assign n41244 = n21278 | n41243 ;
  assign n41245 = n33583 ^ n32009 ^ n20514 ;
  assign n41246 = n10781 | n23282 ;
  assign n41247 = ~n2761 & n3695 ;
  assign n41248 = n41247 ^ n28579 ^ 1'b0 ;
  assign n41249 = ( ~n7578 & n30776 ) | ( ~n7578 & n41248 ) | ( n30776 & n41248 ) ;
  assign n41250 = ( n1090 & n33244 ) | ( n1090 & n39261 ) | ( n33244 & n39261 ) ;
  assign n41251 = ( n4005 & n27550 ) | ( n4005 & ~n41250 ) | ( n27550 & ~n41250 ) ;
  assign n41252 = ( n1000 & n41249 ) | ( n1000 & n41251 ) | ( n41249 & n41251 ) ;
  assign n41253 = ( n2262 & n34879 ) | ( n2262 & ~n37381 ) | ( n34879 & ~n37381 ) ;
  assign n41255 = ( n2755 & n13648 ) | ( n2755 & ~n14965 ) | ( n13648 & ~n14965 ) ;
  assign n41254 = n1784 | n14922 ;
  assign n41256 = n41255 ^ n41254 ^ 1'b0 ;
  assign n41257 = n36132 ^ n34347 ^ n7500 ;
  assign n41258 = n35803 ^ n14422 ^ n11038 ;
  assign n41259 = n41258 ^ n26564 ^ n2423 ;
  assign n41260 = n4093 & ~n39208 ;
  assign n41261 = n37696 ^ n27961 ^ n1909 ;
  assign n41262 = ( n5927 & n24461 ) | ( n5927 & ~n41261 ) | ( n24461 & ~n41261 ) ;
  assign n41263 = n28527 ^ n18769 ^ n3015 ;
  assign n41264 = n40925 ^ n11135 ^ 1'b0 ;
  assign n41265 = n40120 ^ n13217 ^ 1'b0 ;
  assign n41266 = n26479 ^ n14927 ^ n4152 ;
  assign n41267 = n8004 & ~n41266 ;
  assign n41268 = n30230 & n41267 ;
  assign n41269 = n41268 ^ n27113 ^ n17943 ;
  assign n41270 = n40688 & n41269 ;
  assign n41271 = n31164 ^ n12855 ^ 1'b0 ;
  assign n41272 = ~n27594 & n41271 ;
  assign n41273 = n13671 & n32803 ;
  assign n41274 = ( n27462 & ~n32919 ) | ( n27462 & n41273 ) | ( ~n32919 & n41273 ) ;
  assign n41275 = ( n13076 & n24507 ) | ( n13076 & n34090 ) | ( n24507 & n34090 ) ;
  assign n41276 = n12067 ^ n6659 ^ n2260 ;
  assign n41277 = ( ~n7741 & n8432 ) | ( ~n7741 & n16944 ) | ( n8432 & n16944 ) ;
  assign n41278 = n41277 ^ n37035 ^ n4053 ;
  assign n41279 = ( n40828 & n41276 ) | ( n40828 & n41278 ) | ( n41276 & n41278 ) ;
  assign n41280 = n36000 ^ n31693 ^ n7922 ;
  assign n41284 = ( n1096 & n28251 ) | ( n1096 & n30776 ) | ( n28251 & n30776 ) ;
  assign n41282 = n16083 ^ n15632 ^ 1'b0 ;
  assign n41283 = n14941 & n41282 ;
  assign n41281 = ( n505 & n3702 ) | ( n505 & ~n25610 ) | ( n3702 & ~n25610 ) ;
  assign n41285 = n41284 ^ n41283 ^ n41281 ;
  assign n41286 = ( n30519 & n37022 ) | ( n30519 & n41285 ) | ( n37022 & n41285 ) ;
  assign n41287 = n39741 ^ n37232 ^ n28770 ;
  assign n41288 = n14286 ^ n6021 ^ n1436 ;
  assign n41289 = ( ~n4533 & n19252 ) | ( ~n4533 & n41288 ) | ( n19252 & n41288 ) ;
  assign n41290 = ( n1145 & n7823 ) | ( n1145 & n19643 ) | ( n7823 & n19643 ) ;
  assign n41291 = n41290 ^ n17145 ^ n4785 ;
  assign n41292 = n41291 ^ n33250 ^ n658 ;
  assign n41293 = n2954 & n9829 ;
  assign n41294 = n41292 & n41293 ;
  assign n41295 = n33064 ^ n31581 ^ n6596 ;
  assign n41296 = n3607 | n41295 ;
  assign n41297 = n37739 & ~n41296 ;
  assign n41298 = n35605 ^ n18292 ^ n13442 ;
  assign n41299 = ( n9082 & n14234 ) | ( n9082 & n41298 ) | ( n14234 & n41298 ) ;
  assign n41300 = ( n9704 & n32632 ) | ( n9704 & ~n33901 ) | ( n32632 & ~n33901 ) ;
  assign n41301 = n10690 ^ n9253 ^ n8036 ;
  assign n41302 = n38213 ^ n30977 ^ n14505 ;
  assign n41303 = ( ~n21093 & n41301 ) | ( ~n21093 & n41302 ) | ( n41301 & n41302 ) ;
  assign n41304 = ( n11539 & n15213 ) | ( n11539 & n36092 ) | ( n15213 & n36092 ) ;
  assign n41305 = n39196 ^ n12530 ^ n11346 ;
  assign n41306 = ( n35100 & n40476 ) | ( n35100 & n41305 ) | ( n40476 & n41305 ) ;
  assign n41307 = n36604 ^ n27472 ^ n14919 ;
  assign n41308 = ( n1979 & ~n10657 ) | ( n1979 & n28787 ) | ( ~n10657 & n28787 ) ;
  assign n41309 = n41308 ^ n29818 ^ n1232 ;
  assign n41310 = x32 & ~n29800 ;
  assign n41311 = ( ~n2080 & n26048 ) | ( ~n2080 & n41310 ) | ( n26048 & n41310 ) ;
  assign n41312 = n41311 ^ n18787 ^ n5233 ;
  assign n41313 = n3393 & n6333 ;
  assign n41314 = n14764 & n41313 ;
  assign n41315 = n35540 ^ n26184 ^ n3654 ;
  assign n41316 = ( ~n11887 & n32439 ) | ( ~n11887 & n41315 ) | ( n32439 & n41315 ) ;
  assign n41317 = ( n6178 & ~n11996 ) | ( n6178 & n19850 ) | ( ~n11996 & n19850 ) ;
  assign n41318 = ( ~n1522 & n6318 ) | ( ~n1522 & n15519 ) | ( n6318 & n15519 ) ;
  assign n41321 = n22056 ^ n17519 ^ n3259 ;
  assign n41322 = n41321 ^ n5079 ^ 1'b0 ;
  assign n41319 = ~n3794 & n31677 ;
  assign n41320 = n41319 ^ n3365 ^ 1'b0 ;
  assign n41323 = n41322 ^ n41320 ^ n17375 ;
  assign n41324 = n41323 ^ n28016 ^ n22991 ;
  assign n41325 = n22926 ^ n10508 ^ 1'b0 ;
  assign n41327 = ( n537 & n2756 ) | ( n537 & n19393 ) | ( n2756 & n19393 ) ;
  assign n41326 = ( ~n2080 & n10467 ) | ( ~n2080 & n37925 ) | ( n10467 & n37925 ) ;
  assign n41328 = n41327 ^ n41326 ^ n26220 ;
  assign n41329 = n41328 ^ n38465 ^ n35972 ;
  assign n41330 = ( n6254 & n24781 ) | ( n6254 & ~n38674 ) | ( n24781 & ~n38674 ) ;
  assign n41331 = ( n12308 & n38943 ) | ( n12308 & n41330 ) | ( n38943 & n41330 ) ;
  assign n41332 = n11216 ^ n2815 ^ n539 ;
  assign n41333 = n41332 ^ n39714 ^ n7425 ;
  assign n41334 = n29495 ^ n25124 ^ 1'b0 ;
  assign n41335 = n34728 & n41334 ;
  assign n41336 = n9203 & n11821 ;
  assign n41337 = n41336 ^ n4000 ^ 1'b0 ;
  assign n41338 = n41337 ^ n21932 ^ n21180 ;
  assign n41339 = ( n30204 & n34896 ) | ( n30204 & ~n41338 ) | ( n34896 & ~n41338 ) ;
  assign n41340 = ( n1278 & n39259 ) | ( n1278 & ~n41339 ) | ( n39259 & ~n41339 ) ;
  assign n41341 = ( n22294 & n25418 ) | ( n22294 & n41340 ) | ( n25418 & n41340 ) ;
  assign n41342 = ( n1709 & n14817 ) | ( n1709 & ~n41341 ) | ( n14817 & ~n41341 ) ;
  assign n41343 = ( ~n4087 & n6087 ) | ( ~n4087 & n6960 ) | ( n6087 & n6960 ) ;
  assign n41344 = n41343 ^ n14470 ^ n1470 ;
  assign n41345 = n41344 ^ n14219 ^ n3719 ;
  assign n41346 = n31208 ^ n5477 ^ 1'b0 ;
  assign n41347 = n3471 & n41346 ;
  assign n41348 = ~n7926 & n40689 ;
  assign n41349 = ~n41347 & n41348 ;
  assign n41350 = n6684 | n13280 ;
  assign n41351 = n16496 | n41350 ;
  assign n41352 = n29136 ^ n14304 ^ n8382 ;
  assign n41353 = n41352 ^ n23503 ^ n11276 ;
  assign n41354 = ( n9206 & n28732 ) | ( n9206 & n29157 ) | ( n28732 & n29157 ) ;
  assign n41355 = ( ~n9900 & n23880 ) | ( ~n9900 & n41354 ) | ( n23880 & n41354 ) ;
  assign n41356 = ( n7720 & ~n28044 ) | ( n7720 & n31581 ) | ( ~n28044 & n31581 ) ;
  assign n41357 = n30202 ^ n26943 ^ n5270 ;
  assign n41358 = n40207 ^ n35898 ^ n16105 ;
  assign n41359 = n38950 ^ n37643 ^ n5352 ;
  assign n41362 = ~n2378 & n15927 ;
  assign n41360 = ( ~n2899 & n4732 ) | ( ~n2899 & n16047 ) | ( n4732 & n16047 ) ;
  assign n41361 = n41360 ^ n33184 ^ n8191 ;
  assign n41363 = n41362 ^ n41361 ^ 1'b0 ;
  assign n41364 = ( ~n5907 & n9716 ) | ( ~n5907 & n32549 ) | ( n9716 & n32549 ) ;
  assign n41365 = ( n8910 & n16656 ) | ( n8910 & ~n41364 ) | ( n16656 & ~n41364 ) ;
  assign n41366 = n5853 & n37022 ;
  assign n41367 = ~n22531 & n25030 ;
  assign n41368 = n41367 ^ n15069 ^ 1'b0 ;
  assign n41369 = n15871 ^ n12060 ^ 1'b0 ;
  assign n41370 = ( n1771 & ~n14085 ) | ( n1771 & n36154 ) | ( ~n14085 & n36154 ) ;
  assign n41371 = ( n1257 & ~n27490 ) | ( n1257 & n34631 ) | ( ~n27490 & n34631 ) ;
  assign n41372 = ( ~n32816 & n41370 ) | ( ~n32816 & n41371 ) | ( n41370 & n41371 ) ;
  assign n41373 = ~n13031 & n14846 ;
  assign n41374 = n41373 ^ n40795 ^ n5714 ;
  assign n41375 = ( n16947 & n27420 ) | ( n16947 & n41374 ) | ( n27420 & n41374 ) ;
  assign n41376 = ( n8236 & n26220 ) | ( n8236 & n31882 ) | ( n26220 & n31882 ) ;
  assign n41377 = ( n11904 & ~n12163 ) | ( n11904 & n24768 ) | ( ~n12163 & n24768 ) ;
  assign n41378 = ( n13256 & n40956 ) | ( n13256 & n41377 ) | ( n40956 & n41377 ) ;
  assign n41379 = ( n673 & n18018 ) | ( n673 & ~n26972 ) | ( n18018 & ~n26972 ) ;
  assign n41380 = ( n11871 & n33641 ) | ( n11871 & ~n41379 ) | ( n33641 & ~n41379 ) ;
  assign n41381 = ( n12956 & n17875 ) | ( n12956 & ~n41380 ) | ( n17875 & ~n41380 ) ;
  assign n41382 = ( n7542 & ~n19946 ) | ( n7542 & n24981 ) | ( ~n19946 & n24981 ) ;
  assign n41383 = ( ~n13437 & n17670 ) | ( ~n13437 & n41382 ) | ( n17670 & n41382 ) ;
  assign n41384 = ( n14232 & ~n15007 ) | ( n14232 & n41383 ) | ( ~n15007 & n41383 ) ;
  assign n41385 = n15901 ^ n3990 ^ 1'b0 ;
  assign n41386 = ( n3811 & n15504 ) | ( n3811 & n41385 ) | ( n15504 & n41385 ) ;
  assign n41390 = n397 & ~n11776 ;
  assign n41389 = n39109 ^ n37591 ^ n25378 ;
  assign n41387 = ( x34 & n895 ) | ( x34 & ~n37450 ) | ( n895 & ~n37450 ) ;
  assign n41388 = ( n3496 & n30536 ) | ( n3496 & ~n41387 ) | ( n30536 & ~n41387 ) ;
  assign n41391 = n41390 ^ n41389 ^ n41388 ;
  assign n41392 = ( ~n15866 & n41386 ) | ( ~n15866 & n41391 ) | ( n41386 & n41391 ) ;
  assign n41393 = ( n8897 & ~n18781 ) | ( n8897 & n19667 ) | ( ~n18781 & n19667 ) ;
  assign n41394 = n7163 ^ n6901 ^ n760 ;
  assign n41395 = ( n406 & n9528 ) | ( n406 & n21283 ) | ( n9528 & n21283 ) ;
  assign n41396 = n25119 ^ n8587 ^ x68 ;
  assign n41397 = ( n10459 & n14611 ) | ( n10459 & ~n41396 ) | ( n14611 & ~n41396 ) ;
  assign n41398 = n41397 ^ n21702 ^ n17365 ;
  assign n41399 = n41398 ^ n21784 ^ n1686 ;
  assign n41400 = n41399 ^ n7824 ^ n2160 ;
  assign n41401 = ( ~n38546 & n41374 ) | ( ~n38546 & n41400 ) | ( n41374 & n41400 ) ;
  assign n41402 = n36920 ^ n29692 ^ n7968 ;
  assign n41403 = ( n5989 & n33083 ) | ( n5989 & n41402 ) | ( n33083 & n41402 ) ;
  assign n41404 = n35420 ^ n16508 ^ n4533 ;
  assign n41405 = ( n1569 & n12605 ) | ( n1569 & ~n25460 ) | ( n12605 & ~n25460 ) ;
  assign n41406 = ( ~n7201 & n11962 ) | ( ~n7201 & n31153 ) | ( n11962 & n31153 ) ;
  assign n41407 = n6558 | n35027 ;
  assign n41408 = n41407 ^ n7624 ^ 1'b0 ;
  assign n41409 = n41408 ^ n501 ^ 1'b0 ;
  assign n41410 = n41406 & ~n41409 ;
  assign n41411 = ( ~n544 & n13385 ) | ( ~n544 & n21300 ) | ( n13385 & n21300 ) ;
  assign n41412 = n41411 ^ n4455 ^ 1'b0 ;
  assign n41413 = n12129 | n36387 ;
  assign n41414 = n41412 | n41413 ;
  assign n41415 = ( n9885 & n26199 ) | ( n9885 & n32401 ) | ( n26199 & n32401 ) ;
  assign n41417 = ( n20181 & n27644 ) | ( n20181 & ~n32989 ) | ( n27644 & ~n32989 ) ;
  assign n41416 = ( n9958 & ~n17338 ) | ( n9958 & n26997 ) | ( ~n17338 & n26997 ) ;
  assign n41418 = n41417 ^ n41416 ^ n9335 ;
  assign n41419 = n26136 ^ n9937 ^ n8773 ;
  assign n41420 = n41419 ^ n25299 ^ n19977 ;
  assign n41423 = n10720 ^ n10102 ^ n5010 ;
  assign n41424 = n16296 ^ n14950 ^ 1'b0 ;
  assign n41425 = n41423 & ~n41424 ;
  assign n41426 = ( n8975 & n23003 ) | ( n8975 & n41425 ) | ( n23003 & n41425 ) ;
  assign n41421 = ( ~n8186 & n8804 ) | ( ~n8186 & n12735 ) | ( n8804 & n12735 ) ;
  assign n41422 = n41421 ^ n31318 ^ n15817 ;
  assign n41427 = n41426 ^ n41422 ^ n20955 ;
  assign n41428 = n8160 & ~n18716 ;
  assign n41429 = n41428 ^ n35161 ^ 1'b0 ;
  assign n41430 = n31596 ^ n25722 ^ n8809 ;
  assign n41431 = ( n16038 & ~n40926 ) | ( n16038 & n41430 ) | ( ~n40926 & n41430 ) ;
  assign n41432 = ( n1896 & ~n25502 ) | ( n1896 & n25694 ) | ( ~n25502 & n25694 ) ;
  assign n41433 = n41432 ^ n38659 ^ n22978 ;
  assign n41434 = ( n6786 & n20030 ) | ( n6786 & ~n33519 ) | ( n20030 & ~n33519 ) ;
  assign n41436 = n22328 ^ n13436 ^ n4556 ;
  assign n41435 = ( ~n7463 & n14682 ) | ( ~n7463 & n22852 ) | ( n14682 & n22852 ) ;
  assign n41437 = n41436 ^ n41435 ^ n27239 ;
  assign n41438 = ( ~n9555 & n16111 ) | ( ~n9555 & n21951 ) | ( n16111 & n21951 ) ;
  assign n41439 = n41438 ^ n18643 ^ n14417 ;
  assign n41440 = ( n26794 & n28168 ) | ( n26794 & n34308 ) | ( n28168 & n34308 ) ;
  assign n41441 = n41440 ^ n39090 ^ n28784 ;
  assign n41442 = n25944 ^ n12329 ^ n6823 ;
  assign n41443 = n17424 ^ n11569 ^ n2811 ;
  assign n41444 = n38925 ^ n22903 ^ n14843 ;
  assign n41445 = n41444 ^ n28469 ^ n9311 ;
  assign n41450 = n39071 ^ n24993 ^ n15541 ;
  assign n41449 = ~n2820 & n12638 ;
  assign n41451 = n41450 ^ n41449 ^ 1'b0 ;
  assign n41446 = n19830 ^ n11120 ^ n6585 ;
  assign n41447 = n41446 ^ n35230 ^ n2275 ;
  assign n41448 = n5854 & n41447 ;
  assign n41452 = n41451 ^ n41448 ^ 1'b0 ;
  assign n41454 = n26524 ^ n5767 ^ n3482 ;
  assign n41455 = ~n12728 & n22360 ;
  assign n41456 = ~n41454 & n41455 ;
  assign n41453 = n20526 & n33295 ;
  assign n41457 = n41456 ^ n41453 ^ 1'b0 ;
  assign n41460 = n12799 ^ n9070 ^ n5294 ;
  assign n41461 = n41460 ^ n31788 ^ n30528 ;
  assign n41458 = n20094 ^ n10826 ^ n9860 ;
  assign n41459 = n41458 ^ n19819 ^ x22 ;
  assign n41462 = n41461 ^ n41459 ^ n26227 ;
  assign n41463 = n18451 ^ n12546 ^ n8760 ;
  assign n41464 = ~n11106 & n18197 ;
  assign n41465 = n41464 ^ n4767 ^ x50 ;
  assign n41466 = ( n22411 & n41463 ) | ( n22411 & ~n41465 ) | ( n41463 & ~n41465 ) ;
  assign n41467 = ( n13755 & n23825 ) | ( n13755 & n41466 ) | ( n23825 & n41466 ) ;
  assign n41468 = ( n3340 & n3783 ) | ( n3340 & n4015 ) | ( n3783 & n4015 ) ;
  assign n41469 = n41468 ^ n30171 ^ 1'b0 ;
  assign n41470 = ( n3696 & n9747 ) | ( n3696 & ~n30545 ) | ( n9747 & ~n30545 ) ;
  assign n41471 = ( n1708 & n8136 ) | ( n1708 & n29233 ) | ( n8136 & n29233 ) ;
  assign n41472 = n13307 | n16820 ;
  assign n41473 = n7737 | n41472 ;
  assign n41474 = n41473 ^ n28250 ^ n18299 ;
  assign n41475 = n39889 ^ n2344 ^ 1'b0 ;
  assign n41476 = n14568 & ~n41475 ;
  assign n41477 = ( n15700 & n41474 ) | ( n15700 & ~n41476 ) | ( n41474 & ~n41476 ) ;
  assign n41478 = n15747 ^ n7448 ^ n1968 ;
  assign n41479 = n41478 ^ n39030 ^ n16857 ;
  assign n41480 = n30857 ^ n13039 ^ n6644 ;
  assign n41481 = ( n15942 & n31778 ) | ( n15942 & ~n41480 ) | ( n31778 & ~n41480 ) ;
  assign n41482 = ~n2616 & n23676 ;
  assign n41483 = n17754 & n41482 ;
  assign n41484 = x26 & n1015 ;
  assign n41485 = n21759 & n41484 ;
  assign n41486 = ( n5953 & n9693 ) | ( n5953 & n41485 ) | ( n9693 & n41485 ) ;
  assign n41487 = ( n13169 & ~n16168 ) | ( n13169 & n36908 ) | ( ~n16168 & n36908 ) ;
  assign n41488 = ( n4811 & ~n24904 ) | ( n4811 & n41487 ) | ( ~n24904 & n41487 ) ;
  assign n41489 = n36878 & n41488 ;
  assign n41490 = n41486 & n41489 ;
  assign n41491 = n41490 ^ n29146 ^ n16828 ;
  assign n41492 = ( n12682 & n18167 ) | ( n12682 & ~n18534 ) | ( n18167 & ~n18534 ) ;
  assign n41493 = n4433 ^ n4211 ^ 1'b0 ;
  assign n41494 = n41493 ^ n15976 ^ 1'b0 ;
  assign n41495 = n17451 ^ n11175 ^ n9790 ;
  assign n41496 = ( n17226 & n18642 ) | ( n17226 & ~n41495 ) | ( n18642 & ~n41495 ) ;
  assign n41497 = n41496 ^ n25404 ^ n19689 ;
  assign n41498 = ( n6324 & n20098 ) | ( n6324 & n37445 ) | ( n20098 & n37445 ) ;
  assign n41499 = n31794 ^ n26916 ^ 1'b0 ;
  assign n41503 = n6323 ^ n2859 ^ 1'b0 ;
  assign n41504 = ~n515 & n41503 ;
  assign n41500 = n25273 ^ n24717 ^ n1158 ;
  assign n41501 = n41500 ^ n20006 ^ n7430 ;
  assign n41502 = ( n6507 & n30290 ) | ( n6507 & n41501 ) | ( n30290 & n41501 ) ;
  assign n41505 = n41504 ^ n41502 ^ n18342 ;
  assign n41506 = ~n13073 & n33972 ;
  assign n41507 = ~n1570 & n41506 ;
  assign n41508 = n41507 ^ n30093 ^ n29449 ;
  assign n41509 = n33880 ^ n23468 ^ n12883 ;
  assign n41510 = n41509 ^ n23387 ^ n3833 ;
  assign n41511 = ( n1941 & ~n41508 ) | ( n1941 & n41510 ) | ( ~n41508 & n41510 ) ;
  assign n41512 = n24521 ^ n22201 ^ x149 ;
  assign n41513 = ( n25186 & n37666 ) | ( n25186 & n41512 ) | ( n37666 & n41512 ) ;
  assign n41514 = n22392 ^ n18239 ^ n15637 ;
  assign n41515 = n11128 | n20473 ;
  assign n41516 = n41515 ^ n38276 ^ n34914 ;
  assign n41517 = n41516 ^ n40762 ^ n38495 ;
  assign n41518 = n1313 & n10916 ;
  assign n41519 = ( n16010 & n19680 ) | ( n16010 & ~n22786 ) | ( n19680 & ~n22786 ) ;
  assign n41520 = ( n5584 & n23220 ) | ( n5584 & n41519 ) | ( n23220 & n41519 ) ;
  assign n41521 = ( ~n36730 & n41010 ) | ( ~n36730 & n41520 ) | ( n41010 & n41520 ) ;
  assign n41522 = ( n5177 & n8530 ) | ( n5177 & ~n41521 ) | ( n8530 & ~n41521 ) ;
  assign n41524 = n11438 ^ n2068 ^ n962 ;
  assign n41523 = n33092 ^ n11413 ^ n10717 ;
  assign n41525 = n41524 ^ n41523 ^ n39082 ;
  assign n41527 = n14403 ^ n7293 ^ n3206 ;
  assign n41526 = n21348 ^ n15734 ^ 1'b0 ;
  assign n41528 = n41527 ^ n41526 ^ 1'b0 ;
  assign n41529 = n14232 & n37260 ;
  assign n41530 = n41529 ^ n39947 ^ 1'b0 ;
  assign n41531 = n38101 ^ n21220 ^ n19109 ;
  assign n41532 = n4466 & ~n41531 ;
  assign n41533 = n26252 ^ n15483 ^ x207 ;
  assign n41534 = ( ~n1579 & n3773 ) | ( ~n1579 & n41533 ) | ( n3773 & n41533 ) ;
  assign n41535 = ( n1005 & n15370 ) | ( n1005 & ~n26327 ) | ( n15370 & ~n26327 ) ;
  assign n41538 = ( n5656 & n9359 ) | ( n5656 & ~n10718 ) | ( n9359 & ~n10718 ) ;
  assign n41536 = n3841 & ~n27420 ;
  assign n41537 = n36791 & n41536 ;
  assign n41539 = n41538 ^ n41537 ^ n40405 ;
  assign n41540 = ( n3630 & n20185 ) | ( n3630 & n24176 ) | ( n20185 & n24176 ) ;
  assign n41541 = ( n15097 & n26319 ) | ( n15097 & ~n34518 ) | ( n26319 & ~n34518 ) ;
  assign n41542 = n8683 ^ n511 ^ 1'b0 ;
  assign n41543 = n7800 & n41542 ;
  assign n41544 = n21232 ^ n10763 ^ 1'b0 ;
  assign n41545 = n41543 & ~n41544 ;
  assign n41546 = ( n7797 & n13673 ) | ( n7797 & n34939 ) | ( n13673 & n34939 ) ;
  assign n41547 = n6616 | n41546 ;
  assign n41548 = ( n4904 & n23579 ) | ( n4904 & n32357 ) | ( n23579 & n32357 ) ;
  assign n41549 = n34650 ^ n9860 ^ n805 ;
  assign n41550 = n27489 ^ n13688 ^ 1'b0 ;
  assign n41551 = n27657 | n41550 ;
  assign n41556 = ( n23469 & ~n34315 ) | ( n23469 & n40376 ) | ( ~n34315 & n40376 ) ;
  assign n41557 = n41556 ^ n19339 ^ 1'b0 ;
  assign n41552 = ( n4823 & n29403 ) | ( n4823 & ~n29940 ) | ( n29403 & ~n29940 ) ;
  assign n41553 = ( n15416 & n28583 ) | ( n15416 & n41552 ) | ( n28583 & n41552 ) ;
  assign n41554 = n41553 ^ n38767 ^ n10195 ;
  assign n41555 = ( n32976 & ~n40695 ) | ( n32976 & n41554 ) | ( ~n40695 & n41554 ) ;
  assign n41558 = n41557 ^ n41555 ^ n10408 ;
  assign n41559 = n24601 ^ n14243 ^ n13006 ;
  assign n41560 = n35533 ^ n17440 ^ n10307 ;
  assign n41561 = ( n20505 & n41559 ) | ( n20505 & ~n41560 ) | ( n41559 & ~n41560 ) ;
  assign n41562 = n19286 ^ n15292 ^ n10140 ;
  assign n41563 = n3773 & ~n9097 ;
  assign n41564 = ( n1208 & n2982 ) | ( n1208 & ~n6753 ) | ( n2982 & ~n6753 ) ;
  assign n41565 = n41564 ^ n36392 ^ n24171 ;
  assign n41566 = ( n2447 & n36313 ) | ( n2447 & ~n41565 ) | ( n36313 & ~n41565 ) ;
  assign n41567 = ( n1011 & n15830 ) | ( n1011 & n41566 ) | ( n15830 & n41566 ) ;
  assign n41568 = n26914 ^ n24793 ^ n17154 ;
  assign n41569 = n38949 ^ n24751 ^ n3543 ;
  assign n41570 = ( ~n9942 & n22803 ) | ( ~n9942 & n30847 ) | ( n22803 & n30847 ) ;
  assign n41571 = n41570 ^ n13420 ^ n479 ;
  assign n41572 = ( n11464 & n36405 ) | ( n11464 & n37946 ) | ( n36405 & n37946 ) ;
  assign n41573 = n41572 ^ n40178 ^ n13440 ;
  assign n41576 = ~n8307 & n14803 ;
  assign n41575 = n1956 | n17075 ;
  assign n41577 = n41576 ^ n41575 ^ 1'b0 ;
  assign n41574 = ( n4566 & ~n18860 ) | ( n4566 & n19804 ) | ( ~n18860 & n19804 ) ;
  assign n41578 = n41577 ^ n41574 ^ n27846 ;
  assign n41579 = ( n19380 & n28752 ) | ( n19380 & ~n28964 ) | ( n28752 & ~n28964 ) ;
  assign n41580 = ( n1507 & n2630 ) | ( n1507 & ~n3084 ) | ( n2630 & ~n3084 ) ;
  assign n41581 = n41580 ^ n13872 ^ n5132 ;
  assign n41582 = ( ~n25287 & n41579 ) | ( ~n25287 & n41581 ) | ( n41579 & n41581 ) ;
  assign n41584 = n29681 ^ n10575 ^ n8418 ;
  assign n41583 = n28915 ^ n23180 ^ n20226 ;
  assign n41585 = n41584 ^ n41583 ^ n10527 ;
  assign n41586 = ( ~n16954 & n24739 ) | ( ~n16954 & n41585 ) | ( n24739 & n41585 ) ;
  assign n41587 = ( n9180 & n20431 ) | ( n9180 & n41586 ) | ( n20431 & n41586 ) ;
  assign n41588 = n11597 ^ n7884 ^ n1112 ;
  assign n41590 = ( ~n1750 & n25645 ) | ( ~n1750 & n35971 ) | ( n25645 & n35971 ) ;
  assign n41589 = n3860 & ~n18771 ;
  assign n41591 = n41590 ^ n41589 ^ 1'b0 ;
  assign n41592 = n37423 ^ n32579 ^ n17726 ;
  assign n41595 = n6497 | n23216 ;
  assign n41596 = ( n11429 & ~n13068 ) | ( n11429 & n41595 ) | ( ~n13068 & n41595 ) ;
  assign n41597 = n41596 ^ n7044 ^ n1358 ;
  assign n41593 = n20825 ^ n13690 ^ n4528 ;
  assign n41594 = n41593 ^ n28651 ^ n10731 ;
  assign n41598 = n41597 ^ n41594 ^ n36850 ;
  assign n41599 = ( ~n274 & n16623 ) | ( ~n274 & n29044 ) | ( n16623 & n29044 ) ;
  assign n41600 = n41599 ^ n28192 ^ n468 ;
  assign n41601 = n36806 ^ n31324 ^ n8435 ;
  assign n41602 = ( ~n18886 & n27885 ) | ( ~n18886 & n41601 ) | ( n27885 & n41601 ) ;
  assign n41603 = n41602 ^ n29997 ^ n29045 ;
  assign n41604 = n41603 ^ n13513 ^ n13201 ;
  assign n41605 = n3690 & n41604 ;
  assign n41606 = n15006 & n41605 ;
  assign n41607 = n5360 | n32556 ;
  assign n41608 = n41607 ^ n26613 ^ 1'b0 ;
  assign n41609 = n15727 ^ n15490 ^ n11958 ;
  assign n41610 = n41609 ^ n1919 ^ x11 ;
  assign n41611 = ( n11579 & n16861 ) | ( n11579 & ~n23918 ) | ( n16861 & ~n23918 ) ;
  assign n41612 = n41611 ^ n29240 ^ n8393 ;
  assign n41613 = ( ~n3905 & n19080 ) | ( ~n3905 & n41612 ) | ( n19080 & n41612 ) ;
  assign n41614 = n25530 ^ n14547 ^ 1'b0 ;
  assign n41615 = n2754 & n41614 ;
  assign n41616 = n41615 ^ n38903 ^ n18948 ;
  assign n41617 = ( n2910 & ~n4393 ) | ( n2910 & n41616 ) | ( ~n4393 & n41616 ) ;
  assign n41618 = ( n5631 & ~n26263 ) | ( n5631 & n27073 ) | ( ~n26263 & n27073 ) ;
  assign n41619 = n41618 ^ n27545 ^ n26916 ;
  assign n41620 = ( n17841 & ~n17925 ) | ( n17841 & n22666 ) | ( ~n17925 & n22666 ) ;
  assign n41621 = n41620 ^ n32927 ^ n14245 ;
  assign n41622 = ( ~n11948 & n12483 ) | ( ~n11948 & n29364 ) | ( n12483 & n29364 ) ;
  assign n41623 = n33465 ^ n22251 ^ 1'b0 ;
  assign n41624 = n21808 & n41623 ;
  assign n41625 = n19766 & n22843 ;
  assign n41626 = n41625 ^ n15816 ^ 1'b0 ;
  assign n41627 = n37866 ^ n7205 ^ 1'b0 ;
  assign n41628 = ~n41626 & n41627 ;
  assign n41629 = ( n323 & n4543 ) | ( n323 & n6650 ) | ( n4543 & n6650 ) ;
  assign n41630 = n41629 ^ n39907 ^ n36513 ;
  assign n41631 = n35318 ^ n6324 ^ n3723 ;
  assign n41632 = n30974 ^ n21368 ^ 1'b0 ;
  assign n41633 = ( n5911 & n28121 ) | ( n5911 & n36218 ) | ( n28121 & n36218 ) ;
  assign n41634 = n10406 | n30916 ;
  assign n41635 = n14249 & ~n41634 ;
  assign n41636 = n19411 & ~n38048 ;
  assign n41637 = n16514 ^ n8623 ^ n4834 ;
  assign n41638 = ( n1396 & n19619 ) | ( n1396 & ~n41637 ) | ( n19619 & ~n41637 ) ;
  assign n41639 = n16762 & ~n32190 ;
  assign n41640 = ~n41638 & n41639 ;
  assign n41641 = ( n6554 & n41636 ) | ( n6554 & ~n41640 ) | ( n41636 & ~n41640 ) ;
  assign n41642 = n30408 ^ n16623 ^ n1557 ;
  assign n41643 = ( n13242 & n29543 ) | ( n13242 & n41642 ) | ( n29543 & n41642 ) ;
  assign n41647 = n6423 | n16545 ;
  assign n41648 = n41647 ^ n6753 ^ 1'b0 ;
  assign n41644 = n20609 ^ n5081 ^ n3376 ;
  assign n41645 = n41644 ^ n12343 ^ n7544 ;
  assign n41646 = n41645 ^ n18511 ^ 1'b0 ;
  assign n41649 = n41648 ^ n41646 ^ n29086 ;
  assign n41650 = n41649 ^ n30403 ^ n1013 ;
  assign n41651 = ( n4352 & n28915 ) | ( n4352 & n38409 ) | ( n28915 & n38409 ) ;
  assign n41652 = n34267 ^ n19639 ^ n4798 ;
  assign n41653 = n23447 & ~n41652 ;
  assign n41654 = n5940 & n41653 ;
  assign n41655 = n41654 ^ n21920 ^ n1819 ;
  assign n41656 = n24386 ^ n15125 ^ 1'b0 ;
  assign n41657 = ( n8614 & n24508 ) | ( n8614 & n38986 ) | ( n24508 & n38986 ) ;
  assign n41658 = ( n2045 & ~n2217 ) | ( n2045 & n21213 ) | ( ~n2217 & n21213 ) ;
  assign n41659 = n41658 ^ n38096 ^ n13957 ;
  assign n41660 = ( n16085 & n21983 ) | ( n16085 & ~n26366 ) | ( n21983 & ~n26366 ) ;
  assign n41662 = n10795 ^ n1912 ^ 1'b0 ;
  assign n41661 = n34606 ^ n21083 ^ 1'b0 ;
  assign n41663 = n41662 ^ n41661 ^ n19796 ;
  assign n41664 = n41660 & ~n41663 ;
  assign n41665 = ( n8568 & n19416 ) | ( n8568 & n34631 ) | ( n19416 & n34631 ) ;
  assign n41666 = n37229 ^ n21176 ^ n12497 ;
  assign n41667 = n41666 ^ n40713 ^ n988 ;
  assign n41668 = n22075 ^ n16035 ^ n4439 ;
  assign n41669 = ( ~n8680 & n9536 ) | ( ~n8680 & n41668 ) | ( n9536 & n41668 ) ;
  assign n41670 = n41181 ^ n31338 ^ n13842 ;
  assign n41671 = ( ~n19602 & n36318 ) | ( ~n19602 & n41670 ) | ( n36318 & n41670 ) ;
  assign n41672 = n5735 & n19700 ;
  assign n41673 = ~n27169 & n41672 ;
  assign n41674 = ( n482 & n5128 ) | ( n482 & n41225 ) | ( n5128 & n41225 ) ;
  assign n41675 = n27667 ^ n11081 ^ n7565 ;
  assign n41676 = n37158 ^ n6499 ^ n2849 ;
  assign n41677 = n41676 ^ n34843 ^ n9459 ;
  assign n41678 = ( n16184 & n16993 ) | ( n16184 & ~n41677 ) | ( n16993 & ~n41677 ) ;
  assign n41679 = n39561 ^ n2229 ^ 1'b0 ;
  assign n41680 = ( n2007 & ~n19357 ) | ( n2007 & n20353 ) | ( ~n19357 & n20353 ) ;
  assign n41681 = n41680 ^ n24680 ^ n16825 ;
  assign n41682 = n25170 & ~n41681 ;
  assign n41683 = ~n8396 & n41682 ;
  assign n41684 = ( n6721 & n39716 ) | ( n6721 & n41683 ) | ( n39716 & n41683 ) ;
  assign n41685 = ( n9585 & ~n22536 ) | ( n9585 & n41684 ) | ( ~n22536 & n41684 ) ;
  assign n41686 = n23854 ^ n17068 ^ 1'b0 ;
  assign n41687 = ( ~n3199 & n25271 ) | ( ~n3199 & n41686 ) | ( n25271 & n41686 ) ;
  assign n41688 = ( n19162 & n33730 ) | ( n19162 & ~n40452 ) | ( n33730 & ~n40452 ) ;
  assign n41689 = ( n1683 & n27927 ) | ( n1683 & n37741 ) | ( n27927 & n37741 ) ;
  assign n41690 = ( n39858 & ~n41688 ) | ( n39858 & n41689 ) | ( ~n41688 & n41689 ) ;
  assign n41691 = n33051 ^ n16243 ^ n12567 ;
  assign n41692 = n41691 ^ n27990 ^ n12418 ;
  assign n41693 = ~n12764 & n20736 ;
  assign n41694 = n41693 ^ n13386 ^ 1'b0 ;
  assign n41696 = ( n415 & ~n19031 ) | ( n415 & n20848 ) | ( ~n19031 & n20848 ) ;
  assign n41695 = n14374 ^ n6118 ^ n5780 ;
  assign n41697 = n41696 ^ n41695 ^ n11973 ;
  assign n41698 = n26826 ^ n5390 ^ n4668 ;
  assign n41699 = ( n14947 & n18119 ) | ( n14947 & n39123 ) | ( n18119 & n39123 ) ;
  assign n41700 = ( ~n6695 & n10893 ) | ( ~n6695 & n37899 ) | ( n10893 & n37899 ) ;
  assign n41701 = ( ~n17026 & n19995 ) | ( ~n17026 & n40776 ) | ( n19995 & n40776 ) ;
  assign n41702 = ( n609 & n16819 ) | ( n609 & n22785 ) | ( n16819 & n22785 ) ;
  assign n41703 = n41702 ^ n37952 ^ n4970 ;
  assign n41704 = ~n3332 & n21871 ;
  assign n41705 = n17943 & ~n18004 ;
  assign n41706 = n41705 ^ n17823 ^ 1'b0 ;
  assign n41707 = n38178 ^ n26362 ^ n11392 ;
  assign n41714 = ( n5467 & n24435 ) | ( n5467 & ~n25610 ) | ( n24435 & ~n25610 ) ;
  assign n41715 = n41714 ^ n8653 ^ n2970 ;
  assign n41712 = ( ~n10275 & n25056 ) | ( ~n10275 & n26466 ) | ( n25056 & n26466 ) ;
  assign n41713 = n41712 ^ n11013 ^ n10850 ;
  assign n41709 = ( n277 & ~n4575 ) | ( n277 & n16963 ) | ( ~n4575 & n16963 ) ;
  assign n41708 = n20512 ^ n17268 ^ n6387 ;
  assign n41710 = n41709 ^ n41708 ^ n20183 ;
  assign n41711 = n41710 ^ n31162 ^ n27382 ;
  assign n41716 = n41715 ^ n41713 ^ n41711 ;
  assign n41717 = ( n921 & ~n5949 ) | ( n921 & n23473 ) | ( ~n5949 & n23473 ) ;
  assign n41718 = n37825 ^ n36454 ^ n29481 ;
  assign n41719 = ( n20062 & n24269 ) | ( n20062 & n41718 ) | ( n24269 & n41718 ) ;
  assign n41720 = ( x114 & n17924 ) | ( x114 & n19684 ) | ( n17924 & n19684 ) ;
  assign n41721 = n1758 & n7148 ;
  assign n41722 = n11553 & n41721 ;
  assign n41723 = ( n423 & ~n34204 ) | ( n423 & n41722 ) | ( ~n34204 & n41722 ) ;
  assign n41724 = n41723 ^ n16358 ^ n14616 ;
  assign n41725 = ( ~n20536 & n41720 ) | ( ~n20536 & n41724 ) | ( n41720 & n41724 ) ;
  assign n41726 = ( n11580 & n38503 ) | ( n11580 & n39751 ) | ( n38503 & n39751 ) ;
  assign n41727 = n27188 ^ n18304 ^ n12821 ;
  assign n41728 = ~n9548 & n33216 ;
  assign n41729 = ~n30682 & n41728 ;
  assign n41732 = n25776 ^ n21916 ^ 1'b0 ;
  assign n41733 = n12528 & n41732 ;
  assign n41730 = n5271 | n22149 ;
  assign n41731 = n41730 ^ n28771 ^ 1'b0 ;
  assign n41734 = n41733 ^ n41731 ^ n22205 ;
  assign n41739 = ( n2021 & n7751 ) | ( n2021 & ~n7841 ) | ( n7751 & ~n7841 ) ;
  assign n41735 = ( n636 & n7736 ) | ( n636 & n8739 ) | ( n7736 & n8739 ) ;
  assign n41736 = n8894 ^ n5974 ^ 1'b0 ;
  assign n41737 = n41735 | n41736 ;
  assign n41738 = ( n12935 & n22160 ) | ( n12935 & n41737 ) | ( n22160 & n41737 ) ;
  assign n41740 = n41739 ^ n41738 ^ n4380 ;
  assign n41741 = n25880 ^ n14394 ^ n6901 ;
  assign n41742 = n18338 ^ n4693 ^ n399 ;
  assign n41743 = n41742 ^ n28891 ^ n5500 ;
  assign n41744 = ( ~n5946 & n9718 ) | ( ~n5946 & n41743 ) | ( n9718 & n41743 ) ;
  assign n41745 = n41502 ^ n7377 ^ n651 ;
  assign n41746 = ( n897 & n9821 ) | ( n897 & n22196 ) | ( n9821 & n22196 ) ;
  assign n41747 = n41746 ^ n30707 ^ n27282 ;
  assign n41748 = n31614 ^ n21700 ^ 1'b0 ;
  assign n41752 = ( ~n1503 & n11559 ) | ( ~n1503 & n19246 ) | ( n11559 & n19246 ) ;
  assign n41749 = n4925 | n24697 ;
  assign n41750 = n27380 ^ n3724 ^ n1021 ;
  assign n41751 = ( ~n1725 & n41749 ) | ( ~n1725 & n41750 ) | ( n41749 & n41750 ) ;
  assign n41753 = n41752 ^ n41751 ^ n1785 ;
  assign n41754 = n31991 & ~n41019 ;
  assign n41755 = n32852 ^ n15798 ^ n14492 ;
  assign n41756 = n27385 ^ n17909 ^ n3720 ;
  assign n41757 = ( ~n257 & n4737 ) | ( ~n257 & n25214 ) | ( n4737 & n25214 ) ;
  assign n41758 = ( n609 & n41756 ) | ( n609 & n41757 ) | ( n41756 & n41757 ) ;
  assign n41759 = n37983 ^ n26705 ^ n12641 ;
  assign n41760 = n41759 ^ n25138 ^ x196 ;
  assign n41761 = ( n35006 & n36496 ) | ( n35006 & ~n41760 ) | ( n36496 & ~n41760 ) ;
  assign n41762 = n10392 ^ n8025 ^ n6605 ;
  assign n41763 = n41762 ^ n30466 ^ n20249 ;
  assign n41764 = n41763 ^ n9547 ^ 1'b0 ;
  assign n41765 = n13312 ^ n8655 ^ 1'b0 ;
  assign n41766 = ( n8687 & n31915 ) | ( n8687 & ~n34002 ) | ( n31915 & ~n34002 ) ;
  assign n41767 = ( n6463 & n41765 ) | ( n6463 & ~n41766 ) | ( n41765 & ~n41766 ) ;
  assign n41768 = n19170 ^ n3290 ^ 1'b0 ;
  assign n41769 = ~n41767 & n41768 ;
  assign n41770 = n22608 ^ n18481 ^ n14618 ;
  assign n41771 = n41770 ^ n8837 ^ 1'b0 ;
  assign n41772 = n6344 & n41771 ;
  assign n41773 = ( n1424 & ~n7281 ) | ( n1424 & n7383 ) | ( ~n7281 & n7383 ) ;
  assign n41774 = ( n4863 & n19752 ) | ( n4863 & ~n39130 ) | ( n19752 & ~n39130 ) ;
  assign n41775 = ( n34088 & n41773 ) | ( n34088 & ~n41774 ) | ( n41773 & ~n41774 ) ;
  assign n41776 = n24507 ^ n5886 ^ n802 ;
  assign n41777 = n29382 | n41776 ;
  assign n41778 = n41777 ^ n30545 ^ 1'b0 ;
  assign n41779 = n41778 ^ n11406 ^ 1'b0 ;
  assign n41780 = ( n4673 & n5943 ) | ( n4673 & n19534 ) | ( n5943 & n19534 ) ;
  assign n41781 = ( n12097 & ~n22030 ) | ( n12097 & n41780 ) | ( ~n22030 & n41780 ) ;
  assign n41782 = ( n15937 & n25846 ) | ( n15937 & ~n41781 ) | ( n25846 & ~n41781 ) ;
  assign n41783 = ( n19137 & n22505 ) | ( n19137 & n38610 ) | ( n22505 & n38610 ) ;
  assign n41784 = n41783 ^ n25695 ^ n18750 ;
  assign n41785 = n11124 ^ n10241 ^ n1678 ;
  assign n41786 = n41785 ^ n22997 ^ n21438 ;
  assign n41787 = n26897 ^ n12006 ^ n5739 ;
  assign n41788 = n32960 ^ n21989 ^ 1'b0 ;
  assign n41789 = n41787 | n41788 ;
  assign n41790 = n14555 ^ n10756 ^ n8897 ;
  assign n41791 = n25477 ^ n18333 ^ 1'b0 ;
  assign n41792 = ( n22173 & n35709 ) | ( n22173 & n41791 ) | ( n35709 & n41791 ) ;
  assign n41793 = ( n12401 & n14459 ) | ( n12401 & n17414 ) | ( n14459 & n17414 ) ;
  assign n41794 = n17333 ^ n1845 ^ n1431 ;
  assign n41795 = ( x43 & ~n14474 ) | ( x43 & n15982 ) | ( ~n14474 & n15982 ) ;
  assign n41796 = ( n7064 & n13520 ) | ( n7064 & n41795 ) | ( n13520 & n41795 ) ;
  assign n41797 = n3127 & n41215 ;
  assign n41798 = n41797 ^ n30660 ^ n23023 ;
  assign n41799 = n40044 ^ n3056 ^ 1'b0 ;
  assign n41802 = n19818 ^ n6906 ^ n3347 ;
  assign n41803 = ( n15510 & n29917 ) | ( n15510 & n41802 ) | ( n29917 & n41802 ) ;
  assign n41800 = n39562 ^ n473 ^ 1'b0 ;
  assign n41801 = n16103 & n41800 ;
  assign n41804 = n41803 ^ n41801 ^ n28676 ;
  assign n41805 = ( n1752 & ~n19376 ) | ( n1752 & n24032 ) | ( ~n19376 & n24032 ) ;
  assign n41806 = n41805 ^ n27550 ^ n20076 ;
  assign n41807 = n38147 ^ n29521 ^ n3914 ;
  assign n41811 = n12883 & n31547 ;
  assign n41808 = n10374 | n21164 ;
  assign n41809 = n41808 ^ n22741 ^ 1'b0 ;
  assign n41810 = n41809 ^ n38217 ^ n5942 ;
  assign n41812 = n41811 ^ n41810 ^ n36609 ;
  assign n41813 = ( n2865 & ~n4113 ) | ( n2865 & n11773 ) | ( ~n4113 & n11773 ) ;
  assign n41814 = n2392 | n29684 ;
  assign n41815 = n41813 & ~n41814 ;
  assign n41816 = n34568 ^ n12376 ^ n850 ;
  assign n41817 = n41816 ^ n40758 ^ n7513 ;
  assign n41818 = n32755 ^ n29853 ^ n14278 ;
  assign n41819 = ( n661 & n7844 ) | ( n661 & ~n34848 ) | ( n7844 & ~n34848 ) ;
  assign n41820 = n35642 ^ n11314 ^ 1'b0 ;
  assign n41821 = n18882 ^ n6151 ^ 1'b0 ;
  assign n41822 = n41821 ^ n30230 ^ n15201 ;
  assign n41823 = ( n16748 & ~n41820 ) | ( n16748 & n41822 ) | ( ~n41820 & n41822 ) ;
  assign n41824 = n41823 ^ n11043 ^ n6525 ;
  assign n41825 = n41612 ^ n2374 ^ 1'b0 ;
  assign n41826 = ( n9008 & n18584 ) | ( n9008 & n22095 ) | ( n18584 & n22095 ) ;
  assign n41827 = ( n4457 & n37141 ) | ( n4457 & n41826 ) | ( n37141 & n41826 ) ;
  assign n41828 = ( n16271 & n31381 ) | ( n16271 & n41827 ) | ( n31381 & n41827 ) ;
  assign n41829 = n41828 ^ n30936 ^ n18993 ;
  assign n41830 = n5596 & n22691 ;
  assign n41831 = ( n551 & n13301 ) | ( n551 & ~n21063 ) | ( n13301 & ~n21063 ) ;
  assign n41834 = n26371 ^ n12098 ^ n5760 ;
  assign n41832 = ( n14604 & ~n18943 ) | ( n14604 & n29883 ) | ( ~n18943 & n29883 ) ;
  assign n41833 = n41832 ^ n34826 ^ n19039 ;
  assign n41835 = n41834 ^ n41833 ^ n17157 ;
  assign n41836 = n11871 & n12672 ;
  assign n41837 = ~n15886 & n41836 ;
  assign n41838 = n28979 ^ n15144 ^ n3251 ;
  assign n41839 = ( n11448 & n34642 ) | ( n11448 & n41838 ) | ( n34642 & n41838 ) ;
  assign n41840 = n37243 & n39954 ;
  assign n41841 = ( n2071 & ~n14396 ) | ( n2071 & n27868 ) | ( ~n14396 & n27868 ) ;
  assign n41843 = ( n11264 & n16150 ) | ( n11264 & n28550 ) | ( n16150 & n28550 ) ;
  assign n41842 = n5189 & n34437 ;
  assign n41844 = n41843 ^ n41842 ^ 1'b0 ;
  assign n41845 = n23366 & ~n41844 ;
  assign n41847 = n18385 ^ n2777 ^ n990 ;
  assign n41846 = ~n3597 & n18584 ;
  assign n41848 = n41847 ^ n41846 ^ 1'b0 ;
  assign n41849 = n20095 ^ x68 ^ 1'b0 ;
  assign n41850 = n30586 ^ n7283 ^ 1'b0 ;
  assign n41851 = ( n394 & n35786 ) | ( n394 & ~n41850 ) | ( n35786 & ~n41850 ) ;
  assign n41852 = n25966 ^ n12290 ^ n10198 ;
  assign n41853 = ( ~n7824 & n14449 ) | ( ~n7824 & n14783 ) | ( n14449 & n14783 ) ;
  assign n41854 = ( n8463 & n18170 ) | ( n8463 & ~n41853 ) | ( n18170 & ~n41853 ) ;
  assign n41855 = ( ~n24110 & n26306 ) | ( ~n24110 & n41854 ) | ( n26306 & n41854 ) ;
  assign n41856 = n23789 ^ n15561 ^ n4148 ;
  assign n41857 = n41856 ^ n9107 ^ 1'b0 ;
  assign n41860 = ( n4415 & ~n5931 ) | ( n4415 & n9707 ) | ( ~n5931 & n9707 ) ;
  assign n41858 = ( ~n475 & n14551 ) | ( ~n475 & n33668 ) | ( n14551 & n33668 ) ;
  assign n41859 = ( n12535 & n20809 ) | ( n12535 & ~n41858 ) | ( n20809 & ~n41858 ) ;
  assign n41861 = n41860 ^ n41859 ^ n30699 ;
  assign n41867 = n18996 ^ n12551 ^ n7337 ;
  assign n41862 = ( ~n4962 & n11510 ) | ( ~n4962 & n39995 ) | ( n11510 & n39995 ) ;
  assign n41863 = ~n5019 & n16469 ;
  assign n41864 = n13010 | n41863 ;
  assign n41865 = n24220 ^ n16542 ^ n14019 ;
  assign n41866 = ( n41862 & ~n41864 ) | ( n41862 & n41865 ) | ( ~n41864 & n41865 ) ;
  assign n41868 = n41867 ^ n41866 ^ n19796 ;
  assign n41869 = n21030 ^ n20776 ^ 1'b0 ;
  assign n41870 = n30298 ^ n12965 ^ n3372 ;
  assign n41871 = n23631 ^ n10784 ^ n6594 ;
  assign n41872 = ~n28705 & n41871 ;
  assign n41873 = n41872 ^ n40850 ^ 1'b0 ;
  assign n41874 = n17844 | n27309 ;
  assign n41875 = n31373 ^ n14197 ^ n11595 ;
  assign n41876 = ( n11118 & n30329 ) | ( n11118 & n41875 ) | ( n30329 & n41875 ) ;
  assign n41877 = n29506 & ~n41876 ;
  assign n41878 = ( n16101 & ~n33047 ) | ( n16101 & n41877 ) | ( ~n33047 & n41877 ) ;
  assign n41879 = ( ~n11933 & n14174 ) | ( ~n11933 & n16027 ) | ( n14174 & n16027 ) ;
  assign n41880 = ( x35 & ~n5545 ) | ( x35 & n16641 ) | ( ~n5545 & n16641 ) ;
  assign n41881 = n20022 | n41880 ;
  assign n41882 = ~n8726 & n13210 ;
  assign n41883 = n41882 ^ n11037 ^ 1'b0 ;
  assign n41884 = n5806 & n41883 ;
  assign n41885 = n41884 ^ n36913 ^ 1'b0 ;
  assign n41886 = n11333 ^ n1302 ^ 1'b0 ;
  assign n41887 = n15363 | n41886 ;
  assign n41888 = n22730 ^ n18488 ^ n8114 ;
  assign n41889 = ( n16478 & ~n37124 ) | ( n16478 & n41888 ) | ( ~n37124 & n41888 ) ;
  assign n41890 = n30351 ^ n27012 ^ n14262 ;
  assign n41891 = ( n3790 & n26664 ) | ( n3790 & n41890 ) | ( n26664 & n41890 ) ;
  assign n41892 = n24547 ^ n20379 ^ n7150 ;
  assign n41893 = n41892 ^ n31812 ^ n7547 ;
  assign n41895 = n22786 ^ n11003 ^ n10744 ;
  assign n41894 = ( n1880 & n21651 ) | ( n1880 & n22399 ) | ( n21651 & n22399 ) ;
  assign n41896 = n41895 ^ n41894 ^ n2221 ;
  assign n41897 = n16175 ^ n5348 ^ 1'b0 ;
  assign n41898 = n6208 | n41897 ;
  assign n41899 = ( ~n9244 & n41896 ) | ( ~n9244 & n41898 ) | ( n41896 & n41898 ) ;
  assign n41900 = n39086 ^ n23182 ^ n6067 ;
  assign n41901 = ( n12558 & n13926 ) | ( n12558 & n41900 ) | ( n13926 & n41900 ) ;
  assign n41902 = n40566 ^ n38035 ^ n718 ;
  assign n41903 = ( n1396 & n6789 ) | ( n1396 & n38827 ) | ( n6789 & n38827 ) ;
  assign n41904 = n6417 | n7908 ;
  assign n41905 = n31592 ^ n27400 ^ n15314 ;
  assign n41906 = n41905 ^ n20674 ^ n10144 ;
  assign n41907 = n19337 ^ n1570 ^ 1'b0 ;
  assign n41908 = n41907 ^ n14909 ^ n13777 ;
  assign n41909 = n19939 ^ n8857 ^ 1'b0 ;
  assign n41910 = n23650 ^ n17197 ^ 1'b0 ;
  assign n41911 = n24119 ^ n3261 ^ n3234 ;
  assign n41912 = n27691 ^ n14625 ^ n6115 ;
  assign n41913 = n41912 ^ n9109 ^ n1948 ;
  assign n41914 = n5156 & n37439 ;
  assign n41915 = n33759 & n41914 ;
  assign n41916 = n41915 ^ n41425 ^ n4284 ;
  assign n41917 = n41916 ^ n2762 ^ n1866 ;
  assign n41918 = ( n2140 & ~n25390 ) | ( n2140 & n40869 ) | ( ~n25390 & n40869 ) ;
  assign n41920 = n13630 | n13916 ;
  assign n41921 = n8230 & ~n41920 ;
  assign n41922 = n41921 ^ n27478 ^ n20896 ;
  assign n41919 = n13131 & n18735 ;
  assign n41923 = n41922 ^ n41919 ^ n5817 ;
  assign n41924 = n8753 | n32756 ;
  assign n41925 = n41924 ^ n36814 ^ n17902 ;
  assign n41926 = n41923 & ~n41925 ;
  assign n41927 = ~n5643 & n14807 ;
  assign n41928 = ~n31039 & n41927 ;
  assign n41929 = n41928 ^ n21804 ^ n10359 ;
  assign n41930 = n36536 ^ n15115 ^ n10192 ;
  assign n41931 = ( n6150 & n25468 ) | ( n6150 & ~n41930 ) | ( n25468 & ~n41930 ) ;
  assign n41932 = n40426 ^ n21563 ^ n18750 ;
  assign n41933 = n23741 ^ n16188 ^ n10038 ;
  assign n41934 = n23368 ^ n18679 ^ 1'b0 ;
  assign n41935 = ~n41933 & n41934 ;
  assign n41937 = n16965 ^ n6137 ^ n4677 ;
  assign n41938 = n6521 & n14945 ;
  assign n41939 = n41938 ^ n3184 ^ 1'b0 ;
  assign n41940 = n41939 ^ n5314 ^ 1'b0 ;
  assign n41941 = n41937 & ~n41940 ;
  assign n41936 = ~n6238 & n39297 ;
  assign n41942 = n41941 ^ n41936 ^ 1'b0 ;
  assign n41943 = ( n2585 & n6539 ) | ( n2585 & n12264 ) | ( n6539 & n12264 ) ;
  assign n41944 = ( n25303 & n40706 ) | ( n25303 & n41943 ) | ( n40706 & n41943 ) ;
  assign n41945 = n6492 ^ n2155 ^ n1392 ;
  assign n41946 = ( n2599 & n16034 ) | ( n2599 & n41945 ) | ( n16034 & n41945 ) ;
  assign n41947 = n12484 ^ n2976 ^ n1286 ;
  assign n41948 = ( n27372 & n32792 ) | ( n27372 & ~n41947 ) | ( n32792 & ~n41947 ) ;
  assign n41949 = ( n9682 & n41946 ) | ( n9682 & ~n41948 ) | ( n41946 & ~n41948 ) ;
  assign n41950 = ( n13088 & ~n25180 ) | ( n13088 & n31570 ) | ( ~n25180 & n31570 ) ;
  assign n41951 = n41950 ^ n36959 ^ n35733 ;
  assign n41952 = ( n6770 & n13088 ) | ( n6770 & n16984 ) | ( n13088 & n16984 ) ;
  assign n41953 = n21782 ^ n8347 ^ 1'b0 ;
  assign n41954 = ~n13503 & n41953 ;
  assign n41955 = ( n1497 & n14702 ) | ( n1497 & n41954 ) | ( n14702 & n41954 ) ;
  assign n41956 = ( n22345 & n27445 ) | ( n22345 & ~n41955 ) | ( n27445 & ~n41955 ) ;
  assign n41957 = n41956 ^ n16152 ^ n8768 ;
  assign n41958 = n41957 ^ n25207 ^ n12481 ;
  assign n41960 = ~n6476 & n20699 ;
  assign n41961 = n41960 ^ n8157 ^ 1'b0 ;
  assign n41959 = n32093 ^ n13314 ^ n9175 ;
  assign n41962 = n41961 ^ n41959 ^ n30338 ;
  assign n41963 = n2705 | n19875 ;
  assign n41964 = n41963 ^ n25127 ^ n15876 ;
  assign n41967 = n17634 ^ n6767 ^ n2918 ;
  assign n41965 = n33502 ^ n17829 ^ 1'b0 ;
  assign n41966 = n33956 | n41965 ;
  assign n41968 = n41967 ^ n41966 ^ n36356 ;
  assign n41969 = ( n41962 & n41964 ) | ( n41962 & n41968 ) | ( n41964 & n41968 ) ;
  assign n41970 = n16722 & n18442 ;
  assign n41971 = n41970 ^ n7925 ^ 1'b0 ;
  assign n41972 = n29573 ^ n18614 ^ n6242 ;
  assign n41973 = ( n16793 & n25839 ) | ( n16793 & n41972 ) | ( n25839 & n41972 ) ;
  assign n41974 = n41971 | n41973 ;
  assign n41975 = ( n3487 & n22888 ) | ( n3487 & ~n24002 ) | ( n22888 & ~n24002 ) ;
  assign n41976 = ( ~n9833 & n17933 ) | ( ~n9833 & n25952 ) | ( n17933 & n25952 ) ;
  assign n41977 = n8793 & n9392 ;
  assign n41978 = n41977 ^ n6894 ^ 1'b0 ;
  assign n41979 = n41978 ^ n8610 ^ n1615 ;
  assign n41980 = ( n24395 & n28832 ) | ( n24395 & ~n41979 ) | ( n28832 & ~n41979 ) ;
  assign n41981 = ~n41976 & n41980 ;
  assign n41982 = n41975 & n41981 ;
  assign n41983 = ( n3628 & n4068 ) | ( n3628 & n22117 ) | ( n4068 & n22117 ) ;
  assign n41984 = n37752 ^ n13563 ^ n5512 ;
  assign n41985 = ( n4016 & ~n13973 ) | ( n4016 & n17642 ) | ( ~n13973 & n17642 ) ;
  assign n41986 = ( ~n17642 & n41984 ) | ( ~n17642 & n41985 ) | ( n41984 & n41985 ) ;
  assign n41987 = n8616 | n28137 ;
  assign n41988 = n7177 & ~n41987 ;
  assign n41989 = ( n2190 & n9606 ) | ( n2190 & ~n16059 ) | ( n9606 & ~n16059 ) ;
  assign n41990 = ( n1668 & n15932 ) | ( n1668 & n41989 ) | ( n15932 & n41989 ) ;
  assign n41991 = ( n6262 & n41988 ) | ( n6262 & ~n41990 ) | ( n41988 & ~n41990 ) ;
  assign n41992 = n13340 ^ n2082 ^ n618 ;
  assign n41993 = n41992 ^ n19904 ^ n9878 ;
  assign n41996 = ( n3920 & n6464 ) | ( n3920 & n24733 ) | ( n6464 & n24733 ) ;
  assign n41997 = ( n25781 & n37839 ) | ( n25781 & ~n41996 ) | ( n37839 & ~n41996 ) ;
  assign n41994 = ( n732 & ~n14229 ) | ( n732 & n20728 ) | ( ~n14229 & n20728 ) ;
  assign n41995 = ( ~n15374 & n23088 ) | ( ~n15374 & n41994 ) | ( n23088 & n41994 ) ;
  assign n41998 = n41997 ^ n41995 ^ n30220 ;
  assign n41999 = n19076 ^ n8388 ^ 1'b0 ;
  assign n42000 = ( n18584 & n23057 ) | ( n18584 & ~n41999 ) | ( n23057 & ~n41999 ) ;
  assign n42001 = n40525 ^ n20086 ^ n18734 ;
  assign n42002 = n9012 ^ n5540 ^ n1746 ;
  assign n42003 = n42002 ^ n25065 ^ n4897 ;
  assign n42004 = n17629 & ~n42003 ;
  assign n42005 = ( n7000 & n7531 ) | ( n7000 & ~n13617 ) | ( n7531 & ~n13617 ) ;
  assign n42006 = ( n17874 & ~n20690 ) | ( n17874 & n25114 ) | ( ~n20690 & n25114 ) ;
  assign n42007 = ( n619 & ~n42005 ) | ( n619 & n42006 ) | ( ~n42005 & n42006 ) ;
  assign n42009 = n28692 ^ n19650 ^ 1'b0 ;
  assign n42010 = ( ~n1748 & n41191 ) | ( ~n1748 & n42009 ) | ( n41191 & n42009 ) ;
  assign n42008 = n26744 ^ n19806 ^ n10199 ;
  assign n42011 = n42010 ^ n42008 ^ n10449 ;
  assign n42012 = ( n6017 & n13950 ) | ( n6017 & n21449 ) | ( n13950 & n21449 ) ;
  assign n42013 = n21227 ^ n15520 ^ n11315 ;
  assign n42014 = ( ~n4209 & n6842 ) | ( ~n4209 & n9317 ) | ( n6842 & n9317 ) ;
  assign n42015 = ( n6883 & n10067 ) | ( n6883 & n42014 ) | ( n10067 & n42014 ) ;
  assign n42016 = n17010 ^ n10512 ^ n9570 ;
  assign n42017 = n42016 ^ n41967 ^ x89 ;
  assign n42018 = n42017 ^ n9406 ^ 1'b0 ;
  assign n42019 = ( ~n13513 & n16058 ) | ( ~n13513 & n41152 ) | ( n16058 & n41152 ) ;
  assign n42020 = n16326 ^ n8829 ^ n6223 ;
  assign n42021 = ( ~n6715 & n36957 ) | ( ~n6715 & n42020 ) | ( n36957 & n42020 ) ;
  assign n42022 = n40806 ^ n37733 ^ n7707 ;
  assign n42023 = n36191 ^ n17037 ^ n3278 ;
  assign n42024 = n27707 ^ n26498 ^ n12688 ;
  assign n42025 = ( n34405 & n42023 ) | ( n34405 & ~n42024 ) | ( n42023 & ~n42024 ) ;
  assign n42026 = ( n751 & ~n42022 ) | ( n751 & n42025 ) | ( ~n42022 & n42025 ) ;
  assign n42029 = n30398 ^ n9653 ^ n6844 ;
  assign n42027 = n12712 ^ n6413 ^ x185 ;
  assign n42028 = ( ~n3076 & n26902 ) | ( ~n3076 & n42027 ) | ( n26902 & n42027 ) ;
  assign n42030 = n42029 ^ n42028 ^ n24936 ;
  assign n42031 = ( n15805 & n17531 ) | ( n15805 & n31644 ) | ( n17531 & n31644 ) ;
  assign n42032 = n9385 & n19763 ;
  assign n42033 = n8680 & n42032 ;
  assign n42034 = ( n2035 & n42031 ) | ( n2035 & ~n42033 ) | ( n42031 & ~n42033 ) ;
  assign n42037 = x100 & ~n36397 ;
  assign n42038 = n25442 & n42037 ;
  assign n42035 = ( n535 & n13947 ) | ( n535 & n37592 ) | ( n13947 & n37592 ) ;
  assign n42036 = ( x28 & n8918 ) | ( x28 & ~n42035 ) | ( n8918 & ~n42035 ) ;
  assign n42039 = n42038 ^ n42036 ^ n24447 ;
  assign n42040 = ( n1921 & n8431 ) | ( n1921 & n9221 ) | ( n8431 & n9221 ) ;
  assign n42041 = n41168 ^ n15284 ^ 1'b0 ;
  assign n42042 = n14797 & ~n42041 ;
  assign n42043 = n12930 ^ n10524 ^ n487 ;
  assign n42044 = n42043 ^ n27744 ^ n24876 ;
  assign n42045 = n30297 ^ n9646 ^ 1'b0 ;
  assign n42046 = ( n13679 & n19937 ) | ( n13679 & ~n42045 ) | ( n19937 & ~n42045 ) ;
  assign n42047 = n42044 | n42046 ;
  assign n42048 = ( ~n4793 & n16654 ) | ( ~n4793 & n27556 ) | ( n16654 & n27556 ) ;
  assign n42049 = ( n4414 & n12901 ) | ( n4414 & ~n42048 ) | ( n12901 & ~n42048 ) ;
  assign n42050 = ( n28183 & ~n29754 ) | ( n28183 & n36671 ) | ( ~n29754 & n36671 ) ;
  assign n42051 = ( n9186 & n42049 ) | ( n9186 & ~n42050 ) | ( n42049 & ~n42050 ) ;
  assign n42052 = n12571 ^ n12365 ^ n1851 ;
  assign n42053 = n42052 ^ n37967 ^ n726 ;
  assign n42054 = ( n5237 & ~n8869 ) | ( n5237 & n15014 ) | ( ~n8869 & n15014 ) ;
  assign n42055 = ( ~n654 & n30951 ) | ( ~n654 & n42054 ) | ( n30951 & n42054 ) ;
  assign n42056 = n6625 ^ n6034 ^ n5279 ;
  assign n42057 = n42056 ^ n33165 ^ n12435 ;
  assign n42058 = n29908 ^ n13521 ^ n608 ;
  assign n42059 = n25482 ^ n24613 ^ n3339 ;
  assign n42060 = ~n4389 & n42059 ;
  assign n42061 = ( ~n30370 & n34442 ) | ( ~n30370 & n38989 ) | ( n34442 & n38989 ) ;
  assign n42062 = ( n2258 & ~n12204 ) | ( n2258 & n26310 ) | ( ~n12204 & n26310 ) ;
  assign n42063 = ( n30872 & n34264 ) | ( n30872 & n42062 ) | ( n34264 & n42062 ) ;
  assign n42064 = ( n16416 & ~n42061 ) | ( n16416 & n42063 ) | ( ~n42061 & n42063 ) ;
  assign n42065 = n27178 ^ n4854 ^ 1'b0 ;
  assign n42066 = n5095 | n42065 ;
  assign n42067 = n42066 ^ n23463 ^ n16021 ;
  assign n42068 = ( n3920 & n11493 ) | ( n3920 & n42067 ) | ( n11493 & n42067 ) ;
  assign n42069 = n29282 ^ n9449 ^ n3543 ;
  assign n42070 = n3950 & n42069 ;
  assign n42071 = n42070 ^ n6845 ^ 1'b0 ;
  assign n42072 = n31406 ^ n21292 ^ 1'b0 ;
  assign n42073 = n13716 ^ n5754 ^ 1'b0 ;
  assign n42077 = n21097 ^ n7732 ^ n7457 ;
  assign n42075 = ( ~n9896 & n31335 ) | ( ~n9896 & n32889 ) | ( n31335 & n32889 ) ;
  assign n42074 = n7414 & ~n20240 ;
  assign n42076 = n42075 ^ n42074 ^ 1'b0 ;
  assign n42078 = n42077 ^ n42076 ^ 1'b0 ;
  assign n42079 = ( n14966 & n21672 ) | ( n14966 & n42078 ) | ( n21672 & n42078 ) ;
  assign n42080 = ( ~n15665 & n27380 ) | ( ~n15665 & n30346 ) | ( n27380 & n30346 ) ;
  assign n42081 = n42080 ^ n29501 ^ n10230 ;
  assign n42082 = n21044 | n22507 ;
  assign n42083 = ( n9301 & n26461 ) | ( n9301 & n27663 ) | ( n26461 & n27663 ) ;
  assign n42084 = ( n542 & ~n31774 ) | ( n542 & n42083 ) | ( ~n31774 & n42083 ) ;
  assign n42085 = n37797 ^ n12777 ^ x229 ;
  assign n42086 = ( n17989 & ~n28384 ) | ( n17989 & n37816 ) | ( ~n28384 & n37816 ) ;
  assign n42087 = n4288 | n42086 ;
  assign n42088 = n25427 ^ n10548 ^ 1'b0 ;
  assign n42089 = n7287 & n15358 ;
  assign n42090 = n42089 ^ n40305 ^ n10077 ;
  assign n42091 = ( n2157 & n36263 ) | ( n2157 & ~n42090 ) | ( n36263 & ~n42090 ) ;
  assign n42092 = n12616 | n40404 ;
  assign n42093 = n42092 ^ n35832 ^ 1'b0 ;
  assign n42094 = ( n9873 & n27838 ) | ( n9873 & ~n40709 ) | ( n27838 & ~n40709 ) ;
  assign n42095 = ( n14306 & n17872 ) | ( n14306 & ~n21383 ) | ( n17872 & ~n21383 ) ;
  assign n42096 = ( n7786 & ~n16648 ) | ( n7786 & n36450 ) | ( ~n16648 & n36450 ) ;
  assign n42097 = n30962 & n34615 ;
  assign n42101 = n19050 ^ n3515 ^ n1057 ;
  assign n42098 = n13284 ^ n4307 ^ n3134 ;
  assign n42099 = ( n1397 & n11382 ) | ( n1397 & ~n42098 ) | ( n11382 & ~n42098 ) ;
  assign n42100 = ( n8312 & ~n21833 ) | ( n8312 & n42099 ) | ( ~n21833 & n42099 ) ;
  assign n42102 = n42101 ^ n42100 ^ n25273 ;
  assign n42103 = n7706 ^ n6162 ^ n4289 ;
  assign n42104 = ( ~n7483 & n13051 ) | ( ~n7483 & n34422 ) | ( n13051 & n34422 ) ;
  assign n42105 = n26447 ^ n20930 ^ n9469 ;
  assign n42106 = n42105 ^ n40685 ^ n9535 ;
  assign n42107 = n19256 ^ n5013 ^ n613 ;
  assign n42108 = ( n508 & n36941 ) | ( n508 & ~n38054 ) | ( n36941 & ~n38054 ) ;
  assign n42109 = ( n27727 & ~n42003 ) | ( n27727 & n42108 ) | ( ~n42003 & n42108 ) ;
  assign n42110 = n33433 ^ n20268 ^ n10458 ;
  assign n42111 = ~n27172 & n29675 ;
  assign n42112 = ( n3881 & n17044 ) | ( n3881 & n18362 ) | ( n17044 & n18362 ) ;
  assign n42113 = ( ~n11021 & n26836 ) | ( ~n11021 & n31211 ) | ( n26836 & n31211 ) ;
  assign n42114 = ( ~n21025 & n31028 ) | ( ~n21025 & n42113 ) | ( n31028 & n42113 ) ;
  assign n42115 = ( n6293 & n22904 ) | ( n6293 & ~n42114 ) | ( n22904 & ~n42114 ) ;
  assign n42116 = ( n4203 & n36224 ) | ( n4203 & n42115 ) | ( n36224 & n42115 ) ;
  assign n42119 = n19583 ^ n19123 ^ n15126 ;
  assign n42117 = n4449 & n21451 ;
  assign n42118 = ~n21978 & n42117 ;
  assign n42120 = n42119 ^ n42118 ^ n32384 ;
  assign n42121 = n37559 ^ n24468 ^ n12323 ;
  assign n42122 = ( n8822 & n13894 ) | ( n8822 & ~n36083 ) | ( n13894 & ~n36083 ) ;
  assign n42123 = n22222 ^ n22163 ^ n19926 ;
  assign n42124 = ( ~n4223 & n42122 ) | ( ~n4223 & n42123 ) | ( n42122 & n42123 ) ;
  assign n42125 = n2190 & n34157 ;
  assign n42126 = ( n11852 & n27177 ) | ( n11852 & n29131 ) | ( n27177 & n29131 ) ;
  assign n42127 = n21043 ^ n15357 ^ n321 ;
  assign n42128 = ( n42125 & n42126 ) | ( n42125 & ~n42127 ) | ( n42126 & ~n42127 ) ;
  assign n42129 = ( n2243 & ~n11078 ) | ( n2243 & n28837 ) | ( ~n11078 & n28837 ) ;
  assign n42130 = n26144 ^ n9462 ^ 1'b0 ;
  assign n42131 = n38575 ^ n10323 ^ n1368 ;
  assign n42132 = n42131 ^ n38920 ^ n21388 ;
  assign n42133 = n25361 | n40866 ;
  assign n42134 = n5006 | n42133 ;
  assign n42135 = ( n11619 & n16610 ) | ( n11619 & ~n42134 ) | ( n16610 & ~n42134 ) ;
  assign n42136 = n7431 & ~n29181 ;
  assign n42137 = n42135 & n42136 ;
  assign n42138 = ( n42130 & n42132 ) | ( n42130 & n42137 ) | ( n42132 & n42137 ) ;
  assign n42139 = n30767 ^ n24114 ^ n7956 ;
  assign n42140 = ( n6988 & ~n23486 ) | ( n6988 & n37882 ) | ( ~n23486 & n37882 ) ;
  assign n42141 = n25996 ^ n22265 ^ n18665 ;
  assign n42142 = n42140 & ~n42141 ;
  assign n42143 = ( n3035 & ~n11053 ) | ( n3035 & n14820 ) | ( ~n11053 & n14820 ) ;
  assign n42144 = n42143 ^ n25130 ^ 1'b0 ;
  assign n42145 = ( ~n1001 & n4520 ) | ( ~n1001 & n39478 ) | ( n4520 & n39478 ) ;
  assign n42146 = n42145 ^ n31219 ^ n18503 ;
  assign n42147 = ( n5310 & n21714 ) | ( n5310 & n24260 ) | ( n21714 & n24260 ) ;
  assign n42148 = ( n12278 & ~n24994 ) | ( n12278 & n42147 ) | ( ~n24994 & n42147 ) ;
  assign n42149 = ( n21925 & n27287 ) | ( n21925 & n42148 ) | ( n27287 & n42148 ) ;
  assign n42150 = ( ~n17684 & n21636 ) | ( ~n17684 & n42149 ) | ( n21636 & n42149 ) ;
  assign n42151 = n42150 ^ n35741 ^ n11783 ;
  assign n42152 = n20013 & ~n22252 ;
  assign n42153 = ( n3451 & ~n18244 ) | ( n3451 & n24672 ) | ( ~n18244 & n24672 ) ;
  assign n42154 = n42153 ^ n2391 ^ 1'b0 ;
  assign n42155 = n42154 ^ n6589 ^ 1'b0 ;
  assign n42156 = n42152 | n42155 ;
  assign n42157 = ( n1901 & ~n29123 ) | ( n1901 & n34869 ) | ( ~n29123 & n34869 ) ;
  assign n42158 = n27911 ^ n680 ^ 1'b0 ;
  assign n42159 = n10796 & ~n42158 ;
  assign n42160 = ( n5228 & ~n30552 ) | ( n5228 & n42159 ) | ( ~n30552 & n42159 ) ;
  assign n42161 = ( n23184 & ~n23730 ) | ( n23184 & n32527 ) | ( ~n23730 & n32527 ) ;
  assign n42162 = ( ~n9481 & n13368 ) | ( ~n9481 & n36913 ) | ( n13368 & n36913 ) ;
  assign n42163 = ( ~n19315 & n32282 ) | ( ~n19315 & n42162 ) | ( n32282 & n42162 ) ;
  assign n42164 = ( n13740 & ~n42161 ) | ( n13740 & n42163 ) | ( ~n42161 & n42163 ) ;
  assign n42170 = n12111 ^ n9029 ^ n3790 ;
  assign n42167 = ( ~n5746 & n13850 ) | ( ~n5746 & n22070 ) | ( n13850 & n22070 ) ;
  assign n42168 = n42167 ^ n21687 ^ n1334 ;
  assign n42169 = n42168 ^ n34453 ^ n14019 ;
  assign n42165 = n7332 ^ n5896 ^ n4671 ;
  assign n42166 = n42165 ^ n26788 ^ n4954 ;
  assign n42171 = n42170 ^ n42169 ^ n42166 ;
  assign n42172 = n20586 ^ n11130 ^ n2568 ;
  assign n42173 = n30227 ^ n27370 ^ n16158 ;
  assign n42174 = n42173 ^ n9927 ^ n8115 ;
  assign n42175 = ( ~n5302 & n42172 ) | ( ~n5302 & n42174 ) | ( n42172 & n42174 ) ;
  assign n42176 = n42175 ^ n41939 ^ n28538 ;
  assign n42177 = n29242 ^ n4214 ^ x113 ;
  assign n42178 = n22091 ^ n9664 ^ n4128 ;
  assign n42179 = n3982 & n42178 ;
  assign n42180 = ( ~n5787 & n17519 ) | ( ~n5787 & n36646 ) | ( n17519 & n36646 ) ;
  assign n42181 = n25590 & n42180 ;
  assign n42182 = n16271 ^ n9644 ^ n6022 ;
  assign n42183 = n42182 ^ n37438 ^ n4434 ;
  assign n42184 = n42183 ^ n25422 ^ 1'b0 ;
  assign n42185 = n42181 & ~n42184 ;
  assign n42186 = n26471 | n30978 ;
  assign n42187 = n42186 ^ n1746 ^ 1'b0 ;
  assign n42188 = ( n11643 & ~n27374 ) | ( n11643 & n41116 ) | ( ~n27374 & n41116 ) ;
  assign n42189 = ( n8398 & n19566 ) | ( n8398 & n42188 ) | ( n19566 & n42188 ) ;
  assign n42190 = ( n1681 & n2891 ) | ( n1681 & ~n21134 ) | ( n2891 & ~n21134 ) ;
  assign n42191 = ( n1922 & n15203 ) | ( n1922 & ~n23818 ) | ( n15203 & ~n23818 ) ;
  assign n42192 = ( n36720 & n42190 ) | ( n36720 & ~n42191 ) | ( n42190 & ~n42191 ) ;
  assign n42193 = n18946 ^ n11988 ^ 1'b0 ;
  assign n42194 = ( n8668 & n14913 ) | ( n8668 & n16292 ) | ( n14913 & n16292 ) ;
  assign n42195 = n42194 ^ n40278 ^ n29471 ;
  assign n42196 = n39524 ^ n27549 ^ n7886 ;
  assign n42197 = n8685 ^ n6897 ^ x213 ;
  assign n42198 = n38966 ^ n23681 ^ n15022 ;
  assign n42199 = ( n13661 & ~n15101 ) | ( n13661 & n35847 ) | ( ~n15101 & n35847 ) ;
  assign n42200 = ( ~n21676 & n34943 ) | ( ~n21676 & n37149 ) | ( n34943 & n37149 ) ;
  assign n42201 = ( n19965 & ~n20768 ) | ( n19965 & n34761 ) | ( ~n20768 & n34761 ) ;
  assign n42202 = n11218 | n17526 ;
  assign n42203 = n24943 & ~n42202 ;
  assign n42204 = ( n3995 & n25581 ) | ( n3995 & n33896 ) | ( n25581 & n33896 ) ;
  assign n42205 = n18435 ^ n15153 ^ n10022 ;
  assign n42206 = n21893 ^ n16858 ^ n15378 ;
  assign n42207 = ~n20943 & n21483 ;
  assign n42208 = n42207 ^ n39728 ^ 1'b0 ;
  assign n42209 = n31327 ^ x55 ^ 1'b0 ;
  assign n42210 = n33461 & ~n42209 ;
  assign n42211 = n15594 ^ n2107 ^ 1'b0 ;
  assign n42212 = ( n8819 & n16109 ) | ( n8819 & n19658 ) | ( n16109 & n19658 ) ;
  assign n42213 = n30148 ^ n12237 ^ n11771 ;
  assign n42214 = n472 | n789 ;
  assign n42215 = n42214 ^ n27398 ^ n1645 ;
  assign n42216 = n22005 ^ n9599 ^ n4109 ;
  assign n42217 = n42216 ^ n19804 ^ n413 ;
  assign n42218 = ( n10197 & n12142 ) | ( n10197 & n18117 ) | ( n12142 & n18117 ) ;
  assign n42219 = n13862 ^ n13047 ^ n8655 ;
  assign n42220 = n38495 & n42219 ;
  assign n42221 = n25583 & n42220 ;
  assign n42222 = n42218 & ~n42221 ;
  assign n42223 = n24957 & n42222 ;
  assign n42224 = ( n23081 & ~n29741 ) | ( n23081 & n31150 ) | ( ~n29741 & n31150 ) ;
  assign n42225 = ( n4423 & n6408 ) | ( n4423 & ~n10058 ) | ( n6408 & ~n10058 ) ;
  assign n42226 = ( n8726 & ~n14264 ) | ( n8726 & n19488 ) | ( ~n14264 & n19488 ) ;
  assign n42227 = ( n24386 & ~n42225 ) | ( n24386 & n42226 ) | ( ~n42225 & n42226 ) ;
  assign n42228 = n17365 ^ n2406 ^ 1'b0 ;
  assign n42229 = n8031 & ~n42228 ;
  assign n42230 = n42229 ^ n27999 ^ n20370 ;
  assign n42231 = ~n19119 & n42230 ;
  assign n42232 = n42231 ^ n8125 ^ 1'b0 ;
  assign n42233 = ( n8355 & n17599 ) | ( n8355 & n42232 ) | ( n17599 & n42232 ) ;
  assign n42234 = n42233 ^ n7706 ^ 1'b0 ;
  assign n42235 = ~n9082 & n10830 ;
  assign n42236 = n5804 & n42235 ;
  assign n42237 = n22065 ^ n15996 ^ 1'b0 ;
  assign n42238 = ( n12789 & n42236 ) | ( n12789 & n42237 ) | ( n42236 & n42237 ) ;
  assign n42239 = n34349 ^ n15989 ^ n3334 ;
  assign n42240 = n35606 ^ n18886 ^ n10621 ;
  assign n42241 = n42240 ^ n30830 ^ n20618 ;
  assign n42242 = n40226 ^ n20936 ^ 1'b0 ;
  assign n42243 = n26410 | n42242 ;
  assign n42244 = n15940 ^ n8318 ^ n6082 ;
  assign n42245 = n42244 ^ n24885 ^ n445 ;
  assign n42246 = ( n32056 & n42243 ) | ( n32056 & n42245 ) | ( n42243 & n42245 ) ;
  assign n42247 = n33879 ^ n5550 ^ x117 ;
  assign n42248 = ~n5853 & n18129 ;
  assign n42249 = ( ~n8170 & n8184 ) | ( ~n8170 & n25234 ) | ( n8184 & n25234 ) ;
  assign n42250 = ( n31570 & n35533 ) | ( n31570 & ~n42249 ) | ( n35533 & ~n42249 ) ;
  assign n42251 = ( ~n12463 & n18517 ) | ( ~n12463 & n23168 ) | ( n18517 & n23168 ) ;
  assign n42252 = n28283 | n42251 ;
  assign n42253 = n22843 & ~n26231 ;
  assign n42254 = n42253 ^ n22097 ^ 1'b0 ;
  assign n42255 = ( n14698 & n25092 ) | ( n14698 & ~n42254 ) | ( n25092 & ~n42254 ) ;
  assign n42256 = n39351 ^ n38923 ^ 1'b0 ;
  assign n42257 = ~n24939 & n42256 ;
  assign n42258 = ( n18817 & n23091 ) | ( n18817 & ~n42257 ) | ( n23091 & ~n42257 ) ;
  assign n42259 = n21008 & ~n42258 ;
  assign n42260 = ( n3673 & ~n30740 ) | ( n3673 & n42259 ) | ( ~n30740 & n42259 ) ;
  assign n42261 = ( n11511 & n20292 ) | ( n11511 & n27682 ) | ( n20292 & n27682 ) ;
  assign n42265 = n6479 ^ n5938 ^ 1'b0 ;
  assign n42266 = ~n5407 & n42265 ;
  assign n42267 = ( n6911 & ~n38376 ) | ( n6911 & n42266 ) | ( ~n38376 & n42266 ) ;
  assign n42268 = n42267 ^ n28162 ^ n4323 ;
  assign n42262 = n18723 ^ n13218 ^ 1'b0 ;
  assign n42263 = ( n18818 & n28442 ) | ( n18818 & ~n42262 ) | ( n28442 & ~n42262 ) ;
  assign n42264 = n2909 & ~n42263 ;
  assign n42269 = n42268 ^ n42264 ^ 1'b0 ;
  assign n42270 = n42269 ^ n28143 ^ 1'b0 ;
  assign n42271 = n42261 | n42270 ;
  assign n42272 = ( n6389 & ~n26466 ) | ( n6389 & n33870 ) | ( ~n26466 & n33870 ) ;
  assign n42273 = ( n23929 & ~n28264 ) | ( n23929 & n42272 ) | ( ~n28264 & n42272 ) ;
  assign n42274 = ( n5627 & n16693 ) | ( n5627 & n22013 ) | ( n16693 & n22013 ) ;
  assign n42275 = n17780 ^ n1527 ^ n453 ;
  assign n42276 = n42274 | n42275 ;
  assign n42277 = n42276 ^ n14161 ^ n4632 ;
  assign n42278 = n36080 ^ n16049 ^ n4584 ;
  assign n42279 = ( n6321 & n18727 ) | ( n6321 & ~n35136 ) | ( n18727 & ~n35136 ) ;
  assign n42280 = n42279 ^ n34429 ^ n21950 ;
  assign n42281 = n32017 ^ n6767 ^ 1'b0 ;
  assign n42282 = ~n19313 & n42281 ;
  assign n42283 = n42282 ^ n20633 ^ n18875 ;
  assign n42284 = ( n17030 & n19570 ) | ( n17030 & n42283 ) | ( n19570 & n42283 ) ;
  assign n42285 = n42284 ^ n38474 ^ n20975 ;
  assign n42286 = n3573 | n8992 ;
  assign n42287 = ~n318 & n42286 ;
  assign n42288 = ( n22735 & ~n28382 ) | ( n22735 & n40592 ) | ( ~n28382 & n40592 ) ;
  assign n42289 = ( ~n15792 & n31495 ) | ( ~n15792 & n42288 ) | ( n31495 & n42288 ) ;
  assign n42290 = n20753 ^ n17615 ^ n2369 ;
  assign n42291 = ~n20080 & n42290 ;
  assign n42292 = n21312 & n42291 ;
  assign n42293 = n4657 & ~n19882 ;
  assign n42294 = n23316 & n42293 ;
  assign n42296 = n26677 ^ n20802 ^ n4315 ;
  assign n42295 = n6243 & n6825 ;
  assign n42297 = n42296 ^ n42295 ^ 1'b0 ;
  assign n42298 = n42297 ^ n9713 ^ n514 ;
  assign n42299 = n28794 ^ n17708 ^ n17632 ;
  assign n42300 = n42299 ^ n34997 ^ n13347 ;
  assign n42301 = ( n15967 & n37840 ) | ( n15967 & n42300 ) | ( n37840 & n42300 ) ;
  assign n42302 = ~n9053 & n36480 ;
  assign n42303 = ( n8154 & n8731 ) | ( n8154 & n28905 ) | ( n8731 & n28905 ) ;
  assign n42304 = n7918 & ~n13014 ;
  assign n42305 = ( ~n4416 & n5261 ) | ( ~n4416 & n16400 ) | ( n5261 & n16400 ) ;
  assign n42306 = ( ~n11130 & n19119 ) | ( ~n11130 & n19977 ) | ( n19119 & n19977 ) ;
  assign n42307 = ( n5609 & n42305 ) | ( n5609 & n42306 ) | ( n42305 & n42306 ) ;
  assign n42308 = ( n9569 & n15894 ) | ( n9569 & n30178 ) | ( n15894 & n30178 ) ;
  assign n42309 = n42308 ^ n25640 ^ n13354 ;
  assign n42310 = n13955 & n14834 ;
  assign n42311 = n42310 ^ n9008 ^ n422 ;
  assign n42312 = n21647 ^ n4233 ^ n2329 ;
  assign n42313 = ( n18894 & ~n20835 ) | ( n18894 & n42312 ) | ( ~n20835 & n42312 ) ;
  assign n42314 = n42313 ^ n24626 ^ n7964 ;
  assign n42315 = ( n19993 & n42311 ) | ( n19993 & ~n42314 ) | ( n42311 & ~n42314 ) ;
  assign n42317 = ( n11440 & n14616 ) | ( n11440 & ~n32282 ) | ( n14616 & ~n32282 ) ;
  assign n42318 = ( n23882 & n35312 ) | ( n23882 & ~n42317 ) | ( n35312 & ~n42317 ) ;
  assign n42316 = ~n7180 & n7678 ;
  assign n42319 = n42318 ^ n42316 ^ 1'b0 ;
  assign n42320 = n20007 | n23278 ;
  assign n42321 = n24991 & ~n42320 ;
  assign n42322 = n21483 ^ n16998 ^ n4359 ;
  assign n42323 = n31526 ^ n13593 ^ 1'b0 ;
  assign n42324 = n2087 | n42323 ;
  assign n42325 = ( n8073 & ~n29586 ) | ( n8073 & n42324 ) | ( ~n29586 & n42324 ) ;
  assign n42326 = ~n3402 & n6740 ;
  assign n42327 = n42326 ^ n32120 ^ n31407 ;
  assign n42328 = ~n29529 & n42327 ;
  assign n42329 = n42325 & n42328 ;
  assign n42330 = ( n9038 & n19836 ) | ( n9038 & n20883 ) | ( n19836 & n20883 ) ;
  assign n42331 = ( ~n3374 & n42329 ) | ( ~n3374 & n42330 ) | ( n42329 & n42330 ) ;
  assign n42332 = n16137 ^ n7959 ^ n5006 ;
  assign n42333 = ( ~n2274 & n3292 ) | ( ~n2274 & n19063 ) | ( n3292 & n19063 ) ;
  assign n42334 = ( n8718 & n14452 ) | ( n8718 & n42333 ) | ( n14452 & n42333 ) ;
  assign n42335 = n41116 ^ n38910 ^ n8434 ;
  assign n42336 = ( ~n5874 & n34289 ) | ( ~n5874 & n42335 ) | ( n34289 & n42335 ) ;
  assign n42339 = ( n10783 & n31871 ) | ( n10783 & n32606 ) | ( n31871 & n32606 ) ;
  assign n42340 = ( n23010 & n38833 ) | ( n23010 & n42339 ) | ( n38833 & n42339 ) ;
  assign n42338 = n8514 ^ n6375 ^ n3065 ;
  assign n42341 = n42340 ^ n42338 ^ n26824 ;
  assign n42337 = n41962 ^ n32600 ^ n1792 ;
  assign n42342 = n42341 ^ n42337 ^ n36970 ;
  assign n42348 = n2724 | n26250 ;
  assign n42345 = n4965 | n6152 ;
  assign n42346 = n16118 & ~n42345 ;
  assign n42343 = n28415 ^ n7397 ^ n2375 ;
  assign n42344 = n42343 ^ n35502 ^ n31383 ;
  assign n42347 = n42346 ^ n42344 ^ n33068 ;
  assign n42349 = n42348 ^ n42347 ^ x248 ;
  assign n42350 = ( n11770 & n34960 ) | ( n11770 & ~n39712 ) | ( n34960 & ~n39712 ) ;
  assign n42351 = n34904 ^ n24162 ^ 1'b0 ;
  assign n42352 = n15935 | n42351 ;
  assign n42353 = ~n1340 & n36321 ;
  assign n42354 = ( ~n4828 & n13870 ) | ( ~n4828 & n27032 ) | ( n13870 & n27032 ) ;
  assign n42355 = n12613 ^ n5271 ^ n2960 ;
  assign n42356 = n18764 ^ n7830 ^ 1'b0 ;
  assign n42357 = ( n8116 & ~n11376 ) | ( n8116 & n42356 ) | ( ~n11376 & n42356 ) ;
  assign n42358 = ( n975 & n9359 ) | ( n975 & ~n32227 ) | ( n9359 & ~n32227 ) ;
  assign n42359 = ( n42355 & n42357 ) | ( n42355 & n42358 ) | ( n42357 & n42358 ) ;
  assign n42360 = ( n1803 & n2755 ) | ( n1803 & ~n21501 ) | ( n2755 & ~n21501 ) ;
  assign n42361 = n32281 ^ n25719 ^ n6455 ;
  assign n42362 = n42361 ^ n16617 ^ n5305 ;
  assign n42363 = ( ~n29800 & n42360 ) | ( ~n29800 & n42362 ) | ( n42360 & n42362 ) ;
  assign n42364 = ~n14410 & n16957 ;
  assign n42365 = n42364 ^ n8917 ^ 1'b0 ;
  assign n42366 = n42365 ^ n26434 ^ n9352 ;
  assign n42367 = ( n4696 & n6788 ) | ( n4696 & n18244 ) | ( n6788 & n18244 ) ;
  assign n42368 = ( n3140 & n22936 ) | ( n3140 & ~n42367 ) | ( n22936 & ~n42367 ) ;
  assign n42369 = n39296 ^ n29558 ^ n20241 ;
  assign n42370 = ( ~n42366 & n42368 ) | ( ~n42366 & n42369 ) | ( n42368 & n42369 ) ;
  assign n42371 = n22326 ^ n13157 ^ n11792 ;
  assign n42372 = ( n15456 & ~n20811 ) | ( n15456 & n26868 ) | ( ~n20811 & n26868 ) ;
  assign n42373 = n42372 ^ n33616 ^ n14355 ;
  assign n42374 = n42373 ^ n27053 ^ x27 ;
  assign n42375 = ( n14428 & n33484 ) | ( n14428 & ~n42374 ) | ( n33484 & ~n42374 ) ;
  assign n42377 = ~n11501 & n15001 ;
  assign n42378 = n42377 ^ n40700 ^ 1'b0 ;
  assign n42376 = n35679 ^ n13943 ^ n12952 ;
  assign n42379 = n42378 ^ n42376 ^ n41332 ;
  assign n42380 = n42379 ^ n34028 ^ n22091 ;
  assign n42381 = ( n900 & ~n5303 ) | ( n900 & n42025 ) | ( ~n5303 & n42025 ) ;
  assign n42384 = ( n8750 & n25729 ) | ( n8750 & n29162 ) | ( n25729 & n29162 ) ;
  assign n42383 = ( n2311 & n5754 ) | ( n2311 & ~n9308 ) | ( n5754 & ~n9308 ) ;
  assign n42382 = n35942 ^ n23978 ^ n9141 ;
  assign n42385 = n42384 ^ n42383 ^ n42382 ;
  assign n42386 = n23834 ^ n17045 ^ n11205 ;
  assign n42387 = n42386 ^ n20391 ^ n13633 ;
  assign n42388 = ( n17323 & ~n19375 ) | ( n17323 & n42387 ) | ( ~n19375 & n42387 ) ;
  assign n42389 = ( ~n20295 & n21486 ) | ( ~n20295 & n21790 ) | ( n21486 & n21790 ) ;
  assign n42390 = n25224 ^ n11806 ^ n2473 ;
  assign n42391 = n14530 | n28450 ;
  assign n42392 = n42391 ^ n7674 ^ 1'b0 ;
  assign n42393 = n42392 ^ n32435 ^ n9543 ;
  assign n42394 = n21652 ^ n4499 ^ n3392 ;
  assign n42395 = n42394 ^ n34896 ^ 1'b0 ;
  assign n42396 = ( n3807 & n6385 ) | ( n3807 & n42395 ) | ( n6385 & n42395 ) ;
  assign n42397 = n19565 ^ n9112 ^ n2908 ;
  assign n42398 = n14571 | n19446 ;
  assign n42399 = n42397 & ~n42398 ;
  assign n42400 = n34799 ^ n18908 ^ 1'b0 ;
  assign n42401 = ~n9361 & n42400 ;
  assign n42402 = n34728 ^ n21485 ^ n20736 ;
  assign n42403 = n42402 ^ n13347 ^ n3006 ;
  assign n42404 = ( n18352 & n34253 ) | ( n18352 & n42403 ) | ( n34253 & n42403 ) ;
  assign n42405 = n14649 & ~n42404 ;
  assign n42406 = n40370 ^ n26524 ^ n7419 ;
  assign n42407 = ( n14996 & n19812 ) | ( n14996 & ~n42406 ) | ( n19812 & ~n42406 ) ;
  assign n42408 = n39046 ^ n31168 ^ n6361 ;
  assign n42409 = ( n1474 & ~n2509 ) | ( n1474 & n37773 ) | ( ~n2509 & n37773 ) ;
  assign n42410 = n42409 ^ n21232 ^ n6606 ;
  assign n42413 = n20021 | n23268 ;
  assign n42414 = n42413 ^ n1344 ^ 1'b0 ;
  assign n42415 = n24358 & n42414 ;
  assign n42416 = n42415 ^ n10672 ^ 1'b0 ;
  assign n42411 = n16295 ^ n15561 ^ 1'b0 ;
  assign n42412 = n4741 | n42411 ;
  assign n42417 = n42416 ^ n42412 ^ n19671 ;
  assign n42418 = n42410 | n42417 ;
  assign n42419 = n11128 ^ n8849 ^ n482 ;
  assign n42420 = n31562 ^ n30723 ^ n5678 ;
  assign n42421 = ( ~n14190 & n31689 ) | ( ~n14190 & n42420 ) | ( n31689 & n42420 ) ;
  assign n42422 = ( ~n4971 & n39077 ) | ( ~n4971 & n40803 ) | ( n39077 & n40803 ) ;
  assign n42424 = n17356 ^ n11607 ^ n9891 ;
  assign n42423 = n22124 ^ n6154 ^ n4761 ;
  assign n42425 = n42424 ^ n42423 ^ n26401 ;
  assign n42426 = n12281 & ~n42425 ;
  assign n42431 = n4390 | n37696 ;
  assign n42432 = n42431 ^ n5483 ^ 1'b0 ;
  assign n42428 = ~n2943 & n5921 ;
  assign n42429 = n42428 ^ n17639 ^ 1'b0 ;
  assign n42427 = ( ~n1507 & n6927 ) | ( ~n1507 & n19188 ) | ( n6927 & n19188 ) ;
  assign n42430 = n42429 ^ n42427 ^ n37631 ;
  assign n42433 = n42432 ^ n42430 ^ n15579 ;
  assign n42434 = n2590 | n8629 ;
  assign n42435 = ( n6952 & ~n25451 ) | ( n6952 & n33970 ) | ( ~n25451 & n33970 ) ;
  assign n42436 = ( n7863 & n29953 ) | ( n7863 & ~n42435 ) | ( n29953 & ~n42435 ) ;
  assign n42437 = ( ~n11876 & n28680 ) | ( ~n11876 & n41554 ) | ( n28680 & n41554 ) ;
  assign n42438 = ( n42434 & n42436 ) | ( n42434 & n42437 ) | ( n42436 & n42437 ) ;
  assign n42439 = ~n16196 & n40103 ;
  assign n42440 = n26044 ^ n26020 ^ n22365 ;
  assign n42441 = n17414 ^ n11204 ^ n2483 ;
  assign n42442 = n42441 ^ n21330 ^ n17343 ;
  assign n42443 = n40181 ^ n38922 ^ n20943 ;
  assign n42444 = n8383 & n36027 ;
  assign n42445 = n27341 & n42444 ;
  assign n42446 = n32204 & n42445 ;
  assign n42447 = n17191 ^ n6454 ^ 1'b0 ;
  assign n42448 = ~n5140 & n42447 ;
  assign n42450 = n20719 ^ n17629 ^ n17554 ;
  assign n42449 = ( n16763 & n35136 ) | ( n16763 & n39900 ) | ( n35136 & n39900 ) ;
  assign n42451 = n42450 ^ n42449 ^ n26523 ;
  assign n42452 = n41450 ^ n15522 ^ n6599 ;
  assign n42453 = ( n3054 & ~n10700 ) | ( n3054 & n25664 ) | ( ~n10700 & n25664 ) ;
  assign n42454 = ( n7173 & n14022 ) | ( n7173 & ~n42453 ) | ( n14022 & ~n42453 ) ;
  assign n42455 = n32321 ^ n29384 ^ 1'b0 ;
  assign n42456 = ( n1301 & n8007 ) | ( n1301 & n14739 ) | ( n8007 & n14739 ) ;
  assign n42457 = n42456 ^ n24869 ^ n14303 ;
  assign n42458 = n10974 ^ n7934 ^ 1'b0 ;
  assign n42459 = ( n2589 & n20467 ) | ( n2589 & ~n42458 ) | ( n20467 & ~n42458 ) ;
  assign n42460 = ( n12687 & n40436 ) | ( n12687 & n42459 ) | ( n40436 & n42459 ) ;
  assign n42461 = ( n11668 & ~n19036 ) | ( n11668 & n37553 ) | ( ~n19036 & n37553 ) ;
  assign n42462 = ~n17120 & n42461 ;
  assign n42463 = ( n31839 & n32489 ) | ( n31839 & ~n35420 ) | ( n32489 & ~n35420 ) ;
  assign n42464 = n27109 ^ n20989 ^ n11831 ;
  assign n42465 = ( n1490 & n11326 ) | ( n1490 & ~n28506 ) | ( n11326 & ~n28506 ) ;
  assign n42466 = n42465 ^ n14378 ^ n5030 ;
  assign n42467 = n28699 ^ n15309 ^ 1'b0 ;
  assign n42468 = n14392 & n42467 ;
  assign n42469 = n42468 ^ n7203 ^ n3186 ;
  assign n42470 = ( n8102 & n21901 ) | ( n8102 & n42469 ) | ( n21901 & n42469 ) ;
  assign n42471 = ( n6627 & ~n21151 ) | ( n6627 & n39642 ) | ( ~n21151 & n39642 ) ;
  assign n42472 = ( n8704 & n26064 ) | ( n8704 & ~n42471 ) | ( n26064 & ~n42471 ) ;
  assign n42473 = ( n7551 & ~n18670 ) | ( n7551 & n32026 ) | ( ~n18670 & n32026 ) ;
  assign n42474 = n42473 ^ n6240 ^ 1'b0 ;
  assign n42475 = n33125 ^ n6926 ^ 1'b0 ;
  assign n42476 = n26965 | n42475 ;
  assign n42479 = ( n2165 & ~n3601 ) | ( n2165 & n6039 ) | ( ~n3601 & n6039 ) ;
  assign n42477 = n30901 ^ n4104 ^ 1'b0 ;
  assign n42478 = n38541 & ~n42477 ;
  assign n42480 = n42479 ^ n42478 ^ n39153 ;
  assign n42481 = ( ~n2351 & n7833 ) | ( ~n2351 & n21239 ) | ( n7833 & n21239 ) ;
  assign n42482 = n13141 ^ n10695 ^ n2981 ;
  assign n42483 = ~n11803 & n26236 ;
  assign n42484 = n29849 & n42483 ;
  assign n42485 = ( n19329 & ~n30071 ) | ( n19329 & n42484 ) | ( ~n30071 & n42484 ) ;
  assign n42486 = ( ~n6656 & n9806 ) | ( ~n6656 & n18733 ) | ( n9806 & n18733 ) ;
  assign n42487 = n9018 & n27332 ;
  assign n42488 = n13073 | n23221 ;
  assign n42489 = n42488 ^ n7467 ^ 1'b0 ;
  assign n42491 = n22612 ^ n17855 ^ 1'b0 ;
  assign n42492 = ~n5029 & n42491 ;
  assign n42490 = n40230 ^ n38822 ^ n6123 ;
  assign n42493 = n42492 ^ n42490 ^ n36914 ;
  assign n42495 = ( n1471 & n2145 ) | ( n1471 & n9182 ) | ( n2145 & n9182 ) ;
  assign n42496 = n42495 ^ n31616 ^ n5844 ;
  assign n42494 = n27046 & n28591 ;
  assign n42497 = n42496 ^ n42494 ^ n34794 ;
  assign n42498 = n28965 ^ n11478 ^ 1'b0 ;
  assign n42499 = ( n14239 & n34979 ) | ( n14239 & ~n42498 ) | ( n34979 & ~n42498 ) ;
  assign n42500 = n16814 & n35549 ;
  assign n42501 = ( n16222 & ~n42499 ) | ( n16222 & n42500 ) | ( ~n42499 & n42500 ) ;
  assign n42502 = n5650 ^ n2070 ^ 1'b0 ;
  assign n42503 = n42502 ^ n18351 ^ n7806 ;
  assign n42504 = n42503 ^ n23753 ^ n3596 ;
  assign n42505 = n10142 ^ n4153 ^ n779 ;
  assign n42506 = ( ~n9184 & n12609 ) | ( ~n9184 & n42505 ) | ( n12609 & n42505 ) ;
  assign n42507 = ( n5863 & n40341 ) | ( n5863 & n42506 ) | ( n40341 & n42506 ) ;
  assign n42508 = n33700 ^ n11380 ^ n954 ;
  assign n42509 = n7533 ^ n1814 ^ 1'b0 ;
  assign n42510 = ~n8456 & n42509 ;
  assign n42511 = n9535 & n42510 ;
  assign n42512 = n23638 & ~n29528 ;
  assign n42513 = n36697 | n42512 ;
  assign n42514 = n30094 ^ n6497 ^ 1'b0 ;
  assign n42515 = n2908 & n42514 ;
  assign n42516 = n42515 ^ n10513 ^ n1725 ;
  assign n42517 = ( n628 & ~n3173 ) | ( n628 & n42516 ) | ( ~n3173 & n42516 ) ;
  assign n42518 = ( ~n9435 & n20862 ) | ( ~n9435 & n41473 ) | ( n20862 & n41473 ) ;
  assign n42519 = ( ~n12907 & n22550 ) | ( ~n12907 & n42518 ) | ( n22550 & n42518 ) ;
  assign n42520 = ~n608 & n9199 ;
  assign n42521 = ( ~n7537 & n29829 ) | ( ~n7537 & n42520 ) | ( n29829 & n42520 ) ;
  assign n42522 = n42521 ^ n30156 ^ n15044 ;
  assign n42523 = n26535 ^ n23663 ^ n18910 ;
  assign n42524 = n42523 ^ n15295 ^ 1'b0 ;
  assign n42525 = ( n4639 & ~n16969 ) | ( n4639 & n42524 ) | ( ~n16969 & n42524 ) ;
  assign n42526 = n27495 ^ n26972 ^ n3274 ;
  assign n42527 = ( ~n11756 & n39220 ) | ( ~n11756 & n42526 ) | ( n39220 & n42526 ) ;
  assign n42528 = n38625 ^ n23512 ^ n333 ;
  assign n42529 = n11086 & ~n35938 ;
  assign n42530 = n5294 & n42529 ;
  assign n42531 = n33655 ^ n22395 ^ n13883 ;
  assign n42532 = n14167 ^ n1396 ^ 1'b0 ;
  assign n42533 = n13776 | n42532 ;
  assign n42534 = ( n9024 & n33605 ) | ( n9024 & ~n42533 ) | ( n33605 & ~n42533 ) ;
  assign n42535 = ( n9831 & n38486 ) | ( n9831 & ~n42534 ) | ( n38486 & ~n42534 ) ;
  assign n42536 = n7446 ^ n4242 ^ n2006 ;
  assign n42537 = ( ~n2477 & n12494 ) | ( ~n2477 & n13878 ) | ( n12494 & n13878 ) ;
  assign n42538 = n42537 ^ n34044 ^ n23898 ;
  assign n42539 = ( ~n7449 & n32228 ) | ( ~n7449 & n42538 ) | ( n32228 & n42538 ) ;
  assign n42540 = n34760 ^ n27107 ^ n19250 ;
  assign n42541 = n14563 ^ n6528 ^ 1'b0 ;
  assign n42542 = ( ~n301 & n11791 ) | ( ~n301 & n36267 ) | ( n11791 & n36267 ) ;
  assign n42543 = n42542 ^ n30252 ^ n21502 ;
  assign n42544 = ( n2716 & n42541 ) | ( n2716 & n42543 ) | ( n42541 & n42543 ) ;
  assign n42545 = ( ~n1771 & n12836 ) | ( ~n1771 & n42544 ) | ( n12836 & n42544 ) ;
  assign n42546 = ( ~n15410 & n25472 ) | ( ~n15410 & n40179 ) | ( n25472 & n40179 ) ;
  assign n42547 = n15493 ^ n9886 ^ n5304 ;
  assign n42548 = ( n13393 & n28360 ) | ( n13393 & n31973 ) | ( n28360 & n31973 ) ;
  assign n42549 = ( n1509 & ~n18831 ) | ( n1509 & n38526 ) | ( ~n18831 & n38526 ) ;
  assign n42550 = ( n2270 & ~n4635 ) | ( n2270 & n11669 ) | ( ~n4635 & n11669 ) ;
  assign n42551 = n30844 ^ n16879 ^ n1319 ;
  assign n42552 = ( ~n11095 & n20823 ) | ( ~n11095 & n42551 ) | ( n20823 & n42551 ) ;
  assign n42553 = ( ~n22028 & n42550 ) | ( ~n22028 & n42552 ) | ( n42550 & n42552 ) ;
  assign n42554 = n16640 ^ n4718 ^ 1'b0 ;
  assign n42555 = n11895 & ~n42554 ;
  assign n42559 = n18223 & n35509 ;
  assign n42560 = n10381 & n42559 ;
  assign n42558 = n21647 ^ n8872 ^ n6000 ;
  assign n42556 = n9746 ^ n8665 ^ n826 ;
  assign n42557 = n42556 ^ n26781 ^ n9291 ;
  assign n42561 = n42560 ^ n42558 ^ n42557 ;
  assign n42562 = n42561 ^ n36148 ^ n2107 ;
  assign n42563 = n37848 ^ n27903 ^ 1'b0 ;
  assign n42564 = n32728 & n42563 ;
  assign n42565 = n40524 ^ n5220 ^ 1'b0 ;
  assign n42566 = x223 & n42565 ;
  assign n42567 = n42566 ^ n40859 ^ n6281 ;
  assign n42568 = ( n28141 & ~n37218 ) | ( n28141 & n42567 ) | ( ~n37218 & n42567 ) ;
  assign n42569 = ( n1217 & n13311 ) | ( n1217 & ~n15647 ) | ( n13311 & ~n15647 ) ;
  assign n42570 = n25583 ^ n18464 ^ n11539 ;
  assign n42571 = n42570 ^ n30510 ^ n15947 ;
  assign n42572 = n15840 ^ n8586 ^ n372 ;
  assign n42573 = n37025 ^ n34541 ^ n12847 ;
  assign n42574 = n29136 ^ n19937 ^ n11470 ;
  assign n42575 = n6480 ^ n4281 ^ n2643 ;
  assign n42577 = ( n9466 & n9713 ) | ( n9466 & n23929 ) | ( n9713 & n23929 ) ;
  assign n42576 = n25237 | n28461 ;
  assign n42578 = n42577 ^ n42576 ^ 1'b0 ;
  assign n42579 = n1698 & n10124 ;
  assign n42580 = n6977 & n42579 ;
  assign n42581 = n1299 & ~n5314 ;
  assign n42582 = n42581 ^ n16788 ^ 1'b0 ;
  assign n42583 = ( n6072 & n42580 ) | ( n6072 & ~n42582 ) | ( n42580 & ~n42582 ) ;
  assign n42584 = n14843 ^ n1425 ^ 1'b0 ;
  assign n42585 = n259 | n42584 ;
  assign n42586 = n22299 ^ n13640 ^ n7282 ;
  assign n42587 = ( n14006 & n42585 ) | ( n14006 & n42586 ) | ( n42585 & n42586 ) ;
  assign n42588 = ( n23254 & n42583 ) | ( n23254 & n42587 ) | ( n42583 & n42587 ) ;
  assign n42589 = ( n8320 & n11254 ) | ( n8320 & n18531 ) | ( n11254 & n18531 ) ;
  assign n42590 = n42589 ^ n37081 ^ n14871 ;
  assign n42591 = ( n523 & n24904 ) | ( n523 & n42590 ) | ( n24904 & n42590 ) ;
  assign n42592 = n30692 ^ n2506 ^ 1'b0 ;
  assign n42593 = n42592 ^ n25781 ^ n8221 ;
  assign n42594 = ( ~n9433 & n31079 ) | ( ~n9433 & n42593 ) | ( n31079 & n42593 ) ;
  assign n42595 = n42329 ^ n41666 ^ n33267 ;
  assign n42596 = ~n1934 & n5677 ;
  assign n42597 = n42596 ^ n17381 ^ 1'b0 ;
  assign n42598 = n42597 ^ n37740 ^ n2680 ;
  assign n42599 = n28523 ^ n18493 ^ n10386 ;
  assign n42600 = n34617 & ~n42599 ;
  assign n42601 = n31724 ^ n5677 ^ n3911 ;
  assign n42602 = n34475 ^ n24074 ^ n2824 ;
  assign n42603 = n42602 ^ n19393 ^ n4216 ;
  assign n42604 = n42603 ^ n30308 ^ n29242 ;
  assign n42605 = n7666 | n29941 ;
  assign n42606 = n42605 ^ n1339 ^ 1'b0 ;
  assign n42607 = ~n19770 & n42606 ;
  assign n42608 = ( ~n7971 & n11980 ) | ( ~n7971 & n34889 ) | ( n11980 & n34889 ) ;
  assign n42609 = ( ~n13874 & n15792 ) | ( ~n13874 & n42608 ) | ( n15792 & n42608 ) ;
  assign n42610 = n28411 ^ n15147 ^ n5365 ;
  assign n42611 = ( n7097 & ~n24098 ) | ( n7097 & n33353 ) | ( ~n24098 & n33353 ) ;
  assign n42612 = ( n2977 & n42610 ) | ( n2977 & ~n42611 ) | ( n42610 & ~n42611 ) ;
  assign n42613 = ( n8178 & n19322 ) | ( n8178 & ~n36713 ) | ( n19322 & ~n36713 ) ;
  assign n42614 = ( n1993 & ~n16838 ) | ( n1993 & n39782 ) | ( ~n16838 & n39782 ) ;
  assign n42615 = n42614 ^ n10838 ^ n2093 ;
  assign n42616 = n38095 ^ n35938 ^ n2748 ;
  assign n42617 = n42616 ^ n33543 ^ n3360 ;
  assign n42618 = n30856 ^ n4083 ^ 1'b0 ;
  assign n42619 = n30178 | n42618 ;
  assign n42620 = n22686 ^ n20354 ^ n13999 ;
  assign n42621 = ~n27256 & n42620 ;
  assign n42622 = n42621 ^ n36761 ^ 1'b0 ;
  assign n42623 = n16873 ^ n3854 ^ n1714 ;
  assign n42624 = n23901 ^ n16880 ^ n12680 ;
  assign n42625 = n42624 ^ n9091 ^ n1437 ;
  assign n42626 = ( ~n21675 & n29253 ) | ( ~n21675 & n42625 ) | ( n29253 & n42625 ) ;
  assign n42627 = n42582 ^ n7114 ^ n859 ;
  assign n42628 = n32076 ^ n6976 ^ 1'b0 ;
  assign n42629 = n42628 ^ n36082 ^ n33132 ;
  assign n42630 = ( n3740 & n26563 ) | ( n3740 & n41939 ) | ( n26563 & n41939 ) ;
  assign n42631 = n42630 ^ n33422 ^ n9639 ;
  assign n42632 = ( n22292 & ~n38158 ) | ( n22292 & n40911 ) | ( ~n38158 & n40911 ) ;
  assign n42633 = ( n10459 & n39164 ) | ( n10459 & n42632 ) | ( n39164 & n42632 ) ;
  assign n42634 = n2231 & ~n40176 ;
  assign n42635 = n18455 ^ n17214 ^ n2854 ;
  assign n42636 = n7546 & ~n42635 ;
  assign n42637 = ~n42634 & n42636 ;
  assign n42638 = n11275 ^ n10277 ^ n4077 ;
  assign n42639 = ( n4770 & n6626 ) | ( n4770 & n11596 ) | ( n6626 & n11596 ) ;
  assign n42640 = n42639 ^ n14410 ^ n13794 ;
  assign n42641 = n13699 & n42640 ;
  assign n42642 = ~n42638 & n42641 ;
  assign n42643 = n17353 ^ n14077 ^ n11437 ;
  assign n42644 = ( n11312 & n14821 ) | ( n11312 & n24912 ) | ( n14821 & n24912 ) ;
  assign n42645 = n42644 ^ n28212 ^ n16412 ;
  assign n42646 = ~n1327 & n10520 ;
  assign n42647 = ~n28432 & n42646 ;
  assign n42648 = n33983 ^ n30403 ^ n5813 ;
  assign n42649 = ( n39374 & n42647 ) | ( n39374 & ~n42648 ) | ( n42647 & ~n42648 ) ;
  assign n42650 = ( n15281 & ~n37778 ) | ( n15281 & n42649 ) | ( ~n37778 & n42649 ) ;
  assign n42651 = n19583 ^ n7641 ^ n7203 ;
  assign n42652 = n19414 ^ n8393 ^ n623 ;
  assign n42653 = n35100 & ~n42652 ;
  assign n42654 = n26396 ^ n22930 ^ n439 ;
  assign n42655 = n42654 ^ n33302 ^ n16178 ;
  assign n42656 = n37700 ^ n28413 ^ n22911 ;
  assign n42657 = ( n8489 & ~n33221 ) | ( n8489 & n41843 ) | ( ~n33221 & n41843 ) ;
  assign n42658 = ( n6616 & ~n42656 ) | ( n6616 & n42657 ) | ( ~n42656 & n42657 ) ;
  assign n42659 = n10556 | n14822 ;
  assign n42660 = n12988 | n42659 ;
  assign n42661 = n39279 ^ n21027 ^ n2201 ;
  assign n42662 = n40279 | n42661 ;
  assign n42663 = n3508 | n42662 ;
  assign n42664 = n17576 ^ n10658 ^ n4788 ;
  assign n42665 = n39873 & n42664 ;
  assign n42666 = ( n527 & n8554 ) | ( n527 & ~n14423 ) | ( n8554 & ~n14423 ) ;
  assign n42667 = ( n6690 & n9685 ) | ( n6690 & ~n31466 ) | ( n9685 & ~n31466 ) ;
  assign n42668 = n27309 ^ n3151 ^ 1'b0 ;
  assign n42669 = ( n19502 & n31499 ) | ( n19502 & ~n42668 ) | ( n31499 & ~n42668 ) ;
  assign n42670 = n14332 ^ n11195 ^ n6776 ;
  assign n42671 = ( n4678 & n4745 ) | ( n4678 & ~n19244 ) | ( n4745 & ~n19244 ) ;
  assign n42672 = n29869 | n36313 ;
  assign n42673 = n16239 & ~n42672 ;
  assign n42674 = ( ~n15011 & n42671 ) | ( ~n15011 & n42673 ) | ( n42671 & n42673 ) ;
  assign n42675 = ( n671 & n1902 ) | ( n671 & ~n42674 ) | ( n1902 & ~n42674 ) ;
  assign n42676 = ( n19357 & ~n20459 ) | ( n19357 & n25459 ) | ( ~n20459 & n25459 ) ;
  assign n42677 = n27090 ^ n20332 ^ n13087 ;
  assign n42678 = n42677 ^ n11720 ^ n4976 ;
  assign n42679 = ( n1343 & n16160 ) | ( n1343 & n24090 ) | ( n16160 & n24090 ) ;
  assign n42680 = n40382 ^ n23654 ^ n6057 ;
  assign n42685 = ( ~n1977 & n6782 ) | ( ~n1977 & n16805 ) | ( n6782 & n16805 ) ;
  assign n42686 = ( n9632 & n38577 ) | ( n9632 & ~n42685 ) | ( n38577 & ~n42685 ) ;
  assign n42681 = n3132 ^ n3102 ^ 1'b0 ;
  assign n42682 = ~n1031 & n42681 ;
  assign n42683 = ( n8522 & ~n17720 ) | ( n8522 & n42682 ) | ( ~n17720 & n42682 ) ;
  assign n42684 = n37476 & n42683 ;
  assign n42687 = n42686 ^ n42684 ^ 1'b0 ;
  assign n42688 = ( ~n19534 & n23479 ) | ( ~n19534 & n42687 ) | ( n23479 & n42687 ) ;
  assign n42690 = n6636 ^ n6328 ^ n1409 ;
  assign n42689 = ( n12232 & n18663 ) | ( n12232 & n18689 ) | ( n18663 & n18689 ) ;
  assign n42691 = n42690 ^ n42689 ^ n40770 ;
  assign n42692 = n27995 ^ n4018 ^ 1'b0 ;
  assign n42693 = n42692 ^ n30340 ^ n23647 ;
  assign n42694 = ( n935 & n10488 ) | ( n935 & ~n14649 ) | ( n10488 & ~n14649 ) ;
  assign n42695 = ( ~n16911 & n35719 ) | ( ~n16911 & n42694 ) | ( n35719 & n42694 ) ;
  assign n42696 = ( x119 & n272 ) | ( x119 & n35410 ) | ( n272 & n35410 ) ;
  assign n42697 = n18469 ^ n5701 ^ n4429 ;
  assign n42698 = ( n7493 & ~n42696 ) | ( n7493 & n42697 ) | ( ~n42696 & n42697 ) ;
  assign n42699 = n42698 ^ n9902 ^ 1'b0 ;
  assign n42700 = n42695 & ~n42699 ;
  assign n42701 = n41466 ^ n28361 ^ n2028 ;
  assign n42702 = n37611 ^ n26016 ^ n12031 ;
  assign n42703 = n21844 ^ n15675 ^ 1'b0 ;
  assign n42704 = ( n3269 & ~n6958 ) | ( n3269 & n34470 ) | ( ~n6958 & n34470 ) ;
  assign n42705 = ( ~n7525 & n15140 ) | ( ~n7525 & n42704 ) | ( n15140 & n42704 ) ;
  assign n42706 = n20367 ^ n9495 ^ n7029 ;
  assign n42707 = ( ~n11833 & n12048 ) | ( ~n11833 & n14101 ) | ( n12048 & n14101 ) ;
  assign n42708 = n42707 ^ n22860 ^ 1'b0 ;
  assign n42709 = ( n7236 & n42706 ) | ( n7236 & n42708 ) | ( n42706 & n42708 ) ;
  assign n42710 = n24163 ^ n19326 ^ n16116 ;
  assign n42711 = ( n10067 & n12154 ) | ( n10067 & ~n21670 ) | ( n12154 & ~n21670 ) ;
  assign n42712 = n42711 ^ n1176 ^ 1'b0 ;
  assign n42713 = ( n20314 & ~n21241 ) | ( n20314 & n23083 ) | ( ~n21241 & n23083 ) ;
  assign n42714 = n42713 ^ n9422 ^ 1'b0 ;
  assign n42715 = ( n21933 & ~n28782 ) | ( n21933 & n42714 ) | ( ~n28782 & n42714 ) ;
  assign n42716 = n42715 ^ n17707 ^ n12394 ;
  assign n42717 = ( n652 & n21105 ) | ( n652 & ~n33889 ) | ( n21105 & ~n33889 ) ;
  assign n42718 = n8443 & ~n42717 ;
  assign n42719 = n15471 & n42718 ;
  assign n42720 = ( ~n42712 & n42716 ) | ( ~n42712 & n42719 ) | ( n42716 & n42719 ) ;
  assign n42721 = n14732 & n38625 ;
  assign n42722 = n42721 ^ n40956 ^ n38083 ;
  assign n42723 = ~n371 & n23220 ;
  assign n42724 = n42723 ^ n1665 ^ 1'b0 ;
  assign n42725 = n32569 ^ n17199 ^ 1'b0 ;
  assign n42726 = n40186 & ~n42725 ;
  assign n42727 = ( ~n18151 & n24352 ) | ( ~n18151 & n27659 ) | ( n24352 & n27659 ) ;
  assign n42728 = n35518 ^ n16876 ^ n13369 ;
  assign n42729 = ( ~n1481 & n2089 ) | ( ~n1481 & n20508 ) | ( n2089 & n20508 ) ;
  assign n42730 = ( n10578 & ~n42728 ) | ( n10578 & n42729 ) | ( ~n42728 & n42729 ) ;
  assign n42731 = n25283 & ~n32822 ;
  assign n42732 = ( ~n11922 & n19233 ) | ( ~n11922 & n30675 ) | ( n19233 & n30675 ) ;
  assign n42735 = n5474 ^ n4916 ^ n3767 ;
  assign n42733 = n3553 ^ x88 ^ 1'b0 ;
  assign n42734 = ~n30783 & n42733 ;
  assign n42736 = n42735 ^ n42734 ^ n37802 ;
  assign n42737 = ( n13262 & n14720 ) | ( n13262 & n42736 ) | ( n14720 & n42736 ) ;
  assign n42738 = n19764 & ~n26523 ;
  assign n42739 = n42738 ^ n5975 ^ 1'b0 ;
  assign n42740 = ( n2703 & n25636 ) | ( n2703 & ~n39034 ) | ( n25636 & ~n39034 ) ;
  assign n42741 = n32526 ^ n23370 ^ n11582 ;
  assign n42742 = ( n19057 & ~n35668 ) | ( n19057 & n42741 ) | ( ~n35668 & n42741 ) ;
  assign n42743 = ( n11812 & n29818 ) | ( n11812 & n34784 ) | ( n29818 & n34784 ) ;
  assign n42744 = ( n18348 & n42742 ) | ( n18348 & ~n42743 ) | ( n42742 & ~n42743 ) ;
  assign n42745 = n28476 ^ n16434 ^ n6336 ;
  assign n42746 = n9395 ^ n5094 ^ n4371 ;
  assign n42747 = n42746 ^ n17618 ^ n5289 ;
  assign n42748 = n10804 ^ n8324 ^ 1'b0 ;
  assign n42749 = n42230 ^ n12043 ^ 1'b0 ;
  assign n42750 = ~n41500 & n42749 ;
  assign n42751 = ( n14806 & n14913 ) | ( n14806 & n42750 ) | ( n14913 & n42750 ) ;
  assign n42752 = ( ~n7145 & n18713 ) | ( ~n7145 & n41880 ) | ( n18713 & n41880 ) ;
  assign n42753 = n28407 ^ n16538 ^ n658 ;
  assign n42755 = n31397 ^ n10797 ^ n7314 ;
  assign n42754 = n22900 ^ n22372 ^ 1'b0 ;
  assign n42756 = n42755 ^ n42754 ^ n12752 ;
  assign n42762 = n7077 & ~n9245 ;
  assign n42761 = n13926 & n40751 ;
  assign n42757 = n28098 ^ n11503 ^ n10727 ;
  assign n42758 = ( ~n8271 & n15932 ) | ( ~n8271 & n35812 ) | ( n15932 & n35812 ) ;
  assign n42759 = ( n7965 & n27795 ) | ( n7965 & n42758 ) | ( n27795 & n42758 ) ;
  assign n42760 = ( ~n18046 & n42757 ) | ( ~n18046 & n42759 ) | ( n42757 & n42759 ) ;
  assign n42763 = n42762 ^ n42761 ^ n42760 ;
  assign n42764 = n8142 ^ n2762 ^ n2727 ;
  assign n42767 = n20307 ^ n11690 ^ n6684 ;
  assign n42768 = n42767 ^ n17677 ^ n11640 ;
  assign n42765 = n33095 ^ n27981 ^ n26514 ;
  assign n42766 = ( n29941 & n37632 ) | ( n29941 & ~n42765 ) | ( n37632 & ~n42765 ) ;
  assign n42769 = n42768 ^ n42766 ^ n42002 ;
  assign n42770 = ( n664 & n10631 ) | ( n664 & ~n16244 ) | ( n10631 & ~n16244 ) ;
  assign n42772 = n2572 ^ n609 ^ 1'b0 ;
  assign n42771 = n35945 ^ n23121 ^ 1'b0 ;
  assign n42773 = n42772 ^ n42771 ^ n18259 ;
  assign n42774 = ( n38625 & n42770 ) | ( n38625 & n42773 ) | ( n42770 & n42773 ) ;
  assign n42775 = n11269 ^ n2541 ^ n350 ;
  assign n42776 = ~n14076 & n31823 ;
  assign n42777 = ~n16151 & n42776 ;
  assign n42778 = n12962 ^ n5596 ^ 1'b0 ;
  assign n42779 = ~n26538 & n42778 ;
  assign n42780 = n25802 ^ n17790 ^ n11836 ;
  assign n42781 = ( n8699 & n18022 ) | ( n8699 & ~n23184 ) | ( n18022 & ~n23184 ) ;
  assign n42782 = n42781 ^ n41185 ^ n19035 ;
  assign n42784 = n36280 ^ n17411 ^ n5081 ;
  assign n42783 = ( n8701 & ~n24694 ) | ( n8701 & n31761 ) | ( ~n24694 & n31761 ) ;
  assign n42785 = n42784 ^ n42783 ^ n33149 ;
  assign n42786 = n26289 ^ n23313 ^ n5143 ;
  assign n42791 = ( n6626 & ~n6780 ) | ( n6626 & n7166 ) | ( ~n6780 & n7166 ) ;
  assign n42788 = x244 & n9806 ;
  assign n42789 = n6283 & n42788 ;
  assign n42790 = n42789 ^ n12964 ^ n11913 ;
  assign n42787 = n42648 ^ n33254 ^ n2756 ;
  assign n42792 = n42791 ^ n42790 ^ n42787 ;
  assign n42793 = ( n19280 & n31488 ) | ( n19280 & n42792 ) | ( n31488 & n42792 ) ;
  assign n42794 = n10077 & n12140 ;
  assign n42795 = ~n9596 & n42794 ;
  assign n42796 = n29012 ^ n7615 ^ n4654 ;
  assign n42797 = n37629 | n42796 ;
  assign n42798 = ( n2762 & n42795 ) | ( n2762 & n42797 ) | ( n42795 & n42797 ) ;
  assign n42801 = ~n3446 & n4213 ;
  assign n42802 = ~n21209 & n42801 ;
  assign n42799 = n13908 ^ n12153 ^ n1537 ;
  assign n42800 = n42799 ^ n32069 ^ n3853 ;
  assign n42803 = n42802 ^ n42800 ^ n16002 ;
  assign n42804 = ( n4727 & n35039 ) | ( n4727 & ~n42803 ) | ( n35039 & ~n42803 ) ;
  assign n42805 = n21762 ^ n555 ^ 1'b0 ;
  assign n42806 = ( n4751 & ~n34636 ) | ( n4751 & n42805 ) | ( ~n34636 & n42805 ) ;
  assign n42807 = ( n11955 & ~n18922 ) | ( n11955 & n27562 ) | ( ~n18922 & n27562 ) ;
  assign n42808 = n42807 ^ n16242 ^ 1'b0 ;
  assign n42813 = ( ~n8828 & n22770 ) | ( ~n8828 & n35290 ) | ( n22770 & n35290 ) ;
  assign n42809 = n29019 & n30346 ;
  assign n42810 = ~x187 & n42809 ;
  assign n42811 = n36408 ^ n24216 ^ 1'b0 ;
  assign n42812 = n42810 | n42811 ;
  assign n42814 = n42813 ^ n42812 ^ n6384 ;
  assign n42815 = ~n27638 & n42361 ;
  assign n42816 = n19946 ^ n17425 ^ n7444 ;
  assign n42817 = n32766 ^ n23243 ^ n10470 ;
  assign n42818 = n42817 ^ n36132 ^ 1'b0 ;
  assign n42819 = n31991 ^ n28323 ^ n18947 ;
  assign n42820 = ( n9445 & ~n13316 ) | ( n9445 & n26034 ) | ( ~n13316 & n26034 ) ;
  assign n42821 = n5138 ^ n1021 ^ 1'b0 ;
  assign n42822 = ( n2596 & ~n7645 ) | ( n2596 & n35309 ) | ( ~n7645 & n35309 ) ;
  assign n42823 = ( n885 & n21958 ) | ( n885 & ~n42822 ) | ( n21958 & ~n42822 ) ;
  assign n42824 = ( n4292 & n24394 ) | ( n4292 & ~n25158 ) | ( n24394 & ~n25158 ) ;
  assign n42825 = ( n15382 & ~n42823 ) | ( n15382 & n42824 ) | ( ~n42823 & n42824 ) ;
  assign n42826 = ( ~n4467 & n42821 ) | ( ~n4467 & n42825 ) | ( n42821 & n42825 ) ;
  assign n42827 = n32507 ^ n26796 ^ n18886 ;
  assign n42828 = n32343 ^ n22408 ^ n13527 ;
  assign n42829 = n33728 ^ n29013 ^ n9728 ;
  assign n42830 = ( ~n25518 & n29817 ) | ( ~n25518 & n42829 ) | ( n29817 & n42829 ) ;
  assign n42831 = ( n24544 & ~n42828 ) | ( n24544 & n42830 ) | ( ~n42828 & n42830 ) ;
  assign n42832 = n37447 ^ n24197 ^ n8334 ;
  assign n42833 = ( n1105 & n3590 ) | ( n1105 & n8741 ) | ( n3590 & n8741 ) ;
  assign n42834 = ( n15558 & n41963 ) | ( n15558 & n42833 ) | ( n41963 & n42833 ) ;
  assign n42835 = n42834 ^ n11591 ^ n6250 ;
  assign n42836 = n42835 ^ n42105 ^ n12929 ;
  assign n42837 = n42836 ^ n19009 ^ n3115 ;
  assign n42838 = n32572 & ~n41036 ;
  assign n42839 = n37697 ^ n17133 ^ n6831 ;
  assign n42840 = ~n10879 & n16805 ;
  assign n42841 = n11290 & ~n12643 ;
  assign n42842 = n42840 & n42841 ;
  assign n42843 = ( n6040 & n26731 ) | ( n6040 & ~n42842 ) | ( n26731 & ~n42842 ) ;
  assign n42844 = n42638 ^ n31017 ^ n8161 ;
  assign n42845 = ( ~n12290 & n33539 ) | ( ~n12290 & n42844 ) | ( n33539 & n42844 ) ;
  assign n42846 = ( n7033 & n20316 ) | ( n7033 & ~n36546 ) | ( n20316 & ~n36546 ) ;
  assign n42847 = ( n4606 & n20817 ) | ( n4606 & n42846 ) | ( n20817 & n42846 ) ;
  assign n42848 = n19380 ^ n9217 ^ n5188 ;
  assign n42849 = ( ~n31901 & n42847 ) | ( ~n31901 & n42848 ) | ( n42847 & n42848 ) ;
  assign n42850 = n29228 ^ n7106 ^ 1'b0 ;
  assign n42851 = ~n15475 & n42850 ;
  assign n42852 = n33391 ^ n1271 ^ 1'b0 ;
  assign n42853 = n42851 & n42852 ;
  assign n42854 = n35253 ^ n4988 ^ n944 ;
  assign n42855 = ( ~n638 & n3637 ) | ( ~n638 & n17046 ) | ( n3637 & n17046 ) ;
  assign n42856 = ( n37927 & n42597 ) | ( n37927 & ~n42855 ) | ( n42597 & ~n42855 ) ;
  assign n42857 = ( ~n1550 & n2086 ) | ( ~n1550 & n34094 ) | ( n2086 & n34094 ) ;
  assign n42858 = ( n17382 & ~n36742 ) | ( n17382 & n42857 ) | ( ~n36742 & n42857 ) ;
  assign n42859 = ( n3002 & n42856 ) | ( n3002 & n42858 ) | ( n42856 & n42858 ) ;
  assign n42860 = n42859 ^ n27502 ^ 1'b0 ;
  assign n42861 = n42854 & ~n42860 ;
  assign n42864 = ( ~n1971 & n14502 ) | ( ~n1971 & n31728 ) | ( n14502 & n31728 ) ;
  assign n42862 = n5004 ^ n2641 ^ n478 ;
  assign n42863 = n42862 ^ n4182 ^ n2617 ;
  assign n42865 = n42864 ^ n42863 ^ n5706 ;
  assign n42866 = n32438 ^ n4571 ^ x61 ;
  assign n42867 = n29644 ^ n7045 ^ 1'b0 ;
  assign n42868 = n42866 | n42867 ;
  assign n42869 = ( n2675 & n30737 ) | ( n2675 & n33396 ) | ( n30737 & n33396 ) ;
  assign n42870 = ( ~n4619 & n42868 ) | ( ~n4619 & n42869 ) | ( n42868 & n42869 ) ;
  assign n42872 = ( n1104 & n7660 ) | ( n1104 & n8447 ) | ( n7660 & n8447 ) ;
  assign n42871 = ( n15069 & ~n20897 ) | ( n15069 & n34581 ) | ( ~n20897 & n34581 ) ;
  assign n42873 = n42872 ^ n42871 ^ n13572 ;
  assign n42874 = n18799 ^ n17153 ^ n4367 ;
  assign n42875 = n42874 ^ n16062 ^ n10181 ;
  assign n42876 = ( n20486 & ~n24247 ) | ( n20486 & n42875 ) | ( ~n24247 & n42875 ) ;
  assign n42877 = n5406 ^ x105 ^ 1'b0 ;
  assign n42878 = ( n10338 & n18511 ) | ( n10338 & ~n42877 ) | ( n18511 & ~n42877 ) ;
  assign n42879 = n22275 ^ n6751 ^ 1'b0 ;
  assign n42880 = n9821 & ~n42879 ;
  assign n42881 = ( n8277 & ~n33710 ) | ( n8277 & n42880 ) | ( ~n33710 & n42880 ) ;
  assign n42882 = ( n18829 & n29377 ) | ( n18829 & ~n42881 ) | ( n29377 & ~n42881 ) ;
  assign n42883 = ( n1173 & n4042 ) | ( n1173 & n7584 ) | ( n4042 & n7584 ) ;
  assign n42884 = n17191 ^ n14193 ^ n13552 ;
  assign n42885 = ( ~n26999 & n42883 ) | ( ~n26999 & n42884 ) | ( n42883 & n42884 ) ;
  assign n42886 = ( n12815 & ~n26891 ) | ( n12815 & n42885 ) | ( ~n26891 & n42885 ) ;
  assign n42887 = n21076 ^ n14149 ^ n5780 ;
  assign n42888 = n29952 ^ n19090 ^ n3061 ;
  assign n42889 = n10194 | n42888 ;
  assign n42890 = n23734 | n42889 ;
  assign n42891 = n28574 & ~n42890 ;
  assign n42892 = n15760 ^ n13859 ^ n2045 ;
  assign n42893 = ( n42887 & n42891 ) | ( n42887 & ~n42892 ) | ( n42891 & ~n42892 ) ;
  assign n42894 = n40067 ^ n39470 ^ 1'b0 ;
  assign n42895 = n20476 ^ n10146 ^ n6727 ;
  assign n42896 = n26239 ^ n18938 ^ n3428 ;
  assign n42897 = ( ~n9368 & n22117 ) | ( ~n9368 & n42896 ) | ( n22117 & n42896 ) ;
  assign n42898 = ( n4159 & ~n8778 ) | ( n4159 & n15601 ) | ( ~n8778 & n15601 ) ;
  assign n42899 = ( n16375 & n20118 ) | ( n16375 & n42898 ) | ( n20118 & n42898 ) ;
  assign n42900 = n42899 ^ n37063 ^ n15257 ;
  assign n42901 = n18488 ^ n14629 ^ n9458 ;
  assign n42902 = n40635 ^ n21478 ^ n4498 ;
  assign n42903 = n2309 & ~n11834 ;
  assign n42904 = n15717 | n35428 ;
  assign n42905 = n42904 ^ n33488 ^ 1'b0 ;
  assign n42906 = n42903 & ~n42905 ;
  assign n42907 = n6736 | n16818 ;
  assign n42908 = n39073 & ~n42907 ;
  assign n42911 = ( n10546 & n13635 ) | ( n10546 & ~n42167 ) | ( n13635 & ~n42167 ) ;
  assign n42909 = ( n2901 & n21873 ) | ( n2901 & ~n29087 ) | ( n21873 & ~n29087 ) ;
  assign n42910 = ( n30116 & n40224 ) | ( n30116 & ~n42909 ) | ( n40224 & ~n42909 ) ;
  assign n42912 = n42911 ^ n42910 ^ n31666 ;
  assign n42913 = ( n1380 & n2537 ) | ( n1380 & ~n10205 ) | ( n2537 & ~n10205 ) ;
  assign n42919 = n5289 ^ n4043 ^ x61 ;
  assign n42920 = ( n4170 & ~n25760 ) | ( n4170 & n42919 ) | ( ~n25760 & n42919 ) ;
  assign n42921 = ( ~n20188 & n23579 ) | ( ~n20188 & n42920 ) | ( n23579 & n42920 ) ;
  assign n42916 = n2017 & n28514 ;
  assign n42917 = n26678 & n42916 ;
  assign n42914 = n40115 ^ n7238 ^ n4487 ;
  assign n42915 = n42914 ^ n38956 ^ n17481 ;
  assign n42918 = n42917 ^ n42915 ^ 1'b0 ;
  assign n42922 = n42921 ^ n42918 ^ 1'b0 ;
  assign n42923 = ( ~n19483 & n21151 ) | ( ~n19483 & n25421 ) | ( n21151 & n25421 ) ;
  assign n42924 = n39335 ^ n2272 ^ 1'b0 ;
  assign n42925 = n28745 & ~n42924 ;
  assign n42926 = n31040 ^ n29070 ^ n27238 ;
  assign n42929 = ( n1357 & ~n2685 ) | ( n1357 & n12342 ) | ( ~n2685 & n12342 ) ;
  assign n42927 = n31484 ^ n8572 ^ 1'b0 ;
  assign n42928 = n18386 | n42927 ;
  assign n42930 = n42929 ^ n42928 ^ n36860 ;
  assign n42931 = n18177 ^ n16258 ^ n13543 ;
  assign n42932 = ( n38546 & n40618 ) | ( n38546 & n42931 ) | ( n40618 & n42931 ) ;
  assign n42933 = n1775 & n4264 ;
  assign n42934 = ~n42932 & n42933 ;
  assign n42935 = ( n8524 & ~n10495 ) | ( n8524 & n42934 ) | ( ~n10495 & n42934 ) ;
  assign n42936 = n24585 ^ n23908 ^ n21117 ;
  assign n42937 = n42936 ^ n19200 ^ 1'b0 ;
  assign n42938 = n42935 | n42937 ;
  assign n42939 = n11751 ^ n5850 ^ 1'b0 ;
  assign n42940 = ~n13855 & n42939 ;
  assign n42941 = n1282 & ~n4331 ;
  assign n42942 = n42941 ^ n35279 ^ n1710 ;
  assign n42943 = n42942 ^ n38941 ^ n12964 ;
  assign n42944 = ( ~n28356 & n42940 ) | ( ~n28356 & n42943 ) | ( n42940 & n42943 ) ;
  assign n42945 = n24782 ^ n7887 ^ 1'b0 ;
  assign n42946 = n29841 ^ n3689 ^ 1'b0 ;
  assign n42947 = n9339 & n42946 ;
  assign n42948 = ( n23805 & ~n31999 ) | ( n23805 & n42947 ) | ( ~n31999 & n42947 ) ;
  assign n42949 = n42948 ^ n41389 ^ n9165 ;
  assign n42950 = n6545 ^ n5763 ^ 1'b0 ;
  assign n42951 = x38 & n21503 ;
  assign n42952 = n42951 ^ n34340 ^ n4582 ;
  assign n42954 = ( n10389 & ~n11595 ) | ( n10389 & n22917 ) | ( ~n11595 & n22917 ) ;
  assign n42953 = ( n3355 & n10788 ) | ( n3355 & ~n28669 ) | ( n10788 & ~n28669 ) ;
  assign n42955 = n42954 ^ n42953 ^ n18933 ;
  assign n42956 = ( n2765 & n41955 ) | ( n2765 & n42955 ) | ( n41955 & n42955 ) ;
  assign n42957 = n25961 & ~n42956 ;
  assign n42958 = n521 & ~n1079 ;
  assign n42959 = n42958 ^ n14784 ^ 1'b0 ;
  assign n42960 = ( n4922 & ~n35036 ) | ( n4922 & n40278 ) | ( ~n35036 & n40278 ) ;
  assign n42961 = ( n2959 & n37986 ) | ( n2959 & n42960 ) | ( n37986 & n42960 ) ;
  assign n42962 = n27664 & n40984 ;
  assign n42963 = ~n1529 & n18110 ;
  assign n42964 = n30105 & n42963 ;
  assign n42965 = n42964 ^ n38637 ^ n4925 ;
  assign n42966 = n25546 ^ n19643 ^ 1'b0 ;
  assign n42967 = ( n8364 & ~n15029 ) | ( n8364 & n42966 ) | ( ~n15029 & n42966 ) ;
  assign n42968 = n42967 ^ n28143 ^ n2673 ;
  assign n42969 = ( n6832 & ~n14807 ) | ( n6832 & n15156 ) | ( ~n14807 & n15156 ) ;
  assign n42970 = ( n6450 & ~n16425 ) | ( n6450 & n32053 ) | ( ~n16425 & n32053 ) ;
  assign n42971 = n42970 ^ n34001 ^ n2925 ;
  assign n42972 = n10323 ^ n9783 ^ n2656 ;
  assign n42973 = n42972 ^ n31933 ^ n11088 ;
  assign n42976 = n11322 ^ n4761 ^ n1645 ;
  assign n42974 = ( n12119 & n20745 ) | ( n12119 & n24358 ) | ( n20745 & n24358 ) ;
  assign n42975 = n42974 ^ n8861 ^ n1874 ;
  assign n42977 = n42976 ^ n42975 ^ n19048 ;
  assign n42978 = n42518 ^ n23037 ^ n19850 ;
  assign n42979 = ~n14022 & n42978 ;
  assign n42980 = n26615 | n33551 ;
  assign n42981 = n42980 ^ n8929 ^ 1'b0 ;
  assign n42982 = ( n25235 & n40554 ) | ( n25235 & n42981 ) | ( n40554 & n42981 ) ;
  assign n42983 = n16775 ^ n6499 ^ n1600 ;
  assign n42984 = n42983 ^ n19814 ^ n16841 ;
  assign n42985 = ( n2549 & n4261 ) | ( n2549 & n10883 ) | ( n4261 & n10883 ) ;
  assign n42986 = n12448 ^ n10797 ^ n268 ;
  assign n42987 = ( ~n3044 & n30113 ) | ( ~n3044 & n39607 ) | ( n30113 & n39607 ) ;
  assign n42988 = ( ~n42985 & n42986 ) | ( ~n42985 & n42987 ) | ( n42986 & n42987 ) ;
  assign n42989 = n15107 & ~n42988 ;
  assign n42991 = n34352 ^ n30251 ^ n14142 ;
  assign n42990 = n31016 ^ n22317 ^ n18874 ;
  assign n42992 = n42991 ^ n42990 ^ 1'b0 ;
  assign n42993 = ~n22483 & n42992 ;
  assign n42994 = n18313 ^ n6216 ^ n350 ;
  assign n42995 = ( ~n587 & n29843 ) | ( ~n587 & n42994 ) | ( n29843 & n42994 ) ;
  assign n42996 = n31299 & n38443 ;
  assign n42997 = n42996 ^ n35180 ^ n32102 ;
  assign n42998 = ( n25059 & n42995 ) | ( n25059 & n42997 ) | ( n42995 & n42997 ) ;
  assign n42999 = ( ~n398 & n2389 ) | ( ~n398 & n8922 ) | ( n2389 & n8922 ) ;
  assign n43000 = n42999 ^ n37495 ^ n15658 ;
  assign n43001 = n19707 & ~n43000 ;
  assign n43002 = ( n1189 & n5668 ) | ( n1189 & ~n34481 ) | ( n5668 & ~n34481 ) ;
  assign n43003 = n16272 ^ n11286 ^ n2916 ;
  assign n43005 = n18325 & n19081 ;
  assign n43006 = n43005 ^ n8501 ^ 1'b0 ;
  assign n43004 = n25395 ^ n11102 ^ n6285 ;
  assign n43007 = n43006 ^ n43004 ^ n23456 ;
  assign n43008 = n13939 & ~n43007 ;
  assign n43010 = ( ~n379 & n5386 ) | ( ~n379 & n16034 ) | ( n5386 & n16034 ) ;
  assign n43009 = n30168 ^ n10406 ^ n4377 ;
  assign n43011 = n43010 ^ n43009 ^ n22560 ;
  assign n43012 = n43011 ^ n21761 ^ 1'b0 ;
  assign n43017 = ( n11353 & n26658 ) | ( n11353 & ~n32936 ) | ( n26658 & ~n32936 ) ;
  assign n43016 = ( n12997 & n19403 ) | ( n12997 & n31887 ) | ( n19403 & n31887 ) ;
  assign n43013 = ( n13053 & n16263 ) | ( n13053 & n20478 ) | ( n16263 & n20478 ) ;
  assign n43014 = ( n13079 & n28127 ) | ( n13079 & n43013 ) | ( n28127 & n43013 ) ;
  assign n43015 = ( n3400 & n27764 ) | ( n3400 & n43014 ) | ( n27764 & n43014 ) ;
  assign n43018 = n43017 ^ n43016 ^ n43015 ;
  assign n43019 = ( n313 & ~n1268 ) | ( n313 & n2645 ) | ( ~n1268 & n2645 ) ;
  assign n43020 = n32063 ^ n5448 ^ n4824 ;
  assign n43021 = ( ~n16938 & n43019 ) | ( ~n16938 & n43020 ) | ( n43019 & n43020 ) ;
  assign n43022 = ( n6440 & ~n28421 ) | ( n6440 & n42009 ) | ( ~n28421 & n42009 ) ;
  assign n43025 = n3716 | n10203 ;
  assign n43026 = n43025 ^ n19610 ^ 1'b0 ;
  assign n43023 = n21127 ^ n12724 ^ n3533 ;
  assign n43024 = n43023 ^ n35085 ^ n11481 ;
  assign n43027 = n43026 ^ n43024 ^ 1'b0 ;
  assign n43028 = n16468 ^ n14154 ^ n8605 ;
  assign n43029 = ( n6825 & ~n15229 ) | ( n6825 & n39426 ) | ( ~n15229 & n39426 ) ;
  assign n43030 = ( ~n7604 & n43028 ) | ( ~n7604 & n43029 ) | ( n43028 & n43029 ) ;
  assign n43031 = ( n7057 & n19682 ) | ( n7057 & ~n22517 ) | ( n19682 & ~n22517 ) ;
  assign n43032 = ( n27976 & ~n32767 ) | ( n27976 & n43031 ) | ( ~n32767 & n43031 ) ;
  assign n43033 = ( ~n7282 & n19123 ) | ( ~n7282 & n40263 ) | ( n19123 & n40263 ) ;
  assign n43034 = n34921 | n43033 ;
  assign n43035 = n37610 ^ n28784 ^ 1'b0 ;
  assign n43036 = n7989 | n43035 ;
  assign n43037 = n6162 | n16572 ;
  assign n43038 = n42113 ^ n18695 ^ 1'b0 ;
  assign n43039 = n43037 & ~n43038 ;
  assign n43040 = n32630 ^ n8914 ^ n3907 ;
  assign n43041 = ( n11376 & n41854 ) | ( n11376 & ~n43040 ) | ( n41854 & ~n43040 ) ;
  assign n43042 = ( ~n17522 & n24128 ) | ( ~n17522 & n38900 ) | ( n24128 & n38900 ) ;
  assign n43043 = ( n5474 & n37776 ) | ( n5474 & ~n43042 ) | ( n37776 & ~n43042 ) ;
  assign n43044 = n40758 ^ n32215 ^ 1'b0 ;
  assign n43045 = n43044 ^ n38710 ^ n24125 ;
  assign n43046 = n37207 ^ n32947 ^ 1'b0 ;
  assign n43047 = ( n15762 & n31020 ) | ( n15762 & ~n35868 ) | ( n31020 & ~n35868 ) ;
  assign n43048 = ( n2155 & n13248 ) | ( n2155 & n36972 ) | ( n13248 & n36972 ) ;
  assign n43049 = ~n27990 & n43048 ;
  assign n43050 = ~n13040 & n38513 ;
  assign n43051 = ~n9067 & n43050 ;
  assign n43052 = ( n23357 & ~n43049 ) | ( n23357 & n43051 ) | ( ~n43049 & n43051 ) ;
  assign n43053 = ( ~n10983 & n11410 ) | ( ~n10983 & n43052 ) | ( n11410 & n43052 ) ;
  assign n43054 = n21383 ^ n7425 ^ 1'b0 ;
  assign n43055 = n12117 ^ n11611 ^ 1'b0 ;
  assign n43056 = n27744 & ~n43055 ;
  assign n43057 = n22010 & n43056 ;
  assign n43058 = n30202 ^ n5169 ^ 1'b0 ;
  assign n43061 = n10493 & ~n21004 ;
  assign n43062 = n15259 & n43061 ;
  assign n43059 = n38207 ^ n28326 ^ n2781 ;
  assign n43060 = n43059 ^ n17882 ^ n10588 ;
  assign n43063 = n43062 ^ n43060 ^ 1'b0 ;
  assign n43064 = n30392 ^ n14056 ^ n11600 ;
  assign n43065 = ( n7905 & ~n31170 ) | ( n7905 & n43064 ) | ( ~n31170 & n43064 ) ;
  assign n43066 = ( n43058 & ~n43063 ) | ( n43058 & n43065 ) | ( ~n43063 & n43065 ) ;
  assign n43067 = ( ~n14364 & n27384 ) | ( ~n14364 & n32560 ) | ( n27384 & n32560 ) ;
  assign n43068 = n43067 ^ n26366 ^ n1363 ;
  assign n43069 = n33922 ^ n33535 ^ n6267 ;
  assign n43070 = n14749 | n43069 ;
  assign n43071 = n21340 ^ n18349 ^ n8992 ;
  assign n43072 = n29516 & ~n43071 ;
  assign n43073 = n43072 ^ n11864 ^ 1'b0 ;
  assign n43078 = n10428 ^ n7149 ^ n4517 ;
  assign n43074 = n30723 ^ n11211 ^ 1'b0 ;
  assign n43075 = n1426 & n43074 ;
  assign n43076 = n43075 ^ n9379 ^ n6400 ;
  assign n43077 = n43076 ^ n19388 ^ n2279 ;
  assign n43079 = n43078 ^ n43077 ^ n38729 ;
  assign n43080 = ( n1308 & n4665 ) | ( n1308 & n14238 ) | ( n4665 & n14238 ) ;
  assign n43081 = n30987 & n38112 ;
  assign n43082 = n19445 & n43081 ;
  assign n43083 = ( n11069 & ~n43080 ) | ( n11069 & n43082 ) | ( ~n43080 & n43082 ) ;
  assign n43084 = n32735 & n33587 ;
  assign n43085 = n19415 ^ n11038 ^ n3635 ;
  assign n43086 = n43085 ^ n20869 ^ n11795 ;
  assign n43087 = ( n4453 & n22729 ) | ( n4453 & n32767 ) | ( n22729 & n32767 ) ;
  assign n43090 = n28720 ^ n5670 ^ 1'b0 ;
  assign n43091 = n10124 & n43090 ;
  assign n43088 = ( ~n21166 & n21550 ) | ( ~n21166 & n24958 ) | ( n21550 & n24958 ) ;
  assign n43089 = ( n7191 & n27382 ) | ( n7191 & n43088 ) | ( n27382 & n43088 ) ;
  assign n43092 = n43091 ^ n43089 ^ n13617 ;
  assign n43093 = n40750 ^ n26400 ^ 1'b0 ;
  assign n43094 = ( ~n709 & n26011 ) | ( ~n709 & n43093 ) | ( n26011 & n43093 ) ;
  assign n43095 = n43094 ^ n31569 ^ n22844 ;
  assign n43096 = n35398 ^ n23291 ^ 1'b0 ;
  assign n43097 = ( n2431 & ~n23987 ) | ( n2431 & n29002 ) | ( ~n23987 & n29002 ) ;
  assign n43098 = n43097 ^ n13761 ^ n3580 ;
  assign n43099 = ( n33122 & n43096 ) | ( n33122 & ~n43098 ) | ( n43096 & ~n43098 ) ;
  assign n43100 = n31551 ^ n26534 ^ n1301 ;
  assign n43101 = n1548 & ~n43100 ;
  assign n43102 = n11465 & n43101 ;
  assign n43103 = ( n1564 & n15313 ) | ( n1564 & ~n18143 ) | ( n15313 & ~n18143 ) ;
  assign n43104 = n43103 ^ n7736 ^ n5152 ;
  assign n43105 = n43104 ^ n30605 ^ n7802 ;
  assign n43106 = n41860 ^ n32526 ^ n29377 ;
  assign n43107 = n8646 & ~n21379 ;
  assign n43108 = n1003 & ~n7214 ;
  assign n43109 = n43108 ^ n27848 ^ 1'b0 ;
  assign n43110 = ( ~n19308 & n43107 ) | ( ~n19308 & n43109 ) | ( n43107 & n43109 ) ;
  assign n43111 = n31585 ^ n30006 ^ n24226 ;
  assign n43112 = n11058 & n23057 ;
  assign n43113 = n27381 & n43112 ;
  assign n43114 = ( n726 & ~n753 ) | ( n726 & n43113 ) | ( ~n753 & n43113 ) ;
  assign n43115 = ( n9374 & n15046 ) | ( n9374 & n15211 ) | ( n15046 & n15211 ) ;
  assign n43116 = n43115 ^ n18238 ^ n14180 ;
  assign n43117 = ( n10910 & ~n19466 ) | ( n10910 & n26194 ) | ( ~n19466 & n26194 ) ;
  assign n43118 = n43117 ^ n19108 ^ n2444 ;
  assign n43119 = ( n10156 & n16022 ) | ( n10156 & ~n34800 ) | ( n16022 & ~n34800 ) ;
  assign n43120 = n28820 ^ n24568 ^ n8985 ;
  assign n43121 = ( n10434 & n23009 ) | ( n10434 & n38067 ) | ( n23009 & n38067 ) ;
  assign n43122 = n38598 ^ n24460 ^ n825 ;
  assign n43123 = ( ~n11915 & n21919 ) | ( ~n11915 & n41222 ) | ( n21919 & n41222 ) ;
  assign n43124 = n43123 ^ n28844 ^ n11815 ;
  assign n43125 = n25688 ^ n21623 ^ n3523 ;
  assign n43126 = n43125 ^ n14103 ^ n7544 ;
  assign n43127 = n43126 ^ n20730 ^ n17902 ;
  assign n43128 = n38404 ^ n22332 ^ n2670 ;
  assign n43129 = n36852 & ~n41112 ;
  assign n43130 = ~n1996 & n43129 ;
  assign n43131 = n4750 | n5608 ;
  assign n43132 = n5769 & ~n12978 ;
  assign n43133 = ( n5918 & n20551 ) | ( n5918 & ~n43132 ) | ( n20551 & ~n43132 ) ;
  assign n43134 = n43133 ^ n22569 ^ n747 ;
  assign n43135 = n30826 ^ n11279 ^ n2527 ;
  assign n43136 = n20586 ^ n17737 ^ n12986 ;
  assign n43137 = n24730 ^ n23409 ^ n628 ;
  assign n43138 = ( n6579 & n7645 ) | ( n6579 & ~n43137 ) | ( n7645 & ~n43137 ) ;
  assign n43139 = n7605 ^ n5221 ^ n5120 ;
  assign n43140 = n43139 ^ n29544 ^ n16544 ;
  assign n43141 = ( n4500 & n16742 ) | ( n4500 & n43140 ) | ( n16742 & n43140 ) ;
  assign n43142 = n43141 ^ n29309 ^ n5851 ;
  assign n43143 = n43142 ^ n38946 ^ n32923 ;
  assign n43144 = n32991 ^ n27585 ^ n22871 ;
  assign n43145 = ( n7381 & ~n26207 ) | ( n7381 & n40149 ) | ( ~n26207 & n40149 ) ;
  assign n43146 = ( n11929 & n23324 ) | ( n11929 & ~n33972 ) | ( n23324 & ~n33972 ) ;
  assign n43147 = n23471 & ~n43146 ;
  assign n43148 = ~n1220 & n43147 ;
  assign n43149 = n20273 ^ n3106 ^ 1'b0 ;
  assign n43150 = ~n4780 & n9789 ;
  assign n43151 = ( ~n5958 & n20398 ) | ( ~n5958 & n42372 ) | ( n20398 & n42372 ) ;
  assign n43152 = n43151 ^ n40606 ^ n38111 ;
  assign n43153 = ( n11901 & ~n16868 ) | ( n11901 & n30439 ) | ( ~n16868 & n30439 ) ;
  assign n43154 = n26006 ^ n14919 ^ n2394 ;
  assign n43155 = n31097 ^ n879 ^ n792 ;
  assign n43156 = ( n10538 & n43154 ) | ( n10538 & n43155 ) | ( n43154 & n43155 ) ;
  assign n43157 = ( n17468 & n43153 ) | ( n17468 & n43156 ) | ( n43153 & n43156 ) ;
  assign n43158 = n43157 ^ n27751 ^ n13994 ;
  assign n43160 = ( ~n3185 & n14194 ) | ( ~n3185 & n28192 ) | ( n14194 & n28192 ) ;
  assign n43159 = n23958 ^ n16676 ^ n5288 ;
  assign n43161 = n43160 ^ n43159 ^ 1'b0 ;
  assign n43162 = n23930 & ~n43161 ;
  assign n43163 = n43162 ^ n17356 ^ 1'b0 ;
  assign n43164 = n23495 | n26529 ;
  assign n43165 = n536 & ~n43164 ;
  assign n43166 = ( n9357 & ~n23517 ) | ( n9357 & n34836 ) | ( ~n23517 & n34836 ) ;
  assign n43167 = ( n2827 & ~n20112 ) | ( n2827 & n26248 ) | ( ~n20112 & n26248 ) ;
  assign n43168 = ~n14233 & n14592 ;
  assign n43169 = n14824 & n43168 ;
  assign n43170 = ( ~n19359 & n30064 ) | ( ~n19359 & n43169 ) | ( n30064 & n43169 ) ;
  assign n43171 = n43170 ^ n10205 ^ n9659 ;
  assign n43172 = ( n25393 & n30286 ) | ( n25393 & n43171 ) | ( n30286 & n43171 ) ;
  assign n43173 = ( n12408 & ~n43167 ) | ( n12408 & n43172 ) | ( ~n43167 & n43172 ) ;
  assign n43174 = n43173 ^ n939 ^ 1'b0 ;
  assign n43175 = n41192 ^ n13704 ^ n6517 ;
  assign n43176 = n25915 ^ n5229 ^ n3204 ;
  assign n43177 = ( ~n15173 & n35542 ) | ( ~n15173 & n43176 ) | ( n35542 & n43176 ) ;
  assign n43178 = ( ~n7003 & n28931 ) | ( ~n7003 & n43177 ) | ( n28931 & n43177 ) ;
  assign n43179 = n17652 ^ n13429 ^ n865 ;
  assign n43180 = n43179 ^ n38207 ^ n8673 ;
  assign n43181 = n43180 ^ n18598 ^ n11405 ;
  assign n43182 = n31520 ^ n24555 ^ n7047 ;
  assign n43183 = n7090 | n8893 ;
  assign n43184 = n32391 & ~n43183 ;
  assign n43185 = ( n13857 & n36009 ) | ( n13857 & ~n38852 ) | ( n36009 & ~n38852 ) ;
  assign n43186 = n5402 | n43185 ;
  assign n43187 = n43186 ^ n11275 ^ 1'b0 ;
  assign n43188 = ( n14913 & n22410 ) | ( n14913 & ~n23191 ) | ( n22410 & ~n23191 ) ;
  assign n43189 = ( n24174 & ~n34805 ) | ( n24174 & n43188 ) | ( ~n34805 & n43188 ) ;
  assign n43190 = n14914 ^ n6489 ^ n3622 ;
  assign n43191 = ( n3192 & n33633 ) | ( n3192 & ~n43190 ) | ( n33633 & ~n43190 ) ;
  assign n43192 = ( ~n2054 & n7723 ) | ( ~n2054 & n43191 ) | ( n7723 & n43191 ) ;
  assign n43193 = ( n4911 & ~n6480 ) | ( n4911 & n17066 ) | ( ~n6480 & n17066 ) ;
  assign n43194 = n43193 ^ n32416 ^ n7306 ;
  assign n43195 = ( n24061 & ~n28250 ) | ( n24061 & n33720 ) | ( ~n28250 & n33720 ) ;
  assign n43197 = n725 & n6970 ;
  assign n43198 = ~n24517 & n43197 ;
  assign n43196 = ( n8504 & ~n16499 ) | ( n8504 & n25199 ) | ( ~n16499 & n25199 ) ;
  assign n43199 = n43198 ^ n43196 ^ n20291 ;
  assign n43200 = n30904 ^ n22503 ^ n21595 ;
  assign n43201 = ( n9415 & n15972 ) | ( n9415 & ~n32219 ) | ( n15972 & ~n32219 ) ;
  assign n43202 = n43201 ^ n36279 ^ n15754 ;
  assign n43203 = n43202 ^ n25997 ^ n22622 ;
  assign n43204 = ( n5117 & n42126 ) | ( n5117 & ~n43203 ) | ( n42126 & ~n43203 ) ;
  assign n43208 = n24892 ^ n22002 ^ n4877 ;
  assign n43205 = n15564 ^ n5850 ^ n1367 ;
  assign n43206 = n13809 & ~n43205 ;
  assign n43207 = n43206 ^ n3802 ^ 1'b0 ;
  assign n43209 = n43208 ^ n43207 ^ n18257 ;
  assign n43212 = n9721 ^ n5876 ^ 1'b0 ;
  assign n43213 = n7922 & ~n43212 ;
  assign n43210 = ( n2052 & n13353 ) | ( n2052 & n22087 ) | ( n13353 & n22087 ) ;
  assign n43211 = ( x24 & n39067 ) | ( x24 & n43210 ) | ( n39067 & n43210 ) ;
  assign n43214 = n43213 ^ n43211 ^ n9070 ;
  assign n43215 = ( n5649 & ~n8984 ) | ( n5649 & n43049 ) | ( ~n8984 & n43049 ) ;
  assign n43216 = n43215 ^ n37715 ^ n3460 ;
  assign n43217 = n30292 ^ n16668 ^ n9405 ;
  assign n43218 = ( ~n23075 & n26739 ) | ( ~n23075 & n33157 ) | ( n26739 & n33157 ) ;
  assign n43219 = n43217 & ~n43218 ;
  assign n43220 = ( n10158 & n37294 ) | ( n10158 & n42288 ) | ( n37294 & n42288 ) ;
  assign n43221 = n8869 ^ n6618 ^ n3957 ;
  assign n43222 = n43221 ^ n14143 ^ n9429 ;
  assign n43223 = ( ~n14558 & n24654 ) | ( ~n14558 & n43222 ) | ( n24654 & n43222 ) ;
  assign n43224 = n25351 ^ n25233 ^ 1'b0 ;
  assign n43225 = n31499 ^ n6644 ^ n595 ;
  assign n43226 = n1389 & ~n43225 ;
  assign n43227 = n25407 & ~n34829 ;
  assign n43229 = ~n444 & n5051 ;
  assign n43228 = ( ~n13483 & n14808 ) | ( ~n13483 & n29313 ) | ( n14808 & n29313 ) ;
  assign n43230 = n43229 ^ n43228 ^ n39200 ;
  assign n43231 = n34405 ^ n15840 ^ n7089 ;
  assign n43232 = n43231 ^ n32799 ^ n1432 ;
  assign n43233 = n25408 ^ n21167 ^ n17886 ;
  assign n43234 = n7250 ^ n4172 ^ n824 ;
  assign n43235 = n43234 ^ n23544 ^ n13793 ;
  assign n43236 = n43235 ^ n22901 ^ n15049 ;
  assign n43237 = ( ~n14751 & n17131 ) | ( ~n14751 & n43236 ) | ( n17131 & n43236 ) ;
  assign n43238 = ( n18860 & ~n19686 ) | ( n18860 & n30806 ) | ( ~n19686 & n30806 ) ;
  assign n43239 = ( n801 & n40108 ) | ( n801 & n43238 ) | ( n40108 & n43238 ) ;
  assign n43240 = n29835 ^ n20180 ^ n14379 ;
  assign n43241 = n3665 & n43240 ;
  assign n43242 = n30772 ^ n27983 ^ n22098 ;
  assign n43243 = n8828 & ~n43242 ;
  assign n43244 = ~n39938 & n43243 ;
  assign n43245 = n25647 ^ n21168 ^ n1315 ;
  assign n43246 = n20522 ^ n16721 ^ n3475 ;
  assign n43247 = ( n24165 & n30227 ) | ( n24165 & ~n43246 ) | ( n30227 & ~n43246 ) ;
  assign n43248 = n43247 ^ n34858 ^ n1494 ;
  assign n43250 = n18526 ^ n13896 ^ x56 ;
  assign n43249 = n35929 ^ n29516 ^ n22494 ;
  assign n43251 = n43250 ^ n43249 ^ n6546 ;
  assign n43252 = ( ~n1900 & n11672 ) | ( ~n1900 & n17581 ) | ( n11672 & n17581 ) ;
  assign n43253 = n43252 ^ n1501 ^ 1'b0 ;
  assign n43254 = n43253 ^ n42741 ^ n15852 ;
  assign n43255 = n15684 ^ n11963 ^ n2943 ;
  assign n43256 = n43255 ^ n18923 ^ n17526 ;
  assign n43257 = ( n26396 & ~n27575 ) | ( n26396 & n43256 ) | ( ~n27575 & n43256 ) ;
  assign n43258 = ( ~x93 & n27110 ) | ( ~x93 & n36303 ) | ( n27110 & n36303 ) ;
  assign n43259 = ( n20936 & n30205 ) | ( n20936 & n43258 ) | ( n30205 & n43258 ) ;
  assign n43260 = ( n2259 & ~n18901 ) | ( n2259 & n43259 ) | ( ~n18901 & n43259 ) ;
  assign n43261 = ( n1673 & n10753 ) | ( n1673 & ~n43260 ) | ( n10753 & ~n43260 ) ;
  assign n43262 = n6118 | n38045 ;
  assign n43263 = n43262 ^ n39393 ^ 1'b0 ;
  assign n43264 = n21203 | n34132 ;
  assign n43265 = n15423 & ~n43264 ;
  assign n43266 = n33185 ^ n28867 ^ 1'b0 ;
  assign n43270 = n33523 ^ n31960 ^ n13762 ;
  assign n43267 = ( n5909 & n11181 ) | ( n5909 & ~n12344 ) | ( n11181 & ~n12344 ) ;
  assign n43268 = n43267 ^ n30859 ^ n7248 ;
  assign n43269 = n43268 ^ n35555 ^ n19432 ;
  assign n43271 = n43270 ^ n43269 ^ n16258 ;
  assign n43272 = n43271 ^ n27699 ^ n8478 ;
  assign n43277 = n5969 | n36290 ;
  assign n43278 = n43277 ^ n6103 ^ 1'b0 ;
  assign n43273 = n24655 & ~n29758 ;
  assign n43274 = n10206 & n43273 ;
  assign n43275 = n43274 ^ n7884 ^ 1'b0 ;
  assign n43276 = ( n2106 & ~n27249 ) | ( n2106 & n43275 ) | ( ~n27249 & n43275 ) ;
  assign n43279 = n43278 ^ n43276 ^ n1507 ;
  assign n43280 = n43279 ^ n21821 ^ n20875 ;
  assign n43281 = ~n13479 & n35034 ;
  assign n43282 = ( n7606 & n20033 ) | ( n7606 & ~n30615 ) | ( n20033 & ~n30615 ) ;
  assign n43283 = ( n2424 & ~n9729 ) | ( n2424 & n43282 ) | ( ~n9729 & n43282 ) ;
  assign n43284 = ( n6906 & n11809 ) | ( n6906 & n30350 ) | ( n11809 & n30350 ) ;
  assign n43285 = n43284 ^ n22191 ^ n21286 ;
  assign n43286 = n43285 ^ n23638 ^ n18325 ;
  assign n43287 = ( n737 & ~n3674 ) | ( n737 & n13020 ) | ( ~n3674 & n13020 ) ;
  assign n43288 = ( n5625 & n19492 ) | ( n5625 & ~n27868 ) | ( n19492 & ~n27868 ) ;
  assign n43289 = n43288 ^ n40596 ^ n4654 ;
  assign n43290 = ( n6186 & ~n15634 ) | ( n6186 & n43289 ) | ( ~n15634 & n43289 ) ;
  assign n43291 = ( n43160 & n43287 ) | ( n43160 & ~n43290 ) | ( n43287 & ~n43290 ) ;
  assign n43292 = ( n770 & ~n2068 ) | ( n770 & n3849 ) | ( ~n2068 & n3849 ) ;
  assign n43293 = ( ~n2213 & n11834 ) | ( ~n2213 & n43292 ) | ( n11834 & n43292 ) ;
  assign n43294 = n20495 ^ n13235 ^ 1'b0 ;
  assign n43295 = ( x231 & n2687 ) | ( x231 & ~n16252 ) | ( n2687 & ~n16252 ) ;
  assign n43296 = n34287 | n43295 ;
  assign n43297 = ( x28 & n11928 ) | ( x28 & ~n14553 ) | ( n11928 & ~n14553 ) ;
  assign n43298 = n43297 ^ n24665 ^ n508 ;
  assign n43299 = ( n1102 & ~n12124 ) | ( n1102 & n43298 ) | ( ~n12124 & n43298 ) ;
  assign n43300 = ( n6074 & n28236 ) | ( n6074 & n41895 ) | ( n28236 & n41895 ) ;
  assign n43301 = ( n10449 & n28790 ) | ( n10449 & n28826 ) | ( n28790 & n28826 ) ;
  assign n43306 = ( n12167 & ~n16598 ) | ( n12167 & n38338 ) | ( ~n16598 & n38338 ) ;
  assign n43307 = ( n7644 & ~n32018 ) | ( n7644 & n43306 ) | ( ~n32018 & n43306 ) ;
  assign n43308 = ( n1007 & n35664 ) | ( n1007 & ~n43307 ) | ( n35664 & ~n43307 ) ;
  assign n43302 = ( n9533 & ~n10474 ) | ( n9533 & n22887 ) | ( ~n10474 & n22887 ) ;
  assign n43303 = n34929 ^ n265 ^ 1'b0 ;
  assign n43304 = ~n4400 & n43303 ;
  assign n43305 = ( n11149 & ~n43302 ) | ( n11149 & n43304 ) | ( ~n43302 & n43304 ) ;
  assign n43309 = n43308 ^ n43305 ^ n38085 ;
  assign n43310 = n7405 ^ n4888 ^ n1428 ;
  assign n43311 = ( n4286 & ~n37958 ) | ( n4286 & n43310 ) | ( ~n37958 & n43310 ) ;
  assign n43312 = ( n19052 & n20676 ) | ( n19052 & ~n22769 ) | ( n20676 & ~n22769 ) ;
  assign n43313 = n43312 ^ n14050 ^ n3862 ;
  assign n43316 = n35988 ^ n14273 ^ n6472 ;
  assign n43314 = ( n6174 & n7548 ) | ( n6174 & n40163 ) | ( n7548 & n40163 ) ;
  assign n43315 = n43314 ^ n41088 ^ n34520 ;
  assign n43317 = n43316 ^ n43315 ^ n31961 ;
  assign n43318 = n7082 | n14213 ;
  assign n43319 = ( n7470 & n9352 ) | ( n7470 & ~n17438 ) | ( n9352 & ~n17438 ) ;
  assign n43320 = ( ~n4209 & n43318 ) | ( ~n4209 & n43319 ) | ( n43318 & n43319 ) ;
  assign n43321 = n40797 ^ n35433 ^ n9146 ;
  assign n43322 = ( n627 & n38690 ) | ( n627 & ~n38894 ) | ( n38690 & ~n38894 ) ;
  assign n43323 = ( n7047 & n12044 ) | ( n7047 & n43213 ) | ( n12044 & n43213 ) ;
  assign n43324 = n43323 ^ n23383 ^ n5644 ;
  assign n43325 = ( ~n26574 & n43322 ) | ( ~n26574 & n43324 ) | ( n43322 & n43324 ) ;
  assign n43326 = n3422 & ~n12078 ;
  assign n43327 = n43326 ^ n7449 ^ n3178 ;
  assign n43328 = n43327 ^ n31761 ^ n13155 ;
  assign n43329 = n2976 & n19460 ;
  assign n43330 = ~n23817 & n43329 ;
  assign n43331 = n36252 ^ n14629 ^ n7122 ;
  assign n43332 = n4027 ^ n3120 ^ n1044 ;
  assign n43333 = n43332 ^ n20279 ^ n4964 ;
  assign n43334 = ( ~n19250 & n30480 ) | ( ~n19250 & n43333 ) | ( n30480 & n43333 ) ;
  assign n43335 = n43334 ^ n36397 ^ n4791 ;
  assign n43336 = n26539 ^ n710 ^ n371 ;
  assign n43337 = n42299 ^ n17544 ^ n16257 ;
  assign n43338 = ( ~n25148 & n43336 ) | ( ~n25148 & n43337 ) | ( n43336 & n43337 ) ;
  assign n43339 = n35066 ^ n13275 ^ n11282 ;
  assign n43340 = n37097 ^ n19797 ^ n9825 ;
  assign n43341 = ( n3834 & n24881 ) | ( n3834 & n43340 ) | ( n24881 & n43340 ) ;
  assign n43342 = n43341 ^ n14553 ^ n2070 ;
  assign n43345 = n15638 & n17359 ;
  assign n43344 = n26223 ^ n19806 ^ n4370 ;
  assign n43343 = n3375 & ~n29474 ;
  assign n43346 = n43345 ^ n43344 ^ n43343 ;
  assign n43347 = n35906 ^ n27046 ^ n6956 ;
  assign n43348 = ~n4452 & n42624 ;
  assign n43349 = n15063 & n43348 ;
  assign n43350 = n29662 ^ n25361 ^ n14417 ;
  assign n43351 = ~n16264 & n24008 ;
  assign n43352 = ( ~n4493 & n9359 ) | ( ~n4493 & n24797 ) | ( n9359 & n24797 ) ;
  assign n43353 = n43352 ^ n32084 ^ n5027 ;
  assign n43354 = n27901 ^ n3022 ^ x143 ;
  assign n43355 = ( n12914 & n40038 ) | ( n12914 & n43354 ) | ( n40038 & n43354 ) ;
  assign n43360 = ( n17923 & n31492 ) | ( n17923 & n39711 ) | ( n31492 & n39711 ) ;
  assign n43356 = n42268 ^ n7963 ^ n5230 ;
  assign n43357 = n36605 ^ n36172 ^ n9565 ;
  assign n43358 = n43357 ^ n30198 ^ n2543 ;
  assign n43359 = n43356 | n43358 ;
  assign n43361 = n43360 ^ n43359 ^ n32983 ;
  assign n43362 = ( ~n23374 & n25411 ) | ( ~n23374 & n28390 ) | ( n25411 & n28390 ) ;
  assign n43364 = ( n11266 & n37381 ) | ( n11266 & ~n37528 ) | ( n37381 & ~n37528 ) ;
  assign n43363 = n31000 ^ n12718 ^ n5682 ;
  assign n43365 = n43364 ^ n43363 ^ n24620 ;
  assign n43366 = ~n4291 & n37243 ;
  assign n43367 = n6840 & n43366 ;
  assign n43368 = ( n22435 & n27865 ) | ( n22435 & n43367 ) | ( n27865 & n43367 ) ;
  assign n43369 = n5097 & ~n26882 ;
  assign n43370 = ~n16591 & n43369 ;
  assign n43371 = n43370 ^ n21415 ^ n10081 ;
  assign n43372 = n43371 ^ n26368 ^ n7478 ;
  assign n43373 = n2387 & ~n8363 ;
  assign n43374 = ~n30190 & n43373 ;
  assign n43375 = ( x136 & ~n12337 ) | ( x136 & n43374 ) | ( ~n12337 & n43374 ) ;
  assign n43376 = n6058 & n43375 ;
  assign n43377 = ~n43372 & n43376 ;
  assign n43378 = ( n3385 & ~n7359 ) | ( n3385 & n11106 ) | ( ~n7359 & n11106 ) ;
  assign n43379 = n28616 & n43378 ;
  assign n43380 = ( n11279 & n12590 ) | ( n11279 & ~n30004 ) | ( n12590 & ~n30004 ) ;
  assign n43381 = n7531 ^ n7051 ^ n4654 ;
  assign n43382 = n43381 ^ n12868 ^ n8876 ;
  assign n43383 = n43382 ^ n42383 ^ n25427 ;
  assign n43384 = ( n13304 & n43380 ) | ( n13304 & ~n43383 ) | ( n43380 & ~n43383 ) ;
  assign n43385 = n35211 ^ n13755 ^ n9143 ;
  assign n43386 = n43385 ^ n33483 ^ n33092 ;
  assign n43387 = ( n2712 & n5504 ) | ( n2712 & ~n16183 ) | ( n5504 & ~n16183 ) ;
  assign n43388 = ( ~n10459 & n16109 ) | ( ~n10459 & n43387 ) | ( n16109 & n43387 ) ;
  assign n43389 = n43388 ^ n35306 ^ n17886 ;
  assign n43390 = ( n6457 & ~n15659 ) | ( n6457 & n16880 ) | ( ~n15659 & n16880 ) ;
  assign n43392 = ( n1272 & ~n9090 ) | ( n1272 & n15785 ) | ( ~n9090 & n15785 ) ;
  assign n43391 = ~n19262 & n34825 ;
  assign n43393 = n43392 ^ n43391 ^ 1'b0 ;
  assign n43394 = n43393 ^ n24082 ^ n14084 ;
  assign n43395 = ( n12864 & n17053 ) | ( n12864 & ~n43394 ) | ( n17053 & ~n43394 ) ;
  assign n43396 = n16094 ^ n10565 ^ 1'b0 ;
  assign n43397 = ~n14411 & n23545 ;
  assign n43398 = n31958 & n43397 ;
  assign n43399 = n13370 ^ n7146 ^ n2084 ;
  assign n43400 = n12366 ^ n4378 ^ 1'b0 ;
  assign n43401 = n25667 & ~n43400 ;
  assign n43402 = ~n24217 & n43401 ;
  assign n43403 = n11015 & n43402 ;
  assign n43404 = ( ~n22965 & n43399 ) | ( ~n22965 & n43403 ) | ( n43399 & n43403 ) ;
  assign n43405 = ( n8308 & n43398 ) | ( n8308 & n43404 ) | ( n43398 & n43404 ) ;
  assign n43406 = ( n11069 & n16183 ) | ( n11069 & ~n41250 ) | ( n16183 & ~n41250 ) ;
  assign n43407 = n43406 ^ n33508 ^ n26911 ;
  assign n43408 = n33536 ^ n16556 ^ n16226 ;
  assign n43409 = ( n5892 & n38310 ) | ( n5892 & n43408 ) | ( n38310 & n43408 ) ;
  assign n43410 = n13632 ^ n8645 ^ n768 ;
  assign n43411 = n41543 ^ n33275 ^ n20379 ;
  assign n43412 = ( n17840 & n43410 ) | ( n17840 & ~n43411 ) | ( n43410 & ~n43411 ) ;
  assign n43413 = ( n7661 & n19107 ) | ( n7661 & ~n25853 ) | ( n19107 & ~n25853 ) ;
  assign n43414 = n43413 ^ n24350 ^ n7812 ;
  assign n43415 = ~n22531 & n43414 ;
  assign n43416 = n43415 ^ n39570 ^ 1'b0 ;
  assign n43417 = n43416 ^ n20732 ^ n16893 ;
  assign n43418 = n30937 ^ n20928 ^ n17634 ;
  assign n43419 = ( n20307 & ~n26820 ) | ( n20307 & n43418 ) | ( ~n26820 & n43418 ) ;
  assign n43420 = ~n35791 & n43419 ;
  assign n43421 = n22171 ^ n21572 ^ n7170 ;
  assign n43422 = n43421 ^ n36102 ^ n14964 ;
  assign n43423 = ( n1175 & n8011 ) | ( n1175 & n24513 ) | ( n8011 & n24513 ) ;
  assign n43424 = n1639 | n1856 ;
  assign n43425 = n43424 ^ n12371 ^ 1'b0 ;
  assign n43426 = ( n659 & n23702 ) | ( n659 & ~n38740 ) | ( n23702 & ~n38740 ) ;
  assign n43427 = n7274 ^ n1121 ^ 1'b0 ;
  assign n43428 = ( ~n34355 & n36982 ) | ( ~n34355 & n43427 ) | ( n36982 & n43427 ) ;
  assign n43429 = ( x132 & ~n11442 ) | ( x132 & n43428 ) | ( ~n11442 & n43428 ) ;
  assign n43430 = ( ~n21312 & n43426 ) | ( ~n21312 & n43429 ) | ( n43426 & n43429 ) ;
  assign n43431 = n41997 ^ n17406 ^ n12039 ;
  assign n43432 = ( n1014 & n12472 ) | ( n1014 & n43431 ) | ( n12472 & n43431 ) ;
  assign n43433 = n43432 ^ n23080 ^ n9530 ;
  assign n43434 = ( n12011 & ~n19405 ) | ( n12011 & n41490 ) | ( ~n19405 & n41490 ) ;
  assign n43435 = n43434 ^ n15504 ^ n4321 ;
  assign n43436 = n43435 ^ n22263 ^ n6865 ;
  assign n43437 = ( n2818 & ~n9911 ) | ( n2818 & n15985 ) | ( ~n9911 & n15985 ) ;
  assign n43438 = n43437 ^ n2114 ^ n358 ;
  assign n43439 = n43438 ^ n19646 ^ n17074 ;
  assign n43440 = n9819 & ~n23196 ;
  assign n43441 = n43440 ^ n20370 ^ 1'b0 ;
  assign n43442 = ( n2199 & n16303 ) | ( n2199 & ~n43441 ) | ( n16303 & ~n43441 ) ;
  assign n43443 = n43442 ^ n39106 ^ n28615 ;
  assign n43444 = ( n6721 & ~n40212 ) | ( n6721 & n43443 ) | ( ~n40212 & n43443 ) ;
  assign n43445 = n5140 & n16416 ;
  assign n43446 = n43445 ^ n25170 ^ n402 ;
  assign n43447 = ( n13403 & n22282 ) | ( n13403 & n43446 ) | ( n22282 & n43446 ) ;
  assign n43448 = n13760 ^ n3130 ^ 1'b0 ;
  assign n43449 = n33846 & ~n43448 ;
  assign n43450 = n37313 ^ n30161 ^ n15080 ;
  assign n43451 = n11716 ^ n4174 ^ n2869 ;
  assign n43452 = ( ~n18935 & n22230 ) | ( ~n18935 & n36280 ) | ( n22230 & n36280 ) ;
  assign n43453 = ( n3730 & ~n7244 ) | ( n3730 & n8987 ) | ( ~n7244 & n8987 ) ;
  assign n43454 = n30860 ^ n16183 ^ n9119 ;
  assign n43455 = n43454 ^ n16872 ^ n3767 ;
  assign n43456 = ( ~n27445 & n43453 ) | ( ~n27445 & n43455 ) | ( n43453 & n43455 ) ;
  assign n43457 = n17633 & n26107 ;
  assign n43458 = n5599 & n43457 ;
  assign n43459 = ( ~n3675 & n8081 ) | ( ~n3675 & n43458 ) | ( n8081 & n43458 ) ;
  assign n43460 = n42357 ^ n28017 ^ n8872 ;
  assign n43463 = n26220 ^ n10148 ^ 1'b0 ;
  assign n43464 = n43463 ^ n20448 ^ n19827 ;
  assign n43461 = ( ~n547 & n1341 ) | ( ~n547 & n18310 ) | ( n1341 & n18310 ) ;
  assign n43462 = n7535 | n43461 ;
  assign n43465 = n43464 ^ n43462 ^ 1'b0 ;
  assign n43466 = n43465 ^ n2013 ^ n1004 ;
  assign n43467 = n18337 ^ n14386 ^ 1'b0 ;
  assign n43468 = ( n1774 & n6453 ) | ( n1774 & ~n13931 ) | ( n6453 & ~n13931 ) ;
  assign n43469 = ( n13939 & n21568 ) | ( n13939 & n32386 ) | ( n21568 & n32386 ) ;
  assign n43470 = n11598 ^ n1683 ^ 1'b0 ;
  assign n43471 = n25076 | n43470 ;
  assign n43472 = ( n19829 & ~n23998 ) | ( n19829 & n43471 ) | ( ~n23998 & n43471 ) ;
  assign n43473 = ( n9825 & ~n17838 ) | ( n9825 & n43472 ) | ( ~n17838 & n43472 ) ;
  assign n43474 = ( n20002 & n43469 ) | ( n20002 & ~n43473 ) | ( n43469 & ~n43473 ) ;
  assign n43475 = n43474 ^ n21958 ^ n18433 ;
  assign n43476 = ( n6517 & n43468 ) | ( n6517 & ~n43475 ) | ( n43468 & ~n43475 ) ;
  assign n43477 = ( n9448 & n18612 ) | ( n9448 & ~n39016 ) | ( n18612 & ~n39016 ) ;
  assign n43478 = ( n20549 & n27419 ) | ( n20549 & n43477 ) | ( n27419 & n43477 ) ;
  assign n43479 = n11805 ^ n4167 ^ x26 ;
  assign n43480 = n7076 & n43479 ;
  assign n43481 = ( ~n5177 & n6432 ) | ( ~n5177 & n37906 ) | ( n6432 & n37906 ) ;
  assign n43482 = n43481 ^ n37587 ^ n28830 ;
  assign n43483 = n41417 ^ n40042 ^ n27940 ;
  assign n43484 = n11588 ^ n10386 ^ 1'b0 ;
  assign n43485 = n21243 & ~n43484 ;
  assign n43486 = n12576 ^ n8505 ^ n5778 ;
  assign n43487 = n24133 | n32257 ;
  assign n43488 = ( ~n43485 & n43486 ) | ( ~n43485 & n43487 ) | ( n43486 & n43487 ) ;
  assign n43489 = n43488 ^ n31405 ^ n11029 ;
  assign n43490 = n33741 ^ n10929 ^ n6526 ;
  assign n43491 = n43490 ^ n20780 ^ n20721 ;
  assign n43492 = n43491 ^ n32887 ^ n3687 ;
  assign n43493 = n24235 | n25764 ;
  assign n43494 = n43493 ^ n25530 ^ 1'b0 ;
  assign n43495 = ~n9190 & n16881 ;
  assign n43496 = ( n12342 & n13459 ) | ( n12342 & ~n43495 ) | ( n13459 & ~n43495 ) ;
  assign n43497 = ( n18085 & n30715 ) | ( n18085 & n43496 ) | ( n30715 & n43496 ) ;
  assign n43498 = ( n20707 & n30987 ) | ( n20707 & n43497 ) | ( n30987 & n43497 ) ;
  assign n43499 = n43498 ^ n25590 ^ n25222 ;
  assign n43500 = n32745 ^ n16835 ^ n2049 ;
  assign n43501 = ~n24269 & n35307 ;
  assign n43502 = n38386 ^ n28264 ^ n2674 ;
  assign n43503 = n24062 ^ n14735 ^ n9625 ;
  assign n43504 = n43503 ^ n17599 ^ n6400 ;
  assign n43505 = n43504 ^ n35633 ^ n3758 ;
  assign n43506 = n30005 ^ n23776 ^ n15926 ;
  assign n43507 = n2035 | n23206 ;
  assign n43508 = n43507 ^ n6279 ^ 1'b0 ;
  assign n43509 = n20545 ^ n13852 ^ x195 ;
  assign n43510 = n43509 ^ n5128 ^ n2050 ;
  assign n43511 = ( ~n1989 & n17789 ) | ( ~n1989 & n25482 ) | ( n17789 & n25482 ) ;
  assign n43512 = ( ~n5047 & n31167 ) | ( ~n5047 & n43511 ) | ( n31167 & n43511 ) ;
  assign n43513 = n415 & ~n19566 ;
  assign n43514 = n43513 ^ n9969 ^ 1'b0 ;
  assign n43515 = ( n39158 & n41399 ) | ( n39158 & ~n43514 ) | ( n41399 & ~n43514 ) ;
  assign n43516 = n40273 ^ n38620 ^ n12827 ;
  assign n43517 = n13916 ^ n10233 ^ n6823 ;
  assign n43519 = n41157 ^ n28651 ^ n22645 ;
  assign n43518 = n6102 & n14483 ;
  assign n43520 = n43519 ^ n43518 ^ 1'b0 ;
  assign n43521 = n24045 ^ n16137 ^ 1'b0 ;
  assign n43522 = n14915 | n43521 ;
  assign n43523 = n6416 & ~n43522 ;
  assign n43524 = ( n6964 & n17886 ) | ( n6964 & n42976 ) | ( n17886 & n42976 ) ;
  assign n43525 = n10824 | n27234 ;
  assign n43526 = ( n17881 & n43524 ) | ( n17881 & ~n43525 ) | ( n43524 & ~n43525 ) ;
  assign n43527 = ( n16920 & n43523 ) | ( n16920 & ~n43526 ) | ( n43523 & ~n43526 ) ;
  assign n43528 = n18881 ^ n17075 ^ n1779 ;
  assign n43529 = n29800 ^ n21794 ^ n11568 ;
  assign n43530 = n27790 ^ n24604 ^ n20771 ;
  assign n43531 = ( n2575 & n9864 ) | ( n2575 & ~n10255 ) | ( n9864 & ~n10255 ) ;
  assign n43532 = ( n2068 & n3740 ) | ( n2068 & n43531 ) | ( n3740 & n43531 ) ;
  assign n43533 = n14080 & n16861 ;
  assign n43534 = ~n41290 & n43533 ;
  assign n43535 = n43534 ^ n32681 ^ 1'b0 ;
  assign n43536 = ( ~n22544 & n28222 ) | ( ~n22544 & n31236 ) | ( n28222 & n31236 ) ;
  assign n43537 = n43426 ^ n23414 ^ n12775 ;
  assign n43538 = n16602 ^ n9852 ^ n2047 ;
  assign n43539 = n5731 & ~n8653 ;
  assign n43540 = n43539 ^ n2350 ^ 1'b0 ;
  assign n43541 = ( n1949 & n3200 ) | ( n1949 & n43540 ) | ( n3200 & n43540 ) ;
  assign n43542 = n43541 ^ n16494 ^ n7221 ;
  assign n43543 = n37452 & ~n43542 ;
  assign n43544 = ( n36439 & n43538 ) | ( n36439 & ~n43543 ) | ( n43538 & ~n43543 ) ;
  assign n43545 = n32328 ^ n30600 ^ 1'b0 ;
  assign n43546 = n12360 ^ n4834 ^ n4020 ;
  assign n43547 = ( x128 & n18162 ) | ( x128 & ~n43546 ) | ( n18162 & ~n43546 ) ;
  assign n43548 = n24627 ^ n20617 ^ n9169 ;
  assign n43549 = n43548 ^ n24581 ^ n4088 ;
  assign n43550 = ( n16221 & n23665 ) | ( n16221 & n43549 ) | ( n23665 & n43549 ) ;
  assign n43551 = n32026 ^ n5766 ^ 1'b0 ;
  assign n43552 = ~n41172 & n43551 ;
  assign n43553 = ( ~n11029 & n15991 ) | ( ~n11029 & n43552 ) | ( n15991 & n43552 ) ;
  assign n43554 = ( n6022 & n8010 ) | ( n6022 & n19445 ) | ( n8010 & n19445 ) ;
  assign n43555 = ( ~n8949 & n21419 ) | ( ~n8949 & n43554 ) | ( n21419 & n43554 ) ;
  assign n43556 = ( n9510 & n39388 ) | ( n9510 & ~n43555 ) | ( n39388 & ~n43555 ) ;
  assign n43557 = ( n12342 & ~n18868 ) | ( n12342 & n38212 ) | ( ~n18868 & n38212 ) ;
  assign n43558 = n43557 ^ n28145 ^ 1'b0 ;
  assign n43559 = n43558 ^ n34703 ^ n3971 ;
  assign n43560 = n27859 & n43559 ;
  assign n43561 = n41258 ^ n21209 ^ n4663 ;
  assign n43562 = n43561 ^ n19683 ^ n19134 ;
  assign n43563 = n1613 & n7565 ;
  assign n43564 = ( n24950 & n27301 ) | ( n24950 & n43563 ) | ( n27301 & n43563 ) ;
  assign n43565 = ( n4692 & n37792 ) | ( n4692 & ~n43564 ) | ( n37792 & ~n43564 ) ;
  assign n43566 = n18507 ^ n4667 ^ n4393 ;
  assign n43567 = ( n42178 & ~n42929 ) | ( n42178 & n43566 ) | ( ~n42929 & n43566 ) ;
  assign n43568 = n6834 ^ n6630 ^ n1215 ;
  assign n43569 = ( n7476 & n9386 ) | ( n7476 & n14001 ) | ( n9386 & n14001 ) ;
  assign n43570 = ( ~n719 & n35668 ) | ( ~n719 & n43569 ) | ( n35668 & n43569 ) ;
  assign n43571 = n43570 ^ n6795 ^ 1'b0 ;
  assign n43572 = n43568 | n43571 ;
  assign n43573 = n9326 ^ n2673 ^ 1'b0 ;
  assign n43574 = n8945 & ~n43573 ;
  assign n43575 = n7184 | n22599 ;
  assign n43576 = ( ~n8651 & n10508 ) | ( ~n8651 & n11077 ) | ( n10508 & n11077 ) ;
  assign n43577 = ( ~n5829 & n11587 ) | ( ~n5829 & n23707 ) | ( n11587 & n23707 ) ;
  assign n43578 = ( n25834 & n33745 ) | ( n25834 & ~n43577 ) | ( n33745 & ~n43577 ) ;
  assign n43579 = n9939 | n15056 ;
  assign n43580 = n30511 & ~n43579 ;
  assign n43581 = n43580 ^ n39072 ^ n19462 ;
  assign n43582 = ( ~n1716 & n43578 ) | ( ~n1716 & n43581 ) | ( n43578 & n43581 ) ;
  assign n43583 = n41017 ^ n37293 ^ n5834 ;
  assign n43584 = n43583 ^ n15900 ^ n10585 ;
  assign n43585 = n23829 & ~n43584 ;
  assign n43586 = ( n11206 & ~n15807 ) | ( n11206 & n18310 ) | ( ~n15807 & n18310 ) ;
  assign n43587 = ( n2411 & ~n26340 ) | ( n2411 & n43586 ) | ( ~n26340 & n43586 ) ;
  assign n43588 = n11512 & ~n11640 ;
  assign n43589 = n43588 ^ n36533 ^ n11883 ;
  assign n43590 = ( n12120 & n13440 ) | ( n12120 & n29101 ) | ( n13440 & n29101 ) ;
  assign n43591 = n17843 & ~n42713 ;
  assign n43592 = n9147 ^ n8056 ^ n2881 ;
  assign n43593 = n32827 ^ n7706 ^ n1640 ;
  assign n43594 = n16754 ^ n2714 ^ n2437 ;
  assign n43595 = n40300 ^ n15518 ^ n4118 ;
  assign n43596 = n18749 ^ n13494 ^ n8042 ;
  assign n43597 = n43596 ^ n6745 ^ n2813 ;
  assign n43598 = n43597 ^ n40583 ^ n3458 ;
  assign n43600 = ( n5262 & ~n9569 ) | ( n5262 & n22729 ) | ( ~n9569 & n22729 ) ;
  assign n43599 = ( n18188 & n22018 ) | ( n18188 & n43561 ) | ( n22018 & n43561 ) ;
  assign n43601 = n43600 ^ n43599 ^ n23490 ;
  assign n43602 = n30194 | n32357 ;
  assign n43603 = n43602 ^ n19825 ^ 1'b0 ;
  assign n43604 = n24232 & ~n42609 ;
  assign n43605 = ~n1181 & n43604 ;
  assign n43606 = n36857 ^ n31389 ^ n26554 ;
  assign n43612 = n12579 ^ n11453 ^ n10799 ;
  assign n43611 = n10612 ^ n7790 ^ n857 ;
  assign n43607 = ( n13686 & ~n18180 ) | ( n13686 & n26430 ) | ( ~n18180 & n26430 ) ;
  assign n43608 = ( n14259 & n28473 ) | ( n14259 & ~n43607 ) | ( n28473 & ~n43607 ) ;
  assign n43609 = n43608 ^ n22903 ^ n18799 ;
  assign n43610 = n12960 & n43609 ;
  assign n43613 = n43612 ^ n43611 ^ n43610 ;
  assign n43616 = ( n3916 & n6681 ) | ( n3916 & n25343 ) | ( n6681 & n25343 ) ;
  assign n43614 = n19943 & ~n33828 ;
  assign n43615 = n43614 ^ n16915 ^ 1'b0 ;
  assign n43617 = n43616 ^ n43615 ^ n4625 ;
  assign n43618 = n38189 ^ n25798 ^ n10056 ;
  assign n43619 = ( ~n2265 & n25340 ) | ( ~n2265 & n43618 ) | ( n25340 & n43618 ) ;
  assign n43620 = n43619 ^ n16222 ^ n8990 ;
  assign n43621 = ( n2121 & ~n13670 ) | ( n2121 & n30264 ) | ( ~n13670 & n30264 ) ;
  assign n43622 = ( n2278 & n6693 ) | ( n2278 & n9810 ) | ( n6693 & n9810 ) ;
  assign n43623 = n43622 ^ n7578 ^ 1'b0 ;
  assign n43624 = ~n43621 & n43623 ;
  assign n43625 = n8453 ^ n5214 ^ 1'b0 ;
  assign n43626 = n25059 & n43625 ;
  assign n43627 = n36491 ^ n35915 ^ n18041 ;
  assign n43628 = n840 & n43627 ;
  assign n43629 = n30168 ^ n17417 ^ n9829 ;
  assign n43630 = ( ~n9651 & n24173 ) | ( ~n9651 & n30169 ) | ( n24173 & n30169 ) ;
  assign n43631 = ~n5203 & n43630 ;
  assign n43632 = n11775 ^ n1278 ^ 1'b0 ;
  assign n43633 = ( n2290 & ~n6601 ) | ( n2290 & n43632 ) | ( ~n6601 & n43632 ) ;
  assign n43634 = n37740 ^ n36690 ^ n7668 ;
  assign n43635 = n38086 ^ n25514 ^ n1633 ;
  assign n43636 = n30993 ^ n14202 ^ n12483 ;
  assign n43637 = ( n13623 & n23731 ) | ( n13623 & ~n24961 ) | ( n23731 & ~n24961 ) ;
  assign n43638 = ( ~n12151 & n43636 ) | ( ~n12151 & n43637 ) | ( n43636 & n43637 ) ;
  assign n43639 = n20860 ^ n14178 ^ n2430 ;
  assign n43640 = ( ~n9508 & n17584 ) | ( ~n9508 & n43639 ) | ( n17584 & n43639 ) ;
  assign n43641 = ~n19512 & n22564 ;
  assign n43642 = ~n39853 & n43641 ;
  assign n43643 = n43642 ^ n13353 ^ 1'b0 ;
  assign n43644 = n43643 ^ n14563 ^ n2062 ;
  assign n43645 = n38595 ^ n25294 ^ n8133 ;
  assign n43646 = x63 & ~n5714 ;
  assign n43647 = n19618 ^ n8536 ^ 1'b0 ;
  assign n43648 = ( n8442 & ~n14748 ) | ( n8442 & n43647 ) | ( ~n14748 & n43647 ) ;
  assign n43650 = n14687 ^ n8728 ^ n3199 ;
  assign n43649 = n28575 ^ n19813 ^ n6743 ;
  assign n43651 = n43650 ^ n43649 ^ n4302 ;
  assign n43652 = n8672 ^ n7690 ^ n4878 ;
  assign n43653 = ( ~n18489 & n19189 ) | ( ~n18489 & n43652 ) | ( n19189 & n43652 ) ;
  assign n43654 = n10730 & ~n26935 ;
  assign n43655 = n43654 ^ n5239 ^ 1'b0 ;
  assign n43656 = n43655 ^ n39425 ^ n13396 ;
  assign n43657 = n15953 ^ n4283 ^ n934 ;
  assign n43658 = n43657 ^ n37138 ^ n22560 ;
  assign n43659 = n16225 | n17835 ;
  assign n43660 = n17829 | n43659 ;
  assign n43661 = n43660 ^ n24251 ^ n14014 ;
  assign n43662 = n40305 ^ n4746 ^ 1'b0 ;
  assign n43663 = ( n26968 & n43661 ) | ( n26968 & n43662 ) | ( n43661 & n43662 ) ;
  assign n43664 = n30304 ^ n22717 ^ n7155 ;
  assign n43665 = n23081 ^ n6417 ^ 1'b0 ;
  assign n43666 = ( n20280 & n33280 ) | ( n20280 & ~n35454 ) | ( n33280 & ~n35454 ) ;
  assign n43667 = n43666 ^ n37985 ^ n15784 ;
  assign n43668 = n36806 ^ n25343 ^ 1'b0 ;
  assign n43669 = n43668 ^ n38748 ^ n29683 ;
  assign n43670 = ( n10320 & ~n25688 ) | ( n10320 & n43669 ) | ( ~n25688 & n43669 ) ;
  assign n43671 = n43670 ^ n35543 ^ n31059 ;
  assign n43672 = ( ~n450 & n15719 ) | ( ~n450 & n29998 ) | ( n15719 & n29998 ) ;
  assign n43673 = ( ~n499 & n1575 ) | ( ~n499 & n32839 ) | ( n1575 & n32839 ) ;
  assign n43674 = ( n13076 & n33568 ) | ( n13076 & n43673 ) | ( n33568 & n43673 ) ;
  assign n43675 = n31805 ^ n24878 ^ n15477 ;
  assign n43676 = ( n43672 & ~n43674 ) | ( n43672 & n43675 ) | ( ~n43674 & n43675 ) ;
  assign n43677 = n30190 ^ n10399 ^ n833 ;
  assign n43678 = n43677 ^ n1464 ^ 1'b0 ;
  assign n43679 = n8827 & n43678 ;
  assign n43680 = ( n3861 & n13574 ) | ( n3861 & n43679 ) | ( n13574 & n43679 ) ;
  assign n43681 = ( n4433 & ~n8045 ) | ( n4433 & n39302 ) | ( ~n8045 & n39302 ) ;
  assign n43682 = ( n7482 & n16483 ) | ( n7482 & ~n43681 ) | ( n16483 & ~n43681 ) ;
  assign n43683 = n43682 ^ n20427 ^ n3206 ;
  assign n43685 = n37426 ^ n18206 ^ n1396 ;
  assign n43686 = n43685 ^ n11990 ^ 1'b0 ;
  assign n43684 = n24146 ^ n22864 ^ n20654 ;
  assign n43687 = n43686 ^ n43684 ^ n873 ;
  assign n43688 = n43687 ^ n4556 ^ n4483 ;
  assign n43689 = ( n1762 & n1795 ) | ( n1762 & ~n43688 ) | ( n1795 & ~n43688 ) ;
  assign n43690 = ( n12400 & n38005 ) | ( n12400 & n42262 ) | ( n38005 & n42262 ) ;
  assign n43691 = ( n7658 & n11922 ) | ( n7658 & ~n43690 ) | ( n11922 & ~n43690 ) ;
  assign n43692 = ( n29199 & ~n29493 ) | ( n29199 & n43691 ) | ( ~n29493 & n43691 ) ;
  assign n43693 = n43692 ^ n5505 ^ 1'b0 ;
  assign n43694 = ( n9138 & ~n20953 ) | ( n9138 & n36402 ) | ( ~n20953 & n36402 ) ;
  assign n43695 = ( n9636 & n16282 ) | ( n9636 & n33358 ) | ( n16282 & n33358 ) ;
  assign n43696 = ~n16322 & n43695 ;
  assign n43697 = ( ~n9193 & n43694 ) | ( ~n9193 & n43696 ) | ( n43694 & n43696 ) ;
  assign n43698 = n43697 ^ n18687 ^ n1226 ;
  assign n43699 = n26993 ^ n20308 ^ n13417 ;
  assign n43700 = n6344 ^ n5626 ^ n551 ;
  assign n43701 = n43700 ^ n39860 ^ n35936 ;
  assign n43702 = n34111 ^ n9760 ^ n4691 ;
  assign n43703 = ( ~n7441 & n23718 ) | ( ~n7441 & n43702 ) | ( n23718 & n43702 ) ;
  assign n43704 = ( n2782 & ~n17699 ) | ( n2782 & n36373 ) | ( ~n17699 & n36373 ) ;
  assign n43705 = n13700 | n17935 ;
  assign n43706 = n37442 | n43705 ;
  assign n43707 = n497 & n21026 ;
  assign n43708 = n37357 & n43707 ;
  assign n43709 = n8483 | n43708 ;
  assign n43710 = n43709 ^ n13901 ^ 1'b0 ;
  assign n43711 = ( ~n727 & n6173 ) | ( ~n727 & n28887 ) | ( n6173 & n28887 ) ;
  assign n43712 = n43711 ^ n25020 ^ n11244 ;
  assign n43713 = n13136 & ~n43712 ;
  assign n43714 = n43710 & n43713 ;
  assign n43715 = n23873 ^ n4759 ^ 1'b0 ;
  assign n43716 = ( n38952 & n41215 ) | ( n38952 & ~n42244 ) | ( n41215 & ~n42244 ) ;
  assign n43717 = ( ~n19721 & n43715 ) | ( ~n19721 & n43716 ) | ( n43715 & n43716 ) ;
  assign n43718 = n39612 ^ n29558 ^ n4158 ;
  assign n43719 = n13406 | n35780 ;
  assign n43720 = n43719 ^ n4151 ^ 1'b0 ;
  assign n43721 = n43720 ^ n32601 ^ n5990 ;
  assign n43722 = n43496 | n43721 ;
  assign n43723 = n11834 ^ n9366 ^ 1'b0 ;
  assign n43724 = n43723 ^ n19262 ^ 1'b0 ;
  assign n43725 = n26390 & n43724 ;
  assign n43726 = n5228 & n43725 ;
  assign n43727 = ( n658 & n23587 ) | ( n658 & ~n43726 ) | ( n23587 & ~n43726 ) ;
  assign n43728 = n40137 ^ n30960 ^ n10286 ;
  assign n43730 = n23383 ^ n14489 ^ n13183 ;
  assign n43729 = ( n7645 & ~n26182 ) | ( n7645 & n43685 ) | ( ~n26182 & n43685 ) ;
  assign n43731 = n43730 ^ n43729 ^ 1'b0 ;
  assign n43732 = n583 & n8434 ;
  assign n43733 = n23824 | n43732 ;
  assign n43734 = ( n11742 & n15478 ) | ( n11742 & n26705 ) | ( n15478 & n26705 ) ;
  assign n43735 = n23102 & n27536 ;
  assign n43736 = ( n2280 & n11292 ) | ( n2280 & n16962 ) | ( n11292 & n16962 ) ;
  assign n43737 = ( ~n6391 & n22334 ) | ( ~n6391 & n41854 ) | ( n22334 & n41854 ) ;
  assign n43738 = ( n4457 & n11843 ) | ( n4457 & ~n43737 ) | ( n11843 & ~n43737 ) ;
  assign n43739 = ( n469 & n43736 ) | ( n469 & n43738 ) | ( n43736 & n43738 ) ;
  assign n43740 = n19319 | n43739 ;
  assign n43741 = n2463 | n43740 ;
  assign n43744 = n15330 ^ n8024 ^ n7870 ;
  assign n43745 = n43744 ^ n22109 ^ 1'b0 ;
  assign n43742 = n22512 ^ n17845 ^ n2721 ;
  assign n43743 = n43742 ^ n7250 ^ n2159 ;
  assign n43746 = n43745 ^ n43743 ^ n41876 ;
  assign n43747 = n43746 ^ n13248 ^ n2834 ;
  assign n43748 = n33564 ^ n7604 ^ 1'b0 ;
  assign n43749 = n17058 & n18633 ;
  assign n43750 = n43749 ^ n40343 ^ 1'b0 ;
  assign n43751 = n6904 & n14705 ;
  assign n43752 = n34584 & n43751 ;
  assign n43753 = ( n3504 & ~n43750 ) | ( n3504 & n43752 ) | ( ~n43750 & n43752 ) ;
  assign n43754 = n20293 ^ n4839 ^ n4309 ;
  assign n43755 = n2524 & n43754 ;
  assign n43756 = n43755 ^ n25883 ^ 1'b0 ;
  assign n43757 = ( n757 & n32386 ) | ( n757 & ~n43756 ) | ( n32386 & ~n43756 ) ;
  assign n43758 = ( ~n3577 & n16543 ) | ( ~n3577 & n21234 ) | ( n16543 & n21234 ) ;
  assign n43759 = n23321 & ~n23399 ;
  assign n43760 = n43759 ^ n35027 ^ 1'b0 ;
  assign n43761 = ( n19217 & n43758 ) | ( n19217 & n43760 ) | ( n43758 & n43760 ) ;
  assign n43763 = ( ~n607 & n11612 ) | ( ~n607 & n14161 ) | ( n11612 & n14161 ) ;
  assign n43764 = n43763 ^ n31134 ^ 1'b0 ;
  assign n43765 = n4049 & n29658 ;
  assign n43766 = n43764 & n43765 ;
  assign n43762 = ( ~n4723 & n25458 ) | ( ~n4723 & n28903 ) | ( n25458 & n28903 ) ;
  assign n43767 = n43766 ^ n43762 ^ n3477 ;
  assign n43768 = n22567 ^ n17726 ^ n6725 ;
  assign n43769 = ( n29741 & n36380 ) | ( n29741 & ~n43768 ) | ( n36380 & ~n43768 ) ;
  assign n43770 = n24951 ^ n21334 ^ 1'b0 ;
  assign n43771 = n1789 & ~n11765 ;
  assign n43772 = ~n5273 & n43771 ;
  assign n43773 = n1611 & ~n43772 ;
  assign n43774 = ~n11686 & n43773 ;
  assign n43775 = ( ~n19644 & n43770 ) | ( ~n19644 & n43774 ) | ( n43770 & n43774 ) ;
  assign n43776 = ( n7202 & ~n36537 ) | ( n7202 & n43775 ) | ( ~n36537 & n43775 ) ;
  assign n43777 = n32401 ^ n26436 ^ n5603 ;
  assign n43778 = ( ~n13214 & n16722 ) | ( ~n13214 & n43777 ) | ( n16722 & n43777 ) ;
  assign n43779 = n43778 ^ n32006 ^ n10647 ;
  assign n43780 = n24680 ^ n18471 ^ 1'b0 ;
  assign n43781 = n43780 ^ n4142 ^ 1'b0 ;
  assign n43782 = ~n19050 & n43781 ;
  assign n43783 = ( n1549 & n17540 ) | ( n1549 & n23554 ) | ( n17540 & n23554 ) ;
  assign n43784 = ( n17062 & n43343 ) | ( n17062 & ~n43783 ) | ( n43343 & ~n43783 ) ;
  assign n43785 = n12157 & ~n28638 ;
  assign n43786 = n43785 ^ n17830 ^ n11149 ;
  assign n43787 = ( n3540 & n11559 ) | ( n3540 & ~n20373 ) | ( n11559 & ~n20373 ) ;
  assign n43788 = ( n6415 & ~n24706 ) | ( n6415 & n25293 ) | ( ~n24706 & n25293 ) ;
  assign n43789 = ( n8594 & n11816 ) | ( n8594 & ~n43788 ) | ( n11816 & ~n43788 ) ;
  assign n43790 = ( n26658 & n43787 ) | ( n26658 & ~n43789 ) | ( n43787 & ~n43789 ) ;
  assign n43791 = ( n10770 & n43786 ) | ( n10770 & ~n43790 ) | ( n43786 & ~n43790 ) ;
  assign n43792 = ( ~n6418 & n30401 ) | ( ~n6418 & n34736 ) | ( n30401 & n34736 ) ;
  assign n43793 = ( n1830 & ~n25105 ) | ( n1830 & n25530 ) | ( ~n25105 & n25530 ) ;
  assign n43794 = n9404 & ~n12642 ;
  assign n43795 = n43794 ^ n40525 ^ n13337 ;
  assign n43796 = n43795 ^ n9948 ^ n4174 ;
  assign n43797 = ( ~n27566 & n38443 ) | ( ~n27566 & n42172 ) | ( n38443 & n42172 ) ;
  assign n43798 = ( n4433 & n24134 ) | ( n4433 & ~n34710 ) | ( n24134 & ~n34710 ) ;
  assign n43799 = n40255 ^ n15083 ^ n6157 ;
  assign n43800 = n19420 & ~n19956 ;
  assign n43801 = n43800 ^ n3134 ^ 1'b0 ;
  assign n43802 = ( n1546 & n17406 ) | ( n1546 & n18037 ) | ( n17406 & n18037 ) ;
  assign n43803 = ( n14903 & n43801 ) | ( n14903 & ~n43802 ) | ( n43801 & ~n43802 ) ;
  assign n43804 = n43803 ^ n39215 ^ n19727 ;
  assign n43805 = ( ~n43798 & n43799 ) | ( ~n43798 & n43804 ) | ( n43799 & n43804 ) ;
  assign n43806 = n31910 ^ n1502 ^ 1'b0 ;
  assign n43807 = n8610 | n43806 ;
  assign n43808 = n22414 & ~n32616 ;
  assign n43809 = n43808 ^ n28684 ^ 1'b0 ;
  assign n43816 = ( n852 & n21893 ) | ( n852 & n33007 ) | ( n21893 & n33007 ) ;
  assign n43817 = n43816 ^ n33368 ^ n2033 ;
  assign n43813 = ( n10432 & ~n11973 ) | ( n10432 & n13226 ) | ( ~n11973 & n13226 ) ;
  assign n43814 = n43813 ^ n39224 ^ n7997 ;
  assign n43810 = n32273 ^ n15677 ^ n5725 ;
  assign n43811 = ( n1814 & ~n15730 ) | ( n1814 & n29808 ) | ( ~n15730 & n29808 ) ;
  assign n43812 = ( n19700 & ~n43810 ) | ( n19700 & n43811 ) | ( ~n43810 & n43811 ) ;
  assign n43815 = n43814 ^ n43812 ^ 1'b0 ;
  assign n43818 = n43817 ^ n43815 ^ n39871 ;
  assign n43819 = n43818 ^ n15971 ^ n8300 ;
  assign n43820 = ( n1545 & ~n23756 ) | ( n1545 & n25362 ) | ( ~n23756 & n25362 ) ;
  assign n43821 = ( ~n14072 & n15063 ) | ( ~n14072 & n22033 ) | ( n15063 & n22033 ) ;
  assign n43822 = n43821 ^ n31855 ^ n8144 ;
  assign n43830 = n32345 ^ n4940 ^ 1'b0 ;
  assign n43828 = n17136 ^ n9647 ^ n4794 ;
  assign n43829 = n43828 ^ n19462 ^ n16157 ;
  assign n43823 = n38289 ^ n17982 ^ n7842 ;
  assign n43824 = n43823 ^ n10438 ^ n1952 ;
  assign n43825 = n15121 ^ n12420 ^ n2799 ;
  assign n43826 = n43825 ^ n10765 ^ 1'b0 ;
  assign n43827 = n43824 & n43826 ;
  assign n43831 = n43830 ^ n43829 ^ n43827 ;
  assign n43832 = ( ~n4522 & n29773 ) | ( ~n4522 & n31038 ) | ( n29773 & n31038 ) ;
  assign n43833 = n42244 ^ n38074 ^ 1'b0 ;
  assign n43836 = n6431 | n34749 ;
  assign n43837 = n7332 & ~n43836 ;
  assign n43834 = n20839 ^ n18812 ^ n5593 ;
  assign n43835 = ( n404 & n5081 ) | ( n404 & ~n43834 ) | ( n5081 & ~n43834 ) ;
  assign n43838 = n43837 ^ n43835 ^ n20381 ;
  assign n43839 = ( n8136 & ~n21595 ) | ( n8136 & n27231 ) | ( ~n21595 & n27231 ) ;
  assign n43840 = n7978 & n43839 ;
  assign n43841 = ( n13373 & ~n26457 ) | ( n13373 & n36752 ) | ( ~n26457 & n36752 ) ;
  assign n43842 = n916 | n43841 ;
  assign n43843 = n43842 ^ n35225 ^ 1'b0 ;
  assign n43844 = ( n2209 & ~n10326 ) | ( n2209 & n11045 ) | ( ~n10326 & n11045 ) ;
  assign n43845 = ( ~n707 & n10053 ) | ( ~n707 & n10539 ) | ( n10053 & n10539 ) ;
  assign n43846 = n43845 ^ n36754 ^ n16215 ;
  assign n43847 = n28442 ^ n12214 ^ n885 ;
  assign n43848 = n18626 ^ n13046 ^ 1'b0 ;
  assign n43849 = ( ~n4776 & n40147 ) | ( ~n4776 & n43848 ) | ( n40147 & n43848 ) ;
  assign n43850 = n37634 ^ n19723 ^ n1708 ;
  assign n43851 = n34874 ^ n18588 ^ n13466 ;
  assign n43852 = n43851 ^ n21954 ^ n2209 ;
  assign n43853 = ( n277 & n15965 ) | ( n277 & n43852 ) | ( n15965 & n43852 ) ;
  assign n43854 = ( n1952 & n5894 ) | ( n1952 & n33193 ) | ( n5894 & n33193 ) ;
  assign n43855 = n43854 ^ n30129 ^ n10386 ;
  assign n43856 = n43855 ^ n15171 ^ n8383 ;
  assign n43857 = ( n5226 & ~n24979 ) | ( n5226 & n43856 ) | ( ~n24979 & n43856 ) ;
  assign n43858 = ~n20767 & n43857 ;
  assign n43859 = ~n27550 & n43858 ;
  assign n43861 = ( n14286 & n21508 ) | ( n14286 & n22923 ) | ( n21508 & n22923 ) ;
  assign n43860 = ~n26098 & n42883 ;
  assign n43862 = n43861 ^ n43860 ^ n5822 ;
  assign n43863 = n18410 & n34843 ;
  assign n43864 = n22621 ^ n18239 ^ n8810 ;
  assign n43865 = ( n14480 & ~n36422 ) | ( n14480 & n43864 ) | ( ~n36422 & n43864 ) ;
  assign n43866 = n37529 ^ n22221 ^ n8444 ;
  assign n43867 = ( n15558 & ~n30758 ) | ( n15558 & n43866 ) | ( ~n30758 & n43866 ) ;
  assign n43868 = ( n3801 & n26402 ) | ( n3801 & ~n29059 ) | ( n26402 & ~n29059 ) ;
  assign n43869 = n26590 ^ n407 ^ x172 ;
  assign n43870 = n43869 ^ n37285 ^ n19418 ;
  assign n43871 = ( n8044 & n16458 ) | ( n8044 & n33522 ) | ( n16458 & n33522 ) ;
  assign n43872 = ( n14953 & n22486 ) | ( n14953 & n43871 ) | ( n22486 & n43871 ) ;
  assign n43873 = ( n2922 & n6463 ) | ( n2922 & ~n35187 ) | ( n6463 & ~n35187 ) ;
  assign n43874 = n25986 ^ n16389 ^ n7261 ;
  assign n43875 = ( ~n689 & n13812 ) | ( ~n689 & n41178 ) | ( n13812 & n41178 ) ;
  assign n43876 = ( n8498 & n14558 ) | ( n8498 & ~n40591 ) | ( n14558 & ~n40591 ) ;
  assign n43877 = ( ~n19361 & n20635 ) | ( ~n19361 & n29249 ) | ( n20635 & n29249 ) ;
  assign n43878 = ( ~n43875 & n43876 ) | ( ~n43875 & n43877 ) | ( n43876 & n43877 ) ;
  assign n43879 = n37770 ^ n19330 ^ n8273 ;
  assign n43880 = ( n667 & ~n5465 ) | ( n667 & n29295 ) | ( ~n5465 & n29295 ) ;
  assign n43881 = n43880 ^ n16086 ^ n14598 ;
  assign n43882 = n43881 ^ n21929 ^ n16104 ;
  assign n43883 = ( n4042 & ~n18082 ) | ( n4042 & n20292 ) | ( ~n18082 & n20292 ) ;
  assign n43884 = ( n3492 & ~n31415 ) | ( n3492 & n43883 ) | ( ~n31415 & n43883 ) ;
  assign n43885 = n2262 | n42496 ;
  assign n43886 = n26665 | n43885 ;
  assign n43887 = n6312 & n7908 ;
  assign n43888 = n43887 ^ n11896 ^ 1'b0 ;
  assign n43889 = n13792 | n43888 ;
  assign n43890 = n10337 & ~n13579 ;
  assign n43891 = n18770 ^ n18237 ^ n3014 ;
  assign n43892 = n43891 ^ n41209 ^ n17738 ;
  assign n43893 = n43892 ^ n14435 ^ n7225 ;
  assign n43894 = ( n5411 & ~n21666 ) | ( n5411 & n26713 ) | ( ~n21666 & n26713 ) ;
  assign n43895 = ( ~n10846 & n11981 ) | ( ~n10846 & n14418 ) | ( n11981 & n14418 ) ;
  assign n43896 = n43895 ^ n19194 ^ n9081 ;
  assign n43897 = n43896 ^ n25379 ^ x188 ;
  assign n43898 = ( n4381 & ~n27376 ) | ( n4381 & n43319 ) | ( ~n27376 & n43319 ) ;
  assign n43899 = ( n43894 & n43897 ) | ( n43894 & ~n43898 ) | ( n43897 & ~n43898 ) ;
  assign n43900 = n34331 ^ n28032 ^ n6840 ;
  assign n43901 = n43900 ^ n41976 ^ n18975 ;
  assign n43902 = n29199 ^ n8767 ^ n2389 ;
  assign n43903 = n34986 ^ n19799 ^ n8400 ;
  assign n43904 = n7819 ^ n1749 ^ 1'b0 ;
  assign n43905 = n27309 | n43904 ;
  assign n43906 = n43905 ^ n5261 ^ 1'b0 ;
  assign n43907 = n4326 & ~n43906 ;
  assign n43908 = n37359 ^ n12685 ^ n7185 ;
  assign n43909 = n38181 ^ n16861 ^ 1'b0 ;
  assign n43910 = n43908 | n43909 ;
  assign n43911 = n15391 & ~n19160 ;
  assign n43912 = n42534 ^ n11844 ^ n1939 ;
  assign n43913 = n23548 ^ n23032 ^ n22316 ;
  assign n43914 = n39636 ^ n30264 ^ n20700 ;
  assign n43915 = n36405 ^ n30951 ^ n17292 ;
  assign n43916 = ( n36968 & n38702 ) | ( n36968 & ~n40175 ) | ( n38702 & ~n40175 ) ;
  assign n43917 = n27112 ^ n12839 ^ 1'b0 ;
  assign n43918 = n33137 ^ n25892 ^ 1'b0 ;
  assign n43919 = n39468 & ~n43918 ;
  assign n43920 = ( n10445 & ~n14050 ) | ( n10445 & n37300 ) | ( ~n14050 & n37300 ) ;
  assign n43921 = ( n10830 & ~n10897 ) | ( n10830 & n15579 ) | ( ~n10897 & n15579 ) ;
  assign n43922 = ( n12153 & n13103 ) | ( n12153 & ~n43921 ) | ( n13103 & ~n43921 ) ;
  assign n43923 = n43726 ^ n40950 ^ n11679 ;
  assign n43924 = ( n1213 & n3040 ) | ( n1213 & ~n18461 ) | ( n3040 & ~n18461 ) ;
  assign n43926 = ( n1118 & ~n3422 ) | ( n1118 & n8253 ) | ( ~n3422 & n8253 ) ;
  assign n43925 = n27433 ^ n5667 ^ 1'b0 ;
  assign n43927 = n43926 ^ n43925 ^ n13865 ;
  assign n43928 = ( ~n2139 & n9267 ) | ( ~n2139 & n13351 ) | ( n9267 & n13351 ) ;
  assign n43929 = ( n9626 & n17663 ) | ( n9626 & ~n43928 ) | ( n17663 & ~n43928 ) ;
  assign n43930 = n43929 ^ n21968 ^ 1'b0 ;
  assign n43931 = n23959 ^ n11953 ^ n1013 ;
  assign n43932 = ( ~n12962 & n24114 ) | ( ~n12962 & n24944 ) | ( n24114 & n24944 ) ;
  assign n43933 = n43932 ^ n30354 ^ n3028 ;
  assign n43934 = n43933 ^ n31440 ^ n22826 ;
  assign n43936 = n3416 | n18742 ;
  assign n43937 = n43936 ^ n14868 ^ 1'b0 ;
  assign n43935 = ( n5103 & n18381 ) | ( n5103 & ~n19707 ) | ( n18381 & ~n19707 ) ;
  assign n43938 = n43937 ^ n43935 ^ n14613 ;
  assign n43939 = ( n10840 & n39706 ) | ( n10840 & n43938 ) | ( n39706 & n43938 ) ;
  assign n43940 = n38642 & n43939 ;
  assign n43941 = n40722 & n43940 ;
  assign n43942 = ( n3728 & n8505 ) | ( n3728 & ~n10281 ) | ( n8505 & ~n10281 ) ;
  assign n43943 = n43942 ^ n25668 ^ n6375 ;
  assign n43944 = ( n18311 & ~n43137 ) | ( n18311 & n43943 ) | ( ~n43137 & n43943 ) ;
  assign n43945 = n29671 ^ n27085 ^ n19009 ;
  assign n43946 = ( ~n7120 & n13731 ) | ( ~n7120 & n39907 ) | ( n13731 & n39907 ) ;
  assign n43947 = n2685 & ~n43946 ;
  assign n43948 = n20859 & n43947 ;
  assign n43949 = n18597 & n43948 ;
  assign n43950 = n20829 ^ n11792 ^ n1583 ;
  assign n43951 = n43950 ^ n35298 ^ n32754 ;
  assign n43952 = n33236 ^ n12102 ^ n2771 ;
  assign n43953 = n43952 ^ n17167 ^ n5585 ;
  assign n43954 = n39021 ^ n4474 ^ 1'b0 ;
  assign n43955 = n43954 ^ n18804 ^ n8986 ;
  assign n43956 = n12343 & ~n23282 ;
  assign n43957 = ~n26399 & n43956 ;
  assign n43958 = ( n34031 & n43955 ) | ( n34031 & ~n43957 ) | ( n43955 & ~n43957 ) ;
  assign n43959 = ( ~n13528 & n16019 ) | ( ~n13528 & n18038 ) | ( n16019 & n18038 ) ;
  assign n43960 = ( n18026 & n28072 ) | ( n18026 & ~n43959 ) | ( n28072 & ~n43959 ) ;
  assign n43961 = n43926 ^ n21957 ^ n395 ;
  assign n43962 = ( n8565 & n32283 ) | ( n8565 & ~n34182 ) | ( n32283 & ~n34182 ) ;
  assign n43963 = ( n10024 & n16783 ) | ( n10024 & n20505 ) | ( n16783 & n20505 ) ;
  assign n43964 = n43963 ^ n7822 ^ n6581 ;
  assign n43965 = n43964 ^ n20030 ^ n4757 ;
  assign n43966 = n42473 ^ n1872 ^ n1130 ;
  assign n43968 = n19610 ^ n1272 ^ 1'b0 ;
  assign n43967 = n3588 | n9915 ;
  assign n43969 = n43968 ^ n43967 ^ 1'b0 ;
  assign n43970 = ( ~n2752 & n8911 ) | ( ~n2752 & n18745 ) | ( n8911 & n18745 ) ;
  assign n43971 = n43970 ^ n34560 ^ n5477 ;
  assign n43972 = n8589 ^ n5588 ^ n5143 ;
  assign n43973 = ( ~n4341 & n20780 ) | ( ~n4341 & n43972 ) | ( n20780 & n43972 ) ;
  assign n43974 = ( ~n23612 & n37832 ) | ( ~n23612 & n41637 ) | ( n37832 & n41637 ) ;
  assign n43975 = ~n17893 & n43974 ;
  assign n43976 = ( n7984 & n8159 ) | ( n7984 & ~n8639 ) | ( n8159 & ~n8639 ) ;
  assign n43977 = ( n22011 & n26097 ) | ( n22011 & n43976 ) | ( n26097 & n43976 ) ;
  assign n43978 = n42638 ^ n41320 ^ n24180 ;
  assign n43979 = ( ~n36637 & n43977 ) | ( ~n36637 & n43978 ) | ( n43977 & n43978 ) ;
  assign n43980 = n10512 | n33332 ;
  assign n43981 = n27425 ^ n12559 ^ n6726 ;
  assign n43982 = n43981 ^ n15425 ^ n7836 ;
  assign n43983 = n43982 ^ n15729 ^ n14780 ;
  assign n43984 = n13897 ^ n11267 ^ n1683 ;
  assign n43985 = n43984 ^ n42449 ^ n21792 ;
  assign n43986 = n28445 & n38598 ;
  assign n43987 = n43986 ^ n40522 ^ n4765 ;
  assign n43988 = ~n13248 & n43987 ;
  assign n43989 = ( n1484 & n9803 ) | ( n1484 & ~n17967 ) | ( n9803 & ~n17967 ) ;
  assign n43990 = ( ~n18361 & n37683 ) | ( ~n18361 & n43989 ) | ( n37683 & n43989 ) ;
  assign n43991 = n21921 ^ n10522 ^ n2552 ;
  assign n43992 = ( n5876 & n24366 ) | ( n5876 & n43991 ) | ( n24366 & n43991 ) ;
  assign n43994 = n24256 ^ n11752 ^ n7411 ;
  assign n43993 = n35310 ^ n16528 ^ n7287 ;
  assign n43995 = n43994 ^ n43993 ^ n43790 ;
  assign n43997 = n10631 & n14481 ;
  assign n43998 = n378 & n43997 ;
  assign n43999 = n43998 ^ n15663 ^ 1'b0 ;
  assign n43996 = n43115 ^ n11655 ^ n8511 ;
  assign n44000 = n43999 ^ n43996 ^ n932 ;
  assign n44001 = ( n3982 & ~n31616 ) | ( n3982 & n39937 ) | ( ~n31616 & n39937 ) ;
  assign n44002 = ( n6681 & n38227 ) | ( n6681 & n44001 ) | ( n38227 & n44001 ) ;
  assign n44003 = n7231 & n41964 ;
  assign n44004 = n44003 ^ n40734 ^ 1'b0 ;
  assign n44005 = n44004 ^ n23851 ^ n19181 ;
  assign n44006 = ( ~n3977 & n15765 ) | ( ~n3977 & n18053 ) | ( n15765 & n18053 ) ;
  assign n44007 = n10030 & n11734 ;
  assign n44008 = ( n13216 & ~n23170 ) | ( n13216 & n41629 ) | ( ~n23170 & n41629 ) ;
  assign n44009 = n38224 ^ n34884 ^ n7782 ;
  assign n44010 = ( n10673 & n27711 ) | ( n10673 & ~n36600 ) | ( n27711 & ~n36600 ) ;
  assign n44016 = n1888 | n9156 ;
  assign n44015 = ( n8579 & n10957 ) | ( n8579 & ~n28093 ) | ( n10957 & ~n28093 ) ;
  assign n44017 = n44016 ^ n44015 ^ n2511 ;
  assign n44011 = n9889 ^ n6109 ^ 1'b0 ;
  assign n44012 = n13566 | n44011 ;
  assign n44013 = ~n1866 & n19346 ;
  assign n44014 = ( n32039 & ~n44012 ) | ( n32039 & n44013 ) | ( ~n44012 & n44013 ) ;
  assign n44018 = n44017 ^ n44014 ^ n13058 ;
  assign n44019 = n32100 ^ n30459 ^ n15628 ;
  assign n44020 = n44019 ^ n42162 ^ 1'b0 ;
  assign n44021 = n44020 ^ n22512 ^ n14572 ;
  assign n44022 = ( n22887 & ~n36495 ) | ( n22887 & n44021 ) | ( ~n36495 & n44021 ) ;
  assign n44023 = n9564 ^ n6580 ^ n2011 ;
  assign n44024 = n44023 ^ n24167 ^ n16075 ;
  assign n44025 = n14428 ^ n2781 ^ x112 ;
  assign n44026 = n30319 ^ n28814 ^ n18364 ;
  assign n44027 = ( n44024 & n44025 ) | ( n44024 & ~n44026 ) | ( n44025 & ~n44026 ) ;
  assign n44028 = ( ~n14202 & n25254 ) | ( ~n14202 & n30931 ) | ( n25254 & n30931 ) ;
  assign n44029 = ( n15728 & n41844 ) | ( n15728 & ~n44028 ) | ( n41844 & ~n44028 ) ;
  assign n44030 = n44029 ^ n27500 ^ n25496 ;
  assign n44031 = n27957 ^ n7888 ^ n5784 ;
  assign n44032 = ( n7379 & ~n12471 ) | ( n7379 & n23238 ) | ( ~n12471 & n23238 ) ;
  assign n44033 = ( ~n6966 & n44031 ) | ( ~n6966 & n44032 ) | ( n44031 & n44032 ) ;
  assign n44034 = n41746 ^ n17601 ^ 1'b0 ;
  assign n44035 = n37245 | n44034 ;
  assign n44036 = n22388 ^ n3576 ^ n3259 ;
  assign n44037 = ( n3429 & n11795 ) | ( n3429 & n44036 ) | ( n11795 & n44036 ) ;
  assign n44038 = n33991 & n44037 ;
  assign n44039 = ( ~n17539 & n25410 ) | ( ~n17539 & n27323 ) | ( n25410 & n27323 ) ;
  assign n44040 = ( n12120 & n17938 ) | ( n12120 & n34331 ) | ( n17938 & n34331 ) ;
  assign n44041 = ( n11204 & n18822 ) | ( n11204 & ~n44040 ) | ( n18822 & ~n44040 ) ;
  assign n44042 = ( ~n9196 & n31987 ) | ( ~n9196 & n44041 ) | ( n31987 & n44041 ) ;
  assign n44043 = n24698 ^ n16291 ^ n12219 ;
  assign n44044 = n44043 ^ n36779 ^ n8607 ;
  assign n44045 = ( n33114 & n34076 ) | ( n33114 & ~n44044 ) | ( n34076 & ~n44044 ) ;
  assign n44046 = n37553 ^ n36290 ^ n686 ;
  assign n44047 = ( ~n16122 & n24397 ) | ( ~n16122 & n36625 ) | ( n24397 & n36625 ) ;
  assign n44048 = ( n831 & ~n6093 ) | ( n831 & n7009 ) | ( ~n6093 & n7009 ) ;
  assign n44049 = n44048 ^ n38299 ^ n422 ;
  assign n44050 = n43436 ^ n4586 ^ 1'b0 ;
  assign n44051 = n4178 & ~n44050 ;
  assign n44052 = n29629 ^ n17762 ^ n16660 ;
  assign n44053 = ~n7967 & n20429 ;
  assign n44054 = n44053 ^ n15279 ^ 1'b0 ;
  assign n44055 = ( ~n3494 & n28890 ) | ( ~n3494 & n44054 ) | ( n28890 & n44054 ) ;
  assign n44056 = ( ~n5309 & n8646 ) | ( ~n5309 & n39550 ) | ( n8646 & n39550 ) ;
  assign n44057 = ( n5572 & n18892 ) | ( n5572 & ~n25695 ) | ( n18892 & ~n25695 ) ;
  assign n44058 = n44057 ^ n28424 ^ n14857 ;
  assign n44059 = ( ~n478 & n7355 ) | ( ~n478 & n19127 ) | ( n7355 & n19127 ) ;
  assign n44060 = ( n8881 & ~n21359 ) | ( n8881 & n44059 ) | ( ~n21359 & n44059 ) ;
  assign n44061 = n23428 ^ n7986 ^ 1'b0 ;
  assign n44062 = n44060 & n44061 ;
  assign n44063 = n41773 ^ n26235 ^ n19288 ;
  assign n44064 = ( n2608 & n6994 ) | ( n2608 & n44063 ) | ( n6994 & n44063 ) ;
  assign n44065 = n11282 | n14150 ;
  assign n44066 = ( n6126 & n11272 ) | ( n6126 & ~n21898 ) | ( n11272 & ~n21898 ) ;
  assign n44067 = ( n7999 & ~n42126 ) | ( n7999 & n44066 ) | ( ~n42126 & n44066 ) ;
  assign n44068 = n23933 ^ n17252 ^ n3604 ;
  assign n44069 = ( ~n31418 & n43093 ) | ( ~n31418 & n44068 ) | ( n43093 & n44068 ) ;
  assign n44070 = ( n1316 & n2006 ) | ( n1316 & ~n3172 ) | ( n2006 & ~n3172 ) ;
  assign n44071 = ( n27510 & n28098 ) | ( n27510 & n42310 ) | ( n28098 & n42310 ) ;
  assign n44072 = n44071 ^ n21656 ^ 1'b0 ;
  assign n44073 = ( n10169 & n38562 ) | ( n10169 & n44072 ) | ( n38562 & n44072 ) ;
  assign n44074 = n44073 ^ n34541 ^ n20480 ;
  assign n44075 = n33653 ^ n24566 ^ n14975 ;
  assign n44076 = ( ~n44070 & n44074 ) | ( ~n44070 & n44075 ) | ( n44074 & n44075 ) ;
  assign n44077 = ( n9912 & n33480 ) | ( n9912 & ~n36132 ) | ( n33480 & ~n36132 ) ;
  assign n44078 = ( n9100 & n32755 ) | ( n9100 & ~n44077 ) | ( n32755 & ~n44077 ) ;
  assign n44079 = n8726 | n37652 ;
  assign n44080 = n44079 ^ n23184 ^ 1'b0 ;
  assign n44083 = n1856 & ~n20130 ;
  assign n44081 = n43221 ^ n28183 ^ n7284 ;
  assign n44082 = n1398 & n44081 ;
  assign n44084 = n44083 ^ n44082 ^ 1'b0 ;
  assign n44085 = ( n12553 & n17819 ) | ( n12553 & ~n29681 ) | ( n17819 & ~n29681 ) ;
  assign n44086 = ( n8415 & n33199 ) | ( n8415 & n34638 ) | ( n33199 & n34638 ) ;
  assign n44087 = ( ~n10439 & n12335 ) | ( ~n10439 & n34031 ) | ( n12335 & n34031 ) ;
  assign n44088 = n32889 ^ n22966 ^ n1994 ;
  assign n44089 = n21689 ^ n16416 ^ n15834 ;
  assign n44090 = n40876 ^ n21793 ^ 1'b0 ;
  assign n44091 = n42955 & ~n44090 ;
  assign n44092 = n794 | n16927 ;
  assign n44093 = n40292 | n44092 ;
  assign n44094 = ( n7793 & ~n30494 ) | ( n7793 & n38300 ) | ( ~n30494 & n38300 ) ;
  assign n44095 = ( n23729 & ~n24429 ) | ( n23729 & n44094 ) | ( ~n24429 & n44094 ) ;
  assign n44096 = n44095 ^ n4008 ^ 1'b0 ;
  assign n44097 = ( n5957 & n7258 ) | ( n5957 & n30839 ) | ( n7258 & n30839 ) ;
  assign n44098 = n44097 ^ n13813 ^ 1'b0 ;
  assign n44099 = n44098 ^ n16880 ^ n13172 ;
  assign n44101 = n5187 ^ n4509 ^ n614 ;
  assign n44100 = ( n13229 & n27949 ) | ( n13229 & ~n43900 ) | ( n27949 & ~n43900 ) ;
  assign n44102 = n44101 ^ n44100 ^ n41621 ;
  assign n44103 = ~n9655 & n25415 ;
  assign n44104 = n44103 ^ n11068 ^ 1'b0 ;
  assign n44105 = ( n5651 & n26635 ) | ( n5651 & ~n44104 ) | ( n26635 & ~n44104 ) ;
  assign n44106 = ( n8429 & ~n38934 ) | ( n8429 & n44105 ) | ( ~n38934 & n44105 ) ;
  assign n44110 = n19336 ^ n15663 ^ 1'b0 ;
  assign n44111 = ( n27484 & n32990 ) | ( n27484 & n44110 ) | ( n32990 & n44110 ) ;
  assign n44107 = n37497 ^ n32303 ^ n18799 ;
  assign n44108 = ( n9352 & ~n16371 ) | ( n9352 & n42716 ) | ( ~n16371 & n42716 ) ;
  assign n44109 = ( n13036 & n44107 ) | ( n13036 & n44108 ) | ( n44107 & n44108 ) ;
  assign n44112 = n44111 ^ n44109 ^ n8564 ;
  assign n44113 = ( n2209 & n2596 ) | ( n2209 & n8291 ) | ( n2596 & n8291 ) ;
  assign n44114 = n16917 ^ n11708 ^ 1'b0 ;
  assign n44115 = ( ~n17366 & n44113 ) | ( ~n17366 & n44114 ) | ( n44113 & n44114 ) ;
  assign n44117 = n23563 ^ n12543 ^ 1'b0 ;
  assign n44116 = n35866 ^ n29596 ^ n22449 ;
  assign n44118 = n44117 ^ n44116 ^ n16443 ;
  assign n44119 = n12381 ^ n12274 ^ n5704 ;
  assign n44120 = n25722 ^ n9810 ^ n7547 ;
  assign n44121 = n3847 & n42373 ;
  assign n44122 = ~n44120 & n44121 ;
  assign n44123 = ( ~n2224 & n11404 ) | ( ~n2224 & n18352 ) | ( n11404 & n18352 ) ;
  assign n44124 = ( ~n7211 & n13561 ) | ( ~n7211 & n41691 ) | ( n13561 & n41691 ) ;
  assign n44125 = ( n5072 & ~n44123 ) | ( n5072 & n44124 ) | ( ~n44123 & n44124 ) ;
  assign n44126 = n35846 ^ n31294 ^ n8078 ;
  assign n44127 = ( n16927 & ~n20126 ) | ( n16927 & n36768 ) | ( ~n20126 & n36768 ) ;
  assign n44128 = n44127 ^ n15464 ^ n8573 ;
  assign n44129 = ( n1074 & ~n26277 ) | ( n1074 & n44128 ) | ( ~n26277 & n44128 ) ;
  assign n44130 = n9131 | n27104 ;
  assign n44131 = n9751 & ~n43549 ;
  assign n44132 = ~n34941 & n44131 ;
  assign n44133 = n15422 ^ n14372 ^ n7170 ;
  assign n44134 = ( n1648 & n6028 ) | ( n1648 & ~n44133 ) | ( n6028 & ~n44133 ) ;
  assign n44135 = n44134 ^ n19160 ^ x124 ;
  assign n44136 = n44135 ^ n14269 ^ n12223 ;
  assign n44137 = n40919 ^ n31680 ^ 1'b0 ;
  assign n44138 = n2296 & ~n8108 ;
  assign n44139 = ( ~n1039 & n2995 ) | ( ~n1039 & n14616 ) | ( n2995 & n14616 ) ;
  assign n44140 = n24441 ^ n20431 ^ n11140 ;
  assign n44141 = n44140 ^ n22898 ^ n1845 ;
  assign n44142 = n44141 ^ n23079 ^ n16153 ;
  assign n44143 = n10114 ^ n7059 ^ n3911 ;
  assign n44144 = ( n9918 & n13474 ) | ( n9918 & n44143 ) | ( n13474 & n44143 ) ;
  assign n44145 = n4896 ^ n4063 ^ x218 ;
  assign n44146 = n44145 ^ n36511 ^ n16832 ;
  assign n44147 = ( n10827 & n25293 ) | ( n10827 & ~n37098 ) | ( n25293 & ~n37098 ) ;
  assign n44148 = ( n17446 & n22954 ) | ( n17446 & ~n43213 ) | ( n22954 & ~n43213 ) ;
  assign n44149 = ( n19921 & ~n32281 ) | ( n19921 & n44148 ) | ( ~n32281 & n44148 ) ;
  assign n44150 = ( ~n37920 & n44147 ) | ( ~n37920 & n44149 ) | ( n44147 & n44149 ) ;
  assign n44151 = n2564 ^ n1619 ^ 1'b0 ;
  assign n44152 = n15541 & n44151 ;
  assign n44153 = ( n6437 & n16235 ) | ( n6437 & ~n37059 ) | ( n16235 & ~n37059 ) ;
  assign n44154 = ( ~n652 & n28155 ) | ( ~n652 & n44153 ) | ( n28155 & n44153 ) ;
  assign n44155 = ( n15889 & ~n37476 ) | ( n15889 & n44154 ) | ( ~n37476 & n44154 ) ;
  assign n44156 = ( n6681 & n8928 ) | ( n6681 & ~n22073 ) | ( n8928 & ~n22073 ) ;
  assign n44157 = ( n627 & n4029 ) | ( n627 & n20557 ) | ( n4029 & n20557 ) ;
  assign n44158 = ( n8041 & ~n13345 ) | ( n8041 & n44157 ) | ( ~n13345 & n44157 ) ;
  assign n44159 = n7998 | n44158 ;
  assign n44160 = n44156 & n44159 ;
  assign n44161 = ( n3576 & ~n14516 ) | ( n3576 & n35475 ) | ( ~n14516 & n35475 ) ;
  assign n44162 = ( n14200 & n17252 ) | ( n14200 & ~n27681 ) | ( n17252 & ~n27681 ) ;
  assign n44163 = ( ~n16942 & n21079 ) | ( ~n16942 & n44162 ) | ( n21079 & n44162 ) ;
  assign n44164 = n41854 ^ n34807 ^ n27494 ;
  assign n44165 = n40653 ^ n15390 ^ n1139 ;
  assign n44166 = ( n28864 & n44164 ) | ( n28864 & n44165 ) | ( n44164 & n44165 ) ;
  assign n44167 = n9879 ^ n818 ^ 1'b0 ;
  assign n44168 = n11220 ^ n8246 ^ n2452 ;
  assign n44169 = ( ~n28211 & n44167 ) | ( ~n28211 & n44168 ) | ( n44167 & n44168 ) ;
  assign n44170 = ( n4937 & n12815 ) | ( n4937 & n41049 ) | ( n12815 & n41049 ) ;
  assign n44171 = n42873 ^ n17065 ^ 1'b0 ;
  assign n44172 = n15846 | n44171 ;
  assign n44173 = ~n6037 & n17583 ;
  assign n44174 = n14419 | n44173 ;
  assign n44175 = ( n21313 & n21966 ) | ( n21313 & n44174 ) | ( n21966 & n44174 ) ;
  assign n44176 = n33548 ^ n31146 ^ n5547 ;
  assign n44177 = ( x195 & n5918 ) | ( x195 & ~n20257 ) | ( n5918 & ~n20257 ) ;
  assign n44178 = ( ~n1744 & n15738 ) | ( ~n1744 & n44177 ) | ( n15738 & n44177 ) ;
  assign n44179 = n28884 ^ n13219 ^ n6013 ;
  assign n44180 = n44179 ^ n16510 ^ 1'b0 ;
  assign n44181 = n11367 ^ n885 ^ n882 ;
  assign n44182 = ( n8758 & n24041 ) | ( n8758 & ~n36741 ) | ( n24041 & ~n36741 ) ;
  assign n44183 = ~n5586 & n13872 ;
  assign n44184 = ( n16002 & n23894 ) | ( n16002 & n44183 ) | ( n23894 & n44183 ) ;
  assign n44185 = n25810 ^ n18146 ^ n816 ;
  assign n44186 = n16522 ^ n5730 ^ n4465 ;
  assign n44187 = n44186 ^ n37496 ^ n17231 ;
  assign n44188 = ( n44184 & ~n44185 ) | ( n44184 & n44187 ) | ( ~n44185 & n44187 ) ;
  assign n44190 = n25025 ^ n18360 ^ 1'b0 ;
  assign n44189 = ( n8716 & n14127 ) | ( n8716 & n18765 ) | ( n14127 & n18765 ) ;
  assign n44191 = n44190 ^ n44189 ^ n8999 ;
  assign n44192 = n27476 ^ n18022 ^ n14467 ;
  assign n44193 = n21474 | n25379 ;
  assign n44194 = n11501 & ~n44193 ;
  assign n44195 = n44194 ^ n35744 ^ n7573 ;
  assign n44196 = ( ~n26753 & n44192 ) | ( ~n26753 & n44195 ) | ( n44192 & n44195 ) ;
  assign n44199 = n40247 ^ n37585 ^ n12358 ;
  assign n44197 = n8667 ^ n3480 ^ n1711 ;
  assign n44198 = ( ~n7073 & n38642 ) | ( ~n7073 & n44197 ) | ( n38642 & n44197 ) ;
  assign n44200 = n44199 ^ n44198 ^ n14086 ;
  assign n44201 = ( ~n20614 & n26806 ) | ( ~n20614 & n28745 ) | ( n26806 & n28745 ) ;
  assign n44202 = ( n1091 & ~n3689 ) | ( n1091 & n30660 ) | ( ~n3689 & n30660 ) ;
  assign n44203 = n44202 ^ n39729 ^ n25767 ;
  assign n44204 = n44203 ^ n17526 ^ n7405 ;
  assign n44205 = n14446 ^ n4681 ^ n1582 ;
  assign n44206 = n44205 ^ n5197 ^ n2332 ;
  assign n44207 = n18349 ^ n13015 ^ n6214 ;
  assign n44208 = n44207 ^ n36897 ^ n23173 ;
  assign n44211 = ( ~n3709 & n11460 ) | ( ~n3709 & n29978 ) | ( n11460 & n29978 ) ;
  assign n44212 = n15658 | n44211 ;
  assign n44213 = n44212 ^ n34393 ^ 1'b0 ;
  assign n44210 = ( ~n9816 & n26594 ) | ( ~n9816 & n35715 ) | ( n26594 & n35715 ) ;
  assign n44209 = n30730 ^ n22912 ^ n1187 ;
  assign n44214 = n44213 ^ n44210 ^ n44209 ;
  assign n44215 = ( ~n25378 & n27616 ) | ( ~n25378 & n29550 ) | ( n27616 & n29550 ) ;
  assign n44216 = ( n3119 & n31500 ) | ( n3119 & n39761 ) | ( n31500 & n39761 ) ;
  assign n44217 = ( ~n5688 & n24499 ) | ( ~n5688 & n44216 ) | ( n24499 & n44216 ) ;
  assign n44218 = ( n14070 & ~n21220 ) | ( n14070 & n32239 ) | ( ~n21220 & n32239 ) ;
  assign n44219 = n44218 ^ n18193 ^ n4947 ;
  assign n44222 = ( ~n14017 & n19341 ) | ( ~n14017 & n27042 ) | ( n19341 & n27042 ) ;
  assign n44220 = ( ~n19105 & n26818 ) | ( ~n19105 & n42362 ) | ( n26818 & n42362 ) ;
  assign n44221 = ( n11585 & n27833 ) | ( n11585 & n44220 ) | ( n27833 & n44220 ) ;
  assign n44223 = n44222 ^ n44221 ^ n43234 ;
  assign n44224 = ( n1289 & n1357 ) | ( n1289 & n44223 ) | ( n1357 & n44223 ) ;
  assign n44225 = n16702 ^ n16489 ^ n1477 ;
  assign n44226 = n44225 ^ n42884 ^ n19073 ;
  assign n44227 = n40252 ^ n18070 ^ 1'b0 ;
  assign n44228 = n43730 & n44227 ;
  assign n44229 = ( ~n339 & n18836 ) | ( ~n339 & n34344 ) | ( n18836 & n34344 ) ;
  assign n44230 = ( n29749 & n40952 ) | ( n29749 & ~n44229 ) | ( n40952 & ~n44229 ) ;
  assign n44231 = ~n22196 & n25709 ;
  assign n44232 = n44231 ^ n22928 ^ 1'b0 ;
  assign n44233 = ( n17799 & ~n25167 ) | ( n17799 & n44232 ) | ( ~n25167 & n44232 ) ;
  assign n44234 = ( n1928 & n2969 ) | ( n1928 & n8982 ) | ( n2969 & n8982 ) ;
  assign n44236 = n12810 ^ n2186 ^ 1'b0 ;
  assign n44235 = ( ~n6013 & n7506 ) | ( ~n6013 & n31127 ) | ( n7506 & n31127 ) ;
  assign n44237 = n44236 ^ n44235 ^ n36018 ;
  assign n44238 = n32301 ^ n24320 ^ n11992 ;
  assign n44239 = n10433 | n17121 ;
  assign n44240 = n16969 | n44239 ;
  assign n44241 = n35915 & n36227 ;
  assign n44242 = ~n44240 & n44241 ;
  assign n44243 = ( ~n3897 & n5847 ) | ( ~n3897 & n12875 ) | ( n5847 & n12875 ) ;
  assign n44244 = n33265 ^ n30040 ^ 1'b0 ;
  assign n44245 = n13387 & ~n44244 ;
  assign n44246 = n39146 ^ n11975 ^ n5932 ;
  assign n44247 = n44245 & n44246 ;
  assign n44251 = n14101 ^ n7245 ^ n5157 ;
  assign n44248 = ( n6733 & n16497 ) | ( n6733 & ~n18001 ) | ( n16497 & ~n18001 ) ;
  assign n44249 = ( ~n13347 & n38805 ) | ( ~n13347 & n44248 ) | ( n38805 & n44248 ) ;
  assign n44250 = n20591 & ~n44249 ;
  assign n44252 = n44251 ^ n44250 ^ 1'b0 ;
  assign n44253 = ( ~n22554 & n38265 ) | ( ~n22554 & n44252 ) | ( n38265 & n44252 ) ;
  assign n44254 = n44253 ^ n40162 ^ n39100 ;
  assign n44257 = n14914 ^ n7613 ^ 1'b0 ;
  assign n44258 = ~n17530 & n44257 ;
  assign n44255 = n29068 ^ n16852 ^ 1'b0 ;
  assign n44256 = n7591 & n44255 ;
  assign n44259 = n44258 ^ n44256 ^ n10642 ;
  assign n44260 = n14065 & ~n36652 ;
  assign n44261 = n44260 ^ n5520 ^ 1'b0 ;
  assign n44262 = n44261 ^ n33315 ^ n21912 ;
  assign n44263 = ( n20561 & n32546 ) | ( n20561 & n44262 ) | ( n32546 & n44262 ) ;
  assign n44264 = ( ~n8810 & n28229 ) | ( ~n8810 & n40672 ) | ( n28229 & n40672 ) ;
  assign n44265 = n38673 ^ n32865 ^ n9191 ;
  assign n44266 = n44265 ^ n43282 ^ n21481 ;
  assign n44267 = n40556 ^ n39294 ^ n1716 ;
  assign n44268 = n38476 ^ n8068 ^ n4939 ;
  assign n44269 = ( x93 & ~n704 ) | ( x93 & n5286 ) | ( ~n704 & n5286 ) ;
  assign n44270 = n19512 ^ n1347 ^ 1'b0 ;
  assign n44271 = ~n44269 & n44270 ;
  assign n44272 = ( n25114 & n44268 ) | ( n25114 & ~n44271 ) | ( n44268 & ~n44271 ) ;
  assign n44273 = n44272 ^ n11016 ^ n3528 ;
  assign n44274 = n4213 & ~n33517 ;
  assign n44275 = n2508 & ~n3184 ;
  assign n44276 = n44275 ^ n435 ^ 1'b0 ;
  assign n44277 = ~n14968 & n44276 ;
  assign n44278 = n44277 ^ n9784 ^ n7472 ;
  assign n44279 = ( ~n23206 & n27157 ) | ( ~n23206 & n44278 ) | ( n27157 & n44278 ) ;
  assign n44280 = ( n9310 & ~n25897 ) | ( n9310 & n27116 ) | ( ~n25897 & n27116 ) ;
  assign n44281 = n44280 ^ n30350 ^ n805 ;
  assign n44282 = n3235 & n15141 ;
  assign n44283 = n15819 & n44282 ;
  assign n44284 = n42442 ^ n34241 ^ 1'b0 ;
  assign n44285 = n44283 | n44284 ;
  assign n44287 = ( n4656 & n13615 ) | ( n4656 & n14237 ) | ( n13615 & n14237 ) ;
  assign n44288 = n9299 ^ n5684 ^ x7 ;
  assign n44289 = n44288 ^ n30755 ^ n3612 ;
  assign n44290 = ( n3907 & ~n44287 ) | ( n3907 & n44289 ) | ( ~n44287 & n44289 ) ;
  assign n44286 = n15961 | n37163 ;
  assign n44291 = n44290 ^ n44286 ^ 1'b0 ;
  assign n44292 = ( n25191 & n39404 ) | ( n25191 & ~n40626 ) | ( n39404 & ~n40626 ) ;
  assign n44293 = n27441 ^ n11895 ^ n11699 ;
  assign n44294 = ( n4449 & ~n25860 ) | ( n4449 & n37993 ) | ( ~n25860 & n37993 ) ;
  assign n44297 = n32799 ^ x173 ^ 1'b0 ;
  assign n44298 = n31512 & ~n44297 ;
  assign n44295 = n3634 & ~n14098 ;
  assign n44296 = n44295 ^ n30913 ^ n22649 ;
  assign n44299 = n44298 ^ n44296 ^ n7574 ;
  assign n44300 = ( n22495 & ~n23324 ) | ( n22495 & n41240 ) | ( ~n23324 & n41240 ) ;
  assign n44301 = ( n680 & ~n2035 ) | ( n680 & n5391 ) | ( ~n2035 & n5391 ) ;
  assign n44302 = n44301 ^ n30668 ^ n1230 ;
  assign n44303 = n32249 ^ n5196 ^ n2644 ;
  assign n44304 = n44303 ^ n28062 ^ n766 ;
  assign n44305 = n43451 & n44216 ;
  assign n44306 = n3277 & n44305 ;
  assign n44307 = n12038 & n25435 ;
  assign n44308 = n10087 & n44307 ;
  assign n44309 = ~n15279 & n27176 ;
  assign n44310 = n44308 & n44309 ;
  assign n44312 = ( n257 & n8097 ) | ( n257 & ~n8171 ) | ( n8097 & ~n8171 ) ;
  assign n44313 = ~n4941 & n19084 ;
  assign n44314 = ~n44312 & n44313 ;
  assign n44311 = ( n6558 & ~n18819 ) | ( n6558 & n33414 ) | ( ~n18819 & n33414 ) ;
  assign n44315 = n44314 ^ n44311 ^ n30232 ;
  assign n44316 = n26507 ^ n10155 ^ 1'b0 ;
  assign n44317 = ( ~n30074 & n31242 ) | ( ~n30074 & n44316 ) | ( n31242 & n44316 ) ;
  assign n44318 = ( n2407 & n23869 ) | ( n2407 & ~n35739 ) | ( n23869 & ~n35739 ) ;
  assign n44319 = ( ~n26401 & n39987 ) | ( ~n26401 & n44318 ) | ( n39987 & n44318 ) ;
  assign n44320 = ( n8434 & n34183 ) | ( n8434 & n35331 ) | ( n34183 & n35331 ) ;
  assign n44321 = ( n3153 & n43282 ) | ( n3153 & ~n44320 ) | ( n43282 & ~n44320 ) ;
  assign n44327 = n17714 ^ n6985 ^ n566 ;
  assign n44328 = n44327 ^ n18402 ^ 1'b0 ;
  assign n44329 = n15449 | n44328 ;
  assign n44322 = n18237 ^ n301 ^ 1'b0 ;
  assign n44323 = n44322 ^ n13242 ^ n6589 ;
  assign n44324 = n23644 ^ n18522 ^ 1'b0 ;
  assign n44325 = ( ~n24061 & n44323 ) | ( ~n24061 & n44324 ) | ( n44323 & n44324 ) ;
  assign n44326 = n44325 ^ n2585 ^ 1'b0 ;
  assign n44330 = n44329 ^ n44326 ^ n35297 ;
  assign n44331 = n39158 ^ n24416 ^ n4250 ;
  assign n44332 = n27672 ^ n14867 ^ n10883 ;
  assign n44333 = n44332 ^ n15857 ^ n8225 ;
  assign n44334 = n25389 & ~n41128 ;
  assign n44335 = n26018 & n44334 ;
  assign n44336 = n44335 ^ n5894 ^ 1'b0 ;
  assign n44337 = n14246 | n44336 ;
  assign n44340 = n15876 ^ n14602 ^ n10707 ;
  assign n44338 = n12313 ^ x244 ^ 1'b0 ;
  assign n44339 = n13978 & n44338 ;
  assign n44341 = n44340 ^ n44339 ^ n28643 ;
  assign n44342 = n32547 ^ n32215 ^ n8922 ;
  assign n44343 = ( n7939 & n10462 ) | ( n7939 & n10589 ) | ( n10462 & n10589 ) ;
  assign n44344 = n21348 ^ n13893 ^ n11381 ;
  assign n44345 = ( x78 & ~n266 ) | ( x78 & n38295 ) | ( ~n266 & n38295 ) ;
  assign n44346 = n36264 ^ n20421 ^ n2644 ;
  assign n44347 = ( n4374 & n6267 ) | ( n4374 & n44346 ) | ( n6267 & n44346 ) ;
  assign n44348 = n44347 ^ n22568 ^ n5895 ;
  assign n44349 = ( ~n7479 & n34018 ) | ( ~n7479 & n44348 ) | ( n34018 & n44348 ) ;
  assign n44350 = n22131 ^ n2602 ^ 1'b0 ;
  assign n44351 = n44350 ^ n35454 ^ n20222 ;
  assign n44352 = n42582 ^ n8846 ^ n4751 ;
  assign n44353 = ( n17535 & ~n36806 ) | ( n17535 & n44352 ) | ( ~n36806 & n44352 ) ;
  assign n44354 = ( n13894 & n19501 ) | ( n13894 & n43732 ) | ( n19501 & n43732 ) ;
  assign n44355 = ( n1929 & n14410 ) | ( n1929 & n26003 ) | ( n14410 & n26003 ) ;
  assign n44356 = n25081 & ~n44355 ;
  assign n44357 = ( n2877 & n18422 ) | ( n2877 & ~n37592 ) | ( n18422 & ~n37592 ) ;
  assign n44358 = ( ~n25059 & n26482 ) | ( ~n25059 & n44357 ) | ( n26482 & n44357 ) ;
  assign n44359 = n33038 ^ n26445 ^ 1'b0 ;
  assign n44360 = n44359 ^ n31738 ^ n24048 ;
  assign n44361 = n33771 | n36065 ;
  assign n44362 = n26636 ^ n15764 ^ n6248 ;
  assign n44363 = ( n23517 & ~n39154 ) | ( n23517 & n44362 ) | ( ~n39154 & n44362 ) ;
  assign n44364 = n10273 ^ n7814 ^ n5746 ;
  assign n44365 = n17745 ^ n8485 ^ n5267 ;
  assign n44366 = n44365 ^ n8624 ^ n4085 ;
  assign n44367 = n44366 ^ n3194 ^ 1'b0 ;
  assign n44368 = n44367 ^ n36277 ^ 1'b0 ;
  assign n44369 = n19847 & ~n44368 ;
  assign n44370 = ( n16429 & ~n44364 ) | ( n16429 & n44369 ) | ( ~n44364 & n44369 ) ;
  assign n44371 = n31190 ^ n13560 ^ 1'b0 ;
  assign n44372 = ( n25243 & n25584 ) | ( n25243 & n43082 ) | ( n25584 & n43082 ) ;
  assign n44373 = n11742 & ~n27918 ;
  assign n44375 = ( ~n5286 & n26965 ) | ( ~n5286 & n33387 ) | ( n26965 & n33387 ) ;
  assign n44376 = n44375 ^ n6494 ^ n4273 ;
  assign n44374 = n16703 ^ n9796 ^ n4123 ;
  assign n44377 = n44376 ^ n44374 ^ n31403 ;
  assign n44378 = n20892 ^ n16374 ^ n7312 ;
  assign n44379 = ( n2300 & n27342 ) | ( n2300 & ~n44378 ) | ( n27342 & ~n44378 ) ;
  assign n44380 = ( n7463 & n12594 ) | ( n7463 & n44379 ) | ( n12594 & n44379 ) ;
  assign n44381 = n26361 ^ n19673 ^ n6539 ;
  assign n44382 = ( n14334 & n21567 ) | ( n14334 & n35847 ) | ( n21567 & n35847 ) ;
  assign n44383 = n20488 ^ n8062 ^ 1'b0 ;
  assign n44384 = ~n44382 & n44383 ;
  assign n44385 = ( n15762 & n35315 ) | ( n15762 & n41408 ) | ( n35315 & n41408 ) ;
  assign n44386 = n36891 ^ n32046 ^ n30635 ;
  assign n44387 = n14303 ^ n8191 ^ n604 ;
  assign n44388 = ( n11951 & n25008 ) | ( n11951 & ~n44387 ) | ( n25008 & ~n44387 ) ;
  assign n44389 = n7918 ^ n6879 ^ 1'b0 ;
  assign n44390 = n44389 ^ n12357 ^ n1132 ;
  assign n44391 = n21162 ^ n7549 ^ n3305 ;
  assign n44392 = n44391 ^ n12708 ^ n8935 ;
  assign n44393 = ( n11573 & n36553 ) | ( n11573 & ~n38250 ) | ( n36553 & ~n38250 ) ;
  assign n44394 = n16602 ^ n16114 ^ 1'b0 ;
  assign n44395 = ~n29759 & n44394 ;
  assign n44396 = n15434 & n44395 ;
  assign n44397 = n44396 ^ n12831 ^ 1'b0 ;
  assign n44398 = n44397 ^ n31128 ^ n29176 ;
  assign n44399 = n42083 ^ n27759 ^ 1'b0 ;
  assign n44400 = n44399 ^ n23982 ^ n16607 ;
  assign n44401 = n35273 ^ n32589 ^ 1'b0 ;
  assign n44402 = n44401 ^ n21681 ^ n10416 ;
  assign n44403 = n27005 | n44402 ;
  assign n44405 = n9037 ^ n8978 ^ n8020 ;
  assign n44406 = ( n7714 & n23587 ) | ( n7714 & n44405 ) | ( n23587 & n44405 ) ;
  assign n44404 = n38556 ^ n23943 ^ n16386 ;
  assign n44407 = n44406 ^ n44404 ^ n35286 ;
  assign n44408 = ( ~x141 & n10309 ) | ( ~x141 & n16087 ) | ( n10309 & n16087 ) ;
  assign n44409 = ( ~n2877 & n8005 ) | ( ~n2877 & n15269 ) | ( n8005 & n15269 ) ;
  assign n44410 = ( n11915 & n35638 ) | ( n11915 & ~n44409 ) | ( n35638 & ~n44409 ) ;
  assign n44411 = n4430 & ~n6958 ;
  assign n44412 = n25596 ^ n5225 ^ n2891 ;
  assign n44413 = ( ~n33730 & n44411 ) | ( ~n33730 & n44412 ) | ( n44411 & n44412 ) ;
  assign n44414 = n32798 ^ n6579 ^ n4424 ;
  assign n44415 = n31137 ^ n1718 ^ 1'b0 ;
  assign n44416 = ( ~n35962 & n44414 ) | ( ~n35962 & n44415 ) | ( n44414 & n44415 ) ;
  assign n44417 = ( x114 & n19376 ) | ( x114 & ~n20291 ) | ( n19376 & ~n20291 ) ;
  assign n44418 = ( n9523 & n25482 ) | ( n9523 & ~n44417 ) | ( n25482 & ~n44417 ) ;
  assign n44419 = n44418 ^ n19142 ^ n3079 ;
  assign n44420 = n39775 ^ n26440 ^ n13435 ;
  assign n44421 = ( ~n16614 & n16812 ) | ( ~n16614 & n44420 ) | ( n16812 & n44420 ) ;
  assign n44422 = n2540 & ~n34997 ;
  assign n44423 = n20725 & n44422 ;
  assign n44424 = n43037 ^ n16832 ^ n12952 ;
  assign n44425 = ( n12098 & n12455 ) | ( n12098 & ~n12748 ) | ( n12455 & ~n12748 ) ;
  assign n44426 = n44425 ^ n25745 ^ n10511 ;
  assign n44427 = n39888 ^ n37632 ^ n30478 ;
  assign n44428 = n5350 ^ n1783 ^ n838 ;
  assign n44429 = ( ~n15142 & n27955 ) | ( ~n15142 & n44428 ) | ( n27955 & n44428 ) ;
  assign n44430 = n44429 ^ n18438 ^ 1'b0 ;
  assign n44431 = n44430 ^ n41823 ^ n24078 ;
  assign n44432 = n2654 | n25753 ;
  assign n44433 = n3138 | n44432 ;
  assign n44434 = n39767 & n44433 ;
  assign n44435 = n17548 & n22524 ;
  assign n44436 = ( n39300 & n39608 ) | ( n39300 & ~n41136 ) | ( n39608 & ~n41136 ) ;
  assign n44437 = n40995 ^ n21913 ^ n16812 ;
  assign n44438 = ( n4295 & n39066 ) | ( n4295 & n44437 ) | ( n39066 & n44437 ) ;
  assign n44443 = ( n20661 & n25465 ) | ( n20661 & n36528 ) | ( n25465 & n36528 ) ;
  assign n44439 = n17439 ^ n11322 ^ n9485 ;
  assign n44440 = n16198 ^ n6102 ^ n590 ;
  assign n44441 = ( n2171 & ~n44439 ) | ( n2171 & n44440 ) | ( ~n44439 & n44440 ) ;
  assign n44442 = n1594 & n44441 ;
  assign n44444 = n44443 ^ n44442 ^ 1'b0 ;
  assign n44445 = ~n36018 & n40658 ;
  assign n44446 = ( n1991 & ~n7080 ) | ( n1991 & n15664 ) | ( ~n7080 & n15664 ) ;
  assign n44447 = n44446 ^ n22978 ^ 1'b0 ;
  assign n44452 = n6622 & ~n27522 ;
  assign n44448 = n22564 ^ n4646 ^ n2042 ;
  assign n44449 = n17185 & ~n44448 ;
  assign n44450 = ~n15660 & n44449 ;
  assign n44451 = n44450 ^ n39983 ^ n28347 ;
  assign n44453 = n44452 ^ n44451 ^ n7339 ;
  assign n44454 = ( ~n2219 & n24475 ) | ( ~n2219 & n27638 ) | ( n24475 & n27638 ) ;
  assign n44455 = n22624 ^ n20439 ^ n9290 ;
  assign n44456 = n44455 ^ n36745 ^ n8143 ;
  assign n44457 = ~n2026 & n4856 ;
  assign n44458 = n44457 ^ n26901 ^ n16099 ;
  assign n44459 = n11231 & n44458 ;
  assign n44460 = ( n17952 & n18815 ) | ( n17952 & n19953 ) | ( n18815 & n19953 ) ;
  assign n44461 = n44460 ^ n29490 ^ n16419 ;
  assign n44462 = n33747 ^ n32687 ^ 1'b0 ;
  assign n44465 = ( n20943 & n22247 ) | ( n20943 & n37063 ) | ( n22247 & n37063 ) ;
  assign n44463 = n19121 ^ n2201 ^ 1'b0 ;
  assign n44464 = ~n1870 & n44463 ;
  assign n44466 = n44465 ^ n44464 ^ n24329 ;
  assign n44468 = ~n10554 & n20361 ;
  assign n44469 = n44468 ^ n5683 ^ 1'b0 ;
  assign n44467 = ~n15391 & n43743 ;
  assign n44470 = n44469 ^ n44467 ^ n39369 ;
  assign n44471 = n13799 ^ n11943 ^ n1565 ;
  assign n44472 = n44471 ^ n25647 ^ n1777 ;
  assign n44473 = ( n3383 & n22399 ) | ( n3383 & n44472 ) | ( n22399 & n44472 ) ;
  assign n44474 = n24355 ^ n9067 ^ n2647 ;
  assign n44475 = ( ~n10118 & n33688 ) | ( ~n10118 & n44474 ) | ( n33688 & n44474 ) ;
  assign n44476 = n42978 ^ n29347 ^ 1'b0 ;
  assign n44478 = n38213 ^ n23453 ^ n18988 ;
  assign n44479 = n44478 ^ n13771 ^ n8386 ;
  assign n44477 = n28885 ^ n10729 ^ n4484 ;
  assign n44480 = n44479 ^ n44477 ^ n19590 ;
  assign n44481 = n44480 ^ n40625 ^ n3537 ;
  assign n44483 = n35974 ^ n25292 ^ 1'b0 ;
  assign n44482 = ( n8572 & n20027 ) | ( n8572 & n24478 ) | ( n20027 & n24478 ) ;
  assign n44484 = n44483 ^ n44482 ^ n44387 ;
  assign n44485 = ( ~n38035 & n39457 ) | ( ~n38035 & n43060 ) | ( n39457 & n43060 ) ;
  assign n44486 = n44485 ^ n22074 ^ n14811 ;
  assign n44487 = n18976 ^ n18054 ^ n16473 ;
  assign n44488 = ( n16775 & n21641 ) | ( n16775 & ~n22881 ) | ( n21641 & ~n22881 ) ;
  assign n44489 = ( ~n40657 & n44487 ) | ( ~n40657 & n44488 ) | ( n44487 & n44488 ) ;
  assign n44490 = ( n9293 & ~n23645 ) | ( n9293 & n44489 ) | ( ~n23645 & n44489 ) ;
  assign n44491 = n31522 ^ n21961 ^ n18750 ;
  assign n44492 = n30570 ^ n26886 ^ 1'b0 ;
  assign n44493 = ( n7689 & n44491 ) | ( n7689 & n44492 ) | ( n44491 & n44492 ) ;
  assign n44499 = n28345 ^ n16593 ^ n11302 ;
  assign n44498 = ( n572 & n4402 ) | ( n572 & n25931 ) | ( n4402 & n25931 ) ;
  assign n44494 = ( n8833 & ~n9654 ) | ( n8833 & n26897 ) | ( ~n9654 & n26897 ) ;
  assign n44495 = ( n3877 & n12148 ) | ( n3877 & ~n44494 ) | ( n12148 & ~n44494 ) ;
  assign n44496 = n27301 ^ n26284 ^ n3118 ;
  assign n44497 = ( n17356 & ~n44495 ) | ( n17356 & n44496 ) | ( ~n44495 & n44496 ) ;
  assign n44500 = n44499 ^ n44498 ^ n44497 ;
  assign n44501 = ( n3740 & n27097 ) | ( n3740 & ~n30283 ) | ( n27097 & ~n30283 ) ;
  assign n44502 = n42153 ^ n17377 ^ n821 ;
  assign n44506 = ( n8161 & n32875 ) | ( n8161 & n32944 ) | ( n32875 & n32944 ) ;
  assign n44503 = n17572 ^ n12160 ^ n3577 ;
  assign n44504 = n27626 ^ n20092 ^ n12176 ;
  assign n44505 = ( ~n16404 & n44503 ) | ( ~n16404 & n44504 ) | ( n44503 & n44504 ) ;
  assign n44507 = n44506 ^ n44505 ^ n5980 ;
  assign n44508 = ( n44501 & n44502 ) | ( n44501 & ~n44507 ) | ( n44502 & ~n44507 ) ;
  assign n44509 = n23855 ^ n18219 ^ n3682 ;
  assign n44510 = ( n4371 & ~n10708 ) | ( n4371 & n13610 ) | ( ~n10708 & n13610 ) ;
  assign n44511 = n44510 ^ n14791 ^ n2447 ;
  assign n44512 = n24680 ^ n17359 ^ n9948 ;
  assign n44513 = ( n44509 & ~n44511 ) | ( n44509 & n44512 ) | ( ~n44511 & n44512 ) ;
  assign n44514 = ( n7237 & n23910 ) | ( n7237 & ~n31099 ) | ( n23910 & ~n31099 ) ;
  assign n44515 = ~n11790 & n32241 ;
  assign n44516 = ~n11579 & n44515 ;
  assign n44517 = n2528 & ~n40499 ;
  assign n44518 = ~n9542 & n44517 ;
  assign n44519 = n41030 ^ n36182 ^ n9594 ;
  assign n44520 = ( n4595 & n22467 ) | ( n4595 & n35685 ) | ( n22467 & n35685 ) ;
  assign n44521 = ( ~n16598 & n24019 ) | ( ~n16598 & n24296 ) | ( n24019 & n24296 ) ;
  assign n44522 = n44521 ^ n42743 ^ n9850 ;
  assign n44523 = n32438 ^ n24628 ^ n15707 ;
  assign n44524 = ( n16340 & n25806 ) | ( n16340 & ~n44523 ) | ( n25806 & ~n44523 ) ;
  assign n44527 = n302 | n2004 ;
  assign n44528 = n44527 ^ n7849 ^ 1'b0 ;
  assign n44525 = n29555 & ~n31295 ;
  assign n44526 = n44525 ^ n21458 ^ 1'b0 ;
  assign n44529 = n44528 ^ n44526 ^ n8645 ;
  assign n44530 = ( ~n4582 & n6775 ) | ( ~n4582 & n15678 ) | ( n6775 & n15678 ) ;
  assign n44531 = n19785 ^ n16821 ^ n11226 ;
  assign n44532 = ( n5352 & n12727 ) | ( n5352 & n22170 ) | ( n12727 & n22170 ) ;
  assign n44533 = ( ~n4631 & n26896 ) | ( ~n4631 & n44532 ) | ( n26896 & n44532 ) ;
  assign n44534 = ( n9391 & n16666 ) | ( n9391 & n28972 ) | ( n16666 & n28972 ) ;
  assign n44535 = ( n32004 & n44533 ) | ( n32004 & ~n44534 ) | ( n44533 & ~n44534 ) ;
  assign n44536 = ( n31000 & n44531 ) | ( n31000 & ~n44535 ) | ( n44531 & ~n44535 ) ;
  assign n44537 = n41133 ^ n14645 ^ 1'b0 ;
  assign n44538 = n6733 | n44537 ;
  assign n44539 = n17420 ^ n8099 ^ n1224 ;
  assign n44540 = n44539 ^ n39309 ^ n29799 ;
  assign n44544 = n11855 | n17304 ;
  assign n44541 = n38051 ^ n27681 ^ 1'b0 ;
  assign n44542 = n44541 ^ n41000 ^ n27008 ;
  assign n44543 = ( n3852 & ~n17837 ) | ( n3852 & n44542 ) | ( ~n17837 & n44542 ) ;
  assign n44545 = n44544 ^ n44543 ^ 1'b0 ;
  assign n44546 = n24161 ^ n21061 ^ n2592 ;
  assign n44547 = ( n12318 & ~n21129 ) | ( n12318 & n23740 ) | ( ~n21129 & n23740 ) ;
  assign n44548 = ( ~n1321 & n10640 ) | ( ~n1321 & n41387 ) | ( n10640 & n41387 ) ;
  assign n44549 = ( n32666 & n44547 ) | ( n32666 & n44548 ) | ( n44547 & n44548 ) ;
  assign n44550 = n25863 ^ n23575 ^ n18619 ;
  assign n44551 = n26963 ^ n18479 ^ n14894 ;
  assign n44552 = n41776 ^ n41714 ^ n39471 ;
  assign n44553 = ( n22447 & ~n44551 ) | ( n22447 & n44552 ) | ( ~n44551 & n44552 ) ;
  assign n44554 = n13936 ^ n1440 ^ n624 ;
  assign n44555 = n44554 ^ n43616 ^ n34119 ;
  assign n44556 = n21171 & n24795 ;
  assign n44557 = n2463 & n12630 ;
  assign n44558 = n44557 ^ n8117 ^ 1'b0 ;
  assign n44559 = ( n8248 & ~n10067 ) | ( n8248 & n18538 ) | ( ~n10067 & n18538 ) ;
  assign n44560 = ( n2534 & ~n11117 ) | ( n2534 & n44559 ) | ( ~n11117 & n44559 ) ;
  assign n44561 = n17271 ^ n9987 ^ n3816 ;
  assign n44562 = ( ~n28948 & n36703 ) | ( ~n28948 & n44561 ) | ( n36703 & n44561 ) ;
  assign n44563 = n33816 ^ n29917 ^ n18001 ;
  assign n44564 = n29331 ^ n12119 ^ n6898 ;
  assign n44565 = n25547 ^ n23964 ^ n6467 ;
  assign n44566 = n44565 ^ n14288 ^ n14177 ;
  assign n44567 = ( n25106 & n26894 ) | ( n25106 & ~n41964 ) | ( n26894 & ~n41964 ) ;
  assign n44568 = n44567 ^ n10593 ^ n3124 ;
  assign n44569 = n44568 ^ n41466 ^ n5500 ;
  assign n44570 = ( n4731 & n5822 ) | ( n4731 & ~n44569 ) | ( n5822 & ~n44569 ) ;
  assign n44571 = ( n20780 & n21993 ) | ( n20780 & ~n32099 ) | ( n21993 & ~n32099 ) ;
  assign n44572 = ( n12403 & n27501 ) | ( n12403 & ~n44571 ) | ( n27501 & ~n44571 ) ;
  assign n44573 = n44572 ^ n28651 ^ n18001 ;
  assign n44576 = n30629 ^ n21451 ^ n2327 ;
  assign n44574 = n27687 ^ n27221 ^ n12604 ;
  assign n44575 = n23515 & n44574 ;
  assign n44577 = n44576 ^ n44575 ^ 1'b0 ;
  assign n44578 = n10897 & ~n23934 ;
  assign n44579 = n44578 ^ n21786 ^ n18889 ;
  assign n44580 = n14046 ^ n13589 ^ n1683 ;
  assign n44581 = ( n14263 & n44579 ) | ( n14263 & n44580 ) | ( n44579 & n44580 ) ;
  assign n44582 = ( ~n18467 & n19103 ) | ( ~n18467 & n39487 ) | ( n19103 & n39487 ) ;
  assign n44583 = n27515 ^ n26034 ^ 1'b0 ;
  assign n44584 = ( ~n19028 & n28504 ) | ( ~n19028 & n34557 ) | ( n28504 & n34557 ) ;
  assign n44585 = ( x22 & n20398 ) | ( x22 & ~n29602 ) | ( n20398 & ~n29602 ) ;
  assign n44586 = n1717 | n36791 ;
  assign n44587 = ( n3549 & ~n6004 ) | ( n3549 & n17999 ) | ( ~n6004 & n17999 ) ;
  assign n44588 = ( n31614 & ~n44586 ) | ( n31614 & n44587 ) | ( ~n44586 & n44587 ) ;
  assign n44589 = ( n7937 & ~n44585 ) | ( n7937 & n44588 ) | ( ~n44585 & n44588 ) ;
  assign n44590 = ( n4025 & n42975 ) | ( n4025 & ~n44589 ) | ( n42975 & ~n44589 ) ;
  assign n44591 = n27454 ^ n12933 ^ n11484 ;
  assign n44592 = n20163 ^ n10224 ^ n5731 ;
  assign n44593 = n33749 ^ n8413 ^ 1'b0 ;
  assign n44594 = n2911 & n44593 ;
  assign n44595 = ( n18161 & ~n44028 ) | ( n18161 & n44594 ) | ( ~n44028 & n44594 ) ;
  assign n44599 = n37380 ^ n26999 ^ 1'b0 ;
  assign n44600 = n14654 & ~n44599 ;
  assign n44597 = n26036 ^ n7578 ^ n1766 ;
  assign n44598 = n30446 & ~n44597 ;
  assign n44596 = ( n9017 & n28118 ) | ( n9017 & n30016 ) | ( n28118 & n30016 ) ;
  assign n44601 = n44600 ^ n44598 ^ n44596 ;
  assign n44602 = n35202 ^ n31770 ^ 1'b0 ;
  assign n44603 = ~n2922 & n17317 ;
  assign n44604 = n44603 ^ n29992 ^ 1'b0 ;
  assign n44605 = ( n8696 & n44602 ) | ( n8696 & n44604 ) | ( n44602 & n44604 ) ;
  assign n44606 = n14639 & n44605 ;
  assign n44607 = n44606 ^ n3793 ^ 1'b0 ;
  assign n44608 = n9275 | n29347 ;
  assign n44609 = n44608 ^ n25530 ^ 1'b0 ;
  assign n44610 = n40939 ^ n39644 ^ n3172 ;
  assign n44611 = ( n28548 & n29637 ) | ( n28548 & n44610 ) | ( n29637 & n44610 ) ;
  assign n44612 = ( n3223 & ~n9051 ) | ( n3223 & n14617 ) | ( ~n9051 & n14617 ) ;
  assign n44613 = n9190 & ~n44612 ;
  assign n44614 = n44613 ^ n34437 ^ n7320 ;
  assign n44615 = n44614 ^ n30439 ^ n9188 ;
  assign n44620 = n39600 ^ n22096 ^ n9897 ;
  assign n44621 = ( n2627 & n20003 ) | ( n2627 & ~n44620 ) | ( n20003 & ~n44620 ) ;
  assign n44617 = n22503 ^ n10181 ^ n8296 ;
  assign n44618 = n7476 & n44617 ;
  assign n44619 = n8997 & n44618 ;
  assign n44616 = n18695 ^ n9088 ^ 1'b0 ;
  assign n44622 = n44621 ^ n44619 ^ n44616 ;
  assign n44623 = n41765 ^ n30941 ^ n4913 ;
  assign n44624 = n21035 ^ n20512 ^ n16189 ;
  assign n44625 = ( n4137 & ~n9675 ) | ( n4137 & n10884 ) | ( ~n9675 & n10884 ) ;
  assign n44626 = ( n32310 & n44624 ) | ( n32310 & ~n44625 ) | ( n44624 & ~n44625 ) ;
  assign n44627 = ( n9222 & n9775 ) | ( n9222 & n16105 ) | ( n9775 & n16105 ) ;
  assign n44628 = n40534 ^ n30171 ^ n29349 ;
  assign n44629 = ( n13987 & n16068 ) | ( n13987 & ~n44628 ) | ( n16068 & ~n44628 ) ;
  assign n44630 = ( n19265 & n30096 ) | ( n19265 & ~n30375 ) | ( n30096 & ~n30375 ) ;
  assign n44631 = n30692 ^ n27419 ^ 1'b0 ;
  assign n44632 = ( n8789 & n31882 ) | ( n8789 & n44631 ) | ( n31882 & n44631 ) ;
  assign n44633 = n35410 ^ n10056 ^ n667 ;
  assign n44634 = n44633 ^ n15728 ^ n8743 ;
  assign n44635 = ~n11129 & n35201 ;
  assign n44636 = ~n11063 & n44635 ;
  assign n44637 = n44636 ^ n22680 ^ n17940 ;
  assign n44638 = ( n3624 & n17373 ) | ( n3624 & n44637 ) | ( n17373 & n44637 ) ;
  assign n44642 = ~n6279 & n33235 ;
  assign n44640 = n11945 ^ n1987 ^ 1'b0 ;
  assign n44639 = n25536 ^ n23963 ^ n13437 ;
  assign n44641 = n44640 ^ n44639 ^ n14074 ;
  assign n44643 = n44642 ^ n44641 ^ n36321 ;
  assign n44644 = n22780 & n34882 ;
  assign n44645 = ( ~n1354 & n2058 ) | ( ~n1354 & n38208 ) | ( n2058 & n38208 ) ;
  assign n44646 = n32343 ^ n7137 ^ n2254 ;
  assign n44647 = n31014 ^ n9415 ^ 1'b0 ;
  assign n44648 = n18405 | n44647 ;
  assign n44649 = ( n14706 & n19440 ) | ( n14706 & ~n19804 ) | ( n19440 & ~n19804 ) ;
  assign n44650 = ( n677 & n5499 ) | ( n677 & ~n44649 ) | ( n5499 & ~n44649 ) ;
  assign n44651 = ( ~n21198 & n44648 ) | ( ~n21198 & n44650 ) | ( n44648 & n44650 ) ;
  assign n44652 = n15180 ^ n11479 ^ 1'b0 ;
  assign n44653 = n44652 ^ n33424 ^ n18884 ;
  assign n44654 = ( n8935 & ~n32369 ) | ( n8935 & n36712 ) | ( ~n32369 & n36712 ) ;
  assign n44655 = n44654 ^ n42844 ^ n33892 ;
  assign n44656 = n42416 ^ n21801 ^ n18777 ;
  assign n44657 = ( n1958 & n3284 ) | ( n1958 & n44656 ) | ( n3284 & n44656 ) ;
  assign n44658 = ( n20097 & ~n41009 ) | ( n20097 & n44657 ) | ( ~n41009 & n44657 ) ;
  assign n44659 = ( ~n584 & n7167 ) | ( ~n584 & n12456 ) | ( n7167 & n12456 ) ;
  assign n44660 = n44659 ^ n14026 ^ n3479 ;
  assign n44661 = n43146 ^ n18966 ^ n14330 ;
  assign n44662 = ( n13914 & n44660 ) | ( n13914 & n44661 ) | ( n44660 & n44661 ) ;
  assign n44663 = n9107 & n12167 ;
  assign n44664 = n1287 | n32932 ;
  assign n44667 = ( n5899 & n9269 ) | ( n5899 & ~n12716 ) | ( n9269 & ~n12716 ) ;
  assign n44665 = n28432 ^ n26411 ^ n8914 ;
  assign n44666 = ( ~n12285 & n14177 ) | ( ~n12285 & n44665 ) | ( n14177 & n44665 ) ;
  assign n44668 = n44667 ^ n44666 ^ n3753 ;
  assign n44669 = n8598 ^ n4784 ^ n4360 ;
  assign n44670 = ( n3976 & n13887 ) | ( n3976 & ~n44669 ) | ( n13887 & ~n44669 ) ;
  assign n44671 = ( n9380 & ~n12869 ) | ( n9380 & n44670 ) | ( ~n12869 & n44670 ) ;
  assign n44672 = ( ~n5094 & n39737 ) | ( ~n5094 & n44671 ) | ( n39737 & n44671 ) ;
  assign n44673 = n41565 ^ n12022 ^ n4935 ;
  assign n44674 = n40625 | n41444 ;
  assign n44675 = ~n8997 & n12320 ;
  assign n44676 = n16640 ^ n5993 ^ n3013 ;
  assign n44677 = n44676 ^ n13438 ^ 1'b0 ;
  assign n44678 = ~n9081 & n27017 ;
  assign n44679 = n2642 & n44678 ;
  assign n44680 = n44679 ^ n20309 ^ n17378 ;
  assign n44681 = n19659 & n24848 ;
  assign n44682 = ~n7986 & n31670 ;
  assign n44683 = n15032 & ~n27300 ;
  assign n44684 = n39098 ^ n18344 ^ n14420 ;
  assign n44685 = n44684 ^ n26550 ^ n2292 ;
  assign n44686 = ( n15247 & ~n38789 ) | ( n15247 & n44685 ) | ( ~n38789 & n44685 ) ;
  assign n44687 = ( n11439 & n44683 ) | ( n11439 & n44686 ) | ( n44683 & n44686 ) ;
  assign n44688 = n40038 & ~n44687 ;
  assign n44689 = n44682 & n44688 ;
  assign n44690 = n22868 ^ n18509 ^ n505 ;
  assign n44691 = n37035 ^ n22168 ^ n17272 ;
  assign n44692 = ( n12876 & ~n13774 ) | ( n12876 & n44691 ) | ( ~n13774 & n44691 ) ;
  assign n44693 = n1125 | n19315 ;
  assign n44694 = n44693 ^ n26098 ^ 1'b0 ;
  assign n44695 = ( n10972 & n44692 ) | ( n10972 & ~n44694 ) | ( n44692 & ~n44694 ) ;
  assign n44696 = n42840 ^ n12436 ^ 1'b0 ;
  assign n44698 = n10277 & n18165 ;
  assign n44697 = n39680 ^ n25669 ^ n9287 ;
  assign n44699 = n44698 ^ n44697 ^ 1'b0 ;
  assign n44700 = n44696 | n44699 ;
  assign n44701 = n17075 ^ n6294 ^ n2770 ;
  assign n44702 = n34917 ^ n17456 ^ n1827 ;
  assign n44703 = ( n5239 & n15961 ) | ( n5239 & n18732 ) | ( n15961 & n18732 ) ;
  assign n44704 = n40261 ^ n38667 ^ n696 ;
  assign n44705 = ( n9373 & ~n13761 ) | ( n9373 & n15301 ) | ( ~n13761 & n15301 ) ;
  assign n44706 = n44705 ^ n36350 ^ n5521 ;
  assign n44707 = n44706 ^ n32969 ^ n9025 ;
  assign n44708 = n44707 ^ n35778 ^ n17932 ;
  assign n44709 = n44708 ^ n37868 ^ n4698 ;
  assign n44710 = n44709 ^ n28052 ^ n27365 ;
  assign n44711 = ~n25750 & n26016 ;
  assign n44712 = n9704 & n22295 ;
  assign n44713 = n44711 & n44712 ;
  assign n44714 = ( ~n2202 & n2399 ) | ( ~n2202 & n9881 ) | ( n2399 & n9881 ) ;
  assign n44715 = n36019 & ~n44714 ;
  assign n44719 = ~n25154 & n41583 ;
  assign n44717 = ~n5243 & n16032 ;
  assign n44718 = n44717 ^ n10193 ^ 1'b0 ;
  assign n44716 = ( n32531 & n37402 ) | ( n32531 & ~n38217 ) | ( n37402 & ~n38217 ) ;
  assign n44720 = n44719 ^ n44718 ^ n44716 ;
  assign n44721 = ( n3471 & n7140 ) | ( n3471 & n24821 ) | ( n7140 & n24821 ) ;
  assign n44722 = ( n9988 & n23865 ) | ( n9988 & ~n44721 ) | ( n23865 & ~n44721 ) ;
  assign n44723 = n28880 ^ n15089 ^ 1'b0 ;
  assign n44724 = n21762 ^ n2781 ^ n837 ;
  assign n44725 = n44724 ^ n23274 ^ n13805 ;
  assign n44726 = n44725 ^ n41778 ^ n5151 ;
  assign n44727 = n44726 ^ n30052 ^ n13460 ;
  assign n44728 = n36046 ^ n23326 ^ n19505 ;
  assign n44729 = n21972 | n44728 ;
  assign n44733 = ~n12690 & n24253 ;
  assign n44734 = n44733 ^ n41338 ^ 1'b0 ;
  assign n44732 = n37731 ^ n9446 ^ 1'b0 ;
  assign n44730 = n15463 ^ n11502 ^ n1467 ;
  assign n44731 = ~n9416 & n44730 ;
  assign n44735 = n44734 ^ n44732 ^ n44731 ;
  assign n44736 = n36618 & n44016 ;
  assign n44737 = ( n4336 & n14452 ) | ( n4336 & n43657 ) | ( n14452 & n43657 ) ;
  assign n44738 = n44737 ^ n20380 ^ n18790 ;
  assign n44739 = n7820 | n44738 ;
  assign n44740 = n22361 & ~n44739 ;
  assign n44741 = n11555 | n44740 ;
  assign n44742 = n40074 ^ n25328 ^ n12814 ;
  assign n44743 = n44742 ^ n42635 ^ n25387 ;
  assign n44744 = ( n10566 & n17181 ) | ( n10566 & n39013 ) | ( n17181 & n39013 ) ;
  assign n44745 = n5465 & n24495 ;
  assign n44746 = ~n22979 & n44745 ;
  assign n44747 = ( ~n7814 & n10840 ) | ( ~n7814 & n44746 ) | ( n10840 & n44746 ) ;
  assign n44748 = n15879 ^ n11981 ^ n8109 ;
  assign n44749 = n44748 ^ n16045 ^ n14381 ;
  assign n44750 = n44749 ^ n37308 ^ n22007 ;
  assign n44751 = ( ~n11559 & n24854 ) | ( ~n11559 & n41654 ) | ( n24854 & n41654 ) ;
  assign n44752 = n44751 ^ n24827 ^ n20673 ;
  assign n44753 = n21329 ^ n5621 ^ n2628 ;
  assign n44754 = n44753 ^ n17740 ^ n15747 ;
  assign n44755 = ( ~n2727 & n9299 ) | ( ~n2727 & n32125 ) | ( n9299 & n32125 ) ;
  assign n44756 = n11558 | n44659 ;
  assign n44757 = n44756 ^ n8166 ^ 1'b0 ;
  assign n44758 = ( n8699 & n29418 ) | ( n8699 & n44757 ) | ( n29418 & n44757 ) ;
  assign n44759 = ( n13179 & ~n44755 ) | ( n13179 & n44758 ) | ( ~n44755 & n44758 ) ;
  assign n44760 = n44759 ^ n27263 ^ n8231 ;
  assign n44761 = n38811 ^ n37924 ^ 1'b0 ;
  assign n44762 = n34894 ^ n21249 ^ n6664 ;
  assign n44763 = ~n814 & n20851 ;
  assign n44764 = n44763 ^ n1198 ^ 1'b0 ;
  assign n44765 = n44764 ^ n26751 ^ n9024 ;
  assign n44766 = ( ~n23179 & n44762 ) | ( ~n23179 & n44765 ) | ( n44762 & n44765 ) ;
  assign n44767 = n44766 ^ n32819 ^ n15416 ;
  assign n44768 = n32215 ^ n2362 ^ n627 ;
  assign n44769 = ( ~n11696 & n27267 ) | ( ~n11696 & n44768 ) | ( n27267 & n44768 ) ;
  assign n44770 = ( ~n7107 & n9424 ) | ( ~n7107 & n15260 ) | ( n9424 & n15260 ) ;
  assign n44771 = ( n3207 & n7543 ) | ( n3207 & n7937 ) | ( n7543 & n7937 ) ;
  assign n44772 = n44771 ^ n18939 ^ n2478 ;
  assign n44777 = n1432 ^ n706 ^ n396 ;
  assign n44776 = n40820 ^ n23893 ^ n22708 ;
  assign n44773 = n30103 ^ n15632 ^ n13206 ;
  assign n44774 = n36475 ^ n15971 ^ n3081 ;
  assign n44775 = ( n11990 & n44773 ) | ( n11990 & ~n44774 ) | ( n44773 & ~n44774 ) ;
  assign n44778 = n44777 ^ n44776 ^ n44775 ;
  assign n44779 = n44778 ^ n35244 ^ n3509 ;
  assign n44780 = n44779 ^ n2513 ^ 1'b0 ;
  assign n44781 = ~n44772 & n44780 ;
  assign n44782 = n42585 ^ n34812 ^ n16644 ;
  assign n44783 = n16180 ^ n12398 ^ n11200 ;
  assign n44784 = n24295 ^ n9226 ^ n7089 ;
  assign n44785 = n17207 & ~n44784 ;
  assign n44786 = ~n4167 & n44785 ;
  assign n44787 = ( ~n12777 & n20375 ) | ( ~n12777 & n44786 ) | ( n20375 & n44786 ) ;
  assign n44788 = n44787 ^ n7146 ^ n4213 ;
  assign n44789 = n36918 ^ n20563 ^ n17967 ;
  assign n44790 = n9495 | n11664 ;
  assign n44791 = n44790 ^ n20576 ^ 1'b0 ;
  assign n44792 = ( n4903 & n38958 ) | ( n4903 & n44791 ) | ( n38958 & n44791 ) ;
  assign n44793 = ( n25729 & n28013 ) | ( n25729 & ~n29649 ) | ( n28013 & ~n29649 ) ;
  assign n44794 = ( n17735 & n24694 ) | ( n17735 & ~n44793 ) | ( n24694 & ~n44793 ) ;
  assign n44795 = ( n1941 & n6741 ) | ( n1941 & n35605 ) | ( n6741 & n35605 ) ;
  assign n44796 = n44795 ^ n26810 ^ n8370 ;
  assign n44797 = ( ~n11007 & n26011 ) | ( ~n11007 & n44796 ) | ( n26011 & n44796 ) ;
  assign n44798 = n1470 | n4008 ;
  assign n44799 = n44798 ^ n29554 ^ 1'b0 ;
  assign n44800 = ( ~n12446 & n14268 ) | ( ~n12446 & n38708 ) | ( n14268 & n38708 ) ;
  assign n44801 = n44800 ^ n24783 ^ n5063 ;
  assign n44802 = n5844 ^ n2742 ^ 1'b0 ;
  assign n44803 = n44801 | n44802 ;
  assign n44804 = n33871 ^ n11528 ^ n6471 ;
  assign n44805 = n44804 ^ n15188 ^ 1'b0 ;
  assign n44806 = ( n15878 & n18430 ) | ( n15878 & n30169 ) | ( n18430 & n30169 ) ;
  assign n44807 = n25587 ^ n24939 ^ n21144 ;
  assign n44808 = ( n2709 & n8872 ) | ( n2709 & n44807 ) | ( n8872 & n44807 ) ;
  assign n44810 = n41836 ^ n36158 ^ n11530 ;
  assign n44809 = n14254 ^ n5500 ^ n736 ;
  assign n44811 = n44810 ^ n44809 ^ n10567 ;
  assign n44812 = ( n10458 & n26618 ) | ( n10458 & n31349 ) | ( n26618 & n31349 ) ;
  assign n44813 = n11941 ^ n7927 ^ n4865 ;
  assign n44814 = ( n17861 & n18140 ) | ( n17861 & n44813 ) | ( n18140 & n44813 ) ;
  assign n44815 = ( ~n33753 & n36327 ) | ( ~n33753 & n44814 ) | ( n36327 & n44814 ) ;
  assign n44816 = ( n9967 & ~n10255 ) | ( n9967 & n19728 ) | ( ~n10255 & n19728 ) ;
  assign n44817 = n15746 & ~n44816 ;
  assign n44818 = ~n36152 & n44817 ;
  assign n44822 = ( n2627 & n18791 ) | ( n2627 & n40513 ) | ( n18791 & n40513 ) ;
  assign n44819 = n13433 ^ x78 ^ 1'b0 ;
  assign n44820 = ( n8429 & n14616 ) | ( n8429 & n21655 ) | ( n14616 & n21655 ) ;
  assign n44821 = ( n29313 & n44819 ) | ( n29313 & n44820 ) | ( n44819 & n44820 ) ;
  assign n44823 = n44822 ^ n44821 ^ n14321 ;
  assign n44824 = ( n1482 & n6925 ) | ( n1482 & n11152 ) | ( n6925 & n11152 ) ;
  assign n44825 = n7635 ^ n3430 ^ 1'b0 ;
  assign n44826 = n5515 & ~n44825 ;
  assign n44827 = n44824 & n44826 ;
  assign n44828 = ( n25647 & n42692 ) | ( n25647 & ~n44827 ) | ( n42692 & ~n44827 ) ;
  assign n44829 = ( n9763 & ~n29429 ) | ( n9763 & n29799 ) | ( ~n29429 & n29799 ) ;
  assign n44830 = ( n5319 & ~n29861 ) | ( n5319 & n40512 ) | ( ~n29861 & n40512 ) ;
  assign n44831 = n2532 & ~n3650 ;
  assign n44832 = n44831 ^ n43026 ^ 1'b0 ;
  assign n44833 = n44832 ^ n7707 ^ 1'b0 ;
  assign n44834 = ~n18722 & n44833 ;
  assign n44835 = ( n42754 & n44830 ) | ( n42754 & ~n44834 ) | ( n44830 & ~n44834 ) ;
  assign n44836 = n33484 ^ n18810 ^ n2551 ;
  assign n44837 = n15887 | n26292 ;
  assign n44838 = n1751 | n44837 ;
  assign n44839 = ( n6172 & n39510 ) | ( n6172 & ~n44838 ) | ( n39510 & ~n44838 ) ;
  assign n44840 = ( ~n14256 & n44836 ) | ( ~n14256 & n44839 ) | ( n44836 & n44839 ) ;
  assign n44841 = n33260 ^ n31338 ^ n22528 ;
  assign n44842 = ( ~n682 & n1477 ) | ( ~n682 & n3685 ) | ( n1477 & n3685 ) ;
  assign n44843 = ( n8037 & n28348 ) | ( n8037 & n44842 ) | ( n28348 & n44842 ) ;
  assign n44844 = n23089 ^ n11446 ^ n2058 ;
  assign n44845 = n14867 & ~n32475 ;
  assign n44846 = n44845 ^ n1280 ^ 1'b0 ;
  assign n44847 = ( n4834 & n44844 ) | ( n4834 & ~n44846 ) | ( n44844 & ~n44846 ) ;
  assign n44848 = ( n923 & ~n6765 ) | ( n923 & n11152 ) | ( ~n6765 & n11152 ) ;
  assign n44849 = n44848 ^ n26997 ^ n6056 ;
  assign n44850 = ( ~n2114 & n30555 ) | ( ~n2114 & n41833 ) | ( n30555 & n41833 ) ;
  assign n44851 = n400 & ~n12479 ;
  assign n44852 = n9459 & n44851 ;
  assign n44853 = ( n6667 & n11523 ) | ( n6667 & ~n15427 ) | ( n11523 & ~n15427 ) ;
  assign n44854 = n44853 ^ n19196 ^ n17768 ;
  assign n44855 = n44854 ^ n31551 ^ n14612 ;
  assign n44856 = n13986 & n44855 ;
  assign n44857 = n17417 ^ n5101 ^ n2651 ;
  assign n44859 = ( ~n1015 & n1881 ) | ( ~n1015 & n29377 ) | ( n1881 & n29377 ) ;
  assign n44858 = ~n4142 & n19140 ;
  assign n44860 = n44859 ^ n44858 ^ 1'b0 ;
  assign n44861 = ( n38043 & ~n44857 ) | ( n38043 & n44860 ) | ( ~n44857 & n44860 ) ;
  assign n44862 = n44861 ^ n28444 ^ x15 ;
  assign n44863 = ( n2800 & n11125 ) | ( n2800 & ~n12594 ) | ( n11125 & ~n12594 ) ;
  assign n44864 = ( n14060 & ~n15269 ) | ( n14060 & n16562 ) | ( ~n15269 & n16562 ) ;
  assign n44865 = ( n25842 & ~n44863 ) | ( n25842 & n44864 ) | ( ~n44863 & n44864 ) ;
  assign n44866 = n11437 | n12004 ;
  assign n44867 = n9318 & ~n44866 ;
  assign n44868 = n44867 ^ n19871 ^ n19812 ;
  assign n44869 = ~n19337 & n44868 ;
  assign n44870 = n18334 & n44869 ;
  assign n44871 = ( n3992 & n4573 ) | ( n3992 & ~n44870 ) | ( n4573 & ~n44870 ) ;
  assign n44872 = ( n11066 & ~n30240 ) | ( n11066 & n44871 ) | ( ~n30240 & n44871 ) ;
  assign n44873 = n35784 ^ n35382 ^ n17161 ;
  assign n44874 = n44873 ^ n12538 ^ 1'b0 ;
  assign n44875 = n6232 & ~n33606 ;
  assign n44876 = n44875 ^ n24168 ^ 1'b0 ;
  assign n44877 = ( n1450 & n15413 ) | ( n1450 & ~n32988 ) | ( n15413 & ~n32988 ) ;
  assign n44878 = ( n1261 & n38427 ) | ( n1261 & ~n44877 ) | ( n38427 & ~n44877 ) ;
  assign n44879 = n38268 ^ n18612 ^ n17591 ;
  assign n44880 = ( n15328 & ~n25981 ) | ( n15328 & n31879 ) | ( ~n25981 & n31879 ) ;
  assign n44883 = n38048 ^ n29017 ^ 1'b0 ;
  assign n44881 = n2555 ^ n1460 ^ 1'b0 ;
  assign n44882 = n44881 ^ n33389 ^ n11845 ;
  assign n44884 = n44883 ^ n44882 ^ n23860 ;
  assign n44885 = n42560 ^ n28892 ^ 1'b0 ;
  assign n44886 = n31526 ^ n28160 ^ n5048 ;
  assign n44887 = ( ~n1317 & n44885 ) | ( ~n1317 & n44886 ) | ( n44885 & n44886 ) ;
  assign n44892 = ( n6840 & ~n16918 ) | ( n6840 & n37399 ) | ( ~n16918 & n37399 ) ;
  assign n44888 = x220 & ~n1645 ;
  assign n44889 = ~n1518 & n44888 ;
  assign n44890 = ( ~n13436 & n22028 ) | ( ~n13436 & n44889 ) | ( n22028 & n44889 ) ;
  assign n44891 = n44890 ^ n21780 ^ n4297 ;
  assign n44893 = n44892 ^ n44891 ^ n15117 ;
  assign n44894 = ( ~n9577 & n42795 ) | ( ~n9577 & n44893 ) | ( n42795 & n44893 ) ;
  assign n44895 = ( n6023 & ~n8842 ) | ( n6023 & n20550 ) | ( ~n8842 & n20550 ) ;
  assign n44896 = ( n369 & n34386 ) | ( n369 & ~n44895 ) | ( n34386 & ~n44895 ) ;
  assign n44897 = n12612 | n44896 ;
  assign n44898 = n4980 & ~n44897 ;
  assign n44900 = n20240 ^ n5234 ^ 1'b0 ;
  assign n44901 = n12974 ^ n11678 ^ 1'b0 ;
  assign n44902 = ( n17911 & ~n44900 ) | ( n17911 & n44901 ) | ( ~n44900 & n44901 ) ;
  assign n44899 = ( ~n2174 & n19490 ) | ( ~n2174 & n29701 ) | ( n19490 & n29701 ) ;
  assign n44903 = n44902 ^ n44899 ^ n40227 ;
  assign n44904 = n27672 ^ n24701 ^ n16570 ;
  assign n44905 = n9025 | n38119 ;
  assign n44906 = n44905 ^ n19427 ^ n6365 ;
  assign n44907 = n8435 ^ n6927 ^ 1'b0 ;
  assign n44908 = n33864 & ~n44907 ;
  assign n44910 = n21730 ^ n11678 ^ n6515 ;
  assign n44911 = n44910 ^ n15142 ^ n5876 ;
  assign n44909 = n19070 ^ n18222 ^ n985 ;
  assign n44912 = n44911 ^ n44909 ^ n38910 ;
  assign n44915 = ( n2153 & n24141 ) | ( n2153 & n30754 ) | ( n24141 & n30754 ) ;
  assign n44913 = n33926 ^ n5238 ^ n1306 ;
  assign n44914 = n4644 & n44913 ;
  assign n44916 = n44915 ^ n44914 ^ n19845 ;
  assign n44917 = n18621 ^ n12041 ^ n2839 ;
  assign n44918 = n44917 ^ n23605 ^ n7350 ;
  assign n44919 = n44145 ^ n13112 ^ n1877 ;
  assign n44920 = ( n17594 & n35998 ) | ( n17594 & n44919 ) | ( n35998 & n44919 ) ;
  assign n44921 = n31362 ^ n22802 ^ n15903 ;
  assign n44922 = n30884 & n44921 ;
  assign n44923 = ~n16275 & n44922 ;
  assign n44924 = ( ~n6725 & n15867 ) | ( ~n6725 & n20017 ) | ( n15867 & n20017 ) ;
  assign n44925 = ( n2128 & ~n26622 ) | ( n2128 & n44924 ) | ( ~n26622 & n44924 ) ;
  assign n44926 = n40094 ^ n10573 ^ 1'b0 ;
  assign n44928 = n2302 & ~n27221 ;
  assign n44927 = n22529 ^ n21921 ^ n17830 ;
  assign n44929 = n44928 ^ n44927 ^ n16006 ;
  assign n44930 = ( ~n15502 & n23662 ) | ( ~n15502 & n31038 ) | ( n23662 & n31038 ) ;
  assign n44931 = n44930 ^ n36972 ^ n16267 ;
  assign n44932 = ( n6105 & n26424 ) | ( n6105 & ~n44931 ) | ( n26424 & ~n44931 ) ;
  assign n44933 = n44932 ^ n12677 ^ n5670 ;
  assign n44934 = ( n15478 & ~n24161 ) | ( n15478 & n27772 ) | ( ~n24161 & n27772 ) ;
  assign n44937 = ( n3244 & ~n3850 ) | ( n3244 & n8072 ) | ( ~n3850 & n8072 ) ;
  assign n44938 = n44937 ^ n40415 ^ n28838 ;
  assign n44936 = ( n4593 & ~n8104 ) | ( n4593 & n11824 ) | ( ~n8104 & n11824 ) ;
  assign n44935 = n34082 ^ n4009 ^ 1'b0 ;
  assign n44939 = n44938 ^ n44936 ^ n44935 ;
  assign n44940 = n13792 ^ n9892 ^ n6534 ;
  assign n44941 = ( n10646 & n34435 ) | ( n10646 & ~n38529 ) | ( n34435 & ~n38529 ) ;
  assign n44942 = ~n6903 & n35736 ;
  assign n44943 = n44941 & n44942 ;
  assign n44944 = n27097 & ~n39201 ;
  assign n44945 = n44944 ^ n1588 ^ 1'b0 ;
  assign n44946 = n1305 & n44945 ;
  assign n44947 = n9984 ^ n8237 ^ 1'b0 ;
  assign n44948 = n26332 ^ n9069 ^ 1'b0 ;
  assign n44949 = n44947 & ~n44948 ;
  assign n44950 = ( n6951 & n20556 ) | ( n6951 & ~n44949 ) | ( n20556 & ~n44949 ) ;
  assign n44951 = ( n6655 & n23490 ) | ( n6655 & ~n24268 ) | ( n23490 & ~n24268 ) ;
  assign n44952 = ( n8909 & n15464 ) | ( n8909 & ~n18125 ) | ( n15464 & ~n18125 ) ;
  assign n44953 = n44952 ^ n9580 ^ 1'b0 ;
  assign n44954 = n12471 & n44953 ;
  assign n44955 = ( ~n8741 & n10711 ) | ( ~n8741 & n23654 ) | ( n10711 & n23654 ) ;
  assign n44956 = n1555 & n31477 ;
  assign n44957 = n10499 & n44956 ;
  assign n44958 = ( ~n8912 & n44955 ) | ( ~n8912 & n44957 ) | ( n44955 & n44957 ) ;
  assign n44959 = ( ~n33911 & n44954 ) | ( ~n33911 & n44958 ) | ( n44954 & n44958 ) ;
  assign n44960 = ( n6765 & ~n8201 ) | ( n6765 & n10144 ) | ( ~n8201 & n10144 ) ;
  assign n44961 = ( n3214 & n37805 ) | ( n3214 & ~n44960 ) | ( n37805 & ~n44960 ) ;
  assign n44963 = ~n13223 & n20699 ;
  assign n44962 = ( n22393 & n25362 ) | ( n22393 & n40042 ) | ( n25362 & n40042 ) ;
  assign n44964 = n44963 ^ n44962 ^ n7211 ;
  assign n44965 = n21112 ^ n18311 ^ n13974 ;
  assign n44966 = n44965 ^ n36030 ^ n21424 ;
  assign n44967 = n13171 ^ n2923 ^ n554 ;
  assign n44968 = ( n22920 & ~n26619 ) | ( n22920 & n44853 ) | ( ~n26619 & n44853 ) ;
  assign n44969 = ( n17535 & ~n44967 ) | ( n17535 & n44968 ) | ( ~n44967 & n44968 ) ;
  assign n44970 = ( n2053 & ~n18101 ) | ( n2053 & n43431 ) | ( ~n18101 & n43431 ) ;
  assign n44971 = n4324 ^ n332 ^ 1'b0 ;
  assign n44972 = n10054 & n44971 ;
  assign n44973 = ~n32811 & n44972 ;
  assign n44974 = n44973 ^ n6063 ^ 1'b0 ;
  assign n44975 = ( n3232 & ~n22692 ) | ( n3232 & n40452 ) | ( ~n22692 & n40452 ) ;
  assign n44976 = n12835 & n27318 ;
  assign n44977 = n44975 & n44976 ;
  assign n44978 = n27839 & ~n44977 ;
  assign n44979 = ~n23214 & n44978 ;
  assign n44980 = n28212 ^ n21793 ^ n15001 ;
  assign n44981 = n28288 ^ n24264 ^ n22691 ;
  assign n44982 = n43185 ^ n39537 ^ x94 ;
  assign n44983 = n13015 ^ n11945 ^ n7022 ;
  assign n44984 = n44983 ^ n11596 ^ 1'b0 ;
  assign n44985 = n28569 | n44984 ;
  assign n44986 = ~n23825 & n31445 ;
  assign n44987 = ( ~n38789 & n44985 ) | ( ~n38789 & n44986 ) | ( n44985 & n44986 ) ;
  assign n44988 = n11470 | n33592 ;
  assign n44989 = ( n6118 & n21249 ) | ( n6118 & ~n29293 ) | ( n21249 & ~n29293 ) ;
  assign n44990 = n44989 ^ n31240 ^ n22307 ;
  assign n44991 = ( n3152 & ~n32896 ) | ( n3152 & n44990 ) | ( ~n32896 & n44990 ) ;
  assign n44992 = n38449 ^ n11632 ^ n7888 ;
  assign n44993 = ( n13476 & ~n24936 ) | ( n13476 & n44992 ) | ( ~n24936 & n44992 ) ;
  assign n44994 = n44993 ^ n14593 ^ n10123 ;
  assign n44995 = n29536 ^ n23051 ^ n12169 ;
  assign n45002 = n16219 ^ n12168 ^ n10058 ;
  assign n45001 = ( n9537 & n32667 ) | ( n9537 & ~n41995 ) | ( n32667 & ~n41995 ) ;
  assign n44996 = n34848 ^ n27759 ^ 1'b0 ;
  assign n44997 = n19079 ^ n2286 ^ 1'b0 ;
  assign n44998 = ~n30530 & n44997 ;
  assign n44999 = ( n944 & ~n34037 ) | ( n944 & n44998 ) | ( ~n34037 & n44998 ) ;
  assign n45000 = ( ~n5163 & n44996 ) | ( ~n5163 & n44999 ) | ( n44996 & n44999 ) ;
  assign n45003 = n45002 ^ n45001 ^ n45000 ;
  assign n45004 = ( x237 & n17277 ) | ( x237 & ~n45003 ) | ( n17277 & ~n45003 ) ;
  assign n45005 = ( n17490 & n42597 ) | ( n17490 & ~n45004 ) | ( n42597 & ~n45004 ) ;
  assign n45006 = ( n1645 & n20885 ) | ( n1645 & ~n24178 ) | ( n20885 & ~n24178 ) ;
  assign n45007 = ( n12882 & n14791 ) | ( n12882 & ~n23590 ) | ( n14791 & ~n23590 ) ;
  assign n45008 = ( ~n12580 & n43179 ) | ( ~n12580 & n45007 ) | ( n43179 & n45007 ) ;
  assign n45009 = n33651 ^ n33101 ^ n13895 ;
  assign n45010 = ( n21375 & n23014 ) | ( n21375 & ~n38538 ) | ( n23014 & ~n38538 ) ;
  assign n45011 = n45010 ^ n31786 ^ n13122 ;
  assign n45012 = ( n45008 & ~n45009 ) | ( n45008 & n45011 ) | ( ~n45009 & n45011 ) ;
  assign n45013 = n16554 ^ n14950 ^ n2358 ;
  assign n45014 = ( n842 & n21382 ) | ( n842 & n38174 ) | ( n21382 & n38174 ) ;
  assign n45015 = ~n2196 & n45014 ;
  assign n45016 = ( ~n11071 & n11099 ) | ( ~n11071 & n17216 ) | ( n11099 & n17216 ) ;
  assign n45017 = ( ~n45013 & n45015 ) | ( ~n45013 & n45016 ) | ( n45015 & n45016 ) ;
  assign n45021 = ( n13085 & ~n24012 ) | ( n13085 & n43381 ) | ( ~n24012 & n43381 ) ;
  assign n45020 = ( n17345 & n18854 ) | ( n17345 & n28752 ) | ( n18854 & n28752 ) ;
  assign n45018 = ( ~n3063 & n17998 ) | ( ~n3063 & n35937 ) | ( n17998 & n35937 ) ;
  assign n45019 = n45018 ^ n44340 ^ n24262 ;
  assign n45022 = n45021 ^ n45020 ^ n45019 ;
  assign n45023 = n22146 ^ n17974 ^ 1'b0 ;
  assign n45024 = n32268 | n45023 ;
  assign n45025 = n12359 & ~n39685 ;
  assign n45026 = n8451 & n45025 ;
  assign n45027 = n14849 & n45026 ;
  assign n45028 = ( n1255 & ~n4667 ) | ( n1255 & n6857 ) | ( ~n4667 & n6857 ) ;
  assign n45029 = n45028 ^ n22657 ^ n2562 ;
  assign n45030 = ( ~n6625 & n15726 ) | ( ~n6625 & n45029 ) | ( n15726 & n45029 ) ;
  assign n45031 = n45030 ^ n11041 ^ n10405 ;
  assign n45032 = ( ~n45024 & n45027 ) | ( ~n45024 & n45031 ) | ( n45027 & n45031 ) ;
  assign n45037 = n3440 ^ n747 ^ n614 ;
  assign n45038 = ( n2487 & ~n23810 ) | ( n2487 & n45037 ) | ( ~n23810 & n45037 ) ;
  assign n45039 = ~n38626 & n45038 ;
  assign n45040 = n877 & n45039 ;
  assign n45033 = n24620 ^ n20171 ^ n6489 ;
  assign n45034 = n45033 ^ n34305 ^ 1'b0 ;
  assign n45035 = n6910 & n45034 ;
  assign n45036 = ( n11682 & n17542 ) | ( n11682 & n45035 ) | ( n17542 & n45035 ) ;
  assign n45041 = n45040 ^ n45036 ^ n5525 ;
  assign n45042 = n42154 ^ n20408 ^ 1'b0 ;
  assign n45043 = n28091 & ~n45042 ;
  assign n45044 = n29002 ^ n25037 ^ n1548 ;
  assign n45045 = n10199 | n19316 ;
  assign n45046 = n45044 | n45045 ;
  assign n45047 = n27773 & n45046 ;
  assign n45048 = n45047 ^ n10608 ^ 1'b0 ;
  assign n45049 = n27054 ^ n10024 ^ n3338 ;
  assign n45050 = n21438 ^ n17610 ^ n7179 ;
  assign n45055 = n5611 ^ n707 ^ 1'b0 ;
  assign n45056 = n44379 & ~n45055 ;
  assign n45051 = ( n5433 & n33446 ) | ( n5433 & ~n36459 ) | ( n33446 & ~n36459 ) ;
  assign n45052 = n45051 ^ n35228 ^ 1'b0 ;
  assign n45053 = n22478 ^ n21859 ^ 1'b0 ;
  assign n45054 = n45052 & n45053 ;
  assign n45057 = n45056 ^ n45054 ^ n39364 ;
  assign n45058 = n26499 & ~n45057 ;
  assign n45059 = ( n1136 & n5140 ) | ( n1136 & n6168 ) | ( n5140 & n6168 ) ;
  assign n45060 = ~n33300 & n45059 ;
  assign n45061 = n45060 ^ n15185 ^ n9995 ;
  assign n45063 = ~n4507 & n15805 ;
  assign n45062 = ( ~n2041 & n7889 ) | ( ~n2041 & n33170 ) | ( n7889 & n33170 ) ;
  assign n45064 = n45063 ^ n45062 ^ n9266 ;
  assign n45066 = n44439 ^ n16223 ^ n1478 ;
  assign n45065 = ( n3949 & ~n30795 ) | ( n3949 & n35640 ) | ( ~n30795 & n35640 ) ;
  assign n45067 = n45066 ^ n45065 ^ n42059 ;
  assign n45068 = n41397 ^ n28782 ^ n21617 ;
  assign n45069 = ( n36875 & n44830 ) | ( n36875 & ~n45068 ) | ( n44830 & ~n45068 ) ;
  assign n45070 = n4754 | n29710 ;
  assign n45071 = n27284 | n45070 ;
  assign n45072 = ( n8178 & n36372 ) | ( n8178 & ~n41096 ) | ( n36372 & ~n41096 ) ;
  assign n45073 = ( ~n5541 & n28147 ) | ( ~n5541 & n45072 ) | ( n28147 & n45072 ) ;
  assign n45074 = ( n2267 & n24558 ) | ( n2267 & n45073 ) | ( n24558 & n45073 ) ;
  assign n45077 = n30881 ^ n15821 ^ n11847 ;
  assign n45075 = ( ~n5384 & n13984 ) | ( ~n5384 & n20784 ) | ( n13984 & n20784 ) ;
  assign n45076 = n45075 ^ n33076 ^ n12170 ;
  assign n45078 = n45077 ^ n45076 ^ n7730 ;
  assign n45079 = n45078 ^ n30912 ^ 1'b0 ;
  assign n45080 = n45074 | n45079 ;
  assign n45081 = n32610 ^ n22625 ^ n7466 ;
  assign n45082 = n45081 ^ n10251 ^ n3050 ;
  assign n45083 = n17499 ^ n3134 ^ n2388 ;
  assign n45084 = ( n7658 & ~n13842 ) | ( n7658 & n45083 ) | ( ~n13842 & n45083 ) ;
  assign n45085 = ( n11965 & n34786 ) | ( n11965 & n45084 ) | ( n34786 & n45084 ) ;
  assign n45086 = ( n24697 & n25474 ) | ( n24697 & n39065 ) | ( n25474 & n39065 ) ;
  assign n45087 = n30609 & n45086 ;
  assign n45088 = n1330 & n2644 ;
  assign n45089 = ( n4187 & n9715 ) | ( n4187 & n45088 ) | ( n9715 & n45088 ) ;
  assign n45090 = n45089 ^ n8214 ^ n7845 ;
  assign n45091 = ( n23446 & n25996 ) | ( n23446 & n30184 ) | ( n25996 & n30184 ) ;
  assign n45092 = ( n9796 & ~n17296 ) | ( n9796 & n38279 ) | ( ~n17296 & n38279 ) ;
  assign n45093 = ( n11954 & n40861 ) | ( n11954 & n45092 ) | ( n40861 & n45092 ) ;
  assign n45094 = n12540 | n41257 ;
  assign n45095 = n24124 ^ n18531 ^ n8899 ;
  assign n45096 = ( n3355 & n35512 ) | ( n3355 & ~n45095 ) | ( n35512 & ~n45095 ) ;
  assign n45097 = ( n9453 & ~n41382 ) | ( n9453 & n45096 ) | ( ~n41382 & n45096 ) ;
  assign n45098 = n45097 ^ n16459 ^ 1'b0 ;
  assign n45099 = n28837 & ~n37179 ;
  assign n45100 = n45099 ^ n3525 ^ x209 ;
  assign n45101 = n45100 ^ n31693 ^ n27939 ;
  assign n45102 = ( n24850 & ~n45098 ) | ( n24850 & n45101 ) | ( ~n45098 & n45101 ) ;
  assign n45103 = ( n6421 & n27788 ) | ( n6421 & ~n41138 ) | ( n27788 & ~n41138 ) ;
  assign n45104 = n45103 ^ n34016 ^ 1'b0 ;
  assign n45105 = n4206 & ~n45104 ;
  assign n45106 = n1906 & ~n32439 ;
  assign n45107 = n45106 ^ n12036 ^ 1'b0 ;
  assign n45108 = n36302 ^ n27905 ^ n23185 ;
  assign n45109 = n45108 ^ n30129 ^ n11575 ;
  assign n45110 = n13147 & ~n29749 ;
  assign n45111 = n45110 ^ n5880 ^ 1'b0 ;
  assign n45112 = ~n15440 & n45111 ;
  assign n45113 = ~n1337 & n45112 ;
  assign n45114 = n25278 & ~n45113 ;
  assign n45115 = n15735 ^ n5854 ^ 1'b0 ;
  assign n45116 = ( n623 & n18539 ) | ( n623 & n45115 ) | ( n18539 & n45115 ) ;
  assign n45117 = n43586 ^ n26616 ^ n571 ;
  assign n45118 = n45117 ^ n39593 ^ 1'b0 ;
  assign n45119 = ( n2762 & n12175 ) | ( n2762 & ~n45118 ) | ( n12175 & ~n45118 ) ;
  assign n45120 = ( n14816 & n20518 ) | ( n14816 & ~n36970 ) | ( n20518 & ~n36970 ) ;
  assign n45121 = n37851 ^ n544 ^ 1'b0 ;
  assign n45122 = ( ~n5006 & n45120 ) | ( ~n5006 & n45121 ) | ( n45120 & n45121 ) ;
  assign n45123 = n33270 | n43275 ;
  assign n45124 = ( ~n26646 & n27931 ) | ( ~n26646 & n45123 ) | ( n27931 & n45123 ) ;
  assign n45125 = ( ~n2067 & n6981 ) | ( ~n2067 & n24640 ) | ( n6981 & n24640 ) ;
  assign n45126 = ~n18157 & n36303 ;
  assign n45127 = n45125 & n45126 ;
  assign n45128 = ( n6389 & n17874 ) | ( n6389 & ~n45127 ) | ( n17874 & ~n45127 ) ;
  assign n45129 = n45128 ^ n24431 ^ n15035 ;
  assign n45130 = n21617 ^ n18826 ^ 1'b0 ;
  assign n45131 = n15778 & ~n45130 ;
  assign n45132 = ( n20913 & n22801 ) | ( n20913 & ~n43622 ) | ( n22801 & ~n43622 ) ;
  assign n45133 = n24936 & ~n30817 ;
  assign n45134 = ( n22234 & n27349 ) | ( n22234 & ~n45133 ) | ( n27349 & ~n45133 ) ;
  assign n45135 = ( n24012 & n40505 ) | ( n24012 & ~n45134 ) | ( n40505 & ~n45134 ) ;
  assign n45136 = ( ~n17990 & n40466 ) | ( ~n17990 & n43986 ) | ( n40466 & n43986 ) ;
  assign n45137 = n12626 ^ n8318 ^ 1'b0 ;
  assign n45138 = ~n17893 & n45137 ;
  assign n45139 = ( ~n284 & n23214 ) | ( ~n284 & n29326 ) | ( n23214 & n29326 ) ;
  assign n45140 = n45139 ^ n16908 ^ n8903 ;
  assign n45141 = n33908 & n45140 ;
  assign n45142 = n1279 & n45141 ;
  assign n45144 = n9991 ^ x67 ^ 1'b0 ;
  assign n45143 = n32029 ^ n25640 ^ n3515 ;
  assign n45145 = n45144 ^ n45143 ^ n40515 ;
  assign n45146 = ( n45138 & ~n45142 ) | ( n45138 & n45145 ) | ( ~n45142 & n45145 ) ;
  assign n45147 = n29828 ^ n21493 ^ 1'b0 ;
  assign n45148 = ( n959 & n7754 ) | ( n959 & ~n24352 ) | ( n7754 & ~n24352 ) ;
  assign n45149 = n45147 | n45148 ;
  assign n45150 = ( n7487 & ~n12909 ) | ( n7487 & n20897 ) | ( ~n12909 & n20897 ) ;
  assign n45151 = ( n1726 & n6479 ) | ( n1726 & n17706 ) | ( n6479 & n17706 ) ;
  assign n45152 = n15984 ^ n2634 ^ 1'b0 ;
  assign n45153 = n45151 | n45152 ;
  assign n45154 = ( n29539 & ~n45150 ) | ( n29539 & n45153 ) | ( ~n45150 & n45153 ) ;
  assign n45155 = ( n12312 & n20086 ) | ( n12312 & n42577 ) | ( n20086 & n42577 ) ;
  assign n45158 = ( n877 & ~n4796 ) | ( n877 & n26390 ) | ( ~n4796 & n26390 ) ;
  assign n45156 = ( n7042 & n12955 ) | ( n7042 & n27134 ) | ( n12955 & n27134 ) ;
  assign n45157 = ( n11892 & n16788 ) | ( n11892 & n45156 ) | ( n16788 & n45156 ) ;
  assign n45159 = n45158 ^ n45157 ^ x236 ;
  assign n45160 = n45159 ^ n24161 ^ 1'b0 ;
  assign n45161 = n40028 & n45160 ;
  assign n45162 = n11653 ^ n6355 ^ 1'b0 ;
  assign n45163 = ~n8732 & n45162 ;
  assign n45164 = n45163 ^ n17678 ^ 1'b0 ;
  assign n45165 = ( ~n1135 & n6206 ) | ( ~n1135 & n20222 ) | ( n6206 & n20222 ) ;
  assign n45166 = ( ~n10397 & n29766 ) | ( ~n10397 & n45165 ) | ( n29766 & n45165 ) ;
  assign n45167 = ( ~n14073 & n42771 ) | ( ~n14073 & n45166 ) | ( n42771 & n45166 ) ;
  assign n45169 = n19092 ^ n10346 ^ n4781 ;
  assign n45170 = n20844 ^ n13828 ^ 1'b0 ;
  assign n45171 = n45169 & ~n45170 ;
  assign n45168 = n27413 ^ n12082 ^ 1'b0 ;
  assign n45172 = n45171 ^ n45168 ^ n28261 ;
  assign n45173 = ( n2784 & ~n7893 ) | ( n2784 & n13127 ) | ( ~n7893 & n13127 ) ;
  assign n45174 = ( n12313 & n40641 ) | ( n12313 & n45173 ) | ( n40641 & n45173 ) ;
  assign n45175 = ( n8830 & ~n19791 ) | ( n8830 & n27675 ) | ( ~n19791 & n27675 ) ;
  assign n45176 = n40836 ^ n12544 ^ 1'b0 ;
  assign n45177 = n43270 ^ n23660 ^ n20605 ;
  assign n45178 = n37486 ^ n21131 ^ n4522 ;
  assign n45179 = n9437 ^ n3649 ^ 1'b0 ;
  assign n45180 = ~n37836 & n45179 ;
  assign n45181 = ( ~n6863 & n45178 ) | ( ~n6863 & n45180 ) | ( n45178 & n45180 ) ;
  assign n45182 = n29734 ^ n22577 ^ 1'b0 ;
  assign n45183 = n9932 & n45182 ;
  assign n45184 = ~n28011 & n31068 ;
  assign n45185 = n45184 ^ n6694 ^ 1'b0 ;
  assign n45186 = ( n22294 & n31439 ) | ( n22294 & ~n35093 ) | ( n31439 & ~n35093 ) ;
  assign n45187 = n1435 | n19042 ;
  assign n45188 = n45186 & ~n45187 ;
  assign n45189 = n16999 ^ n10267 ^ n4765 ;
  assign n45190 = n10722 | n14045 ;
  assign n45191 = n45190 ^ n26893 ^ n6765 ;
  assign n45192 = ( n8946 & n25977 ) | ( n8946 & n26114 ) | ( n25977 & n26114 ) ;
  assign n45193 = n45192 ^ n10567 ^ n5411 ;
  assign n45194 = n26897 ^ n10564 ^ 1'b0 ;
  assign n45195 = n15157 | n45194 ;
  assign n45196 = ( n13648 & ~n21240 ) | ( n13648 & n31822 ) | ( ~n21240 & n31822 ) ;
  assign n45197 = ( n4032 & n37686 ) | ( n4032 & ~n45196 ) | ( n37686 & ~n45196 ) ;
  assign n45198 = ( n22727 & ~n45195 ) | ( n22727 & n45197 ) | ( ~n45195 & n45197 ) ;
  assign n45199 = ( n15505 & n25385 ) | ( n15505 & n38678 ) | ( n25385 & n38678 ) ;
  assign n45200 = n45199 ^ n2695 ^ n2511 ;
  assign n45201 = ( n2248 & n13719 ) | ( n2248 & ~n45200 ) | ( n13719 & ~n45200 ) ;
  assign n45202 = n7463 | n24815 ;
  assign n45203 = n2781 | n45202 ;
  assign n45204 = ( ~n14076 & n18243 ) | ( ~n14076 & n27224 ) | ( n18243 & n27224 ) ;
  assign n45205 = n45204 ^ n17107 ^ n7232 ;
  assign n45206 = ( n23130 & ~n45203 ) | ( n23130 & n45205 ) | ( ~n45203 & n45205 ) ;
  assign n45207 = n45206 ^ n38361 ^ n28810 ;
  assign n45208 = n32328 ^ n13683 ^ x17 ;
  assign n45209 = n35815 ^ n12461 ^ 1'b0 ;
  assign n45210 = n35580 ^ n16611 ^ n13517 ;
  assign n45211 = n599 & n45210 ;
  assign n45212 = n45211 ^ n7110 ^ 1'b0 ;
  assign n45216 = ( n5237 & n10848 ) | ( n5237 & ~n28247 ) | ( n10848 & ~n28247 ) ;
  assign n45214 = ( ~n2157 & n27469 ) | ( ~n2157 & n27777 ) | ( n27469 & n27777 ) ;
  assign n45215 = ( n4810 & n17115 ) | ( n4810 & ~n45214 ) | ( n17115 & ~n45214 ) ;
  assign n45213 = n42899 ^ n26700 ^ n21340 ;
  assign n45217 = n45216 ^ n45215 ^ n45213 ;
  assign n45218 = n34342 ^ n33497 ^ n32572 ;
  assign n45219 = ( n5072 & n28805 ) | ( n5072 & n29019 ) | ( n28805 & n29019 ) ;
  assign n45220 = ( n4071 & n40325 ) | ( n4071 & ~n42161 ) | ( n40325 & ~n42161 ) ;
  assign n45221 = ( n35435 & n38417 ) | ( n35435 & ~n45220 ) | ( n38417 & ~n45220 ) ;
  assign n45222 = ( n6224 & n19729 ) | ( n6224 & n27051 ) | ( n19729 & n27051 ) ;
  assign n45224 = ( ~n5801 & n16658 ) | ( ~n5801 & n20937 ) | ( n16658 & n20937 ) ;
  assign n45223 = n34836 ^ n24738 ^ n1720 ;
  assign n45225 = n45224 ^ n45223 ^ n14575 ;
  assign n45226 = n15178 ^ n7891 ^ x156 ;
  assign n45227 = n37124 ^ n21826 ^ n5635 ;
  assign n45228 = ~n11606 & n34952 ;
  assign n45229 = n9981 & n28412 ;
  assign n45230 = n45229 ^ n2001 ^ 1'b0 ;
  assign n45231 = n18594 ^ n17854 ^ n5464 ;
  assign n45232 = n25722 ^ n12400 ^ n4129 ;
  assign n45233 = ( n3498 & n32525 ) | ( n3498 & n45232 ) | ( n32525 & n45232 ) ;
  assign n45235 = n2732 & ~n5010 ;
  assign n45236 = ~n2087 & n14285 ;
  assign n45237 = n8831 & n45236 ;
  assign n45238 = n45237 ^ n32328 ^ n2713 ;
  assign n45239 = n45235 & n45238 ;
  assign n45234 = n36335 ^ n26523 ^ n7010 ;
  assign n45240 = n45239 ^ n45234 ^ n18162 ;
  assign n45241 = ( ~x52 & n29345 ) | ( ~x52 & n43162 ) | ( n29345 & n43162 ) ;
  assign n45242 = n32560 ^ n9570 ^ 1'b0 ;
  assign n45243 = ~n16208 & n45242 ;
  assign n45244 = ( ~n3432 & n31810 ) | ( ~n3432 & n38220 ) | ( n31810 & n38220 ) ;
  assign n45245 = n17652 & ~n38252 ;
  assign n45246 = n31398 & n45245 ;
  assign n45247 = ( n26517 & n45244 ) | ( n26517 & n45246 ) | ( n45244 & n45246 ) ;
  assign n45248 = ( n6238 & n10707 ) | ( n6238 & ~n20723 ) | ( n10707 & ~n20723 ) ;
  assign n45249 = ( ~n20214 & n22831 ) | ( ~n20214 & n23914 ) | ( n22831 & n23914 ) ;
  assign n45250 = ( n18972 & n45248 ) | ( n18972 & n45249 ) | ( n45248 & n45249 ) ;
  assign n45251 = n45076 ^ n31011 ^ n7107 ;
  assign n45252 = ( n2968 & n7024 ) | ( n2968 & n43861 ) | ( n7024 & n43861 ) ;
  assign n45253 = n31168 ^ n19818 ^ n14884 ;
  assign n45254 = ( n10779 & n37381 ) | ( n10779 & ~n45253 ) | ( n37381 & ~n45253 ) ;
  assign n45255 = n43825 ^ n21200 ^ n4261 ;
  assign n45256 = ( ~n2517 & n2661 ) | ( ~n2517 & n28247 ) | ( n2661 & n28247 ) ;
  assign n45257 = n11574 | n23365 ;
  assign n45258 = n45257 ^ n9680 ^ 1'b0 ;
  assign n45259 = ( n8960 & ~n15119 ) | ( n8960 & n30503 ) | ( ~n15119 & n30503 ) ;
  assign n45260 = n45259 ^ n13157 ^ n9939 ;
  assign n45261 = ( ~n2674 & n37189 ) | ( ~n2674 & n39264 ) | ( n37189 & n39264 ) ;
  assign n45262 = n31126 ^ n23188 ^ n4003 ;
  assign n45263 = n30075 ^ n15654 ^ n12493 ;
  assign n45264 = ( n23223 & ~n45262 ) | ( n23223 & n45263 ) | ( ~n45262 & n45263 ) ;
  assign n45265 = n19726 ^ n10082 ^ n1000 ;
  assign n45266 = n45265 ^ n38858 ^ n23445 ;
  assign n45267 = n15470 ^ n13292 ^ n1528 ;
  assign n45273 = ( n11765 & ~n30618 ) | ( n11765 & n41232 ) | ( ~n30618 & n41232 ) ;
  assign n45271 = ( n1762 & n9707 ) | ( n1762 & n25501 ) | ( n9707 & n25501 ) ;
  assign n45268 = n19393 ^ n5916 ^ 1'b0 ;
  assign n45269 = n45268 ^ n37562 ^ n1092 ;
  assign n45270 = ~n12746 & n45269 ;
  assign n45272 = n45271 ^ n45270 ^ 1'b0 ;
  assign n45274 = n45273 ^ n45272 ^ n26534 ;
  assign n45275 = ( n1424 & ~n45267 ) | ( n1424 & n45274 ) | ( ~n45267 & n45274 ) ;
  assign n45282 = ~n27419 & n35430 ;
  assign n45283 = n44541 & n45282 ;
  assign n45276 = ( ~n2573 & n7610 ) | ( ~n2573 & n17046 ) | ( n7610 & n17046 ) ;
  assign n45277 = n45276 ^ n28692 ^ n14044 ;
  assign n45278 = n45277 ^ n6020 ^ 1'b0 ;
  assign n45279 = ~n23216 & n45278 ;
  assign n45280 = n42167 ^ n37394 ^ n11410 ;
  assign n45281 = ( ~n41715 & n45279 ) | ( ~n41715 & n45280 ) | ( n45279 & n45280 ) ;
  assign n45284 = n45283 ^ n45281 ^ n25360 ;
  assign n45288 = n38215 ^ n16878 ^ n7909 ;
  assign n45285 = n44083 ^ n36074 ^ n16110 ;
  assign n45286 = ( n24735 & n33732 ) | ( n24735 & ~n35843 ) | ( n33732 & ~n35843 ) ;
  assign n45287 = ( n16198 & n45285 ) | ( n16198 & ~n45286 ) | ( n45285 & ~n45286 ) ;
  assign n45289 = n45288 ^ n45287 ^ n8971 ;
  assign n45290 = ( n15521 & n17307 ) | ( n15521 & n31084 ) | ( n17307 & n31084 ) ;
  assign n45291 = n3624 & n45290 ;
  assign n45292 = ~n14026 & n45291 ;
  assign n45293 = n24461 ^ n16831 ^ n4233 ;
  assign n45294 = n40312 ^ n26277 ^ n8856 ;
  assign n45295 = ( n23446 & ~n45293 ) | ( n23446 & n45294 ) | ( ~n45293 & n45294 ) ;
  assign n45296 = ~n8129 & n22769 ;
  assign n45297 = n12224 ^ n1191 ^ n632 ;
  assign n45298 = n45297 ^ n41122 ^ n10164 ;
  assign n45299 = n16275 ^ n13599 ^ n13519 ;
  assign n45300 = ( ~n2675 & n3081 ) | ( ~n2675 & n24072 ) | ( n3081 & n24072 ) ;
  assign n45301 = n45300 ^ n26632 ^ n17075 ;
  assign n45302 = n45301 ^ n36059 ^ n17315 ;
  assign n45303 = n45302 ^ n24384 ^ n3242 ;
  assign n45304 = n45303 ^ n28695 ^ n27817 ;
  assign n45305 = n38244 ^ n35571 ^ n12060 ;
  assign n45306 = ( ~n11654 & n43895 ) | ( ~n11654 & n45305 ) | ( n43895 & n45305 ) ;
  assign n45307 = ( ~n9079 & n24397 ) | ( ~n9079 & n31142 ) | ( n24397 & n31142 ) ;
  assign n45308 = n21481 & n22312 ;
  assign n45309 = n22529 & n45308 ;
  assign n45312 = ( n1795 & n30261 ) | ( n1795 & ~n39008 ) | ( n30261 & ~n39008 ) ;
  assign n45310 = n34331 ^ n16173 ^ n9497 ;
  assign n45311 = n45310 ^ n31190 ^ n575 ;
  assign n45313 = n45312 ^ n45311 ^ n21253 ;
  assign n45314 = n41149 ^ n22961 ^ n7626 ;
  assign n45315 = n45314 ^ n5783 ^ n4523 ;
  assign n45316 = ( n5902 & n17286 ) | ( n5902 & n37108 ) | ( n17286 & n37108 ) ;
  assign n45317 = n13601 ^ n9070 ^ n1464 ;
  assign n45318 = ( n3543 & ~n43287 ) | ( n3543 & n45317 ) | ( ~n43287 & n45317 ) ;
  assign n45319 = ( n2124 & n23340 ) | ( n2124 & n45318 ) | ( n23340 & n45318 ) ;
  assign n45320 = n17231 & n45319 ;
  assign n45321 = n45320 ^ n38918 ^ 1'b0 ;
  assign n45322 = n45321 ^ n32676 ^ n24391 ;
  assign n45323 = n38351 ^ n28333 ^ n12735 ;
  assign n45324 = n37390 ^ n14917 ^ n12340 ;
  assign n45325 = n579 & n25122 ;
  assign n45326 = n45325 ^ n20894 ^ 1'b0 ;
  assign n45327 = ( ~n21844 & n23305 ) | ( ~n21844 & n35694 ) | ( n23305 & n35694 ) ;
  assign n45328 = ( n19506 & n30656 ) | ( n19506 & ~n45327 ) | ( n30656 & ~n45327 ) ;
  assign n45329 = n45328 ^ n29559 ^ n28965 ;
  assign n45330 = ( ~n22973 & n25274 ) | ( ~n22973 & n31687 ) | ( n25274 & n31687 ) ;
  assign n45331 = n38373 ^ n2550 ^ 1'b0 ;
  assign n45332 = n23274 | n45331 ;
  assign n45333 = ( n11905 & n42966 ) | ( n11905 & n45332 ) | ( n42966 & n45332 ) ;
  assign n45334 = ( ~n7212 & n27245 ) | ( ~n7212 & n45333 ) | ( n27245 & n45333 ) ;
  assign n45335 = ~n8114 & n45334 ;
  assign n45336 = ( n3325 & n23740 ) | ( n3325 & n44348 ) | ( n23740 & n44348 ) ;
  assign n45337 = ( n11539 & n39088 ) | ( n11539 & n41465 ) | ( n39088 & n41465 ) ;
  assign n45338 = n28925 ^ n11612 ^ n10434 ;
  assign n45339 = n45337 & ~n45338 ;
  assign n45340 = n36926 ^ n28157 ^ n13020 ;
  assign n45341 = n33537 ^ n22641 ^ n20109 ;
  assign n45342 = n45341 ^ n10390 ^ n5845 ;
  assign n45346 = n11326 ^ n9451 ^ 1'b0 ;
  assign n45347 = n45346 ^ n14887 ^ n14145 ;
  assign n45343 = n10068 | n19179 ;
  assign n45344 = n45343 ^ n3863 ^ 1'b0 ;
  assign n45345 = n38933 | n45344 ;
  assign n45348 = n45347 ^ n45345 ^ 1'b0 ;
  assign n45349 = n7737 & n8001 ;
  assign n45350 = n30978 & n45349 ;
  assign n45351 = ( ~n1076 & n10451 ) | ( ~n1076 & n34928 ) | ( n10451 & n34928 ) ;
  assign n45352 = ( n5728 & n14907 ) | ( n5728 & n45351 ) | ( n14907 & n45351 ) ;
  assign n45353 = n19262 ^ n18325 ^ n10025 ;
  assign n45354 = n45353 ^ n5918 ^ 1'b0 ;
  assign n45355 = n45354 ^ n25790 ^ n2452 ;
  assign n45359 = ( n1340 & ~n25668 ) | ( n1340 & n37551 ) | ( ~n25668 & n37551 ) ;
  assign n45356 = n15226 ^ n6536 ^ n909 ;
  assign n45357 = ( n2019 & n9605 ) | ( n2019 & n45356 ) | ( n9605 & n45356 ) ;
  assign n45358 = ( n6847 & n15775 ) | ( n6847 & n45357 ) | ( n15775 & n45357 ) ;
  assign n45360 = n45359 ^ n45358 ^ n44882 ;
  assign n45361 = n41626 ^ n11488 ^ n11416 ;
  assign n45362 = ( n542 & n11878 ) | ( n542 & n21154 ) | ( n11878 & n21154 ) ;
  assign n45363 = n45362 ^ n29828 ^ n19641 ;
  assign n45364 = n12215 ^ n7833 ^ n6017 ;
  assign n45365 = ~n24980 & n28168 ;
  assign n45366 = ( ~n1330 & n6359 ) | ( ~n1330 & n11299 ) | ( n6359 & n11299 ) ;
  assign n45368 = ( n2167 & n14673 ) | ( n2167 & ~n21602 ) | ( n14673 & ~n21602 ) ;
  assign n45369 = n45368 ^ n6512 ^ n2468 ;
  assign n45367 = x125 & n40133 ;
  assign n45370 = n45369 ^ n45367 ^ 1'b0 ;
  assign n45371 = ( n4142 & ~n11069 ) | ( n4142 & n14852 ) | ( ~n11069 & n14852 ) ;
  assign n45372 = ( n1739 & n45370 ) | ( n1739 & n45371 ) | ( n45370 & n45371 ) ;
  assign n45373 = n25333 ^ n10250 ^ n3480 ;
  assign n45374 = ( n291 & n2919 ) | ( n291 & n45373 ) | ( n2919 & n45373 ) ;
  assign n45375 = ( n8666 & ~n12593 ) | ( n8666 & n14435 ) | ( ~n12593 & n14435 ) ;
  assign n45376 = n45375 ^ n26662 ^ n20657 ;
  assign n45377 = ( n23310 & n45374 ) | ( n23310 & n45376 ) | ( n45374 & n45376 ) ;
  assign n45378 = ( ~n12403 & n17611 ) | ( ~n12403 & n34889 ) | ( n17611 & n34889 ) ;
  assign n45379 = ( n4725 & ~n7929 ) | ( n4725 & n30824 ) | ( ~n7929 & n30824 ) ;
  assign n45380 = n45379 ^ n10390 ^ n8134 ;
  assign n45381 = ( n2363 & n45378 ) | ( n2363 & ~n45380 ) | ( n45378 & ~n45380 ) ;
  assign n45382 = ( ~n1116 & n12125 ) | ( ~n1116 & n18549 ) | ( n12125 & n18549 ) ;
  assign n45383 = ( n5515 & n10602 ) | ( n5515 & ~n45382 ) | ( n10602 & ~n45382 ) ;
  assign n45384 = n27990 ^ n20777 ^ n15404 ;
  assign n45385 = ( n12890 & ~n40974 ) | ( n12890 & n45384 ) | ( ~n40974 & n45384 ) ;
  assign n45388 = n31600 ^ n8376 ^ n5444 ;
  assign n45386 = n13752 | n27249 ;
  assign n45387 = n45386 ^ n38807 ^ n14225 ;
  assign n45389 = n45388 ^ n45387 ^ n29385 ;
  assign n45390 = n45389 ^ n42716 ^ n27376 ;
  assign n45391 = n19840 ^ n13660 ^ n1514 ;
  assign n45392 = n28940 | n45391 ;
  assign n45393 = n45120 ^ n15551 ^ n8201 ;
  assign n45394 = n30505 ^ n23393 ^ 1'b0 ;
  assign n45395 = ~n45393 & n45394 ;
  assign n45397 = ( n7978 & n22852 ) | ( n7978 & ~n28877 ) | ( n22852 & ~n28877 ) ;
  assign n45396 = ( ~n10758 & n15215 ) | ( ~n10758 & n27311 ) | ( n15215 & n27311 ) ;
  assign n45398 = n45397 ^ n45396 ^ n29881 ;
  assign n45401 = ( n4288 & ~n5192 ) | ( n4288 & n6208 ) | ( ~n5192 & n6208 ) ;
  assign n45400 = n32489 ^ n15564 ^ n332 ;
  assign n45399 = n11910 & n37128 ;
  assign n45402 = n45401 ^ n45400 ^ n45399 ;
  assign n45404 = ( n7409 & n19747 ) | ( n7409 & n33889 ) | ( n19747 & n33889 ) ;
  assign n45403 = ( n19630 & n30089 ) | ( n19630 & ~n36351 ) | ( n30089 & ~n36351 ) ;
  assign n45405 = n45404 ^ n45403 ^ n24953 ;
  assign n45406 = n45405 ^ n34177 ^ 1'b0 ;
  assign n45407 = ( ~n7173 & n29953 ) | ( ~n7173 & n45406 ) | ( n29953 & n45406 ) ;
  assign n45408 = n30305 ^ n12498 ^ n3242 ;
  assign n45409 = n12126 & n14886 ;
  assign n45410 = ( n9789 & n18799 ) | ( n9789 & n21760 ) | ( n18799 & n21760 ) ;
  assign n45411 = n45410 ^ n43360 ^ n12607 ;
  assign n45412 = ( n12587 & n17609 ) | ( n12587 & n18078 ) | ( n17609 & n18078 ) ;
  assign n45413 = n21125 & n45412 ;
  assign n45414 = ( n7114 & n8468 ) | ( n7114 & n45413 ) | ( n8468 & n45413 ) ;
  assign n45415 = ( n26277 & ~n39154 ) | ( n26277 & n45414 ) | ( ~n39154 & n45414 ) ;
  assign n45416 = n982 & ~n28081 ;
  assign n45417 = ~n3380 & n18330 ;
  assign n45418 = n27186 & n45417 ;
  assign n45419 = n16146 & n18805 ;
  assign n45420 = ~n21806 & n45419 ;
  assign n45421 = n45420 ^ n1907 ^ 1'b0 ;
  assign n45422 = n22310 | n45421 ;
  assign n45423 = n43203 ^ n31660 ^ n7774 ;
  assign n45424 = n38533 ^ n28576 ^ n7251 ;
  assign n45425 = ( ~n7791 & n36598 ) | ( ~n7791 & n45424 ) | ( n36598 & n45424 ) ;
  assign n45426 = n40859 ^ n13523 ^ n4974 ;
  assign n45427 = n45426 ^ n18785 ^ 1'b0 ;
  assign n45428 = n45427 ^ n36759 ^ 1'b0 ;
  assign n45429 = ( n1975 & ~n2056 ) | ( n1975 & n34431 ) | ( ~n2056 & n34431 ) ;
  assign n45431 = n27900 ^ n13864 ^ n10416 ;
  assign n45432 = ( n39635 & ~n41435 ) | ( n39635 & n45431 ) | ( ~n41435 & n45431 ) ;
  assign n45433 = n45432 ^ n30911 ^ 1'b0 ;
  assign n45430 = n28600 ^ n23477 ^ n9733 ;
  assign n45434 = n45433 ^ n45430 ^ n30824 ;
  assign n45437 = n9805 ^ n5552 ^ 1'b0 ;
  assign n45438 = n45437 ^ n15551 ^ n9677 ;
  assign n45439 = ( n6926 & ~n9114 ) | ( n6926 & n45438 ) | ( ~n9114 & n45438 ) ;
  assign n45436 = ( n5923 & n30214 ) | ( n5923 & ~n42898 ) | ( n30214 & ~n42898 ) ;
  assign n45435 = ( n14978 & ~n18881 ) | ( n14978 & n36399 ) | ( ~n18881 & n36399 ) ;
  assign n45440 = n45439 ^ n45436 ^ n45435 ;
  assign n45441 = ( ~n4027 & n25843 ) | ( ~n4027 & n45440 ) | ( n25843 & n45440 ) ;
  assign n45442 = ~n4346 & n17056 ;
  assign n45443 = n45442 ^ n34963 ^ 1'b0 ;
  assign n45444 = ( x73 & ~n6765 ) | ( x73 & n8298 ) | ( ~n6765 & n8298 ) ;
  assign n45445 = n18204 & n22355 ;
  assign n45446 = n45444 & n45445 ;
  assign n45448 = n30978 ^ n11195 ^ 1'b0 ;
  assign n45447 = n13635 ^ n6527 ^ n914 ;
  assign n45449 = n45448 ^ n45447 ^ n17211 ;
  assign n45450 = n38005 ^ n15282 ^ n3310 ;
  assign n45451 = ~n4128 & n45450 ;
  assign n45452 = ( n29423 & ~n30400 ) | ( n29423 & n45451 ) | ( ~n30400 & n45451 ) ;
  assign n45453 = ( n6287 & n40685 ) | ( n6287 & n44001 ) | ( n40685 & n44001 ) ;
  assign n45454 = ( ~n773 & n15848 ) | ( ~n773 & n45453 ) | ( n15848 & n45453 ) ;
  assign n45455 = n21817 ^ n9092 ^ 1'b0 ;
  assign n45456 = ( ~n5629 & n8557 ) | ( ~n5629 & n34373 ) | ( n8557 & n34373 ) ;
  assign n45457 = ( x176 & ~n17866 ) | ( x176 & n34052 ) | ( ~n17866 & n34052 ) ;
  assign n45460 = n22097 ^ n20875 ^ n7863 ;
  assign n45458 = n17937 & n23002 ;
  assign n45459 = n36148 & n45458 ;
  assign n45461 = n45460 ^ n45459 ^ n1286 ;
  assign n45462 = ( n5739 & ~n45457 ) | ( n5739 & n45461 ) | ( ~n45457 & n45461 ) ;
  assign n45463 = n25206 ^ n23005 ^ n21312 ;
  assign n45464 = ( n554 & n955 ) | ( n554 & n3532 ) | ( n955 & n3532 ) ;
  assign n45465 = n15996 & n45464 ;
  assign n45466 = ~n38594 & n45465 ;
  assign n45467 = ~n28899 & n42638 ;
  assign n45468 = x213 & ~n33445 ;
  assign n45469 = n45467 & n45468 ;
  assign n45470 = n26859 ^ n23154 ^ n17366 ;
  assign n45471 = n45470 ^ n40556 ^ n26564 ;
  assign n45472 = ( n7905 & n17332 ) | ( n7905 & ~n37077 ) | ( n17332 & ~n37077 ) ;
  assign n45473 = ( n1742 & ~n11338 ) | ( n1742 & n20144 ) | ( ~n11338 & n20144 ) ;
  assign n45474 = ~n13381 & n45473 ;
  assign n45475 = ~n4289 & n45474 ;
  assign n45476 = n45475 ^ n31727 ^ n22511 ;
  assign n45477 = ( n3138 & n15715 ) | ( n3138 & n26836 ) | ( n15715 & n26836 ) ;
  assign n45478 = ( n3342 & n3859 ) | ( n3342 & ~n14738 ) | ( n3859 & ~n14738 ) ;
  assign n45479 = n45478 ^ n23529 ^ n7430 ;
  assign n45480 = ( n4650 & n18362 ) | ( n4650 & n35761 ) | ( n18362 & n35761 ) ;
  assign n45482 = n27799 ^ n19665 ^ n308 ;
  assign n45483 = n45482 ^ n15357 ^ 1'b0 ;
  assign n45481 = ( n7329 & ~n15052 ) | ( n7329 & n37885 ) | ( ~n15052 & n37885 ) ;
  assign n45484 = n45483 ^ n45481 ^ n10991 ;
  assign n45485 = ~n11840 & n37719 ;
  assign n45486 = n45485 ^ n30967 ^ 1'b0 ;
  assign n45487 = n20200 ^ n1325 ^ 1'b0 ;
  assign n45488 = n6464 & n45487 ;
  assign n45489 = n45488 ^ n21019 ^ 1'b0 ;
  assign n45490 = n1670 & ~n7824 ;
  assign n45491 = ( ~n2341 & n19712 ) | ( ~n2341 & n45490 ) | ( n19712 & n45490 ) ;
  assign n45492 = ( n5087 & n39805 ) | ( n5087 & n42038 ) | ( n39805 & n42038 ) ;
  assign n45493 = n12030 ^ n10715 ^ 1'b0 ;
  assign n45494 = ~n34877 & n45493 ;
  assign n45495 = n30343 | n42616 ;
  assign n45498 = ( n10430 & ~n13342 ) | ( n10430 & n16007 ) | ( ~n13342 & n16007 ) ;
  assign n45499 = n45498 ^ n42762 ^ n6216 ;
  assign n45496 = ~n2662 & n6304 ;
  assign n45497 = ( n3223 & ~n3255 ) | ( n3223 & n45496 ) | ( ~n3255 & n45496 ) ;
  assign n45500 = n45499 ^ n45497 ^ n19646 ;
  assign n45502 = ( n5053 & ~n7227 ) | ( n5053 & n23223 ) | ( ~n7227 & n23223 ) ;
  assign n45501 = n30347 ^ n17004 ^ n2140 ;
  assign n45503 = n45502 ^ n45501 ^ n36030 ;
  assign n45504 = n45503 ^ n1687 ^ 1'b0 ;
  assign n45505 = n45500 & n45504 ;
  assign n45506 = ( ~n45494 & n45495 ) | ( ~n45494 & n45505 ) | ( n45495 & n45505 ) ;
  assign n45507 = ( n25079 & ~n29747 ) | ( n25079 & n32154 ) | ( ~n29747 & n32154 ) ;
  assign n45509 = ( n7035 & ~n12275 ) | ( n7035 & n28043 ) | ( ~n12275 & n28043 ) ;
  assign n45508 = ( n11317 & n15132 ) | ( n11317 & ~n38521 ) | ( n15132 & ~n38521 ) ;
  assign n45510 = n45509 ^ n45508 ^ n31699 ;
  assign n45511 = n19084 ^ n4404 ^ n3296 ;
  assign n45512 = ( n9679 & n27500 ) | ( n9679 & ~n45511 ) | ( n27500 & ~n45511 ) ;
  assign n45513 = n42647 ^ n26362 ^ n7240 ;
  assign n45514 = n45513 ^ n26470 ^ n724 ;
  assign n45515 = n8446 & n15406 ;
  assign n45516 = n45515 ^ n12654 ^ 1'b0 ;
  assign n45518 = ( ~n1435 & n8541 ) | ( ~n1435 & n12388 ) | ( n8541 & n12388 ) ;
  assign n45519 = ( n26286 & n28096 ) | ( n26286 & n45518 ) | ( n28096 & n45518 ) ;
  assign n45517 = n43712 ^ n22604 ^ n15329 ;
  assign n45520 = n45519 ^ n45517 ^ n11669 ;
  assign n45521 = n45520 ^ n37744 ^ 1'b0 ;
  assign n45522 = n45516 | n45521 ;
  assign n45523 = n35835 ^ n25273 ^ n14162 ;
  assign n45524 = n36511 ^ n16802 ^ n417 ;
  assign n45525 = ( n12849 & n41683 ) | ( n12849 & n45524 ) | ( n41683 & n45524 ) ;
  assign n45526 = n23167 ^ n22001 ^ 1'b0 ;
  assign n45527 = ( n7772 & n8400 ) | ( n7772 & ~n18539 ) | ( n8400 & ~n18539 ) ;
  assign n45528 = ( n7862 & n25228 ) | ( n7862 & ~n42781 ) | ( n25228 & ~n42781 ) ;
  assign n45529 = n34517 ^ n18688 ^ n7183 ;
  assign n45530 = ( ~n18563 & n45528 ) | ( ~n18563 & n45529 ) | ( n45528 & n45529 ) ;
  assign n45531 = ( n9568 & ~n12866 ) | ( n9568 & n17308 ) | ( ~n12866 & n17308 ) ;
  assign n45532 = ( n16554 & n33316 ) | ( n16554 & n45531 ) | ( n33316 & n45531 ) ;
  assign n45533 = n24993 ^ n15589 ^ n8700 ;
  assign n45534 = ( n3831 & n27854 ) | ( n3831 & ~n45533 ) | ( n27854 & ~n45533 ) ;
  assign n45535 = n45534 ^ n11535 ^ n6100 ;
  assign n45536 = n28915 ^ n12867 ^ n9968 ;
  assign n45537 = n17713 ^ n5306 ^ 1'b0 ;
  assign n45538 = n16429 | n45537 ;
  assign n45539 = n25558 ^ n14878 ^ n8476 ;
  assign n45540 = ( n10364 & n14156 ) | ( n10364 & n45539 ) | ( n14156 & n45539 ) ;
  assign n45541 = ( ~n20243 & n44698 ) | ( ~n20243 & n45540 ) | ( n44698 & n45540 ) ;
  assign n45543 = n31983 ^ n11614 ^ n4526 ;
  assign n45544 = n45543 ^ n32487 ^ n3462 ;
  assign n45542 = ( n4886 & n16462 ) | ( n4886 & ~n37585 ) | ( n16462 & ~n37585 ) ;
  assign n45545 = n45544 ^ n45542 ^ n38103 ;
  assign n45551 = n31424 ^ n23529 ^ n22708 ;
  assign n45546 = ( ~n881 & n11415 ) | ( ~n881 & n39511 ) | ( n11415 & n39511 ) ;
  assign n45547 = n23282 | n33113 ;
  assign n45548 = n45547 ^ n27085 ^ 1'b0 ;
  assign n45549 = ( ~n3917 & n38823 ) | ( ~n3917 & n45548 ) | ( n38823 & n45548 ) ;
  assign n45550 = ( n13619 & n45546 ) | ( n13619 & ~n45549 ) | ( n45546 & ~n45549 ) ;
  assign n45552 = n45551 ^ n45550 ^ n27738 ;
  assign n45553 = ( ~n1106 & n34879 ) | ( ~n1106 & n37773 ) | ( n34879 & n37773 ) ;
  assign n45554 = n45553 ^ n26664 ^ n22920 ;
  assign n45555 = ~n12231 & n28718 ;
  assign n45556 = n45555 ^ n4321 ^ 1'b0 ;
  assign n45557 = ( n15537 & ~n25326 ) | ( n15537 & n45556 ) | ( ~n25326 & n45556 ) ;
  assign n45558 = n41458 ^ n30055 ^ n15678 ;
  assign n45559 = ( n40264 & ~n45557 ) | ( n40264 & n45558 ) | ( ~n45557 & n45558 ) ;
  assign n45560 = n32689 ^ n22183 ^ 1'b0 ;
  assign n45561 = ( n1119 & n39041 ) | ( n1119 & ~n45560 ) | ( n39041 & ~n45560 ) ;
  assign n45562 = n13282 & n27761 ;
  assign n45563 = ~x195 & n45562 ;
  assign n45564 = ( n10901 & n23779 ) | ( n10901 & ~n45563 ) | ( n23779 & ~n45563 ) ;
  assign n45565 = x85 & ~n31331 ;
  assign n45566 = n45565 ^ n357 ^ 1'b0 ;
  assign n45567 = n4236 & ~n33316 ;
  assign n45568 = n12648 & n45567 ;
  assign n45569 = n45568 ^ n26865 ^ n4434 ;
  assign n45570 = ( ~n15881 & n28537 ) | ( ~n15881 & n45569 ) | ( n28537 & n45569 ) ;
  assign n45571 = ( ~n13908 & n18962 ) | ( ~n13908 & n24642 ) | ( n18962 & n24642 ) ;
  assign n45572 = ( ~n24282 & n35732 ) | ( ~n24282 & n36456 ) | ( n35732 & n36456 ) ;
  assign n45573 = ( n42754 & n45571 ) | ( n42754 & n45572 ) | ( n45571 & n45572 ) ;
  assign n45574 = n28345 ^ n22302 ^ n19618 ;
  assign n45575 = n45574 ^ n24821 ^ n24033 ;
  assign n45576 = n1543 & ~n45575 ;
  assign n45577 = ( n5249 & n8584 ) | ( n5249 & n21871 ) | ( n8584 & n21871 ) ;
  assign n45578 = n45577 ^ n33861 ^ 1'b0 ;
  assign n45579 = n22225 ^ n11237 ^ n5351 ;
  assign n45580 = n45579 ^ n36884 ^ n5949 ;
  assign n45581 = n45580 ^ n11528 ^ n2423 ;
  assign n45582 = ~n3619 & n22461 ;
  assign n45583 = n45582 ^ n1318 ^ 1'b0 ;
  assign n45584 = ( n7741 & n8306 ) | ( n7741 & n45583 ) | ( n8306 & n45583 ) ;
  assign n45585 = n45584 ^ n25161 ^ n24016 ;
  assign n45586 = n45585 ^ n20432 ^ 1'b0 ;
  assign n45587 = n22992 ^ n21881 ^ n5044 ;
  assign n45588 = n45587 ^ n13493 ^ n4640 ;
  assign n45589 = ( n2792 & n11703 ) | ( n2792 & ~n45588 ) | ( n11703 & ~n45588 ) ;
  assign n45590 = ( ~n2744 & n21166 ) | ( ~n2744 & n45589 ) | ( n21166 & n45589 ) ;
  assign n45591 = ( ~n7764 & n16306 ) | ( ~n7764 & n45590 ) | ( n16306 & n45590 ) ;
  assign n45592 = n33773 ^ n29739 ^ 1'b0 ;
  assign n45593 = ~n15898 & n45592 ;
  assign n45594 = n14453 | n24325 ;
  assign n45595 = n18121 & ~n45594 ;
  assign n45596 = n45595 ^ n10657 ^ n3663 ;
  assign n45597 = n10301 ^ n2233 ^ 1'b0 ;
  assign n45598 = ( n662 & n10301 ) | ( n662 & n45597 ) | ( n10301 & n45597 ) ;
  assign n45599 = n45598 ^ n24727 ^ n4740 ;
  assign n45600 = n45599 ^ n22802 ^ n9560 ;
  assign n45601 = n45600 ^ n24284 ^ n14973 ;
  assign n45602 = n45601 ^ n41594 ^ n41538 ;
  assign n45603 = ( n12869 & ~n17430 ) | ( n12869 & n45602 ) | ( ~n17430 & n45602 ) ;
  assign n45604 = n9280 ^ n5914 ^ n1078 ;
  assign n45605 = n45604 ^ n30171 ^ n26593 ;
  assign n45606 = n26493 ^ n19806 ^ n15262 ;
  assign n45607 = n11374 ^ n5737 ^ 1'b0 ;
  assign n45608 = ~n1112 & n45607 ;
  assign n45609 = ~n15685 & n40834 ;
  assign n45610 = n45608 | n45609 ;
  assign n45611 = n41907 ^ n41228 ^ n27669 ;
  assign n45612 = n45611 ^ n36249 ^ n32523 ;
  assign n45613 = n1349 | n17208 ;
  assign n45614 = n45613 ^ n42664 ^ n37895 ;
  assign n45620 = n24965 ^ n7572 ^ n2627 ;
  assign n45615 = n1356 & ~n4852 ;
  assign n45616 = n45615 ^ n9035 ^ 1'b0 ;
  assign n45617 = n11451 & n32549 ;
  assign n45618 = n45617 ^ n34355 ^ 1'b0 ;
  assign n45619 = ( ~n31516 & n45616 ) | ( ~n31516 & n45618 ) | ( n45616 & n45618 ) ;
  assign n45621 = n45620 ^ n45619 ^ 1'b0 ;
  assign n45622 = n4356 | n33253 ;
  assign n45623 = n3320 | n45622 ;
  assign n45624 = ( ~n13632 & n25222 ) | ( ~n13632 & n45318 ) | ( n25222 & n45318 ) ;
  assign n45625 = ( n8976 & n40709 ) | ( n8976 & ~n45624 ) | ( n40709 & ~n45624 ) ;
  assign n45629 = ( n1665 & ~n8903 ) | ( n1665 & n10717 ) | ( ~n8903 & n10717 ) ;
  assign n45626 = ( n2328 & n5631 ) | ( n2328 & n24179 ) | ( n5631 & n24179 ) ;
  assign n45627 = n45626 ^ n29568 ^ n1171 ;
  assign n45628 = ( ~n27224 & n29179 ) | ( ~n27224 & n45627 ) | ( n29179 & n45627 ) ;
  assign n45630 = n45629 ^ n45628 ^ n41500 ;
  assign n45631 = ( n9451 & ~n33857 ) | ( n9451 & n42634 ) | ( ~n33857 & n42634 ) ;
  assign n45632 = ( ~n15808 & n45630 ) | ( ~n15808 & n45631 ) | ( n45630 & n45631 ) ;
  assign n45633 = ( n34480 & n42098 ) | ( n34480 & ~n45618 ) | ( n42098 & ~n45618 ) ;
  assign n45634 = n45401 ^ n23446 ^ 1'b0 ;
  assign n45635 = n45634 ^ n15430 ^ n427 ;
  assign n45636 = ~n28061 & n45635 ;
  assign n45637 = n45636 ^ n38754 ^ n16099 ;
  assign n45638 = ( ~n10675 & n37136 ) | ( ~n10675 & n45520 ) | ( n37136 & n45520 ) ;
  assign n45642 = ( n13602 & n25316 ) | ( n13602 & ~n31229 ) | ( n25316 & ~n31229 ) ;
  assign n45640 = n548 | n21320 ;
  assign n45641 = n45640 ^ n5025 ^ 1'b0 ;
  assign n45639 = n40131 ^ n16850 ^ n12607 ;
  assign n45643 = n45642 ^ n45641 ^ n45639 ;
  assign n45644 = ( n11655 & ~n22766 ) | ( n11655 & n45643 ) | ( ~n22766 & n45643 ) ;
  assign n45645 = ( ~n10910 & n16738 ) | ( ~n10910 & n17052 ) | ( n16738 & n17052 ) ;
  assign n45646 = ( n15708 & ~n35966 ) | ( n15708 & n45645 ) | ( ~n35966 & n45645 ) ;
  assign n45647 = n26363 | n33449 ;
  assign n45648 = n13481 & ~n17377 ;
  assign n45649 = n15879 & n45648 ;
  assign n45650 = ( n17610 & n36221 ) | ( n17610 & n45649 ) | ( n36221 & n45649 ) ;
  assign n45651 = ( n6785 & ~n11507 ) | ( n6785 & n19675 ) | ( ~n11507 & n19675 ) ;
  assign n45652 = ( n20272 & n45650 ) | ( n20272 & n45651 ) | ( n45650 & n45651 ) ;
  assign n45653 = ( n4099 & n27003 ) | ( n4099 & ~n31025 ) | ( n27003 & ~n31025 ) ;
  assign n45654 = n45653 ^ n26914 ^ n15533 ;
  assign n45655 = n30364 ^ n1760 ^ 1'b0 ;
  assign n45656 = n27556 ^ n23682 ^ n21734 ;
  assign n45657 = ( ~n31937 & n38917 ) | ( ~n31937 & n45656 ) | ( n38917 & n45656 ) ;
  assign n45658 = n45657 ^ n29857 ^ n1686 ;
  assign n45659 = ( n2193 & n17584 ) | ( n2193 & n45658 ) | ( n17584 & n45658 ) ;
  assign n45660 = ( n16548 & ~n18390 ) | ( n16548 & n21797 ) | ( ~n18390 & n21797 ) ;
  assign n45661 = ( ~n9219 & n19983 ) | ( ~n9219 & n43708 ) | ( n19983 & n43708 ) ;
  assign n45663 = n25234 ^ n11563 ^ n2068 ;
  assign n45662 = n17337 ^ n15678 ^ 1'b0 ;
  assign n45664 = n45663 ^ n45662 ^ n365 ;
  assign n45665 = ( n980 & n2833 ) | ( n980 & n11645 ) | ( n2833 & n11645 ) ;
  assign n45666 = n2139 & ~n45665 ;
  assign n45667 = n45664 & n45666 ;
  assign n45668 = ( n7937 & n19721 ) | ( n7937 & n37009 ) | ( n19721 & n37009 ) ;
  assign n45669 = n29179 ^ n688 ^ x225 ;
  assign n45670 = n45668 | n45669 ;
  assign n45675 = n29162 ^ n26949 ^ n843 ;
  assign n45671 = ( n1818 & n10422 ) | ( n1818 & n27660 ) | ( n10422 & n27660 ) ;
  assign n45672 = n18903 ^ n1154 ^ 1'b0 ;
  assign n45673 = n45671 | n45672 ;
  assign n45674 = ( n11590 & ~n35422 ) | ( n11590 & n45673 ) | ( ~n35422 & n45673 ) ;
  assign n45676 = n45675 ^ n45674 ^ n5201 ;
  assign n45677 = ( ~n2784 & n7608 ) | ( ~n2784 & n9359 ) | ( n7608 & n9359 ) ;
  assign n45678 = n5140 ^ n2039 ^ 1'b0 ;
  assign n45679 = ( n23268 & n45677 ) | ( n23268 & ~n45678 ) | ( n45677 & ~n45678 ) ;
  assign n45680 = ( n16208 & n24043 ) | ( n16208 & n45679 ) | ( n24043 & n45679 ) ;
  assign n45681 = n7277 | n7593 ;
  assign n45682 = ( ~n2985 & n4464 ) | ( ~n2985 & n24467 ) | ( n4464 & n24467 ) ;
  assign n45683 = ( ~n5917 & n9710 ) | ( ~n5917 & n32999 ) | ( n9710 & n32999 ) ;
  assign n45684 = n22808 ^ n4648 ^ 1'b0 ;
  assign n45685 = n17689 ^ n4266 ^ 1'b0 ;
  assign n45686 = ~n42728 & n45685 ;
  assign n45687 = ( n1803 & ~n2319 ) | ( n1803 & n19276 ) | ( ~n2319 & n19276 ) ;
  assign n45688 = n20344 | n45687 ;
  assign n45689 = ~n20014 & n45688 ;
  assign n45690 = ( n21997 & n25148 ) | ( n21997 & ~n26769 ) | ( n25148 & ~n26769 ) ;
  assign n45691 = ( n9926 & ~n31062 ) | ( n9926 & n45690 ) | ( ~n31062 & n45690 ) ;
  assign n45692 = n23514 ^ n10068 ^ n4520 ;
  assign n45693 = n45692 ^ n31158 ^ n4402 ;
  assign n45700 = n22714 ^ n14098 ^ n13212 ;
  assign n45698 = ~n12247 & n29213 ;
  assign n45699 = n12852 & n45698 ;
  assign n45694 = n4588 ^ n1315 ^ 1'b0 ;
  assign n45695 = n16094 & n45694 ;
  assign n45696 = n45695 ^ n30220 ^ n10094 ;
  assign n45697 = n45696 ^ n17823 ^ n11695 ;
  assign n45701 = n45700 ^ n45699 ^ n45697 ;
  assign n45704 = n16442 ^ n4677 ^ 1'b0 ;
  assign n45705 = ~n21665 & n45704 ;
  assign n45706 = n38357 & n45705 ;
  assign n45707 = ~n21938 & n45706 ;
  assign n45702 = n43738 ^ n25145 ^ n3579 ;
  assign n45703 = n45702 ^ n40382 ^ n12505 ;
  assign n45708 = n45707 ^ n45703 ^ n29992 ;
  assign n45709 = n21144 ^ n13164 ^ n1496 ;
  assign n45710 = n18994 ^ n8628 ^ n4593 ;
  assign n45711 = n30129 | n45710 ;
  assign n45712 = n24817 ^ n13993 ^ 1'b0 ;
  assign n45713 = n2765 | n45712 ;
  assign n45714 = ( ~n45709 & n45711 ) | ( ~n45709 & n45713 ) | ( n45711 & n45713 ) ;
  assign n45716 = n34510 ^ n14540 ^ n7537 ;
  assign n45715 = n44844 ^ n20480 ^ n11347 ;
  assign n45717 = n45716 ^ n45715 ^ n4445 ;
  assign n45718 = ( n18749 & ~n29695 ) | ( n18749 & n45717 ) | ( ~n29695 & n45717 ) ;
  assign n45719 = n9779 ^ n7251 ^ 1'b0 ;
  assign n45720 = n45719 ^ n35337 ^ n6972 ;
  assign n45721 = ( n1804 & n6589 ) | ( n1804 & n13400 ) | ( n6589 & n13400 ) ;
  assign n45722 = n45721 ^ n24984 ^ n10614 ;
  assign n45723 = n40805 ^ n26684 ^ 1'b0 ;
  assign n45724 = n32580 & n45723 ;
  assign n45725 = n39533 ^ n25387 ^ n682 ;
  assign n45726 = ( n8881 & ~n45724 ) | ( n8881 & n45725 ) | ( ~n45724 & n45725 ) ;
  assign n45727 = n42031 ^ n19501 ^ 1'b0 ;
  assign n45728 = ( n13578 & ~n43770 ) | ( n13578 & n45727 ) | ( ~n43770 & n45727 ) ;
  assign n45730 = n9323 ^ n8196 ^ n8181 ;
  assign n45729 = n15012 & ~n15440 ;
  assign n45731 = n45730 ^ n45729 ^ 1'b0 ;
  assign n45732 = ( n36054 & n43485 ) | ( n36054 & n45731 ) | ( n43485 & n45731 ) ;
  assign n45733 = ( n4151 & ~n16842 ) | ( n4151 & n44732 ) | ( ~n16842 & n44732 ) ;
  assign n45734 = n18076 & n35157 ;
  assign n45735 = n45734 ^ n38497 ^ 1'b0 ;
  assign n45736 = ( ~n45732 & n45733 ) | ( ~n45732 & n45735 ) | ( n45733 & n45735 ) ;
  assign n45737 = n27529 ^ n24760 ^ 1'b0 ;
  assign n45738 = n28541 & ~n32225 ;
  assign n45739 = n45738 ^ n6135 ^ 1'b0 ;
  assign n45740 = ( n13729 & n15311 ) | ( n13729 & ~n24015 ) | ( n15311 & ~n24015 ) ;
  assign n45741 = n4496 ^ n1262 ^ n904 ;
  assign n45742 = ( n29212 & n45740 ) | ( n29212 & n45741 ) | ( n45740 & n45741 ) ;
  assign n45743 = n21680 ^ n11834 ^ n8323 ;
  assign n45744 = n32131 ^ n2545 ^ n324 ;
  assign n45745 = ( n5184 & ~n10310 ) | ( n5184 & n45744 ) | ( ~n10310 & n45744 ) ;
  assign n45746 = ( n7218 & n45743 ) | ( n7218 & n45745 ) | ( n45743 & n45745 ) ;
  assign n45747 = n45746 ^ n36158 ^ n35784 ;
  assign n45748 = n20847 ^ n9147 ^ n3616 ;
  assign n45753 = n1268 & ~n18752 ;
  assign n45750 = ( n16227 & n30848 ) | ( n16227 & ~n33780 ) | ( n30848 & ~n33780 ) ;
  assign n45751 = n45750 ^ n7628 ^ n894 ;
  assign n45752 = n45751 ^ n40977 ^ n19393 ;
  assign n45749 = ( n15631 & ~n27795 ) | ( n15631 & n28413 ) | ( ~n27795 & n28413 ) ;
  assign n45754 = n45753 ^ n45752 ^ n45749 ;
  assign n45755 = ( ~n4209 & n8856 ) | ( ~n4209 & n12792 ) | ( n8856 & n12792 ) ;
  assign n45756 = ( ~n21403 & n24544 ) | ( ~n21403 & n39936 ) | ( n24544 & n39936 ) ;
  assign n45757 = n29036 ^ n6922 ^ n439 ;
  assign n45758 = ( n10969 & n26702 ) | ( n10969 & n45757 ) | ( n26702 & n45757 ) ;
  assign n45759 = n16310 & n30916 ;
  assign n45760 = ( n8880 & n21837 ) | ( n8880 & n45759 ) | ( n21837 & n45759 ) ;
  assign n45761 = n38090 ^ n20289 ^ n13440 ;
  assign n45762 = ( n1683 & n37639 ) | ( n1683 & ~n45761 ) | ( n37639 & ~n45761 ) ;
  assign n45763 = n45762 ^ n28890 ^ n11725 ;
  assign n45764 = n32391 ^ n20722 ^ n9708 ;
  assign n45765 = n45764 ^ n524 ^ 1'b0 ;
  assign n45766 = ~n9270 & n29964 ;
  assign n45767 = n45766 ^ n12654 ^ 1'b0 ;
  assign n45768 = n39626 | n45767 ;
  assign n45769 = n45768 ^ n19393 ^ 1'b0 ;
  assign n45770 = n45769 ^ n10784 ^ n5206 ;
  assign n45772 = n2601 | n4433 ;
  assign n45773 = n45772 ^ n16535 ^ 1'b0 ;
  assign n45771 = n27425 ^ n11546 ^ n7556 ;
  assign n45774 = n45773 ^ n45771 ^ n27489 ;
  assign n45775 = ~n3084 & n45774 ;
  assign n45776 = n23145 & ~n35288 ;
  assign n45777 = ~n42098 & n45776 ;
  assign n45778 = n33825 ^ n9015 ^ n7995 ;
  assign n45779 = n45778 ^ n38850 ^ 1'b0 ;
  assign n45780 = ~n45777 & n45779 ;
  assign n45782 = n8523 ^ n2498 ^ n719 ;
  assign n45781 = n34241 ^ n29462 ^ n25714 ;
  assign n45783 = n45782 ^ n45781 ^ n30161 ;
  assign n45784 = ( n7715 & ~n11013 ) | ( n7715 & n23079 ) | ( ~n11013 & n23079 ) ;
  assign n45785 = n11311 | n34350 ;
  assign n45786 = n31982 & ~n45785 ;
  assign n45787 = ( n1053 & ~n18888 ) | ( n1053 & n26701 ) | ( ~n18888 & n26701 ) ;
  assign n45788 = n45602 ^ n37327 ^ n30902 ;
  assign n45790 = ( ~n3194 & n20961 ) | ( ~n3194 & n30317 ) | ( n20961 & n30317 ) ;
  assign n45789 = ( n11274 & n13370 ) | ( n11274 & ~n24936 ) | ( n13370 & ~n24936 ) ;
  assign n45791 = n45790 ^ n45789 ^ n9970 ;
  assign n45792 = n45791 ^ n17284 ^ n10498 ;
  assign n45793 = n25749 ^ n10673 ^ 1'b0 ;
  assign n45794 = ( ~n13369 & n17942 ) | ( ~n13369 & n31382 ) | ( n17942 & n31382 ) ;
  assign n45795 = ( n685 & n2597 ) | ( n685 & n26701 ) | ( n2597 & n26701 ) ;
  assign n45796 = n45795 ^ n36290 ^ 1'b0 ;
  assign n45797 = n45796 ^ n28230 ^ n24360 ;
  assign n45798 = n3925 & ~n6489 ;
  assign n45799 = ~n27770 & n41708 ;
  assign n45800 = n45056 ^ n3456 ^ 1'b0 ;
  assign n45801 = ~n21482 & n45800 ;
  assign n45802 = ( n5025 & ~n45799 ) | ( n5025 & n45801 ) | ( ~n45799 & n45801 ) ;
  assign n45803 = n16155 ^ n15286 ^ n402 ;
  assign n45804 = n39516 ^ n29212 ^ n8201 ;
  assign n45805 = n23287 ^ n12667 ^ 1'b0 ;
  assign n45806 = ( n45803 & ~n45804 ) | ( n45803 & n45805 ) | ( ~n45804 & n45805 ) ;
  assign n45807 = ( n11500 & n23651 ) | ( n11500 & n27789 ) | ( n23651 & n27789 ) ;
  assign n45808 = n45807 ^ n37676 ^ n31015 ;
  assign n45809 = ( n6780 & n34848 ) | ( n6780 & n45808 ) | ( n34848 & n45808 ) ;
  assign n45810 = ( n18251 & ~n23505 ) | ( n18251 & n29362 ) | ( ~n23505 & n29362 ) ;
  assign n45811 = n35223 ^ n25081 ^ n24820 ;
  assign n45812 = n45811 ^ n41586 ^ n20329 ;
  assign n45813 = n3828 & ~n8477 ;
  assign n45814 = n45813 ^ n24206 ^ n17877 ;
  assign n45815 = ( n2926 & ~n45812 ) | ( n2926 & n45814 ) | ( ~n45812 & n45814 ) ;
  assign n45816 = ( n7325 & n14000 ) | ( n7325 & ~n22885 ) | ( n14000 & ~n22885 ) ;
  assign n45817 = ( n5536 & ~n6602 ) | ( n5536 & n10826 ) | ( ~n6602 & n10826 ) ;
  assign n45818 = n16016 ^ n14381 ^ x3 ;
  assign n45819 = n802 & n5922 ;
  assign n45820 = n45819 ^ n2880 ^ 1'b0 ;
  assign n45821 = ( n6287 & ~n35065 ) | ( n6287 & n45820 ) | ( ~n35065 & n45820 ) ;
  assign n45822 = n9200 ^ n1813 ^ n552 ;
  assign n45824 = n30092 ^ n13850 ^ n7771 ;
  assign n45823 = n39641 ^ n38756 ^ n8472 ;
  assign n45825 = n45824 ^ n45823 ^ n13004 ;
  assign n45826 = ( n1111 & n45822 ) | ( n1111 & n45825 ) | ( n45822 & n45825 ) ;
  assign n45827 = n43065 ^ n39200 ^ n11802 ;
  assign n45828 = n37169 ^ n21497 ^ n18897 ;
  assign n45829 = x8 & ~n45828 ;
  assign n45830 = n40311 ^ n33750 ^ n2761 ;
  assign n45831 = n14345 & ~n45830 ;
  assign n45832 = ~n13113 & n45831 ;
  assign n45833 = n43742 ^ n35423 ^ n14126 ;
  assign n45834 = n45833 ^ n18371 ^ 1'b0 ;
  assign n45835 = n25543 ^ n17414 ^ n7944 ;
  assign n45836 = ~n4317 & n33015 ;
  assign n45837 = n41765 ^ n35389 ^ n32219 ;
  assign n45838 = n8821 & ~n17963 ;
  assign n45839 = n19226 | n45838 ;
  assign n45840 = x227 | n45839 ;
  assign n45841 = ( n6737 & ~n14483 ) | ( n6737 & n45840 ) | ( ~n14483 & n45840 ) ;
  assign n45842 = ( ~n14362 & n17052 ) | ( ~n14362 & n38403 ) | ( n17052 & n38403 ) ;
  assign n45843 = n23074 ^ n9167 ^ n2855 ;
  assign n45844 = ( n6018 & n12266 ) | ( n6018 & n45843 ) | ( n12266 & n45843 ) ;
  assign n45848 = n35868 ^ n29560 ^ n23770 ;
  assign n45845 = n32529 ^ n18076 ^ n1848 ;
  assign n45846 = ~n26157 & n45845 ;
  assign n45847 = n13035 & n45846 ;
  assign n45849 = n45848 ^ n45847 ^ n29288 ;
  assign n45850 = ( n4390 & n15060 ) | ( n4390 & n32542 ) | ( n15060 & n32542 ) ;
  assign n45851 = n18199 ^ n10865 ^ x89 ;
  assign n45852 = ( n17181 & n20957 ) | ( n17181 & n45851 ) | ( n20957 & n45851 ) ;
  assign n45853 = n40101 ^ n40019 ^ n3983 ;
  assign n45854 = n45853 ^ n17907 ^ n2080 ;
  assign n45855 = n45852 & ~n45854 ;
  assign n45856 = n45855 ^ n28601 ^ 1'b0 ;
  assign n45857 = ( n9654 & n13180 ) | ( n9654 & ~n45856 ) | ( n13180 & ~n45856 ) ;
  assign n45858 = n45857 ^ n40207 ^ n29366 ;
  assign n45859 = n44022 & n45858 ;
  assign n45860 = ~n10548 & n45859 ;
  assign n45861 = ( n13694 & n16895 ) | ( n13694 & n17931 ) | ( n16895 & n17931 ) ;
  assign n45862 = n45861 ^ n17111 ^ n7078 ;
  assign n45863 = ( ~n7170 & n38200 ) | ( ~n7170 & n45862 ) | ( n38200 & n45862 ) ;
  assign n45864 = n21220 ^ n6018 ^ 1'b0 ;
  assign n45865 = n45864 ^ n19762 ^ 1'b0 ;
  assign n45866 = n45865 ^ n44499 ^ n41821 ;
  assign n45867 = ( n29825 & ~n33971 ) | ( n29825 & n45866 ) | ( ~n33971 & n45866 ) ;
  assign n45872 = n38436 ^ n17738 ^ n14948 ;
  assign n45868 = ( n14616 & ~n20508 ) | ( n14616 & n34552 ) | ( ~n20508 & n34552 ) ;
  assign n45869 = n15923 ^ n11279 ^ n5723 ;
  assign n45870 = ( n28915 & n45868 ) | ( n28915 & n45869 ) | ( n45868 & n45869 ) ;
  assign n45871 = n45870 ^ n28845 ^ n7978 ;
  assign n45873 = n45872 ^ n45871 ^ n37394 ;
  assign n45874 = n22312 ^ n13528 ^ n4364 ;
  assign n45875 = n25547 ^ n15128 ^ n2765 ;
  assign n45876 = ( ~n1284 & n8558 ) | ( ~n1284 & n44610 ) | ( n8558 & n44610 ) ;
  assign n45877 = n26666 ^ n11667 ^ n2949 ;
  assign n45878 = n45877 ^ n32598 ^ n15801 ;
  assign n45879 = ( n45875 & n45876 ) | ( n45875 & ~n45878 ) | ( n45876 & ~n45878 ) ;
  assign n45880 = n21242 & ~n34018 ;
  assign n45881 = n45880 ^ n6532 ^ 1'b0 ;
  assign n45882 = n7740 & n30961 ;
  assign n45883 = ~n45881 & n45882 ;
  assign n45884 = n13116 ^ n13044 ^ 1'b0 ;
  assign n45889 = n39733 ^ n31822 ^ n7442 ;
  assign n45886 = n12360 ^ n10991 ^ n4277 ;
  assign n45885 = ( n8706 & n13843 ) | ( n8706 & ~n17848 ) | ( n13843 & ~n17848 ) ;
  assign n45887 = n45886 ^ n45885 ^ n18936 ;
  assign n45888 = n45887 ^ n34917 ^ n32664 ;
  assign n45890 = n45889 ^ n45888 ^ n2748 ;
  assign n45891 = n45890 ^ n35714 ^ n14937 ;
  assign n45892 = n45891 ^ n20309 ^ n10277 ;
  assign n45893 = n4290 & ~n34435 ;
  assign n45894 = ( n25840 & n38852 ) | ( n25840 & ~n45893 ) | ( n38852 & ~n45893 ) ;
  assign n45895 = n45894 ^ n30917 ^ n28877 ;
  assign n45896 = ( n2044 & n3207 ) | ( n2044 & n7667 ) | ( n3207 & n7667 ) ;
  assign n45897 = ( x221 & n22591 ) | ( x221 & ~n45896 ) | ( n22591 & ~n45896 ) ;
  assign n45898 = n21193 ^ n16861 ^ n1481 ;
  assign n45899 = ( n19985 & ~n38945 ) | ( n19985 & n45898 ) | ( ~n38945 & n45898 ) ;
  assign n45900 = ( ~n17604 & n45897 ) | ( ~n17604 & n45899 ) | ( n45897 & n45899 ) ;
  assign n45901 = n11714 ^ n2246 ^ 1'b0 ;
  assign n45902 = n45901 ^ n33584 ^ n11692 ;
  assign n45903 = n4417 & ~n12929 ;
  assign n45904 = n29816 ^ n10127 ^ n3601 ;
  assign n45905 = n4468 ^ n427 ^ 1'b0 ;
  assign n45906 = n4458 & ~n45905 ;
  assign n45907 = n45710 ^ n25848 ^ n10233 ;
  assign n45908 = ( ~n7125 & n45906 ) | ( ~n7125 & n45907 ) | ( n45906 & n45907 ) ;
  assign n45909 = ( ~n4463 & n14231 ) | ( ~n4463 & n44409 ) | ( n14231 & n44409 ) ;
  assign n45910 = ~n14575 & n23721 ;
  assign n45911 = n1145 & n35058 ;
  assign n45912 = ~n7725 & n45911 ;
  assign n45913 = n45912 ^ n41354 ^ n31563 ;
  assign n45914 = n20740 ^ n15185 ^ n15170 ;
  assign n45915 = ( n6341 & ~n7853 ) | ( n6341 & n45914 ) | ( ~n7853 & n45914 ) ;
  assign n45916 = n45915 ^ n28838 ^ n22952 ;
  assign n45917 = ( n2381 & ~n10266 ) | ( n2381 & n40134 ) | ( ~n10266 & n40134 ) ;
  assign n45918 = n24168 | n45917 ;
  assign n45919 = n17155 & n25540 ;
  assign n45920 = n45919 ^ n6924 ^ 1'b0 ;
  assign n45921 = n17478 | n45920 ;
  assign n45922 = ( ~n12514 & n42240 ) | ( ~n12514 & n45921 ) | ( n42240 & n45921 ) ;
  assign n45923 = n41088 ^ n18709 ^ n10937 ;
  assign n45924 = ( ~n2310 & n6605 ) | ( ~n2310 & n38035 ) | ( n6605 & n38035 ) ;
  assign n45925 = ( n26864 & n31011 ) | ( n26864 & n34722 ) | ( n31011 & n34722 ) ;
  assign n45926 = n22400 & n45925 ;
  assign n45927 = n1341 & n45926 ;
  assign n45928 = ( n33800 & n45924 ) | ( n33800 & ~n45927 ) | ( n45924 & ~n45927 ) ;
  assign n45929 = ( n27918 & ~n33730 ) | ( n27918 & n45928 ) | ( ~n33730 & n45928 ) ;
  assign n45930 = ( n6115 & n6273 ) | ( n6115 & n12713 ) | ( n6273 & n12713 ) ;
  assign n45931 = n31699 ^ n21104 ^ n12360 ;
  assign n45932 = ( n12566 & n21883 ) | ( n12566 & n45931 ) | ( n21883 & n45931 ) ;
  assign n45933 = n45932 ^ n8878 ^ n5544 ;
  assign n45934 = n41912 ^ n10718 ^ 1'b0 ;
  assign n45935 = ( n45930 & n45933 ) | ( n45930 & ~n45934 ) | ( n45933 & ~n45934 ) ;
  assign n45936 = n38660 ^ n35850 ^ n21182 ;
  assign n45937 = ( n7702 & n14675 ) | ( n7702 & n25780 ) | ( n14675 & n25780 ) ;
  assign n45938 = n45937 ^ n8891 ^ n8254 ;
  assign n45939 = ( n9605 & n10857 ) | ( n9605 & ~n41709 ) | ( n10857 & ~n41709 ) ;
  assign n45940 = ( n15195 & n45938 ) | ( n15195 & n45939 ) | ( n45938 & n45939 ) ;
  assign n45941 = ( n5312 & n45936 ) | ( n5312 & ~n45940 ) | ( n45936 & ~n45940 ) ;
  assign n45942 = ( ~x108 & n659 ) | ( ~x108 & n45941 ) | ( n659 & n45941 ) ;
  assign n45943 = n20644 & n29766 ;
  assign n45944 = n42366 ^ n13136 ^ n4605 ;
  assign n45945 = n42229 ^ n39763 ^ n27553 ;
  assign n45946 = n12640 ^ n782 ^ n706 ;
  assign n45947 = n34621 ^ n22588 ^ n5731 ;
  assign n45948 = n20118 & ~n45947 ;
  assign n45949 = ( x109 & n14487 ) | ( x109 & n45948 ) | ( n14487 & n45948 ) ;
  assign n45950 = ( n5909 & n6382 ) | ( n5909 & ~n9280 ) | ( n6382 & ~n9280 ) ;
  assign n45951 = n45950 ^ n24459 ^ n14093 ;
  assign n45952 = ( n8506 & n13146 ) | ( n8506 & ~n23759 ) | ( n13146 & ~n23759 ) ;
  assign n45953 = n26757 & n33374 ;
  assign n45954 = ( n3067 & ~n36097 ) | ( n3067 & n45953 ) | ( ~n36097 & n45953 ) ;
  assign n45955 = n26643 ^ n11341 ^ 1'b0 ;
  assign n45956 = ( n27413 & ~n42386 ) | ( n27413 & n45955 ) | ( ~n42386 & n45955 ) ;
  assign n45957 = ( n26843 & ~n43172 ) | ( n26843 & n45956 ) | ( ~n43172 & n45956 ) ;
  assign n45958 = n3813 & ~n17504 ;
  assign n45959 = n4012 & n45958 ;
  assign n45960 = n4246 | n7698 ;
  assign n45961 = n45959 & ~n45960 ;
  assign n45962 = n45961 ^ n20238 ^ n3185 ;
  assign n45964 = n42067 ^ n30375 ^ n3537 ;
  assign n45963 = n39796 & ~n39990 ;
  assign n45965 = n45964 ^ n45963 ^ 1'b0 ;
  assign n45966 = n26550 ^ n11614 ^ x174 ;
  assign n45967 = ( n2064 & ~n7078 ) | ( n2064 & n25970 ) | ( ~n7078 & n25970 ) ;
  assign n45968 = n45967 ^ n15152 ^ n8701 ;
  assign n45969 = ( ~n32140 & n39268 ) | ( ~n32140 & n45968 ) | ( n39268 & n45968 ) ;
  assign n45970 = ( ~n13240 & n35510 ) | ( ~n13240 & n45969 ) | ( n35510 & n45969 ) ;
  assign n45971 = ( n452 & ~n8708 ) | ( n452 & n45803 ) | ( ~n8708 & n45803 ) ;
  assign n45972 = n18954 ^ n12798 ^ n10101 ;
  assign n45973 = n45972 ^ n16090 ^ n401 ;
  assign n45974 = ( n1076 & n28550 ) | ( n1076 & n44177 ) | ( n28550 & n44177 ) ;
  assign n45975 = n11589 ^ n6477 ^ n1193 ;
  assign n45976 = ( n1172 & ~n4663 ) | ( n1172 & n45975 ) | ( ~n4663 & n45975 ) ;
  assign n45977 = ( n8040 & n31475 ) | ( n8040 & ~n38220 ) | ( n31475 & ~n38220 ) ;
  assign n45978 = ( n11405 & ~n45976 ) | ( n11405 & n45977 ) | ( ~n45976 & n45977 ) ;
  assign n45979 = ( n32163 & n45974 ) | ( n32163 & n45978 ) | ( n45974 & n45978 ) ;
  assign n45980 = n18051 ^ n3235 ^ n3198 ;
  assign n45981 = n45980 ^ n26933 ^ n8157 ;
  assign n45982 = n28639 ^ n27976 ^ n2184 ;
  assign n45983 = n7629 ^ n1153 ^ 1'b0 ;
  assign n45984 = n26729 & ~n45983 ;
  assign n45985 = ( n732 & n24922 ) | ( n732 & ~n31545 ) | ( n24922 & ~n31545 ) ;
  assign n45986 = n5050 | n43960 ;
  assign n45987 = n45985 & ~n45986 ;
  assign n45988 = n42891 ^ n25208 ^ n7546 ;
  assign n45989 = ( ~n930 & n25226 ) | ( ~n930 & n45988 ) | ( n25226 & n45988 ) ;
  assign n45990 = n19752 ^ n17043 ^ n15695 ;
  assign n45991 = n45989 & ~n45990 ;
  assign n45992 = ( n22895 & n42023 ) | ( n22895 & ~n45991 ) | ( n42023 & ~n45991 ) ;
  assign n45993 = n7566 & ~n45992 ;
  assign n45994 = ( ~n14276 & n16919 ) | ( ~n14276 & n40628 ) | ( n16919 & n40628 ) ;
  assign n45996 = ( n1428 & n4231 ) | ( n1428 & ~n37513 ) | ( n4231 & ~n37513 ) ;
  assign n45995 = n27240 ^ n22263 ^ 1'b0 ;
  assign n45997 = n45996 ^ n45995 ^ n11008 ;
  assign n45998 = n45997 ^ n42909 ^ n9090 ;
  assign n45999 = ( n2413 & n10253 ) | ( n2413 & n45705 ) | ( n10253 & n45705 ) ;
  assign n46000 = n16135 ^ n2029 ^ 1'b0 ;
  assign n46001 = ~n45999 & n46000 ;
  assign n46002 = ( ~n20031 & n37474 ) | ( ~n20031 & n46001 ) | ( n37474 & n46001 ) ;
  assign n46003 = n34810 ^ n22098 ^ n9199 ;
  assign n46004 = ( n6350 & n15665 ) | ( n6350 & n46003 ) | ( n15665 & n46003 ) ;
  assign n46005 = n44501 ^ n37671 ^ n24985 ;
  assign n46010 = n38974 ^ n22395 ^ x143 ;
  assign n46011 = ( ~n25170 & n32841 ) | ( ~n25170 & n46010 ) | ( n32841 & n46010 ) ;
  assign n46009 = n4981 & n6366 ;
  assign n46006 = n1594 ^ n1583 ^ x234 ;
  assign n46007 = n36286 ^ n2561 ^ n867 ;
  assign n46008 = ( n7196 & n46006 ) | ( n7196 & ~n46007 ) | ( n46006 & ~n46007 ) ;
  assign n46012 = n46011 ^ n46009 ^ n46008 ;
  assign n46013 = n45508 ^ n29829 ^ n3949 ;
  assign n46014 = n11770 ^ n7960 ^ 1'b0 ;
  assign n46015 = n36086 ^ n25408 ^ n9801 ;
  assign n46016 = n34031 ^ n13887 ^ n8265 ;
  assign n46017 = ( n20226 & n24498 ) | ( n20226 & ~n46016 ) | ( n24498 & ~n46016 ) ;
  assign n46018 = ( n13837 & ~n27568 ) | ( n13837 & n46017 ) | ( ~n27568 & n46017 ) ;
  assign n46019 = n28038 ^ n19660 ^ n2405 ;
  assign n46021 = ( ~n14244 & n17941 ) | ( ~n14244 & n31546 ) | ( n17941 & n31546 ) ;
  assign n46020 = n2480 | n37555 ;
  assign n46022 = n46021 ^ n46020 ^ n1489 ;
  assign n46023 = ( n11758 & ~n41749 ) | ( n11758 & n46022 ) | ( ~n41749 & n46022 ) ;
  assign n46024 = ( n10326 & n19562 ) | ( n10326 & ~n46023 ) | ( n19562 & ~n46023 ) ;
  assign n46025 = ( n5859 & n9204 ) | ( n5859 & ~n22968 ) | ( n9204 & ~n22968 ) ;
  assign n46026 = ( n19035 & n25539 ) | ( n19035 & ~n42403 ) | ( n25539 & ~n42403 ) ;
  assign n46027 = n947 & ~n36368 ;
  assign n46029 = n20958 & ~n23409 ;
  assign n46030 = ~n19491 & n46029 ;
  assign n46031 = n46030 ^ n29389 ^ n901 ;
  assign n46028 = n12973 | n27986 ;
  assign n46032 = n46031 ^ n46028 ^ 1'b0 ;
  assign n46035 = n22996 ^ n4952 ^ n4922 ;
  assign n46033 = n40169 ^ n5317 ^ 1'b0 ;
  assign n46034 = n46033 ^ n40255 ^ 1'b0 ;
  assign n46036 = n46035 ^ n46034 ^ n20602 ;
  assign n46037 = ~n2840 & n29749 ;
  assign n46038 = n31418 ^ n18483 ^ n16495 ;
  assign n46039 = n46038 ^ n31177 ^ n12278 ;
  assign n46040 = n28748 ^ n23259 ^ n21853 ;
  assign n46041 = n46040 ^ n39725 ^ n2704 ;
  assign n46042 = ( n8014 & ~n46039 ) | ( n8014 & n46041 ) | ( ~n46039 & n46041 ) ;
  assign n46043 = n28170 ^ n23523 ^ n10800 ;
  assign n46044 = n46043 ^ n30629 ^ n20400 ;
  assign n46045 = n25466 ^ n24501 ^ n5824 ;
  assign n46046 = n21735 ^ n19108 ^ 1'b0 ;
  assign n46047 = n18462 & ~n46046 ;
  assign n46048 = ~n45585 & n46047 ;
  assign n46049 = ( n28781 & n46045 ) | ( n28781 & n46048 ) | ( n46045 & n46048 ) ;
  assign n46050 = ( n18916 & ~n19434 ) | ( n18916 & n27976 ) | ( ~n19434 & n27976 ) ;
  assign n46051 = n30985 ^ n19169 ^ n2624 ;
  assign n46053 = ( n14724 & ~n28090 ) | ( n14724 & n29417 ) | ( ~n28090 & n29417 ) ;
  assign n46052 = n12232 ^ n4721 ^ n2180 ;
  assign n46054 = n46053 ^ n46052 ^ n37942 ;
  assign n46055 = n12452 & ~n43205 ;
  assign n46056 = ~n46054 & n46055 ;
  assign n46057 = n7191 ^ n3852 ^ 1'b0 ;
  assign n46058 = ( n2565 & n9697 ) | ( n2565 & ~n39163 ) | ( n9697 & ~n39163 ) ;
  assign n46059 = n14025 ^ n13909 ^ 1'b0 ;
  assign n46060 = n32812 & ~n46059 ;
  assign n46061 = n46060 ^ n5914 ^ 1'b0 ;
  assign n46062 = n37832 ^ n32294 ^ n10451 ;
  assign n46063 = n19084 ^ n18574 ^ 1'b0 ;
  assign n46064 = ( n10249 & n10587 ) | ( n10249 & n27669 ) | ( n10587 & n27669 ) ;
  assign n46065 = n46064 ^ n31144 ^ n4036 ;
  assign n46066 = ( n13904 & n40251 ) | ( n13904 & n46065 ) | ( n40251 & n46065 ) ;
  assign n46067 = n14261 ^ n6621 ^ 1'b0 ;
  assign n46068 = n46067 ^ n2134 ^ 1'b0 ;
  assign n46069 = n18965 & n46068 ;
  assign n46072 = n38616 ^ n25232 ^ n22161 ;
  assign n46073 = ( n43825 & n45086 ) | ( n43825 & n46072 ) | ( n45086 & n46072 ) ;
  assign n46070 = n15076 ^ n14242 ^ 1'b0 ;
  assign n46071 = n11282 & ~n46070 ;
  assign n46074 = n46073 ^ n46071 ^ n6367 ;
  assign n46075 = n46074 ^ n21618 ^ n17987 ;
  assign n46076 = ( n16291 & n22290 ) | ( n16291 & n39234 ) | ( n22290 & n39234 ) ;
  assign n46077 = ( ~n30371 & n34759 ) | ( ~n30371 & n46076 ) | ( n34759 & n46076 ) ;
  assign n46078 = n42955 ^ n19854 ^ n4435 ;
  assign n46079 = ( n5705 & ~n19258 ) | ( n5705 & n46078 ) | ( ~n19258 & n46078 ) ;
  assign n46084 = n13654 & ~n42341 ;
  assign n46080 = n21454 ^ n2858 ^ 1'b0 ;
  assign n46081 = n46080 ^ n40305 ^ n9542 ;
  assign n46082 = ( n5025 & n19162 ) | ( n5025 & n46081 ) | ( n19162 & n46081 ) ;
  assign n46083 = n46082 ^ n36508 ^ n36241 ;
  assign n46085 = n46084 ^ n46083 ^ 1'b0 ;
  assign n46087 = n26153 | n27810 ;
  assign n46086 = ( n16647 & n25225 ) | ( n16647 & n35188 ) | ( n25225 & n35188 ) ;
  assign n46088 = n46087 ^ n46086 ^ n15845 ;
  assign n46093 = ( n13123 & n15367 ) | ( n13123 & n30090 ) | ( n15367 & n30090 ) ;
  assign n46094 = n46093 ^ n22458 ^ n7313 ;
  assign n46090 = n7681 ^ n2538 ^ n481 ;
  assign n46091 = ( ~n3475 & n4892 ) | ( ~n3475 & n46090 ) | ( n4892 & n46090 ) ;
  assign n46092 = n46091 ^ n19076 ^ n14344 ;
  assign n46095 = n46094 ^ n46092 ^ n24649 ;
  assign n46089 = ( n9849 & n9855 ) | ( n9849 & ~n42736 ) | ( n9855 & ~n42736 ) ;
  assign n46096 = n46095 ^ n46089 ^ 1'b0 ;
  assign n46097 = ( n33405 & n39058 ) | ( n33405 & ~n46096 ) | ( n39058 & ~n46096 ) ;
  assign n46098 = n25006 ^ n23915 ^ n8709 ;
  assign n46099 = n32863 ^ n3604 ^ 1'b0 ;
  assign n46100 = n23478 | n39314 ;
  assign n46101 = n39297 | n46100 ;
  assign n46102 = ( n3771 & ~n4163 ) | ( n3771 & n13159 ) | ( ~n4163 & n13159 ) ;
  assign n46103 = n46102 ^ n20031 ^ n5918 ;
  assign n46104 = ( n35358 & n45499 ) | ( n35358 & ~n46103 ) | ( n45499 & ~n46103 ) ;
  assign n46105 = ( ~n30916 & n37115 ) | ( ~n30916 & n46104 ) | ( n37115 & n46104 ) ;
  assign n46106 = n32250 ^ n25853 ^ n972 ;
  assign n46107 = ( n7272 & n16222 ) | ( n7272 & n16718 ) | ( n16222 & n16718 ) ;
  assign n46108 = n46107 ^ n42172 ^ n16702 ;
  assign n46109 = ( n16656 & n25982 ) | ( n16656 & ~n43987 ) | ( n25982 & ~n43987 ) ;
  assign n46110 = n42590 ^ n16826 ^ 1'b0 ;
  assign n46111 = n46110 ^ n7066 ^ 1'b0 ;
  assign n46112 = n29883 ^ n6322 ^ n5438 ;
  assign n46113 = n16695 & n46112 ;
  assign n46114 = n46113 ^ n7358 ^ 1'b0 ;
  assign n46116 = n33508 ^ n283 ^ 1'b0 ;
  assign n46115 = ( n12153 & ~n14803 ) | ( n12153 & n39500 ) | ( ~n14803 & n39500 ) ;
  assign n46117 = n46116 ^ n46115 ^ 1'b0 ;
  assign n46118 = n14455 ^ n5813 ^ 1'b0 ;
  assign n46119 = ( n20593 & ~n33083 ) | ( n20593 & n46118 ) | ( ~n33083 & n46118 ) ;
  assign n46120 = n46119 ^ n38574 ^ n715 ;
  assign n46121 = n40195 ^ n14114 ^ n1751 ;
  assign n46123 = n20162 ^ n8897 ^ n5563 ;
  assign n46122 = ( n9905 & n14136 ) | ( n9905 & n43026 ) | ( n14136 & n43026 ) ;
  assign n46124 = n46123 ^ n46122 ^ n2331 ;
  assign n46132 = n9129 | n9717 ;
  assign n46133 = n17303 & ~n46132 ;
  assign n46125 = ( n5938 & n9044 ) | ( n5938 & ~n40734 ) | ( n9044 & ~n40734 ) ;
  assign n46128 = ( n7692 & n8773 ) | ( n7692 & n35433 ) | ( n8773 & n35433 ) ;
  assign n46127 = n35854 ^ n24828 ^ n2735 ;
  assign n46129 = n46128 ^ n46127 ^ n10068 ;
  assign n46126 = ~n4229 & n21590 ;
  assign n46130 = n46129 ^ n46126 ^ 1'b0 ;
  assign n46131 = ( n38019 & ~n46125 ) | ( n38019 & n46130 ) | ( ~n46125 & n46130 ) ;
  assign n46134 = n46133 ^ n46131 ^ n26894 ;
  assign n46135 = ( n10152 & n16520 ) | ( n10152 & ~n27307 ) | ( n16520 & ~n27307 ) ;
  assign n46136 = n10917 & ~n14817 ;
  assign n46137 = n46136 ^ n9855 ^ 1'b0 ;
  assign n46138 = n46137 ^ n34672 ^ n10963 ;
  assign n46139 = ( ~n946 & n46135 ) | ( ~n946 & n46138 ) | ( n46135 & n46138 ) ;
  assign n46140 = n14787 ^ n11450 ^ n10132 ;
  assign n46141 = n46140 ^ n39012 ^ n2880 ;
  assign n46142 = ( n7057 & ~n7463 ) | ( n7057 & n46141 ) | ( ~n7463 & n46141 ) ;
  assign n46143 = n12185 ^ n2840 ^ n1413 ;
  assign n46144 = n46143 ^ n17996 ^ n16335 ;
  assign n46145 = ( n6011 & ~n46142 ) | ( n6011 & n46144 ) | ( ~n46142 & n46144 ) ;
  assign n46146 = n46145 ^ n19948 ^ n3023 ;
  assign n46147 = ( n19683 & ~n27854 ) | ( n19683 & n39164 ) | ( ~n27854 & n39164 ) ;
  assign n46148 = n34529 ^ n23575 ^ n20215 ;
  assign n46149 = ( n694 & ~n7877 ) | ( n694 & n16504 ) | ( ~n7877 & n16504 ) ;
  assign n46150 = n46149 ^ n31236 ^ n13973 ;
  assign n46151 = ( n11159 & n20018 ) | ( n11159 & n27777 ) | ( n20018 & n27777 ) ;
  assign n46152 = n5276 ^ n4173 ^ n2004 ;
  assign n46153 = n43981 ^ n21893 ^ n19010 ;
  assign n46154 = ( n44020 & ~n46152 ) | ( n44020 & n46153 ) | ( ~n46152 & n46153 ) ;
  assign n46155 = n13780 ^ n2278 ^ 1'b0 ;
  assign n46156 = ~n16946 & n27852 ;
  assign n46157 = ~n17748 & n46156 ;
  assign n46158 = n31090 ^ n21752 ^ n5784 ;
  assign n46159 = ( ~n29612 & n29782 ) | ( ~n29612 & n46158 ) | ( n29782 & n46158 ) ;
  assign n46160 = ( ~n20198 & n46157 ) | ( ~n20198 & n46159 ) | ( n46157 & n46159 ) ;
  assign n46162 = ( n24506 & n33346 ) | ( n24506 & ~n33507 ) | ( n33346 & ~n33507 ) ;
  assign n46161 = n6978 & ~n22888 ;
  assign n46163 = n46162 ^ n46161 ^ 1'b0 ;
  assign n46164 = ~n23176 & n25231 ;
  assign n46165 = n34972 ^ n22473 ^ 1'b0 ;
  assign n46166 = ( n2592 & n35476 ) | ( n2592 & ~n39920 ) | ( n35476 & ~n39920 ) ;
  assign n46167 = n33101 ^ n3014 ^ n1595 ;
  assign n46168 = n46167 ^ n20305 ^ 1'b0 ;
  assign n46169 = n33257 ^ n12370 ^ n2855 ;
  assign n46170 = ( ~n6046 & n44891 ) | ( ~n6046 & n46169 ) | ( n44891 & n46169 ) ;
  assign n46173 = n15634 ^ n15176 ^ n14914 ;
  assign n46171 = ( n2035 & n12268 ) | ( n2035 & n18064 ) | ( n12268 & n18064 ) ;
  assign n46172 = n46171 ^ n24713 ^ n11169 ;
  assign n46174 = n46173 ^ n46172 ^ 1'b0 ;
  assign n46175 = ( n7292 & ~n46170 ) | ( n7292 & n46174 ) | ( ~n46170 & n46174 ) ;
  assign n46176 = n23238 ^ n9429 ^ n3088 ;
  assign n46177 = ( n10260 & n35518 ) | ( n10260 & n46176 ) | ( n35518 & n46176 ) ;
  assign n46178 = n46177 ^ n30761 ^ 1'b0 ;
  assign n46179 = ~n7730 & n26759 ;
  assign n46180 = n23023 & n46179 ;
  assign n46181 = n22058 | n43334 ;
  assign n46182 = n46181 ^ n36404 ^ 1'b0 ;
  assign n46187 = ( n8810 & ~n11981 ) | ( n8810 & n21514 ) | ( ~n11981 & n21514 ) ;
  assign n46185 = n18422 ^ n9604 ^ 1'b0 ;
  assign n46186 = n9483 & n46185 ;
  assign n46183 = n29737 ^ n15313 ^ n3162 ;
  assign n46184 = ( n28377 & n36181 ) | ( n28377 & ~n46183 ) | ( n36181 & ~n46183 ) ;
  assign n46188 = n46187 ^ n46186 ^ n46184 ;
  assign n46189 = n36154 ^ n24791 ^ n11899 ;
  assign n46190 = ( n19993 & ~n41486 ) | ( n19993 & n46189 ) | ( ~n41486 & n46189 ) ;
  assign n46191 = ( ~n3862 & n9825 ) | ( ~n3862 & n18675 ) | ( n9825 & n18675 ) ;
  assign n46192 = n46191 ^ n12612 ^ n7193 ;
  assign n46193 = n43881 ^ n16130 ^ n5066 ;
  assign n46194 = ( n9555 & n35398 ) | ( n9555 & ~n39130 ) | ( n35398 & ~n39130 ) ;
  assign n46195 = ( n21017 & n31753 ) | ( n21017 & ~n46194 ) | ( n31753 & ~n46194 ) ;
  assign n46197 = n43410 ^ n10418 ^ n1902 ;
  assign n46196 = n30824 ^ n14264 ^ n2925 ;
  assign n46198 = n46197 ^ n46196 ^ n19513 ;
  assign n46199 = ( n13484 & n39909 ) | ( n13484 & n43207 ) | ( n39909 & n43207 ) ;
  assign n46200 = ( n10897 & n19021 ) | ( n10897 & n46199 ) | ( n19021 & n46199 ) ;
  assign n46201 = ( n12347 & n16624 ) | ( n12347 & n39305 ) | ( n16624 & n39305 ) ;
  assign n46202 = n41399 ^ n37817 ^ n2342 ;
  assign n46203 = n46202 ^ n8207 ^ 1'b0 ;
  assign n46204 = n39419 ^ n35134 ^ n13261 ;
  assign n46205 = ( n10300 & n15104 ) | ( n10300 & ~n25703 ) | ( n15104 & ~n25703 ) ;
  assign n46206 = n46205 ^ n37473 ^ n855 ;
  assign n46207 = n46206 ^ n29779 ^ n10165 ;
  assign n46208 = ( ~n4262 & n4876 ) | ( ~n4262 & n19213 ) | ( n4876 & n19213 ) ;
  assign n46209 = n46208 ^ n13627 ^ n4481 ;
  assign n46215 = n16408 ^ n6815 ^ n3348 ;
  assign n46214 = n31983 ^ n23452 ^ x103 ;
  assign n46216 = n46215 ^ n46214 ^ n41696 ;
  assign n46213 = n26111 ^ n24033 ^ 1'b0 ;
  assign n46210 = n15768 ^ x116 ^ 1'b0 ;
  assign n46211 = ~n22810 & n39069 ;
  assign n46212 = n46210 & n46211 ;
  assign n46217 = n46216 ^ n46213 ^ n46212 ;
  assign n46219 = n31837 ^ n14159 ^ n13593 ;
  assign n46220 = x63 & n1489 ;
  assign n46221 = n46220 ^ n11126 ^ 1'b0 ;
  assign n46222 = n46221 ^ n16039 ^ n5863 ;
  assign n46223 = ( n28940 & n46219 ) | ( n28940 & ~n46222 ) | ( n46219 & ~n46222 ) ;
  assign n46218 = n33298 ^ n19586 ^ 1'b0 ;
  assign n46224 = n46223 ^ n46218 ^ n11632 ;
  assign n46225 = n2498 & ~n30127 ;
  assign n46226 = n37683 ^ n10967 ^ n3542 ;
  assign n46230 = n39726 ^ n27419 ^ 1'b0 ;
  assign n46231 = n40602 | n46230 ;
  assign n46227 = n8341 ^ n4082 ^ n1848 ;
  assign n46228 = ( n3954 & ~n39887 ) | ( n3954 & n46227 ) | ( ~n39887 & n46227 ) ;
  assign n46229 = ( n9924 & n18660 ) | ( n9924 & ~n46228 ) | ( n18660 & ~n46228 ) ;
  assign n46232 = n46231 ^ n46229 ^ n43470 ;
  assign n46234 = ( ~n6871 & n13117 ) | ( ~n6871 & n14647 ) | ( n13117 & n14647 ) ;
  assign n46233 = n22547 ^ n16626 ^ n7160 ;
  assign n46235 = n46234 ^ n46233 ^ n22806 ;
  assign n46236 = n15089 & ~n46235 ;
  assign n46237 = ( n12965 & ~n38025 ) | ( n12965 & n43071 ) | ( ~n38025 & n43071 ) ;
  assign n46238 = ( n8386 & ~n8913 ) | ( n8386 & n11442 ) | ( ~n8913 & n11442 ) ;
  assign n46239 = ( n6016 & n9984 ) | ( n6016 & n46238 ) | ( n9984 & n46238 ) ;
  assign n46240 = ( n20625 & n35963 ) | ( n20625 & ~n46239 ) | ( n35963 & ~n46239 ) ;
  assign n46241 = ( n6007 & n11832 ) | ( n6007 & n19005 ) | ( n11832 & n19005 ) ;
  assign n46242 = n46241 ^ n19201 ^ n5597 ;
  assign n46243 = ( ~n3971 & n14254 ) | ( ~n3971 & n46242 ) | ( n14254 & n46242 ) ;
  assign n46244 = ( n46237 & ~n46240 ) | ( n46237 & n46243 ) | ( ~n46240 & n46243 ) ;
  assign n46245 = ( n8984 & n10891 ) | ( n8984 & ~n36296 ) | ( n10891 & ~n36296 ) ;
  assign n46246 = n29311 ^ n20549 ^ n7332 ;
  assign n46247 = n46246 ^ n33792 ^ n29366 ;
  assign n46248 = n25335 ^ n14879 ^ 1'b0 ;
  assign n46249 = ( n23795 & n32637 ) | ( n23795 & ~n46248 ) | ( n32637 & ~n46248 ) ;
  assign n46252 = n15892 ^ n5896 ^ n1267 ;
  assign n46251 = ( n8784 & ~n15620 ) | ( n8784 & n21402 ) | ( ~n15620 & n21402 ) ;
  assign n46250 = n30044 ^ n20886 ^ 1'b0 ;
  assign n46253 = n46252 ^ n46251 ^ n46250 ;
  assign n46254 = n30772 ^ n7640 ^ n4309 ;
  assign n46255 = n34773 ^ n13014 ^ 1'b0 ;
  assign n46256 = n907 & n46255 ;
  assign n46257 = n46256 ^ n590 ^ 1'b0 ;
  assign n46258 = ( ~n10775 & n46254 ) | ( ~n10775 & n46257 ) | ( n46254 & n46257 ) ;
  assign n46259 = n43160 ^ n18072 ^ 1'b0 ;
  assign n46260 = n34910 & ~n46259 ;
  assign n46261 = ( n1432 & ~n22063 ) | ( n1432 & n37179 ) | ( ~n22063 & n37179 ) ;
  assign n46262 = n46261 ^ n8588 ^ n3923 ;
  assign n46263 = ~n9092 & n24182 ;
  assign n46264 = ~n8862 & n46263 ;
  assign n46265 = ( ~n18185 & n30896 ) | ( ~n18185 & n35950 ) | ( n30896 & n35950 ) ;
  assign n46266 = ( n46262 & ~n46264 ) | ( n46262 & n46265 ) | ( ~n46264 & n46265 ) ;
  assign n46267 = n35043 ^ n25546 ^ 1'b0 ;
  assign n46268 = ~n46266 & n46267 ;
  assign n46269 = n2566 & ~n27343 ;
  assign n46270 = n46269 ^ n31472 ^ n15259 ;
  assign n46271 = ( n4835 & n8420 ) | ( n4835 & ~n40524 ) | ( n8420 & ~n40524 ) ;
  assign n46272 = n46271 ^ n35310 ^ n14401 ;
  assign n46273 = ( n10252 & n30215 ) | ( n10252 & n46272 ) | ( n30215 & n46272 ) ;
  assign n46274 = ( n1971 & ~n44248 ) | ( n1971 & n45639 ) | ( ~n44248 & n45639 ) ;
  assign n46275 = ( n7496 & n29227 ) | ( n7496 & n46274 ) | ( n29227 & n46274 ) ;
  assign n46277 = ( n2421 & n7585 ) | ( n2421 & n41875 ) | ( n7585 & n41875 ) ;
  assign n46278 = ( n16581 & n26247 ) | ( n16581 & n46277 ) | ( n26247 & n46277 ) ;
  assign n46279 = ( n34113 & ~n35419 ) | ( n34113 & n46278 ) | ( ~n35419 & n46278 ) ;
  assign n46276 = n20975 ^ n2673 ^ 1'b0 ;
  assign n46280 = n46279 ^ n46276 ^ n30957 ;
  assign n46281 = n35868 | n44760 ;
  assign n46282 = ~n9533 & n14506 ;
  assign n46283 = n13985 | n46282 ;
  assign n46284 = n46283 ^ n6552 ^ 1'b0 ;
  assign n46285 = ~n25798 & n31784 ;
  assign n46286 = ( n15113 & n36158 ) | ( n15113 & ~n43738 ) | ( n36158 & ~n43738 ) ;
  assign n46287 = ~n435 & n28513 ;
  assign n46288 = n44868 ^ n20447 ^ 1'b0 ;
  assign n46289 = ( ~n5489 & n8849 ) | ( ~n5489 & n11354 ) | ( n8849 & n11354 ) ;
  assign n46290 = ( ~n12540 & n14317 ) | ( ~n12540 & n46289 ) | ( n14317 & n46289 ) ;
  assign n46291 = n46290 ^ n37041 ^ x160 ;
  assign n46292 = ( n28778 & n36264 ) | ( n28778 & ~n45557 ) | ( n36264 & ~n45557 ) ;
  assign n46293 = ( x60 & n31253 ) | ( x60 & n46292 ) | ( n31253 & n46292 ) ;
  assign n46294 = ( ~n8178 & n19426 ) | ( ~n8178 & n46293 ) | ( n19426 & n46293 ) ;
  assign n46295 = n2029 ^ n487 ^ 1'b0 ;
  assign n46296 = ~n10385 & n46295 ;
  assign n46297 = ( n8738 & n26246 ) | ( n8738 & ~n46296 ) | ( n26246 & ~n46296 ) ;
  assign n46298 = ( n3333 & n19284 ) | ( n3333 & ~n46297 ) | ( n19284 & ~n46297 ) ;
  assign n46299 = n34050 ^ n12275 ^ n5345 ;
  assign n46300 = n46299 ^ n5336 ^ n1024 ;
  assign n46301 = n46300 ^ n32478 ^ n6650 ;
  assign n46302 = ( ~n11951 & n30609 ) | ( ~n11951 & n33430 ) | ( n30609 & n33430 ) ;
  assign n46304 = n29836 ^ n5395 ^ n3826 ;
  assign n46303 = ~n14085 & n39249 ;
  assign n46305 = n46304 ^ n46303 ^ 1'b0 ;
  assign n46306 = ( ~n2564 & n16094 ) | ( ~n2564 & n35756 ) | ( n16094 & n35756 ) ;
  assign n46307 = n35832 ^ n33042 ^ n16945 ;
  assign n46308 = n35062 ^ n3957 ^ n1492 ;
  assign n46309 = ( n5013 & ~n5603 ) | ( n5013 & n12103 ) | ( ~n5603 & n12103 ) ;
  assign n46310 = n46309 ^ n10073 ^ n6742 ;
  assign n46311 = ( n5757 & ~n46308 ) | ( n5757 & n46310 ) | ( ~n46308 & n46310 ) ;
  assign n46312 = ( ~n1645 & n4168 ) | ( ~n1645 & n36027 ) | ( n4168 & n36027 ) ;
  assign n46313 = ( ~n1759 & n6353 ) | ( ~n1759 & n16305 ) | ( n6353 & n16305 ) ;
  assign n46314 = ( x243 & ~n7212 ) | ( x243 & n13198 ) | ( ~n7212 & n13198 ) ;
  assign n46315 = n3189 | n3340 ;
  assign n46316 = n15658 & ~n46315 ;
  assign n46317 = n46316 ^ n32714 ^ n21494 ;
  assign n46321 = ( n7146 & n23617 ) | ( n7146 & ~n45868 ) | ( n23617 & ~n45868 ) ;
  assign n46318 = ( n25781 & ~n28891 ) | ( n25781 & n29759 ) | ( ~n28891 & n29759 ) ;
  assign n46319 = n33876 ^ n30670 ^ n26366 ;
  assign n46320 = n46318 | n46319 ;
  assign n46322 = n46321 ^ n46320 ^ 1'b0 ;
  assign n46323 = n22400 ^ n12042 ^ n10477 ;
  assign n46324 = n46323 ^ n40685 ^ n39642 ;
  assign n46325 = n24562 ^ n23237 ^ n7684 ;
  assign n46326 = ( n27858 & n38174 ) | ( n27858 & n46325 ) | ( n38174 & n46325 ) ;
  assign n46327 = n1378 | n13123 ;
  assign n46328 = n21636 | n46327 ;
  assign n46329 = n46328 ^ n31713 ^ n5441 ;
  assign n46330 = n17048 ^ n12259 ^ n10105 ;
  assign n46331 = n39058 & n46330 ;
  assign n46332 = n46331 ^ n39665 ^ n6192 ;
  assign n46335 = n44585 ^ n4096 ^ 1'b0 ;
  assign n46336 = ~n40612 & n46335 ;
  assign n46333 = n19802 ^ n11353 ^ n2748 ;
  assign n46334 = ( n21502 & n24615 ) | ( n21502 & n46333 ) | ( n24615 & n46333 ) ;
  assign n46337 = n46336 ^ n46334 ^ n24835 ;
  assign n46338 = n35218 ^ n24873 ^ n19042 ;
  assign n46339 = n46338 ^ n44379 ^ 1'b0 ;
  assign n46340 = ( n9181 & ~n20530 ) | ( n9181 & n29608 ) | ( ~n20530 & n29608 ) ;
  assign n46341 = n44568 ^ n44223 ^ n38414 ;
  assign n46342 = ( n2159 & n13766 ) | ( n2159 & ~n13886 ) | ( n13766 & ~n13886 ) ;
  assign n46343 = n46342 ^ n26450 ^ n8746 ;
  assign n46346 = ( n10643 & n12108 ) | ( n10643 & ~n41446 ) | ( n12108 & ~n41446 ) ;
  assign n46344 = ( n10489 & n17084 ) | ( n10489 & ~n30529 ) | ( n17084 & ~n30529 ) ;
  assign n46345 = ( n7554 & ~n22972 ) | ( n7554 & n46344 ) | ( ~n22972 & n46344 ) ;
  assign n46347 = n46346 ^ n46345 ^ n31563 ;
  assign n46348 = ( n3889 & ~n4816 ) | ( n3889 & n36112 ) | ( ~n4816 & n36112 ) ;
  assign n46349 = n46348 ^ n7703 ^ n6829 ;
  assign n46350 = ( n31736 & n45626 ) | ( n31736 & ~n46349 ) | ( n45626 & ~n46349 ) ;
  assign n46351 = ( ~n5808 & n12732 ) | ( ~n5808 & n32350 ) | ( n12732 & n32350 ) ;
  assign n46352 = ( n3465 & n46344 ) | ( n3465 & ~n46351 ) | ( n46344 & ~n46351 ) ;
  assign n46353 = ( n38373 & ~n46350 ) | ( n38373 & n46352 ) | ( ~n46350 & n46352 ) ;
  assign n46354 = n2214 | n22722 ;
  assign n46355 = n46354 ^ n10261 ^ n9422 ;
  assign n46356 = n34602 ^ n2000 ^ 1'b0 ;
  assign n46357 = ~n2538 & n46356 ;
  assign n46358 = ( n26357 & ~n46355 ) | ( n26357 & n46357 ) | ( ~n46355 & n46357 ) ;
  assign n46359 = n27534 ^ n12366 ^ n1531 ;
  assign n46360 = n46359 ^ n42757 ^ n19334 ;
  assign n46361 = ( n15188 & n21232 ) | ( n15188 & ~n46360 ) | ( n21232 & ~n46360 ) ;
  assign n46362 = ( n11651 & n17998 ) | ( n11651 & ~n46361 ) | ( n17998 & ~n46361 ) ;
  assign n46363 = n37138 ^ n26943 ^ 1'b0 ;
  assign n46364 = n15234 | n46363 ;
  assign n46365 = ( n24500 & n25142 ) | ( n24500 & ~n46364 ) | ( n25142 & ~n46364 ) ;
  assign n46366 = n8228 ^ n448 ^ 1'b0 ;
  assign n46367 = ~n12803 & n46366 ;
  assign n46368 = n29302 ^ n10488 ^ n4282 ;
  assign n46369 = n24476 ^ n13007 ^ n9406 ;
  assign n46370 = n32973 ^ n30783 ^ n28375 ;
  assign n46371 = n17411 ^ n7554 ^ n6156 ;
  assign n46372 = n46371 ^ n39003 ^ n589 ;
  assign n46376 = n898 & n19730 ;
  assign n46377 = n14918 ^ n1247 ^ 1'b0 ;
  assign n46378 = n46376 & n46377 ;
  assign n46373 = ( n2775 & n3520 ) | ( n2775 & n25741 ) | ( n3520 & n25741 ) ;
  assign n46374 = ( ~x157 & x204 ) | ( ~x157 & n46373 ) | ( x204 & n46373 ) ;
  assign n46375 = n46374 ^ n33935 ^ n9690 ;
  assign n46379 = n46378 ^ n46375 ^ n39708 ;
  assign n46381 = n9265 & n10252 ;
  assign n46382 = ~n32505 & n46381 ;
  assign n46380 = n16255 & ~n34841 ;
  assign n46383 = n46382 ^ n46380 ^ 1'b0 ;
  assign n46384 = n31461 ^ n9066 ^ n6285 ;
  assign n46385 = n46384 ^ n23775 ^ n8118 ;
  assign n46386 = n44147 ^ n23431 ^ n15088 ;
  assign n46387 = ( n18318 & n33029 ) | ( n18318 & ~n46130 ) | ( n33029 & ~n46130 ) ;
  assign n46388 = n39106 ^ n26039 ^ n3359 ;
  assign n46389 = n18259 ^ n4941 ^ n2037 ;
  assign n46390 = n13978 & ~n36304 ;
  assign n46391 = n46389 & n46390 ;
  assign n46392 = n46391 ^ n7145 ^ n5612 ;
  assign n46393 = ( n20817 & n30022 ) | ( n20817 & n46392 ) | ( n30022 & n46392 ) ;
  assign n46394 = n38566 ^ n32439 ^ n31403 ;
  assign n46395 = ( n2445 & n6260 ) | ( n2445 & ~n37786 ) | ( n6260 & ~n37786 ) ;
  assign n46396 = ( n15174 & n21511 ) | ( n15174 & n46395 ) | ( n21511 & n46395 ) ;
  assign n46397 = n19258 ^ n6444 ^ 1'b0 ;
  assign n46398 = ( n3976 & ~n15435 ) | ( n3976 & n26430 ) | ( ~n15435 & n26430 ) ;
  assign n46399 = ( n26665 & ~n46397 ) | ( n26665 & n46398 ) | ( ~n46397 & n46398 ) ;
  assign n46400 = n35356 ^ n23313 ^ n6347 ;
  assign n46401 = n45205 | n46400 ;
  assign n46402 = ( n6494 & ~n17545 ) | ( n6494 & n26199 ) | ( ~n17545 & n26199 ) ;
  assign n46403 = n46402 ^ n8428 ^ 1'b0 ;
  assign n46404 = n14883 ^ n12507 ^ n5566 ;
  assign n46405 = n46404 ^ n36294 ^ n26322 ;
  assign n46406 = n41616 ^ n32098 ^ n6846 ;
  assign n46407 = ~n37710 & n39370 ;
  assign n46408 = n40635 ^ n17425 ^ n369 ;
  assign n46409 = ( ~n4931 & n13458 ) | ( ~n4931 & n18660 ) | ( n13458 & n18660 ) ;
  assign n46410 = ( ~n28437 & n32416 ) | ( ~n28437 & n43696 ) | ( n32416 & n43696 ) ;
  assign n46411 = n22368 ^ n3813 ^ 1'b0 ;
  assign n46412 = n11119 & ~n46411 ;
  assign n46413 = n45531 ^ n26430 ^ n11244 ;
  assign n46414 = n46413 ^ n4445 ^ 1'b0 ;
  assign n46415 = n1681 & ~n46414 ;
  assign n46416 = n20717 ^ n8440 ^ n3062 ;
  assign n46417 = n46416 ^ n21758 ^ n867 ;
  assign n46418 = n46417 ^ n35105 ^ 1'b0 ;
  assign n46419 = ~n9606 & n46418 ;
  assign n46420 = ( n1903 & n22252 ) | ( n1903 & ~n46419 ) | ( n22252 & ~n46419 ) ;
  assign n46421 = ( n3646 & n21984 ) | ( n3646 & n46420 ) | ( n21984 & n46420 ) ;
  assign n46422 = ~n35527 & n40019 ;
  assign n46423 = n4426 | n18313 ;
  assign n46424 = n27876 ^ n6854 ^ n1492 ;
  assign n46425 = n33263 ^ n20464 ^ n3657 ;
  assign n46426 = n5068 & n15088 ;
  assign n46427 = n46426 ^ n17777 ^ 1'b0 ;
  assign n46428 = n46427 ^ n45310 ^ n9164 ;
  assign n46429 = ( n46424 & n46425 ) | ( n46424 & n46428 ) | ( n46425 & n46428 ) ;
  assign n46430 = n32041 | n34226 ;
  assign n46431 = n46430 ^ n21196 ^ 1'b0 ;
  assign n46432 = ( n5872 & ~n7690 ) | ( n5872 & n16617 ) | ( ~n7690 & n16617 ) ;
  assign n46433 = ( n7947 & n15336 ) | ( n7947 & n46432 ) | ( n15336 & n46432 ) ;
  assign n46434 = ( n2214 & n3905 ) | ( n2214 & n46433 ) | ( n3905 & n46433 ) ;
  assign n46435 = ( n13773 & n46431 ) | ( n13773 & ~n46434 ) | ( n46431 & ~n46434 ) ;
  assign n46436 = n38370 ^ n7837 ^ n6109 ;
  assign n46437 = ( n2018 & n29154 ) | ( n2018 & ~n46436 ) | ( n29154 & ~n46436 ) ;
  assign n46438 = n28069 ^ n13100 ^ n295 ;
  assign n46439 = n26546 & n36086 ;
  assign n46440 = n46439 ^ n19723 ^ n11840 ;
  assign n46441 = n46440 ^ n44617 ^ n32611 ;
  assign n46442 = n13760 & n22113 ;
  assign n46443 = n46442 ^ n42997 ^ 1'b0 ;
  assign n46444 = n7403 & ~n9204 ;
  assign n46445 = n46444 ^ n45076 ^ 1'b0 ;
  assign n46446 = n35494 ^ n24574 ^ n2303 ;
  assign n46447 = n46446 ^ n15802 ^ 1'b0 ;
  assign n46448 = ~n2449 & n46447 ;
  assign n46449 = ( ~n21409 & n23059 ) | ( ~n21409 & n46448 ) | ( n23059 & n46448 ) ;
  assign n46450 = ( n899 & n1964 ) | ( n899 & n46449 ) | ( n1964 & n46449 ) ;
  assign n46451 = ( ~n4250 & n17398 ) | ( ~n4250 & n29218 ) | ( n17398 & n29218 ) ;
  assign n46452 = ( n7502 & n12348 ) | ( n7502 & ~n46451 ) | ( n12348 & ~n46451 ) ;
  assign n46453 = ( ~n21280 & n22830 ) | ( ~n21280 & n28597 ) | ( n22830 & n28597 ) ;
  assign n46454 = n2189 & n46453 ;
  assign n46455 = ( n11364 & n22996 ) | ( n11364 & ~n23166 ) | ( n22996 & ~n23166 ) ;
  assign n46456 = n39341 ^ n11284 ^ n5505 ;
  assign n46457 = ( n22643 & n25065 ) | ( n22643 & ~n46456 ) | ( n25065 & ~n46456 ) ;
  assign n46458 = ( n31145 & ~n46455 ) | ( n31145 & n46457 ) | ( ~n46455 & n46457 ) ;
  assign n46459 = n8885 ^ n7163 ^ n5298 ;
  assign n46460 = ( n12969 & ~n38625 ) | ( n12969 & n46090 ) | ( ~n38625 & n46090 ) ;
  assign n46461 = ( n22979 & n38806 ) | ( n22979 & ~n46460 ) | ( n38806 & ~n46460 ) ;
  assign n46462 = ( ~n7674 & n42929 ) | ( ~n7674 & n46461 ) | ( n42929 & n46461 ) ;
  assign n46463 = ( n20930 & n46459 ) | ( n20930 & n46462 ) | ( n46459 & n46462 ) ;
  assign n46464 = n11291 | n20181 ;
  assign n46465 = n24018 | n46464 ;
  assign n46466 = ( n3777 & n12748 ) | ( n3777 & ~n46465 ) | ( n12748 & ~n46465 ) ;
  assign n46467 = ( ~n1884 & n6639 ) | ( ~n1884 & n46466 ) | ( n6639 & n46466 ) ;
  assign n46468 = x108 & n3349 ;
  assign n46469 = n3786 & n29250 ;
  assign n46470 = ( n35472 & n46468 ) | ( n35472 & n46469 ) | ( n46468 & n46469 ) ;
  assign n46473 = n23855 ^ n6250 ^ n2854 ;
  assign n46471 = n14378 | n32678 ;
  assign n46472 = n46471 ^ n3694 ^ 1'b0 ;
  assign n46474 = n46473 ^ n46472 ^ n31467 ;
  assign n46475 = ( n3921 & n10411 ) | ( n3921 & ~n46474 ) | ( n10411 & ~n46474 ) ;
  assign n46476 = n46475 ^ n42604 ^ 1'b0 ;
  assign n46477 = n46103 | n46476 ;
  assign n46478 = n25957 ^ n16790 ^ 1'b0 ;
  assign n46479 = ( n7977 & ~n11425 ) | ( n7977 & n13440 ) | ( ~n11425 & n13440 ) ;
  assign n46480 = ( n3832 & n33806 ) | ( n3832 & ~n46479 ) | ( n33806 & ~n46479 ) ;
  assign n46481 = ( ~n10098 & n22078 ) | ( ~n10098 & n42677 ) | ( n22078 & n42677 ) ;
  assign n46482 = n42288 ^ n19752 ^ n13612 ;
  assign n46483 = ( ~n12288 & n16370 ) | ( ~n12288 & n28897 ) | ( n16370 & n28897 ) ;
  assign n46484 = n5027 & ~n46483 ;
  assign n46485 = ( ~n23234 & n28987 ) | ( ~n23234 & n46484 ) | ( n28987 & n46484 ) ;
  assign n46486 = ( ~n10474 & n11948 ) | ( ~n10474 & n25234 ) | ( n11948 & n25234 ) ;
  assign n46487 = n46486 ^ n21560 ^ n6849 ;
  assign n46491 = n28096 ^ n7257 ^ n3597 ;
  assign n46488 = n11125 ^ n9017 ^ n4997 ;
  assign n46489 = n24608 & ~n39088 ;
  assign n46490 = n46488 & n46489 ;
  assign n46492 = n46491 ^ n46490 ^ n8290 ;
  assign n46493 = ( n23313 & n39457 ) | ( n23313 & ~n46492 ) | ( n39457 & ~n46492 ) ;
  assign n46494 = ( n14589 & n46487 ) | ( n14589 & ~n46493 ) | ( n46487 & ~n46493 ) ;
  assign n46495 = ( ~n24717 & n29452 ) | ( ~n24717 & n30084 ) | ( n29452 & n30084 ) ;
  assign n46496 = ( ~n21112 & n22190 ) | ( ~n21112 & n46495 ) | ( n22190 & n46495 ) ;
  assign n46497 = ( n378 & n26470 ) | ( n378 & n46496 ) | ( n26470 & n46496 ) ;
  assign n46498 = ~n19534 & n23315 ;
  assign n46499 = n46074 ^ n34278 ^ n31692 ;
  assign n46500 = n37785 ^ n6096 ^ x61 ;
  assign n46504 = n21066 & n25667 ;
  assign n46505 = n2840 & n46504 ;
  assign n46503 = n40247 ^ n24568 ^ n13892 ;
  assign n46501 = ( n2509 & ~n12447 ) | ( n2509 & n22808 ) | ( ~n12447 & n22808 ) ;
  assign n46502 = n46501 ^ n12044 ^ n8271 ;
  assign n46506 = n46505 ^ n46503 ^ n46502 ;
  assign n46507 = ( n10442 & n46500 ) | ( n10442 & n46506 ) | ( n46500 & n46506 ) ;
  assign n46508 = ( n25220 & ~n33321 ) | ( n25220 & n46507 ) | ( ~n33321 & n46507 ) ;
  assign n46509 = n3781 ^ n3194 ^ 1'b0 ;
  assign n46510 = n46509 ^ n17821 ^ n13605 ;
  assign n46513 = n10401 ^ n1390 ^ 1'b0 ;
  assign n46514 = n1323 | n46513 ;
  assign n46512 = n8227 ^ n3025 ^ n1362 ;
  assign n46511 = n29577 ^ n12551 ^ n7939 ;
  assign n46515 = n46514 ^ n46512 ^ n46511 ;
  assign n46516 = n15694 ^ n4275 ^ 1'b0 ;
  assign n46517 = n46516 ^ n33449 ^ n28475 ;
  assign n46518 = n11275 ^ n8546 ^ n4888 ;
  assign n46519 = n33420 | n46518 ;
  assign n46520 = n19917 ^ n2188 ^ n1932 ;
  assign n46521 = ( n8101 & n12967 ) | ( n8101 & n25966 ) | ( n12967 & n25966 ) ;
  assign n46522 = n45732 ^ n25587 ^ n11833 ;
  assign n46524 = n24372 ^ n11164 ^ n9962 ;
  assign n46523 = n12406 & ~n42550 ;
  assign n46525 = n46524 ^ n46523 ^ 1'b0 ;
  assign n46526 = n40905 ^ n22839 ^ 1'b0 ;
  assign n46527 = n11618 & ~n46526 ;
  assign n46528 = n25274 ^ n9073 ^ n4856 ;
  assign n46529 = n46528 ^ n9261 ^ 1'b0 ;
  assign n46530 = n8923 ^ n6414 ^ n3523 ;
  assign n46531 = ( n15602 & ~n29284 ) | ( n15602 & n40285 ) | ( ~n29284 & n40285 ) ;
  assign n46534 = ( n6736 & n30050 ) | ( n6736 & ~n38784 ) | ( n30050 & ~n38784 ) ;
  assign n46532 = n8761 ^ n7663 ^ n1539 ;
  assign n46533 = n46532 ^ n25428 ^ n1578 ;
  assign n46535 = n46534 ^ n46533 ^ n35250 ;
  assign n46536 = ( n24541 & n31418 ) | ( n24541 & n46413 ) | ( n31418 & n46413 ) ;
  assign n46537 = n20522 ^ n19127 ^ n16574 ;
  assign n46539 = n21200 ^ n16173 ^ 1'b0 ;
  assign n46538 = n46459 ^ n37305 ^ n10885 ;
  assign n46540 = n46539 ^ n46538 ^ n7692 ;
  assign n46545 = n3402 & n13048 ;
  assign n46546 = n46545 ^ n40893 ^ n943 ;
  assign n46541 = n6710 & n13553 ;
  assign n46542 = n46541 ^ n10419 ^ n1322 ;
  assign n46543 = n46542 ^ n42123 ^ n3613 ;
  assign n46544 = n22265 | n46543 ;
  assign n46547 = n46546 ^ n46544 ^ 1'b0 ;
  assign n46548 = n31604 ^ n9965 ^ n2041 ;
  assign n46549 = n46548 ^ n46223 ^ n13155 ;
  assign n46552 = n14724 ^ n11566 ^ n5387 ;
  assign n46550 = n10036 & n28799 ;
  assign n46551 = ~n840 & n46550 ;
  assign n46553 = n46552 ^ n46551 ^ n6532 ;
  assign n46554 = ( n4189 & n6124 ) | ( n4189 & n23138 ) | ( n6124 & n23138 ) ;
  assign n46555 = ( n547 & ~n22632 ) | ( n547 & n46554 ) | ( ~n22632 & n46554 ) ;
  assign n46556 = n38543 ^ n14624 ^ 1'b0 ;
  assign n46557 = ~n11155 & n46556 ;
  assign n46558 = n46557 ^ n14321 ^ n12672 ;
  assign n46559 = n46558 ^ n35071 ^ n3631 ;
  assign n46560 = n13984 ^ n12528 ^ n9741 ;
  assign n46561 = n32611 ^ n4869 ^ 1'b0 ;
  assign n46562 = ( ~n8156 & n15872 ) | ( ~n8156 & n42225 ) | ( n15872 & n42225 ) ;
  assign n46563 = ( ~n20332 & n46561 ) | ( ~n20332 & n46562 ) | ( n46561 & n46562 ) ;
  assign n46564 = n22236 | n40967 ;
  assign n46565 = n17135 & n34937 ;
  assign n46566 = n28127 ^ n22926 ^ n8793 ;
  assign n46567 = ( n4801 & n14417 ) | ( n4801 & n17734 ) | ( n14417 & n17734 ) ;
  assign n46568 = ( n6311 & n31219 ) | ( n6311 & ~n46567 ) | ( n31219 & ~n46567 ) ;
  assign n46569 = n7937 & ~n46568 ;
  assign n46570 = ~n46566 & n46569 ;
  assign n46571 = n24388 & ~n28641 ;
  assign n46572 = n46571 ^ n10304 ^ 1'b0 ;
  assign n46573 = ~n46022 & n46572 ;
  assign n46574 = n14172 ^ n6917 ^ 1'b0 ;
  assign n46575 = n19809 ^ n7167 ^ n7140 ;
  assign n46576 = n44148 ^ n39938 ^ n15339 ;
  assign n46577 = n44378 ^ n12506 ^ n6118 ;
  assign n46578 = ( n25216 & n34155 ) | ( n25216 & n46577 ) | ( n34155 & n46577 ) ;
  assign n46579 = ( ~n5245 & n39342 ) | ( ~n5245 & n45724 ) | ( n39342 & n45724 ) ;
  assign n46580 = n42365 ^ n5076 ^ 1'b0 ;
  assign n46581 = n41360 | n46580 ;
  assign n46582 = n9190 ^ n8259 ^ 1'b0 ;
  assign n46583 = n17432 | n46582 ;
  assign n46584 = ( n15292 & ~n15717 ) | ( n15292 & n46583 ) | ( ~n15717 & n46583 ) ;
  assign n46585 = ~n44821 & n46584 ;
  assign n46586 = n44153 ^ n39308 ^ 1'b0 ;
  assign n46587 = ~n46585 & n46586 ;
  assign n46588 = n32806 ^ n29720 ^ n13735 ;
  assign n46589 = n7173 ^ n3068 ^ n1134 ;
  assign n46591 = n19578 ^ n11734 ^ n2617 ;
  assign n46590 = n15617 ^ n12114 ^ n6795 ;
  assign n46592 = n46591 ^ n46590 ^ n38117 ;
  assign n46593 = ( n7098 & n14386 ) | ( n7098 & n29305 ) | ( n14386 & n29305 ) ;
  assign n46594 = n46593 ^ n15116 ^ 1'b0 ;
  assign n46595 = ( ~n46589 & n46592 ) | ( ~n46589 & n46594 ) | ( n46592 & n46594 ) ;
  assign n46596 = n42070 ^ n41412 ^ n15377 ;
  assign n46597 = n29435 ^ n17997 ^ n14084 ;
  assign n46598 = n37013 ^ n24969 ^ n1153 ;
  assign n46599 = ( n669 & n40311 ) | ( n669 & n46598 ) | ( n40311 & n46598 ) ;
  assign n46600 = ( n15422 & ~n44057 ) | ( n15422 & n46599 ) | ( ~n44057 & n46599 ) ;
  assign n46601 = ( n3491 & ~n7808 ) | ( n3491 & n21383 ) | ( ~n7808 & n21383 ) ;
  assign n46602 = n46601 ^ n15358 ^ 1'b0 ;
  assign n46603 = n17179 & n46602 ;
  assign n46604 = ( n6462 & ~n12626 ) | ( n6462 & n15188 ) | ( ~n12626 & n15188 ) ;
  assign n46605 = ( n26678 & n33539 ) | ( n26678 & ~n46604 ) | ( n33539 & ~n46604 ) ;
  assign n46606 = ( ~n8679 & n24405 ) | ( ~n8679 & n46605 ) | ( n24405 & n46605 ) ;
  assign n46607 = n37913 ^ n24801 ^ n1971 ;
  assign n46608 = n3461 & n6917 ;
  assign n46609 = n46608 ^ n9190 ^ 1'b0 ;
  assign n46610 = n46609 ^ n44327 ^ n1078 ;
  assign n46611 = n46610 ^ n13515 ^ 1'b0 ;
  assign n46612 = ( n6169 & n7362 ) | ( n6169 & n17547 ) | ( n7362 & n17547 ) ;
  assign n46613 = n1356 & n46612 ;
  assign n46614 = ( n2809 & n39346 ) | ( n2809 & ~n46613 ) | ( n39346 & ~n46613 ) ;
  assign n46615 = n38770 ^ n36712 ^ n27655 ;
  assign n46616 = n46615 ^ n36937 ^ n35933 ;
  assign n46617 = ( n355 & n1588 ) | ( n355 & ~n36459 ) | ( n1588 & ~n36459 ) ;
  assign n46618 = ( n13508 & n45925 ) | ( n13508 & n46617 ) | ( n45925 & n46617 ) ;
  assign n46619 = ( n2337 & n6559 ) | ( n2337 & ~n18702 ) | ( n6559 & ~n18702 ) ;
  assign n46620 = ( n365 & n9720 ) | ( n365 & ~n44469 ) | ( n9720 & ~n44469 ) ;
  assign n46621 = ( ~n18771 & n46619 ) | ( ~n18771 & n46620 ) | ( n46619 & n46620 ) ;
  assign n46622 = n9725 ^ n3391 ^ 1'b0 ;
  assign n46623 = n23556 | n46622 ;
  assign n46624 = n42652 ^ n31639 ^ n20241 ;
  assign n46625 = ( n14690 & n19009 ) | ( n14690 & n46624 ) | ( n19009 & n46624 ) ;
  assign n46626 = n46625 ^ n10997 ^ n4623 ;
  assign n46627 = n8911 ^ x248 ^ 1'b0 ;
  assign n46630 = ( n19982 & n27307 ) | ( n19982 & n27896 ) | ( n27307 & n27896 ) ;
  assign n46628 = ~n3561 & n32447 ;
  assign n46629 = n46628 ^ n22874 ^ 1'b0 ;
  assign n46631 = n46630 ^ n46629 ^ n23918 ;
  assign n46635 = ( n10826 & n16500 ) | ( n10826 & n33365 ) | ( n16500 & n33365 ) ;
  assign n46632 = x200 & ~n453 ;
  assign n46633 = n46632 ^ n1733 ^ 1'b0 ;
  assign n46634 = ( ~n2747 & n30604 ) | ( ~n2747 & n46633 ) | ( n30604 & n46633 ) ;
  assign n46636 = n46635 ^ n46634 ^ n6077 ;
  assign n46637 = n46636 ^ n42166 ^ n1396 ;
  assign n46638 = ( n1367 & n11171 ) | ( n1367 & ~n17640 ) | ( n11171 & ~n17640 ) ;
  assign n46639 = ( n6506 & ~n34562 ) | ( n6506 & n46638 ) | ( ~n34562 & n46638 ) ;
  assign n46640 = n46639 ^ n14094 ^ n1566 ;
  assign n46644 = n39747 ^ n19828 ^ n889 ;
  assign n46642 = n39105 ^ n21062 ^ n12977 ;
  assign n46643 = ( n7997 & n15532 ) | ( n7997 & n46642 ) | ( n15532 & n46642 ) ;
  assign n46641 = n25793 ^ n15117 ^ n317 ;
  assign n46645 = n46644 ^ n46643 ^ n46641 ;
  assign n46646 = ( n11237 & n27662 ) | ( n11237 & ~n45645 ) | ( n27662 & ~n45645 ) ;
  assign n46647 = n40632 ^ n15246 ^ n7851 ;
  assign n46648 = ( n7734 & n46646 ) | ( n7734 & n46647 ) | ( n46646 & n46647 ) ;
  assign n46650 = n20954 ^ n17912 ^ n9931 ;
  assign n46649 = n1258 & n11442 ;
  assign n46651 = n46650 ^ n46649 ^ 1'b0 ;
  assign n46652 = n36179 ^ n23752 ^ n16192 ;
  assign n46653 = n36022 ^ n24009 ^ n4636 ;
  assign n46654 = ( n5654 & n41360 ) | ( n5654 & n46653 ) | ( n41360 & n46653 ) ;
  assign n46655 = n12640 ^ n9664 ^ 1'b0 ;
  assign n46656 = n46655 ^ n21996 ^ n15340 ;
  assign n46657 = ( x63 & n27797 ) | ( x63 & n44642 ) | ( n27797 & n44642 ) ;
  assign n46658 = ~n22736 & n46657 ;
  assign n46659 = n46067 ^ n8473 ^ n3479 ;
  assign n46660 = n35383 & n42941 ;
  assign n46661 = n770 & n46660 ;
  assign n46662 = ( n6734 & n14224 ) | ( n6734 & n46661 ) | ( n14224 & n46661 ) ;
  assign n46663 = ( n384 & n46659 ) | ( n384 & ~n46662 ) | ( n46659 & ~n46662 ) ;
  assign n46664 = n2311 & n43886 ;
  assign n46665 = ~x13 & n46664 ;
  assign n46668 = n28716 ^ n16573 ^ n9000 ;
  assign n46667 = ( n6198 & ~n32662 ) | ( n6198 & n39232 ) | ( ~n32662 & n39232 ) ;
  assign n46666 = ( ~n10024 & n24666 ) | ( ~n10024 & n27256 ) | ( n24666 & n27256 ) ;
  assign n46669 = n46668 ^ n46667 ^ n46666 ;
  assign n46670 = n19544 ^ n15156 ^ n1950 ;
  assign n46673 = ( ~n7272 & n40235 ) | ( ~n7272 & n43685 ) | ( n40235 & n43685 ) ;
  assign n46671 = ~n18258 & n24031 ;
  assign n46672 = n46671 ^ n21853 ^ 1'b0 ;
  assign n46674 = n46673 ^ n46672 ^ n26693 ;
  assign n46675 = ( ~n6552 & n9715 ) | ( ~n6552 & n26987 ) | ( n9715 & n26987 ) ;
  assign n46676 = n14220 & n28399 ;
  assign n46677 = n46676 ^ n10765 ^ 1'b0 ;
  assign n46678 = n414 & n46677 ;
  assign n46679 = n27902 & ~n44083 ;
  assign n46680 = n968 | n11552 ;
  assign n46681 = n46680 ^ n17376 ^ 1'b0 ;
  assign n46682 = n46681 ^ n38107 ^ n11604 ;
  assign n46684 = ( n4446 & n22181 ) | ( n4446 & n25593 ) | ( n22181 & n25593 ) ;
  assign n46685 = n46684 ^ n37285 ^ n21125 ;
  assign n46683 = ~n1492 & n35104 ;
  assign n46686 = n46685 ^ n46683 ^ 1'b0 ;
  assign n46687 = n12668 ^ n10865 ^ 1'b0 ;
  assign n46688 = n46687 ^ n11216 ^ n5550 ;
  assign n46689 = ( ~n17366 & n32816 ) | ( ~n17366 & n46688 ) | ( n32816 & n46688 ) ;
  assign n46690 = n46689 ^ n46346 ^ n2777 ;
  assign n46691 = n34139 ^ n20148 ^ n11912 ;
  assign n46692 = ( ~n8811 & n18535 ) | ( ~n8811 & n25257 ) | ( n18535 & n25257 ) ;
  assign n46693 = n46692 ^ n21599 ^ n11314 ;
  assign n46694 = n46693 ^ n24246 ^ n19397 ;
  assign n46695 = n46694 ^ n26829 ^ n14410 ;
  assign n46696 = n46695 ^ n44387 ^ n13075 ;
  assign n46699 = ( n7199 & n17743 ) | ( n7199 & ~n21207 ) | ( n17743 & ~n21207 ) ;
  assign n46700 = n32328 ^ n4688 ^ n1406 ;
  assign n46701 = ( n18199 & ~n46699 ) | ( n18199 & n46700 ) | ( ~n46699 & n46700 ) ;
  assign n46697 = ~n16965 & n19650 ;
  assign n46698 = n46697 ^ n22581 ^ 1'b0 ;
  assign n46702 = n46701 ^ n46698 ^ n38685 ;
  assign n46703 = ( ~n9748 & n13631 ) | ( ~n9748 & n29665 ) | ( n13631 & n29665 ) ;
  assign n46704 = ( ~n2966 & n42552 ) | ( ~n2966 & n46703 ) | ( n42552 & n46703 ) ;
  assign n46706 = n13828 & n19501 ;
  assign n46707 = n17526 & n46706 ;
  assign n46705 = ( n14802 & n20016 ) | ( n14802 & n30295 ) | ( n20016 & n30295 ) ;
  assign n46708 = n46707 ^ n46705 ^ n44778 ;
  assign n46709 = n17294 & n29985 ;
  assign n46713 = n5674 & ~n14540 ;
  assign n46710 = n30504 ^ n27788 ^ n5772 ;
  assign n46711 = n46710 ^ n39906 ^ n19614 ;
  assign n46712 = n27229 & ~n46711 ;
  assign n46714 = n46713 ^ n46712 ^ 1'b0 ;
  assign n46715 = n27862 ^ n12931 ^ 1'b0 ;
  assign n46716 = n41396 ^ n33371 ^ 1'b0 ;
  assign n46717 = n33001 & ~n46716 ;
  assign n46718 = n45866 ^ n17737 ^ n16497 ;
  assign n46719 = ( ~n3848 & n19483 ) | ( ~n3848 & n33527 ) | ( n19483 & n33527 ) ;
  assign n46720 = n46719 ^ n45732 ^ n42276 ;
  assign n46721 = n13218 & ~n45111 ;
  assign n46722 = n46721 ^ n39708 ^ 1'b0 ;
  assign n46723 = n23592 & ~n29578 ;
  assign n46724 = n46723 ^ n18766 ^ 1'b0 ;
  assign n46725 = ( n12769 & ~n38490 ) | ( n12769 & n46724 ) | ( ~n38490 & n46724 ) ;
  assign n46726 = n46725 ^ n39692 ^ n27785 ;
  assign n46727 = n46726 ^ n32607 ^ n4159 ;
  assign n46728 = n40026 ^ n25942 ^ n748 ;
  assign n46729 = n46728 ^ n35019 ^ n20860 ;
  assign n46730 = n6757 & ~n11420 ;
  assign n46731 = n46730 ^ n26288 ^ 1'b0 ;
  assign n46732 = ( ~n3375 & n5512 ) | ( ~n3375 & n28497 ) | ( n5512 & n28497 ) ;
  assign n46733 = n39711 ^ n15603 ^ 1'b0 ;
  assign n46734 = n46733 ^ n42566 ^ n32170 ;
  assign n46735 = n38175 ^ n23970 ^ n10718 ;
  assign n46736 = n38742 ^ n19258 ^ n7514 ;
  assign n46737 = ( n17983 & ~n46735 ) | ( n17983 & n46736 ) | ( ~n46735 & n46736 ) ;
  assign n46738 = n35319 ^ n34052 ^ n20991 ;
  assign n46739 = ( n29517 & n42715 ) | ( n29517 & n43093 ) | ( n42715 & n43093 ) ;
  assign n46740 = n46739 ^ n10786 ^ n6602 ;
  assign n46741 = ~n4315 & n30866 ;
  assign n46742 = n46741 ^ n13276 ^ 1'b0 ;
  assign n46743 = ( n9073 & ~n23713 ) | ( n9073 & n39214 ) | ( ~n23713 & n39214 ) ;
  assign n46744 = n37528 ^ n22210 ^ n7278 ;
  assign n46745 = ( n5889 & ~n46743 ) | ( n5889 & n46744 ) | ( ~n46743 & n46744 ) ;
  assign n46746 = ( n310 & n26532 ) | ( n310 & n46745 ) | ( n26532 & n46745 ) ;
  assign n46747 = ( n14360 & n19731 ) | ( n14360 & n29956 ) | ( n19731 & n29956 ) ;
  assign n46748 = ( n2659 & ~n28094 ) | ( n2659 & n29374 ) | ( ~n28094 & n29374 ) ;
  assign n46749 = n27500 ^ n25303 ^ n8003 ;
  assign n46750 = n46749 ^ n11156 ^ 1'b0 ;
  assign n46751 = n46750 ^ n45396 ^ n30283 ;
  assign n46753 = ( ~n19754 & n20586 ) | ( ~n19754 & n26644 ) | ( n20586 & n26644 ) ;
  assign n46754 = n46753 ^ x75 ^ 1'b0 ;
  assign n46755 = n19735 & n46754 ;
  assign n46752 = n30016 ^ n924 ^ 1'b0 ;
  assign n46756 = n46755 ^ n46752 ^ n16106 ;
  assign n46757 = ( ~n7457 & n8090 ) | ( ~n7457 & n46756 ) | ( n8090 & n46756 ) ;
  assign n46759 = n30643 ^ n21859 ^ n17408 ;
  assign n46758 = ( ~n12407 & n21790 ) | ( ~n12407 & n41956 ) | ( n21790 & n41956 ) ;
  assign n46760 = n46759 ^ n46758 ^ n13989 ;
  assign n46762 = ( n816 & n5234 ) | ( n816 & ~n12470 ) | ( n5234 & ~n12470 ) ;
  assign n46763 = n46762 ^ n31434 ^ n11647 ;
  assign n46761 = n37083 ^ n31082 ^ n14423 ;
  assign n46764 = n46763 ^ n46761 ^ n26926 ;
  assign n46765 = n283 & ~n12099 ;
  assign n46766 = ~n39853 & n46765 ;
  assign n46771 = ( n9162 & n19923 ) | ( n9162 & ~n44786 ) | ( n19923 & ~n44786 ) ;
  assign n46767 = ( n1534 & ~n8721 ) | ( n1534 & n14829 ) | ( ~n8721 & n14829 ) ;
  assign n46768 = n46767 ^ n1099 ^ 1'b0 ;
  assign n46769 = n37637 & n46768 ;
  assign n46770 = ~n25187 & n46769 ;
  assign n46772 = n46771 ^ n46770 ^ 1'b0 ;
  assign n46774 = n40656 ^ n34148 ^ 1'b0 ;
  assign n46775 = n32452 & ~n46774 ;
  assign n46773 = ~n8384 & n22065 ;
  assign n46776 = n46775 ^ n46773 ^ n12067 ;
  assign n46777 = n20348 ^ n7367 ^ 1'b0 ;
  assign n46778 = n46777 ^ n40540 ^ n18645 ;
  assign n46779 = ( n3093 & ~n26843 ) | ( n3093 & n33732 ) | ( ~n26843 & n33732 ) ;
  assign n46780 = n45627 ^ n27650 ^ n5174 ;
  assign n46781 = n46780 ^ n16893 ^ n452 ;
  assign n46782 = n46781 ^ n34986 ^ n3184 ;
  assign n46783 = n23795 ^ n21574 ^ n9412 ;
  assign n46784 = n46783 ^ n35838 ^ n30579 ;
  assign n46785 = n38443 ^ n10822 ^ n1471 ;
  assign n46786 = n40363 & ~n46785 ;
  assign n46787 = n24416 ^ n16028 ^ 1'b0 ;
  assign n46788 = n17788 | n46787 ;
  assign n46789 = ( ~n2757 & n8348 ) | ( ~n2757 & n46788 ) | ( n8348 & n46788 ) ;
  assign n46790 = ( n14549 & ~n16003 ) | ( n14549 & n39367 ) | ( ~n16003 & n39367 ) ;
  assign n46791 = n46790 ^ n18848 ^ n16570 ;
  assign n46792 = n15455 | n31862 ;
  assign n46794 = n44962 ^ n17481 ^ n4224 ;
  assign n46793 = n28695 & ~n38913 ;
  assign n46795 = n46794 ^ n46793 ^ 1'b0 ;
  assign n46796 = ( n4305 & n12682 ) | ( n4305 & n45886 ) | ( n12682 & n45886 ) ;
  assign n46797 = n46796 ^ n21735 ^ 1'b0 ;
  assign n46798 = n28091 ^ n20817 ^ n9570 ;
  assign n46799 = ( n15530 & ~n20995 ) | ( n15530 & n46798 ) | ( ~n20995 & n46798 ) ;
  assign n46800 = n46799 ^ n41654 ^ n2362 ;
  assign n46801 = n34921 ^ n27316 ^ n23274 ;
  assign n46802 = ~n1111 & n13827 ;
  assign n46803 = n46802 ^ n44572 ^ n31720 ;
  assign n46804 = ( n5039 & n8452 ) | ( n5039 & ~n46803 ) | ( n8452 & ~n46803 ) ;
  assign n46805 = ( n6257 & ~n12462 ) | ( n6257 & n41616 ) | ( ~n12462 & n41616 ) ;
  assign n46806 = n26184 ^ n25267 ^ n9178 ;
  assign n46807 = ( n3988 & n10257 ) | ( n3988 & ~n36988 ) | ( n10257 & ~n36988 ) ;
  assign n46808 = ( n3671 & n42099 ) | ( n3671 & ~n46807 ) | ( n42099 & ~n46807 ) ;
  assign n46809 = ( n19717 & n39108 ) | ( n19717 & n46808 ) | ( n39108 & n46808 ) ;
  assign n46810 = ( n3065 & ~n21374 ) | ( n3065 & n26661 ) | ( ~n21374 & n26661 ) ;
  assign n46811 = ( x46 & ~n40643 ) | ( x46 & n46810 ) | ( ~n40643 & n46810 ) ;
  assign n46812 = n25118 ^ n10557 ^ 1'b0 ;
  assign n46813 = n35840 & n46812 ;
  assign n46814 = n14250 | n25872 ;
  assign n46815 = ( n1109 & n6626 ) | ( n1109 & ~n30784 ) | ( n6626 & ~n30784 ) ;
  assign n46816 = ( n17451 & ~n27852 ) | ( n17451 & n38189 ) | ( ~n27852 & n38189 ) ;
  assign n46817 = n15969 ^ n8454 ^ n6328 ;
  assign n46818 = n46817 ^ n15793 ^ n4588 ;
  assign n46819 = n38764 & n46818 ;
  assign n46820 = n46819 ^ n16573 ^ 1'b0 ;
  assign n46821 = ( n13779 & ~n24400 ) | ( n13779 & n46820 ) | ( ~n24400 & n46820 ) ;
  assign n46822 = ( n30869 & n46816 ) | ( n30869 & n46821 ) | ( n46816 & n46821 ) ;
  assign n46823 = n26069 & n43357 ;
  assign n46824 = n35310 ^ n23173 ^ n18723 ;
  assign n46825 = ( n17267 & n44075 ) | ( n17267 & n46824 ) | ( n44075 & n46824 ) ;
  assign n46827 = ( n16309 & n22065 ) | ( n16309 & ~n27638 ) | ( n22065 & ~n27638 ) ;
  assign n46826 = n2773 | n13808 ;
  assign n46828 = n46827 ^ n46826 ^ 1'b0 ;
  assign n46829 = n14894 ^ n5844 ^ n1252 ;
  assign n46830 = ( n12232 & n46828 ) | ( n12232 & n46829 ) | ( n46828 & n46829 ) ;
  assign n46831 = ( n3398 & n41961 ) | ( n3398 & n46830 ) | ( n41961 & n46830 ) ;
  assign n46834 = ( ~n26374 & n26880 ) | ( ~n26374 & n41389 ) | ( n26880 & n41389 ) ;
  assign n46832 = ( n14825 & n17561 ) | ( n14825 & n30027 ) | ( n17561 & n30027 ) ;
  assign n46833 = n46832 ^ n16762 ^ n6952 ;
  assign n46835 = n46834 ^ n46833 ^ n34362 ;
  assign n46836 = n17699 ^ n5473 ^ 1'b0 ;
  assign n46837 = ( n4371 & ~n5539 ) | ( n4371 & n46836 ) | ( ~n5539 & n46836 ) ;
  assign n46838 = n46837 ^ n33981 ^ 1'b0 ;
  assign n46839 = n3450 & n3620 ;
  assign n46840 = n46838 & n46839 ;
  assign n46841 = n46840 ^ n24059 ^ n1648 ;
  assign n46843 = ( n1638 & ~n18502 ) | ( n1638 & n41688 ) | ( ~n18502 & n41688 ) ;
  assign n46842 = n19766 & ~n31552 ;
  assign n46844 = n46843 ^ n46842 ^ 1'b0 ;
  assign n46845 = ~n26594 & n41259 ;
  assign n46846 = n46844 & n46845 ;
  assign n46847 = n39495 ^ n18562 ^ n9541 ;
  assign n46848 = n46847 ^ n34458 ^ n4041 ;
  assign n46849 = n22682 ^ n14941 ^ n9375 ;
  assign n46850 = ( ~n3873 & n18280 ) | ( ~n3873 & n18580 ) | ( n18280 & n18580 ) ;
  assign n46851 = ( n42009 & n46849 ) | ( n42009 & ~n46850 ) | ( n46849 & ~n46850 ) ;
  assign n46852 = ( ~n23767 & n46848 ) | ( ~n23767 & n46851 ) | ( n46848 & n46851 ) ;
  assign n46853 = n32486 ^ n20397 ^ n14281 ;
  assign n46854 = n46853 ^ n20360 ^ n17161 ;
  assign n46855 = ( n27374 & n44753 ) | ( n27374 & ~n46089 ) | ( n44753 & ~n46089 ) ;
  assign n46856 = n10438 ^ n3303 ^ 1'b0 ;
  assign n46857 = n8483 | n46856 ;
  assign n46858 = n46857 ^ n12725 ^ 1'b0 ;
  assign n46859 = n20220 & ~n22294 ;
  assign n46860 = n46859 ^ n27477 ^ 1'b0 ;
  assign n46861 = n46860 ^ n39067 ^ n8162 ;
  assign n46862 = ( ~n28632 & n39173 ) | ( ~n28632 & n41478 ) | ( n39173 & n41478 ) ;
  assign n46863 = ( n8115 & n16345 ) | ( n8115 & ~n18245 ) | ( n16345 & ~n18245 ) ;
  assign n46864 = ~n8306 & n46863 ;
  assign n46865 = ~n28718 & n46864 ;
  assign n46866 = n20617 ^ n20223 ^ n12471 ;
  assign n46867 = n46866 ^ n45021 ^ n28916 ;
  assign n46868 = n46867 ^ n46599 ^ n34429 ;
  assign n46869 = ( n12283 & n16815 ) | ( n12283 & ~n21946 ) | ( n16815 & ~n21946 ) ;
  assign n46870 = n27368 | n38903 ;
  assign n46871 = n46870 ^ n25581 ^ 1'b0 ;
  assign n46872 = ( n8848 & ~n22637 ) | ( n8848 & n35778 ) | ( ~n22637 & n35778 ) ;
  assign n46873 = ( ~n46869 & n46871 ) | ( ~n46869 & n46872 ) | ( n46871 & n46872 ) ;
  assign n46874 = ( n6259 & ~n20676 ) | ( n6259 & n24904 ) | ( ~n20676 & n24904 ) ;
  assign n46876 = ( n11214 & n13680 ) | ( n11214 & ~n33880 ) | ( n13680 & ~n33880 ) ;
  assign n46875 = n42799 ^ n37083 ^ n9146 ;
  assign n46877 = n46876 ^ n46875 ^ n38873 ;
  assign n46878 = ( ~n15867 & n46874 ) | ( ~n15867 & n46877 ) | ( n46874 & n46877 ) ;
  assign n46879 = ~n24424 & n30071 ;
  assign n46880 = ( ~x222 & n3047 ) | ( ~x222 & n14807 ) | ( n3047 & n14807 ) ;
  assign n46881 = ( n12724 & ~n21018 ) | ( n12724 & n24321 ) | ( ~n21018 & n24321 ) ;
  assign n46882 = ( ~n37866 & n44568 ) | ( ~n37866 & n46881 ) | ( n44568 & n46881 ) ;
  assign n46883 = n42753 ^ n21610 ^ 1'b0 ;
  assign n46884 = n2298 | n46883 ;
  assign n46885 = n46884 ^ n11701 ^ n10903 ;
  assign n46886 = n18428 & ~n36547 ;
  assign n46887 = n7960 & n46886 ;
  assign n46888 = n6069 & n40626 ;
  assign n46889 = n46888 ^ n15081 ^ 1'b0 ;
  assign n46890 = n41722 ^ n34054 ^ n24699 ;
  assign n46891 = n36267 ^ n20511 ^ n11317 ;
  assign n46892 = ( n356 & ~n9059 ) | ( n356 & n46891 ) | ( ~n9059 & n46891 ) ;
  assign n46893 = n11982 ^ n1161 ^ 1'b0 ;
  assign n46894 = ( n18987 & ~n46892 ) | ( n18987 & n46893 ) | ( ~n46892 & n46893 ) ;
  assign n46897 = ( n12590 & n29521 ) | ( n12590 & n37971 ) | ( n29521 & n37971 ) ;
  assign n46895 = n40922 ^ n8288 ^ n2935 ;
  assign n46896 = ( ~n2395 & n18557 ) | ( ~n2395 & n46895 ) | ( n18557 & n46895 ) ;
  assign n46898 = n46897 ^ n46896 ^ 1'b0 ;
  assign n46899 = n11801 ^ n8394 ^ 1'b0 ;
  assign n46900 = ( n3803 & n13960 ) | ( n3803 & n37881 ) | ( n13960 & n37881 ) ;
  assign n46901 = ( n30105 & n46899 ) | ( n30105 & ~n46900 ) | ( n46899 & ~n46900 ) ;
  assign n46905 = n17204 ^ n6044 ^ 1'b0 ;
  assign n46906 = ~n6827 & n46905 ;
  assign n46904 = n20517 ^ n16535 ^ n1397 ;
  assign n46907 = n46906 ^ n46904 ^ n4082 ;
  assign n46902 = n22263 ^ n4959 ^ x128 ;
  assign n46903 = ( n21140 & n25855 ) | ( n21140 & ~n46902 ) | ( n25855 & ~n46902 ) ;
  assign n46908 = n46907 ^ n46903 ^ n19324 ;
  assign n46910 = ( n3149 & ~n15561 ) | ( n3149 & n28184 ) | ( ~n15561 & n28184 ) ;
  assign n46911 = ( n3631 & n11715 ) | ( n3631 & n46910 ) | ( n11715 & n46910 ) ;
  assign n46909 = n5198 & ~n41988 ;
  assign n46912 = n46911 ^ n46909 ^ 1'b0 ;
  assign n46913 = ( n5768 & n20104 ) | ( n5768 & n34609 ) | ( n20104 & n34609 ) ;
  assign n46914 = n24514 ^ n6511 ^ n1208 ;
  assign n46915 = n46914 ^ n27564 ^ n446 ;
  assign n46916 = ( n31734 & n33730 ) | ( n31734 & n45074 ) | ( n33730 & n45074 ) ;
  assign n46917 = n46916 ^ n43642 ^ n1075 ;
  assign n46918 = n31857 ^ n18719 ^ n17567 ;
  assign n46920 = n11795 ^ n6993 ^ n2662 ;
  assign n46921 = ( n9217 & ~n22871 ) | ( n9217 & n46920 ) | ( ~n22871 & n46920 ) ;
  assign n46919 = ( n1678 & ~n8121 ) | ( n1678 & n26792 ) | ( ~n8121 & n26792 ) ;
  assign n46922 = n46921 ^ n46919 ^ n4589 ;
  assign n46923 = n2967 & ~n13660 ;
  assign n46924 = n46923 ^ n14089 ^ 1'b0 ;
  assign n46925 = n21278 | n46924 ;
  assign n46926 = n46925 ^ n12302 ^ 1'b0 ;
  assign n46927 = n46926 ^ n28612 ^ n19820 ;
  assign n46928 = ( ~n13375 & n27863 ) | ( ~n13375 & n40252 ) | ( n27863 & n40252 ) ;
  assign n46929 = ( n16050 & ~n21190 ) | ( n16050 & n46928 ) | ( ~n21190 & n46928 ) ;
  assign n46930 = n45368 ^ n7615 ^ 1'b0 ;
  assign n46931 = n14250 ^ n7786 ^ n2033 ;
  assign n46932 = n15269 ^ n4038 ^ n1416 ;
  assign n46933 = ( n6454 & n10024 ) | ( n6454 & n10952 ) | ( n10024 & n10952 ) ;
  assign n46934 = n46933 ^ n32834 ^ n17975 ;
  assign n46935 = ( n433 & n2380 ) | ( n433 & n5599 ) | ( n2380 & n5599 ) ;
  assign n46936 = n40893 ^ n29366 ^ n11693 ;
  assign n46937 = ( ~n22961 & n46935 ) | ( ~n22961 & n46936 ) | ( n46935 & n46936 ) ;
  assign n46938 = ( ~n7800 & n41956 ) | ( ~n7800 & n46937 ) | ( n41956 & n46937 ) ;
  assign n46939 = ( n46932 & n46934 ) | ( n46932 & ~n46938 ) | ( n46934 & ~n46938 ) ;
  assign n46940 = ( n904 & n2479 ) | ( n904 & n18714 ) | ( n2479 & n18714 ) ;
  assign n46941 = n41691 & n46940 ;
  assign n46942 = ~n4149 & n18727 ;
  assign n46943 = ( n4858 & n25348 ) | ( n4858 & ~n46942 ) | ( n25348 & ~n46942 ) ;
  assign n46944 = n46943 ^ n43723 ^ n42891 ;
  assign n46945 = ( n2893 & ~n19527 ) | ( n2893 & n19541 ) | ( ~n19527 & n19541 ) ;
  assign n46946 = n46945 ^ n13119 ^ n4287 ;
  assign n46947 = ( ~n22927 & n27014 ) | ( ~n22927 & n43375 ) | ( n27014 & n43375 ) ;
  assign n46948 = n5472 & ~n46947 ;
  assign n46949 = n14681 & n46948 ;
  assign n46950 = n24857 & ~n46949 ;
  assign n46951 = n4312 & ~n26147 ;
  assign n46952 = ~n29788 & n46951 ;
  assign n46953 = ( n8535 & n17887 ) | ( n8535 & n21412 ) | ( n17887 & n21412 ) ;
  assign n46954 = n16099 & ~n46953 ;
  assign n46955 = n46952 & n46954 ;
  assign n46956 = ~n10970 & n21953 ;
  assign n46957 = n46956 ^ n8785 ^ 1'b0 ;
  assign n46958 = n46957 ^ n1288 ^ 1'b0 ;
  assign n46959 = ( n4368 & n4457 ) | ( n4368 & ~n34217 ) | ( n4457 & ~n34217 ) ;
  assign n46960 = n5685 & ~n26303 ;
  assign n46961 = n46960 ^ n1277 ^ 1'b0 ;
  assign n46962 = n46961 ^ n4155 ^ 1'b0 ;
  assign n46963 = n46962 ^ n21017 ^ n15720 ;
  assign n46964 = n42805 ^ n21703 ^ n4020 ;
  assign n46965 = ~n11133 & n28268 ;
  assign n46966 = n42943 ^ n23280 ^ n11134 ;
  assign n46967 = n7955 & ~n12491 ;
  assign n46968 = ~n6787 & n20260 ;
  assign n46969 = ~n46967 & n46968 ;
  assign n46970 = n23399 ^ n5447 ^ 1'b0 ;
  assign n46971 = ( n5056 & n18110 ) | ( n5056 & n29471 ) | ( n18110 & n29471 ) ;
  assign n46972 = ( ~n36305 & n42614 ) | ( ~n36305 & n46971 ) | ( n42614 & n46971 ) ;
  assign n46977 = n14238 ^ n10407 ^ 1'b0 ;
  assign n46978 = n1969 & n46977 ;
  assign n46976 = ~n11558 & n22062 ;
  assign n46979 = n46978 ^ n46976 ^ 1'b0 ;
  assign n46973 = ( ~n11655 & n14984 ) | ( ~n11655 & n21157 ) | ( n14984 & n21157 ) ;
  assign n46974 = n46973 ^ n23321 ^ n16226 ;
  assign n46975 = ( ~n10378 & n19578 ) | ( ~n10378 & n46974 ) | ( n19578 & n46974 ) ;
  assign n46980 = n46979 ^ n46975 ^ n9233 ;
  assign n46981 = n18259 ^ n15612 ^ n11481 ;
  assign n46982 = n41564 ^ n9782 ^ n8012 ;
  assign n46983 = n46982 ^ n23772 ^ n756 ;
  assign n46984 = ( n8217 & n39408 ) | ( n8217 & ~n46983 ) | ( n39408 & ~n46983 ) ;
  assign n46985 = n46984 ^ n26140 ^ 1'b0 ;
  assign n46986 = n19663 ^ n9797 ^ n4680 ;
  assign n46987 = ( ~n4393 & n13603 ) | ( ~n4393 & n33216 ) | ( n13603 & n33216 ) ;
  assign n46988 = n32443 ^ n22230 ^ 1'b0 ;
  assign n46989 = n46988 ^ n46373 ^ n14147 ;
  assign n46990 = ( ~n3721 & n36112 ) | ( ~n3721 & n37858 ) | ( n36112 & n37858 ) ;
  assign n46991 = n31135 ^ n17241 ^ n4662 ;
  assign n46992 = ( n2190 & n8253 ) | ( n2190 & ~n46991 ) | ( n8253 & ~n46991 ) ;
  assign n46993 = n14235 & ~n37107 ;
  assign n46994 = ~n46992 & n46993 ;
  assign n46998 = ( n16583 & n31234 ) | ( n16583 & n40351 ) | ( n31234 & n40351 ) ;
  assign n46995 = ( n840 & n1174 ) | ( n840 & ~n11598 ) | ( n1174 & ~n11598 ) ;
  assign n46996 = n46995 ^ n41739 ^ n5880 ;
  assign n46997 = ( n23206 & ~n32860 ) | ( n23206 & n46996 ) | ( ~n32860 & n46996 ) ;
  assign n46999 = n46998 ^ n46997 ^ n26538 ;
  assign n47000 = ( n33494 & n45346 ) | ( n33494 & n46999 ) | ( n45346 & n46999 ) ;
  assign n47001 = ( n6100 & n6168 ) | ( n6100 & n28213 ) | ( n6168 & n28213 ) ;
  assign n47002 = n47001 ^ n15955 ^ n5725 ;
  assign n47003 = ( n2774 & ~n40758 ) | ( n2774 & n47002 ) | ( ~n40758 & n47002 ) ;
  assign n47004 = n4789 & n19123 ;
  assign n47005 = ~n21486 & n47004 ;
  assign n47006 = n47005 ^ n15486 ^ n8425 ;
  assign n47007 = n33315 ^ n10676 ^ n5660 ;
  assign n47008 = n47007 ^ n26239 ^ n17519 ;
  assign n47009 = ( ~n4681 & n10013 ) | ( ~n4681 & n22671 ) | ( n10013 & n22671 ) ;
  assign n47010 = ( n3508 & n16092 ) | ( n3508 & n47009 ) | ( n16092 & n47009 ) ;
  assign n47011 = ( ~n9079 & n10118 ) | ( ~n9079 & n25148 ) | ( n10118 & n25148 ) ;
  assign n47012 = n31339 ^ n19373 ^ n3265 ;
  assign n47013 = ( n28021 & n35043 ) | ( n28021 & n47012 ) | ( n35043 & n47012 ) ;
  assign n47014 = n14511 ^ n6734 ^ 1'b0 ;
  assign n47015 = n21252 | n47014 ;
  assign n47016 = ( n7467 & n15319 ) | ( n7467 & ~n16572 ) | ( n15319 & ~n16572 ) ;
  assign n47017 = ( n7783 & ~n24928 ) | ( n7783 & n36290 ) | ( ~n24928 & n36290 ) ;
  assign n47018 = n47017 ^ n41665 ^ 1'b0 ;
  assign n47019 = n47016 & n47018 ;
  assign n47023 = ( n5156 & n10976 ) | ( n5156 & ~n44417 ) | ( n10976 & ~n44417 ) ;
  assign n47022 = ( n15197 & n30583 ) | ( n15197 & n35422 ) | ( n30583 & n35422 ) ;
  assign n47020 = n38095 ^ n30050 ^ n12011 ;
  assign n47021 = n47020 ^ n31802 ^ n25472 ;
  assign n47024 = n47023 ^ n47022 ^ n47021 ;
  assign n47025 = n4564 ^ n2477 ^ n1515 ;
  assign n47026 = n47025 ^ n22953 ^ 1'b0 ;
  assign n47027 = n43044 ^ n12097 ^ n9258 ;
  assign n47028 = n24815 ^ n20084 ^ n1528 ;
  assign n47029 = ( n5136 & n29973 ) | ( n5136 & n35978 ) | ( n29973 & n35978 ) ;
  assign n47030 = ~n11440 & n19981 ;
  assign n47031 = ~n12343 & n47030 ;
  assign n47032 = n16341 ^ n14944 ^ n10752 ;
  assign n47033 = ( x134 & n27079 ) | ( x134 & ~n47032 ) | ( n27079 & ~n47032 ) ;
  assign n47034 = ( n1337 & n40127 ) | ( n1337 & ~n47033 ) | ( n40127 & ~n47033 ) ;
  assign n47035 = n47034 ^ n45237 ^ n40314 ;
  assign n47036 = n44565 ^ n25465 ^ n17143 ;
  assign n47037 = ( n8460 & ~n38019 ) | ( n8460 & n47036 ) | ( ~n38019 & n47036 ) ;
  assign n47038 = n3103 & n6933 ;
  assign n47039 = ( n3500 & n18724 ) | ( n3500 & ~n47038 ) | ( n18724 & ~n47038 ) ;
  assign n47040 = n47039 ^ n10440 ^ n6715 ;
  assign n47041 = n41276 ^ n25861 ^ n11494 ;
  assign n47042 = n37733 ^ n5118 ^ n4872 ;
  assign n47043 = n47042 ^ n22988 ^ 1'b0 ;
  assign n47044 = ( n7306 & n23977 ) | ( n7306 & ~n44666 ) | ( n23977 & ~n44666 ) ;
  assign n47045 = ( n12308 & ~n13919 ) | ( n12308 & n35946 ) | ( ~n13919 & n35946 ) ;
  assign n47046 = n3499 | n11191 ;
  assign n47047 = n47046 ^ n12542 ^ 1'b0 ;
  assign n47048 = ( ~n12767 & n14653 ) | ( ~n12767 & n38700 ) | ( n14653 & n38700 ) ;
  assign n47049 = n15445 | n47048 ;
  assign n47050 = n42813 | n47049 ;
  assign n47051 = n42044 ^ n23167 ^ n12376 ;
  assign n47052 = ( n14237 & n19877 ) | ( n14237 & n47051 ) | ( n19877 & n47051 ) ;
  assign n47053 = n34520 ^ n32019 ^ n7249 ;
  assign n47054 = ( n12979 & n12993 ) | ( n12979 & n34143 ) | ( n12993 & n34143 ) ;
  assign n47055 = n43372 ^ n41168 ^ n10070 ;
  assign n47056 = n47055 ^ n35815 ^ n24282 ;
  assign n47057 = n10321 & ~n37158 ;
  assign n47058 = n47057 ^ n4463 ^ 1'b0 ;
  assign n47059 = n47058 ^ n24606 ^ n5573 ;
  assign n47060 = n41223 ^ n16460 ^ n8511 ;
  assign n47061 = n28058 ^ n20610 ^ 1'b0 ;
  assign n47062 = ~n47060 & n47061 ;
  assign n47063 = n47062 ^ n4453 ^ 1'b0 ;
  assign n47064 = ( n1021 & n5791 ) | ( n1021 & n17989 ) | ( n5791 & n17989 ) ;
  assign n47065 = n47064 ^ n4182 ^ 1'b0 ;
  assign n47066 = n9169 | n45478 ;
  assign n47067 = ( n3781 & n11354 ) | ( n3781 & n18934 ) | ( n11354 & n18934 ) ;
  assign n47068 = n27567 ^ n13708 ^ n7390 ;
  assign n47069 = ( ~n12673 & n47067 ) | ( ~n12673 & n47068 ) | ( n47067 & n47068 ) ;
  assign n47070 = n44707 ^ n650 ^ 1'b0 ;
  assign n47071 = ~n29212 & n47070 ;
  assign n47072 = ( ~n2657 & n17463 ) | ( ~n2657 & n31437 ) | ( n17463 & n31437 ) ;
  assign n47073 = n47072 ^ n44746 ^ 1'b0 ;
  assign n47074 = ( n31771 & ~n47071 ) | ( n31771 & n47073 ) | ( ~n47071 & n47073 ) ;
  assign n47075 = n18741 ^ n12279 ^ n7012 ;
  assign n47076 = ( n11346 & n42119 ) | ( n11346 & ~n47075 ) | ( n42119 & ~n47075 ) ;
  assign n47077 = n47076 ^ n31338 ^ n15593 ;
  assign n47078 = ( n2859 & ~n9953 ) | ( n2859 & n47077 ) | ( ~n9953 & n47077 ) ;
  assign n47079 = n14643 ^ n12094 ^ 1'b0 ;
  assign n47080 = n47079 ^ n46866 ^ n40658 ;
  assign n47081 = n34168 ^ n29661 ^ n3269 ;
  assign n47082 = ( n8334 & n16926 ) | ( n8334 & ~n42365 ) | ( n16926 & ~n42365 ) ;
  assign n47084 = n9324 ^ n4696 ^ n1783 ;
  assign n47085 = n47084 ^ n28397 ^ n1236 ;
  assign n47083 = n38796 ^ n19961 ^ 1'b0 ;
  assign n47086 = n47085 ^ n47083 ^ n28293 ;
  assign n47088 = n19714 ^ n3244 ^ n599 ;
  assign n47089 = n47088 ^ n20503 ^ n6038 ;
  assign n47090 = ( n17635 & ~n34211 ) | ( n17635 & n47089 ) | ( ~n34211 & n47089 ) ;
  assign n47091 = n47090 ^ n28531 ^ n2492 ;
  assign n47087 = n5820 & n19146 ;
  assign n47092 = n47091 ^ n47087 ^ 1'b0 ;
  assign n47093 = ( n3171 & n17787 ) | ( n3171 & n21434 ) | ( n17787 & n21434 ) ;
  assign n47094 = n47093 ^ n7755 ^ n7202 ;
  assign n47095 = n47094 ^ n45387 ^ n34511 ;
  assign n47096 = n7049 & n32931 ;
  assign n47097 = n47096 ^ n11262 ^ 1'b0 ;
  assign n47098 = ( n19421 & n33303 ) | ( n19421 & ~n47097 ) | ( n33303 & ~n47097 ) ;
  assign n47099 = ( ~n12749 & n26425 ) | ( ~n12749 & n37132 ) | ( n26425 & n37132 ) ;
  assign n47100 = ( n7422 & n30855 ) | ( n7422 & n47099 ) | ( n30855 & n47099 ) ;
  assign n47101 = ( n3920 & n12213 ) | ( n3920 & ~n36840 ) | ( n12213 & ~n36840 ) ;
  assign n47102 = n47101 ^ n25540 ^ n12523 ;
  assign n47103 = n6733 ^ n5858 ^ n518 ;
  assign n47104 = n16933 & ~n38155 ;
  assign n47105 = n47104 ^ n26694 ^ 1'b0 ;
  assign n47106 = ~n12715 & n33422 ;
  assign n47107 = n47106 ^ n10042 ^ 1'b0 ;
  assign n47108 = ( x224 & ~n2825 ) | ( x224 & n5243 ) | ( ~n2825 & n5243 ) ;
  assign n47109 = ( n19103 & n23969 ) | ( n19103 & n47108 ) | ( n23969 & n47108 ) ;
  assign n47110 = ( n4904 & n14073 ) | ( n4904 & n17844 ) | ( n14073 & n17844 ) ;
  assign n47111 = n17333 ^ n9402 ^ 1'b0 ;
  assign n47112 = n23756 | n47111 ;
  assign n47113 = ( n8011 & n47110 ) | ( n8011 & n47112 ) | ( n47110 & n47112 ) ;
  assign n47114 = ( n20947 & n27272 ) | ( n20947 & ~n40042 ) | ( n27272 & ~n40042 ) ;
  assign n47115 = n14234 ^ n5366 ^ n4551 ;
  assign n47116 = n25010 ^ n24474 ^ n5189 ;
  assign n47117 = ( n5605 & n47115 ) | ( n5605 & ~n47116 ) | ( n47115 & ~n47116 ) ;
  assign n47118 = ( ~n21275 & n25553 ) | ( ~n21275 & n42858 ) | ( n25553 & n42858 ) ;
  assign n47119 = n41330 ^ n16865 ^ 1'b0 ;
  assign n47120 = n47119 ^ n32230 ^ n22998 ;
  assign n47121 = ( n13157 & ~n14528 ) | ( n13157 & n31513 ) | ( ~n14528 & n31513 ) ;
  assign n47122 = ( ~n1334 & n8945 ) | ( ~n1334 & n36267 ) | ( n8945 & n36267 ) ;
  assign n47123 = n20017 & n45483 ;
  assign n47131 = ( n18533 & ~n38319 ) | ( n18533 & n46650 ) | ( ~n38319 & n46650 ) ;
  assign n47132 = ( n9493 & n19532 ) | ( n9493 & n47131 ) | ( n19532 & n47131 ) ;
  assign n47124 = n5235 ^ n4531 ^ n3331 ;
  assign n47125 = n47124 ^ n44755 ^ n29766 ;
  assign n47128 = n25042 ^ n5947 ^ n591 ;
  assign n47127 = ( n10530 & n26738 ) | ( n10530 & n35978 ) | ( n26738 & n35978 ) ;
  assign n47126 = ( n13508 & n16732 ) | ( n13508 & ~n42999 ) | ( n16732 & ~n42999 ) ;
  assign n47129 = n47128 ^ n47127 ^ n47126 ;
  assign n47130 = ~n47125 & n47129 ;
  assign n47133 = n47132 ^ n47130 ^ 1'b0 ;
  assign n47136 = n27949 ^ n4945 ^ x49 ;
  assign n47134 = n18275 ^ n17461 ^ n12818 ;
  assign n47135 = n47134 ^ n40873 ^ n4310 ;
  assign n47137 = n47136 ^ n47135 ^ n19140 ;
  assign n47138 = n47137 ^ n42118 ^ n38903 ;
  assign n47139 = ( ~n25321 & n33323 ) | ( ~n25321 & n47138 ) | ( n33323 & n47138 ) ;
  assign n47140 = n47139 ^ n16251 ^ n12911 ;
  assign n47141 = n36234 ^ n4560 ^ 1'b0 ;
  assign n47142 = ( n2359 & n15970 ) | ( n2359 & n21755 ) | ( n15970 & n21755 ) ;
  assign n47143 = n47142 ^ n12648 ^ n8244 ;
  assign n47144 = n36375 ^ n33686 ^ n7451 ;
  assign n47145 = ( n24232 & n40639 ) | ( n24232 & ~n47144 ) | ( n40639 & ~n47144 ) ;
  assign n47149 = ( n2107 & ~n6052 ) | ( n2107 & n41609 ) | ( ~n6052 & n41609 ) ;
  assign n47150 = ( n13523 & n33686 ) | ( n13523 & n47149 ) | ( n33686 & n47149 ) ;
  assign n47147 = n38868 ^ n14191 ^ n7024 ;
  assign n47146 = ( n9506 & ~n27901 ) | ( n9506 & n31084 ) | ( ~n27901 & n31084 ) ;
  assign n47148 = n47147 ^ n47146 ^ n6298 ;
  assign n47151 = n47150 ^ n47148 ^ n4420 ;
  assign n47152 = n42044 ^ n27937 ^ n15572 ;
  assign n47153 = ( n5117 & n9619 ) | ( n5117 & ~n12757 ) | ( n9619 & ~n12757 ) ;
  assign n47154 = ( n16319 & n42550 ) | ( n16319 & n47153 ) | ( n42550 & n47153 ) ;
  assign n47155 = ( n8377 & n18509 ) | ( n8377 & ~n39314 ) | ( n18509 & ~n39314 ) ;
  assign n47157 = ( n10127 & n30795 ) | ( n10127 & ~n46227 ) | ( n30795 & ~n46227 ) ;
  assign n47158 = n7436 | n47157 ;
  assign n47156 = ~n11751 & n31939 ;
  assign n47159 = n47158 ^ n47156 ^ 1'b0 ;
  assign n47161 = n18397 | n29127 ;
  assign n47162 = n11460 & ~n47161 ;
  assign n47160 = ( n4402 & n16158 ) | ( n4402 & n16204 ) | ( n16158 & n16204 ) ;
  assign n47163 = n47162 ^ n47160 ^ n14768 ;
  assign n47164 = n47163 ^ n36282 ^ n25593 ;
  assign n47165 = n28245 ^ n22567 ^ n17594 ;
  assign n47166 = n47165 ^ n5069 ^ n4863 ;
  assign n47168 = n36986 ^ n27808 ^ n9692 ;
  assign n47167 = ( n6410 & n15128 ) | ( n6410 & n15970 ) | ( n15128 & n15970 ) ;
  assign n47169 = n47168 ^ n47167 ^ n37863 ;
  assign n47170 = n30761 ^ n13628 ^ n5991 ;
  assign n47171 = n47170 ^ n35956 ^ n1621 ;
  assign n47172 = ( n7478 & n43344 ) | ( n7478 & ~n47171 ) | ( n43344 & ~n47171 ) ;
  assign n47173 = n11531 ^ n10663 ^ n7039 ;
  assign n47174 = ~n6238 & n19542 ;
  assign n47175 = n47174 ^ n3323 ^ 1'b0 ;
  assign n47176 = n47175 ^ n33147 ^ 1'b0 ;
  assign n47177 = n28191 ^ n21180 ^ n14532 ;
  assign n47178 = ~n2865 & n24076 ;
  assign n47179 = n47178 ^ n26598 ^ 1'b0 ;
  assign n47180 = ( n6397 & n25597 ) | ( n6397 & n46693 ) | ( n25597 & n46693 ) ;
  assign n47181 = n16957 & n40509 ;
  assign n47182 = n38970 ^ n33633 ^ n23647 ;
  assign n47185 = ( n24776 & n25399 ) | ( n24776 & ~n32971 ) | ( n25399 & ~n32971 ) ;
  assign n47183 = n2220 | n45951 ;
  assign n47184 = n47183 ^ n2007 ^ 1'b0 ;
  assign n47186 = n47185 ^ n47184 ^ 1'b0 ;
  assign n47187 = ( ~n4049 & n13797 ) | ( ~n4049 & n26859 ) | ( n13797 & n26859 ) ;
  assign n47188 = n18107 & ~n22454 ;
  assign n47189 = n1183 & n47188 ;
  assign n47190 = n47189 ^ n16351 ^ n14322 ;
  assign n47191 = n22233 | n22835 ;
  assign n47192 = n47191 ^ n42329 ^ n41714 ;
  assign n47193 = ( n26884 & n28242 ) | ( n26884 & n47192 ) | ( n28242 & n47192 ) ;
  assign n47194 = n24733 ^ n8989 ^ 1'b0 ;
  assign n47195 = n2871 | n47194 ;
  assign n47196 = n11567 ^ n5599 ^ n1055 ;
  assign n47197 = ( n23617 & ~n45702 ) | ( n23617 & n47196 ) | ( ~n45702 & n47196 ) ;
  assign n47198 = n29897 ^ n29031 ^ n4682 ;
  assign n47199 = n47198 ^ n15917 ^ n1327 ;
  assign n47200 = n47199 ^ n20403 ^ n465 ;
  assign n47201 = n35167 ^ n13789 ^ n6558 ;
  assign n47202 = n47201 ^ n32483 ^ n1711 ;
  assign n47203 = n779 & n17687 ;
  assign n47204 = n47203 ^ n12244 ^ 1'b0 ;
  assign n47205 = n45898 ^ n20431 ^ n12035 ;
  assign n47206 = n26695 ^ n15068 ^ n10529 ;
  assign n47207 = n24234 ^ n22022 ^ n17487 ;
  assign n47208 = n34905 ^ n16670 ^ 1'b0 ;
  assign n47209 = n43632 | n47208 ;
  assign n47210 = n47209 ^ n19997 ^ 1'b0 ;
  assign n47211 = ( n11963 & ~n47207 ) | ( n11963 & n47210 ) | ( ~n47207 & n47210 ) ;
  assign n47212 = n12824 ^ n2890 ^ n1807 ;
  assign n47213 = n47212 ^ n30670 ^ n7669 ;
  assign n47214 = n45646 & n47213 ;
  assign n47215 = n47214 ^ n38799 ^ 1'b0 ;
  assign n47218 = n28868 ^ n21212 ^ n13589 ;
  assign n47216 = n30095 ^ n23322 ^ 1'b0 ;
  assign n47217 = n2296 & n47216 ;
  assign n47219 = n47218 ^ n47217 ^ n43616 ;
  assign n47220 = n4047 & ~n8640 ;
  assign n47221 = n47220 ^ n44759 ^ 1'b0 ;
  assign n47222 = ( ~n29058 & n32891 ) | ( ~n29058 & n47221 ) | ( n32891 & n47221 ) ;
  assign n47223 = ( n36074 & ~n39762 ) | ( n36074 & n47222 ) | ( ~n39762 & n47222 ) ;
  assign n47224 = n41032 ^ n280 ^ 1'b0 ;
  assign n47225 = ( n10293 & ~n16915 ) | ( n10293 & n47224 ) | ( ~n16915 & n47224 ) ;
  assign n47226 = n42602 ^ n6957 ^ 1'b0 ;
  assign n47227 = n4339 & ~n6866 ;
  assign n47228 = n1007 | n47227 ;
  assign n47229 = n47228 ^ n41995 ^ n22816 ;
  assign n47230 = n39620 ^ n1824 ^ 1'b0 ;
  assign n47231 = n47230 ^ n25400 ^ n22578 ;
  assign n47232 = n14455 ^ n13359 ^ 1'b0 ;
  assign n47233 = n17991 & ~n44097 ;
  assign n47234 = ( n14639 & n20414 ) | ( n14639 & ~n47233 ) | ( n20414 & ~n47233 ) ;
  assign n47235 = n47234 ^ n14643 ^ 1'b0 ;
  assign n47236 = n39752 ^ n7891 ^ n1534 ;
  assign n47237 = ( n28443 & n46115 ) | ( n28443 & n47236 ) | ( n46115 & n47236 ) ;
  assign n47238 = n15529 ^ n6470 ^ n5413 ;
  assign n47239 = n47238 ^ n12022 ^ n11749 ;
  assign n47241 = n24581 ^ n13425 ^ n12089 ;
  assign n47240 = ( n6502 & n7549 ) | ( n6502 & ~n9555 ) | ( n7549 & ~n9555 ) ;
  assign n47242 = n47241 ^ n47240 ^ n13455 ;
  assign n47245 = n39321 ^ n14100 ^ n2642 ;
  assign n47243 = n33360 ^ n10642 ^ n6227 ;
  assign n47244 = ( n15837 & ~n32526 ) | ( n15837 & n47243 ) | ( ~n32526 & n47243 ) ;
  assign n47246 = n47245 ^ n47244 ^ n5401 ;
  assign n47247 = n28048 ^ n26068 ^ 1'b0 ;
  assign n47248 = n42800 ^ n38225 ^ n2173 ;
  assign n47249 = x51 & n6854 ;
  assign n47250 = n47249 ^ n11716 ^ 1'b0 ;
  assign n47251 = ( n33038 & n39044 ) | ( n33038 & ~n47250 ) | ( n39044 & ~n47250 ) ;
  assign n47252 = n26298 ^ n23803 ^ 1'b0 ;
  assign n47253 = n24968 ^ n15867 ^ 1'b0 ;
  assign n47254 = n36582 | n47253 ;
  assign n47256 = ( n3920 & ~n19183 ) | ( n3920 & n29716 ) | ( ~n19183 & n29716 ) ;
  assign n47255 = n24947 ^ n20826 ^ n9465 ;
  assign n47257 = n47256 ^ n47255 ^ n14509 ;
  assign n47258 = ( ~n20492 & n25738 ) | ( ~n20492 & n47257 ) | ( n25738 & n47257 ) ;
  assign n47259 = n28091 ^ n19836 ^ n16578 ;
  assign n47260 = ( n6488 & n16707 ) | ( n6488 & ~n32440 ) | ( n16707 & ~n32440 ) ;
  assign n47261 = n47260 ^ n14222 ^ n9311 ;
  assign n47262 = ( ~n32003 & n47259 ) | ( ~n32003 & n47261 ) | ( n47259 & n47261 ) ;
  assign n47263 = ( n15037 & ~n40238 ) | ( n15037 & n41919 ) | ( ~n40238 & n41919 ) ;
  assign n47264 = ( n23357 & ~n30335 ) | ( n23357 & n41261 ) | ( ~n30335 & n41261 ) ;
  assign n47265 = ( ~n33919 & n47263 ) | ( ~n33919 & n47264 ) | ( n47263 & n47264 ) ;
  assign n47266 = n750 & n3885 ;
  assign n47267 = n47266 ^ n4315 ^ 1'b0 ;
  assign n47268 = n47267 ^ n33347 ^ n11938 ;
  assign n47269 = ( n28240 & n30954 ) | ( n28240 & n40579 ) | ( n30954 & n40579 ) ;
  assign n47270 = n38415 ^ n33793 ^ n23962 ;
  assign n47271 = n35725 ^ n11914 ^ 1'b0 ;
  assign n47272 = n47271 ^ n33685 ^ n2260 ;
  assign n47273 = n47272 ^ n14138 ^ 1'b0 ;
  assign n47275 = ( n17268 & n24293 ) | ( n17268 & n36636 ) | ( n24293 & n36636 ) ;
  assign n47276 = n47275 ^ n14960 ^ n980 ;
  assign n47274 = n18056 & ~n25137 ;
  assign n47277 = n47276 ^ n47274 ^ 1'b0 ;
  assign n47280 = ( ~n9440 & n10861 ) | ( ~n9440 & n20508 ) | ( n10861 & n20508 ) ;
  assign n47278 = n29866 ^ n20600 ^ 1'b0 ;
  assign n47279 = n41116 | n47278 ;
  assign n47281 = n47280 ^ n47279 ^ n17793 ;
  assign n47282 = n8886 & ~n13687 ;
  assign n47283 = n4074 & n47282 ;
  assign n47284 = ( ~n20987 & n21169 ) | ( ~n20987 & n47283 ) | ( n21169 & n47283 ) ;
  assign n47285 = n8861 ^ n5659 ^ n3672 ;
  assign n47286 = n45478 ^ n13076 ^ 1'b0 ;
  assign n47287 = ~n20929 & n47286 ;
  assign n47288 = ( n7766 & n47285 ) | ( n7766 & ~n47287 ) | ( n47285 & ~n47287 ) ;
  assign n47289 = n43388 ^ n16984 ^ n8325 ;
  assign n47290 = ( n7457 & ~n16819 ) | ( n7457 & n28475 ) | ( ~n16819 & n28475 ) ;
  assign n47291 = ( ~n8475 & n29221 ) | ( ~n8475 & n47290 ) | ( n29221 & n47290 ) ;
  assign n47292 = n12649 ^ n11196 ^ n3914 ;
  assign n47293 = n29932 | n42432 ;
  assign n47294 = ( n38546 & n47292 ) | ( n38546 & n47293 ) | ( n47292 & n47293 ) ;
  assign n47295 = n44637 ^ n5429 ^ n696 ;
  assign n47296 = ( ~n20208 & n46514 ) | ( ~n20208 & n47295 ) | ( n46514 & n47295 ) ;
  assign n47297 = n23422 ^ n13395 ^ 1'b0 ;
  assign n47298 = ~n1757 & n47297 ;
  assign n47299 = n24915 & ~n27966 ;
  assign n47300 = n47299 ^ n7544 ^ 1'b0 ;
  assign n47301 = n30004 ^ n15546 ^ n6166 ;
  assign n47302 = n28018 ^ n19307 ^ n2278 ;
  assign n47303 = ( n13182 & n18286 ) | ( n13182 & n40531 ) | ( n18286 & n40531 ) ;
  assign n47304 = ( n28713 & n36996 ) | ( n28713 & ~n47303 ) | ( n36996 & ~n47303 ) ;
  assign n47305 = n35773 ^ n23294 ^ n21412 ;
  assign n47306 = ~n24223 & n36690 ;
  assign n47307 = n47306 ^ n41658 ^ n12758 ;
  assign n47308 = n24503 ^ n22306 ^ 1'b0 ;
  assign n47309 = ( n13184 & ~n20305 ) | ( n13184 & n47308 ) | ( ~n20305 & n47308 ) ;
  assign n47310 = n47309 ^ n23274 ^ n12277 ;
  assign n47311 = ( n10327 & n15004 ) | ( n10327 & ~n16122 ) | ( n15004 & ~n16122 ) ;
  assign n47312 = ( n20962 & n22672 ) | ( n20962 & n47311 ) | ( n22672 & n47311 ) ;
  assign n47313 = ( n3631 & ~n45432 ) | ( n3631 & n47312 ) | ( ~n45432 & n47312 ) ;
  assign n47314 = ( n47307 & n47310 ) | ( n47307 & ~n47313 ) | ( n47310 & ~n47313 ) ;
  assign n47315 = n11117 & n39341 ;
  assign n47316 = n17097 ^ n7466 ^ 1'b0 ;
  assign n47317 = n36270 ^ n33263 ^ n25919 ;
  assign n47318 = n25468 | n38662 ;
  assign n47319 = ( ~n17874 & n47317 ) | ( ~n17874 & n47318 ) | ( n47317 & n47318 ) ;
  assign n47320 = ( ~n10162 & n14463 ) | ( ~n10162 & n43438 ) | ( n14463 & n43438 ) ;
  assign n47321 = n47320 ^ n45750 ^ 1'b0 ;
  assign n47322 = ( ~n6775 & n42551 ) | ( ~n6775 & n47321 ) | ( n42551 & n47321 ) ;
  assign n47323 = n16821 ^ n13356 ^ n1434 ;
  assign n47324 = n47323 ^ n16680 ^ n4371 ;
  assign n47325 = n40797 ^ n32258 ^ n22145 ;
  assign n47326 = n34473 ^ n23295 ^ n4018 ;
  assign n47327 = n24171 ^ n10116 ^ n9622 ;
  assign n47328 = n1727 & ~n37789 ;
  assign n47329 = n7253 & n47328 ;
  assign n47330 = n8409 ^ n284 ^ 1'b0 ;
  assign n47331 = n25708 & n47330 ;
  assign n47332 = n33175 ^ n8030 ^ 1'b0 ;
  assign n47333 = ( n9015 & ~n12535 ) | ( n9015 & n33552 ) | ( ~n12535 & n33552 ) ;
  assign n47334 = n47333 ^ n21568 ^ n419 ;
  assign n47335 = n12499 & ~n36017 ;
  assign n47336 = n47335 ^ n25187 ^ 1'b0 ;
  assign n47337 = n34284 ^ n22350 ^ n13995 ;
  assign n47338 = n47337 ^ n46534 ^ n14160 ;
  assign n47339 = n47336 & ~n47338 ;
  assign n47340 = ( n6579 & ~n38198 ) | ( n6579 & n45147 ) | ( ~n38198 & n45147 ) ;
  assign n47344 = n12036 & n13597 ;
  assign n47345 = ( n7967 & n8159 ) | ( n7967 & ~n47344 ) | ( n8159 & ~n47344 ) ;
  assign n47341 = ( n16738 & ~n18682 ) | ( n16738 & n45280 ) | ( ~n18682 & n45280 ) ;
  assign n47342 = ( n16417 & ~n35245 ) | ( n16417 & n39755 ) | ( ~n35245 & n39755 ) ;
  assign n47343 = ( n32370 & ~n47341 ) | ( n32370 & n47342 ) | ( ~n47341 & n47342 ) ;
  assign n47346 = n47345 ^ n47343 ^ n30487 ;
  assign n47347 = n29131 ^ n20232 ^ n3246 ;
  assign n47348 = n13690 ^ n7132 ^ 1'b0 ;
  assign n47349 = n28515 & n47348 ;
  assign n47350 = ( n24976 & n46488 ) | ( n24976 & n47349 ) | ( n46488 & n47349 ) ;
  assign n47351 = ( n10949 & n47347 ) | ( n10949 & n47350 ) | ( n47347 & n47350 ) ;
  assign n47352 = n17469 ^ n16223 ^ n2011 ;
  assign n47353 = n47352 ^ n26296 ^ n8396 ;
  assign n47354 = ~n16440 & n28279 ;
  assign n47355 = n29403 & ~n29730 ;
  assign n47356 = n47140 & n47355 ;
  assign n47357 = n7162 ^ n4485 ^ n3272 ;
  assign n47358 = ~n5042 & n20128 ;
  assign n47359 = n47357 & n47358 ;
  assign n47360 = n42025 ^ n25855 ^ n3689 ;
  assign n47361 = n43524 ^ n23985 ^ n5515 ;
  assign n47362 = n47361 ^ n41032 ^ n15030 ;
  assign n47364 = n22568 ^ n15097 ^ n4315 ;
  assign n47363 = ( ~n1288 & n2029 ) | ( ~n1288 & n46541 ) | ( n2029 & n46541 ) ;
  assign n47365 = n47364 ^ n47363 ^ 1'b0 ;
  assign n47366 = n11635 ^ n11006 ^ n10769 ;
  assign n47368 = ( n7539 & ~n7923 ) | ( n7539 & n10252 ) | ( ~n7923 & n10252 ) ;
  assign n47367 = ~n294 & n2762 ;
  assign n47369 = n47368 ^ n47367 ^ 1'b0 ;
  assign n47370 = n47369 ^ n40185 ^ n11962 ;
  assign n47371 = n47370 ^ n14507 ^ n7166 ;
  assign n47372 = ( n16528 & ~n22311 ) | ( n16528 & n30719 ) | ( ~n22311 & n30719 ) ;
  assign n47373 = n47372 ^ n15422 ^ 1'b0 ;
  assign n47374 = ( ~n3117 & n11063 ) | ( ~n3117 & n47373 ) | ( n11063 & n47373 ) ;
  assign n47375 = ~n5959 & n32055 ;
  assign n47376 = n47375 ^ n7288 ^ n6544 ;
  assign n47377 = n2304 ^ n877 ^ 1'b0 ;
  assign n47378 = n47377 ^ n4647 ^ n810 ;
  assign n47379 = ( n13724 & n29087 ) | ( n13724 & n47378 ) | ( n29087 & n47378 ) ;
  assign n47380 = ( x19 & n10896 ) | ( x19 & ~n47379 ) | ( n10896 & ~n47379 ) ;
  assign n47381 = n22796 ^ n11809 ^ n10262 ;
  assign n47382 = n47381 ^ n18481 ^ 1'b0 ;
  assign n47383 = n14090 & ~n47382 ;
  assign n47384 = ( n657 & n11052 ) | ( n657 & ~n19829 ) | ( n11052 & ~n19829 ) ;
  assign n47386 = n2338 & n3739 ;
  assign n47387 = ( n16420 & n27568 ) | ( n16420 & ~n47386 ) | ( n27568 & ~n47386 ) ;
  assign n47385 = ( ~n1391 & n5577 ) | ( ~n1391 & n5911 ) | ( n5577 & n5911 ) ;
  assign n47388 = n47387 ^ n47385 ^ n15108 ;
  assign n47389 = ( n27351 & ~n47384 ) | ( n27351 & n47388 ) | ( ~n47384 & n47388 ) ;
  assign n47390 = n33437 ^ n12310 ^ n10775 ;
  assign n47391 = ( n4738 & n40728 ) | ( n4738 & n47390 ) | ( n40728 & n47390 ) ;
  assign n47392 = n1546 & ~n18185 ;
  assign n47393 = n47392 ^ n7842 ^ 1'b0 ;
  assign n47394 = ( ~n10148 & n21870 ) | ( ~n10148 & n47393 ) | ( n21870 & n47393 ) ;
  assign n47395 = n4347 & ~n37645 ;
  assign n47396 = ~n22780 & n47395 ;
  assign n47397 = ( n34001 & n43238 ) | ( n34001 & ~n47396 ) | ( n43238 & ~n47396 ) ;
  assign n47399 = n26742 ^ n16230 ^ n14572 ;
  assign n47398 = n8124 & ~n30203 ;
  assign n47400 = n47399 ^ n47398 ^ 1'b0 ;
  assign n47401 = ~n25231 & n47400 ;
  assign n47402 = n15052 & ~n18679 ;
  assign n47403 = n47402 ^ n13649 ^ 1'b0 ;
  assign n47404 = n11404 & ~n42872 ;
  assign n47405 = ( n2181 & n26202 ) | ( n2181 & ~n40657 ) | ( n26202 & ~n40657 ) ;
  assign n47406 = n10847 & ~n47405 ;
  assign n47407 = n47404 & n47406 ;
  assign n47408 = n19308 ^ n5925 ^ n5284 ;
  assign n47409 = ( n15492 & ~n32234 ) | ( n15492 & n32676 ) | ( ~n32234 & n32676 ) ;
  assign n47410 = n24227 ^ n5781 ^ n559 ;
  assign n47411 = ( n23376 & ~n35735 ) | ( n23376 & n43925 ) | ( ~n35735 & n43925 ) ;
  assign n47412 = ( n35588 & n47410 ) | ( n35588 & n47411 ) | ( n47410 & n47411 ) ;
  assign n47413 = ( n1379 & n1872 ) | ( n1379 & n5993 ) | ( n1872 & n5993 ) ;
  assign n47414 = ( ~n32864 & n42161 ) | ( ~n32864 & n47413 ) | ( n42161 & n47413 ) ;
  assign n47415 = n47414 ^ n6517 ^ n1662 ;
  assign n47416 = ( ~n912 & n19356 ) | ( ~n912 & n28810 ) | ( n19356 & n28810 ) ;
  assign n47417 = n17305 ^ n10242 ^ 1'b0 ;
  assign n47418 = ( n32520 & n46300 ) | ( n32520 & n47417 ) | ( n46300 & n47417 ) ;
  assign n47419 = n25710 ^ n13855 ^ n10542 ;
  assign n47420 = ( ~n9619 & n27501 ) | ( ~n9619 & n47419 ) | ( n27501 & n47419 ) ;
  assign n47421 = n20181 ^ n7981 ^ n925 ;
  assign n47422 = n5451 & n47421 ;
  assign n47423 = n47420 & n47422 ;
  assign n47424 = n44639 ^ n14489 ^ 1'b0 ;
  assign n47425 = n47424 ^ n691 ^ n362 ;
  assign n47426 = ( ~n21288 & n26661 ) | ( ~n21288 & n47425 ) | ( n26661 & n47425 ) ;
  assign n47427 = n47426 ^ n44026 ^ n40749 ;
  assign n47428 = n31953 ^ n28604 ^ n21834 ;
  assign n47429 = n47428 ^ n38564 ^ n1259 ;
  assign n47430 = ( n11961 & n14903 ) | ( n11961 & ~n43188 ) | ( n14903 & ~n43188 ) ;
  assign n47431 = n21826 ^ n19401 ^ n5374 ;
  assign n47432 = ( ~n3185 & n5970 ) | ( ~n3185 & n17592 ) | ( n5970 & n17592 ) ;
  assign n47433 = ( ~n921 & n35719 ) | ( ~n921 & n45400 ) | ( n35719 & n45400 ) ;
  assign n47434 = n47433 ^ n16709 ^ n15128 ;
  assign n47435 = ( ~n34427 & n47432 ) | ( ~n34427 & n47434 ) | ( n47432 & n47434 ) ;
  assign n47436 = ( n2140 & n19953 ) | ( n2140 & ~n25490 ) | ( n19953 & ~n25490 ) ;
  assign n47437 = n47436 ^ n15351 ^ n15140 ;
  assign n47438 = ( n9688 & n10502 ) | ( n9688 & ~n11300 ) | ( n10502 & ~n11300 ) ;
  assign n47439 = n47438 ^ n17029 ^ 1'b0 ;
  assign n47440 = n47439 ^ n46639 ^ n10616 ;
  assign n47441 = ( n8553 & n47437 ) | ( n8553 & n47440 ) | ( n47437 & n47440 ) ;
  assign n47443 = n5851 ^ n4064 ^ n2609 ;
  assign n47442 = n25219 ^ n13919 ^ n2436 ;
  assign n47444 = n47443 ^ n47442 ^ n2062 ;
  assign n47445 = ( n5306 & ~n42970 ) | ( n5306 & n47444 ) | ( ~n42970 & n47444 ) ;
  assign n47446 = n47445 ^ n44915 ^ n4849 ;
  assign n47447 = ( n6018 & n15046 ) | ( n6018 & ~n16538 ) | ( n15046 & ~n16538 ) ;
  assign n47448 = ( n11065 & n42062 ) | ( n11065 & n47447 ) | ( n42062 & n47447 ) ;
  assign n47449 = n2426 & n25132 ;
  assign n47450 = ~n47448 & n47449 ;
  assign n47451 = n45894 ^ n9861 ^ n4419 ;
  assign n47452 = ( n965 & ~n23456 ) | ( n965 & n47451 ) | ( ~n23456 & n47451 ) ;
  assign n47453 = n47452 ^ n27825 ^ n21622 ;
  assign n47454 = ( n6748 & n18641 ) | ( n6748 & ~n28456 ) | ( n18641 & ~n28456 ) ;
  assign n47455 = n1840 & ~n47454 ;
  assign n47456 = ( n7867 & n18102 ) | ( n7867 & n47455 ) | ( n18102 & n47455 ) ;
  assign n47457 = ( ~n15691 & n32152 ) | ( ~n15691 & n47456 ) | ( n32152 & n47456 ) ;
  assign n47458 = n47457 ^ n10738 ^ x146 ;
  assign n47459 = ( n2845 & ~n38317 ) | ( n2845 & n39539 ) | ( ~n38317 & n39539 ) ;
  assign n47460 = n47459 ^ n43670 ^ n40577 ;
  assign n47461 = n21684 ^ n16262 ^ n1009 ;
  assign n47462 = n12442 | n30861 ;
  assign n47465 = ( n5210 & n27229 ) | ( n5210 & ~n28036 ) | ( n27229 & ~n28036 ) ;
  assign n47466 = n47465 ^ n44639 ^ n6853 ;
  assign n47463 = n25381 ^ n5460 ^ n1972 ;
  assign n47464 = n47463 ^ n38595 ^ n36270 ;
  assign n47467 = n47466 ^ n47464 ^ n40626 ;
  assign n47468 = n29110 ^ n8767 ^ 1'b0 ;
  assign n47469 = n20339 ^ n15051 ^ n3856 ;
  assign n47470 = n17367 & n24060 ;
  assign n47471 = n47470 ^ n11321 ^ 1'b0 ;
  assign n47472 = n31027 ^ n22406 ^ n3539 ;
  assign n47473 = n27949 & ~n40776 ;
  assign n47474 = n20995 ^ n14387 ^ n5560 ;
  assign n47475 = ( n9340 & ~n16217 ) | ( n9340 & n47474 ) | ( ~n16217 & n47474 ) ;
  assign n47476 = ( n12915 & n13269 ) | ( n12915 & ~n34377 ) | ( n13269 & ~n34377 ) ;
  assign n47477 = ( n9482 & n10179 ) | ( n9482 & ~n47476 ) | ( n10179 & ~n47476 ) ;
  assign n47478 = ( n16051 & ~n18633 ) | ( n16051 & n42538 ) | ( ~n18633 & n42538 ) ;
  assign n47479 = n39128 ^ x135 ^ 1'b0 ;
  assign n47480 = n18714 ^ n5085 ^ n2131 ;
  assign n47481 = ( n26688 & ~n33037 ) | ( n26688 & n34024 ) | ( ~n33037 & n34024 ) ;
  assign n47482 = ( ~n1553 & n46875 ) | ( ~n1553 & n47481 ) | ( n46875 & n47481 ) ;
  assign n47483 = n39007 ^ n22011 ^ 1'b0 ;
  assign n47484 = ~n35584 & n47483 ;
  assign n47485 = n10692 | n35165 ;
  assign n47486 = n36188 ^ n26861 ^ n12084 ;
  assign n47488 = n7136 ^ n6224 ^ n2523 ;
  assign n47489 = n47488 ^ n18711 ^ n8269 ;
  assign n47490 = n47489 ^ n34560 ^ 1'b0 ;
  assign n47491 = n47124 & n47490 ;
  assign n47487 = n39384 ^ n19561 ^ x244 ;
  assign n47492 = n47491 ^ n47487 ^ n11845 ;
  assign n47493 = n24845 ^ n18963 ^ 1'b0 ;
  assign n47494 = ~n7012 & n47493 ;
  assign n47495 = n47494 ^ n36208 ^ n26331 ;
  assign n47496 = ( n3430 & ~n6824 ) | ( n3430 & n8955 ) | ( ~n6824 & n8955 ) ;
  assign n47497 = n5944 & ~n41228 ;
  assign n47498 = ~n36774 & n47497 ;
  assign n47499 = ( n22896 & n24222 ) | ( n22896 & ~n47498 ) | ( n24222 & ~n47498 ) ;
  assign n47500 = ( n14027 & n23236 ) | ( n14027 & n47499 ) | ( n23236 & n47499 ) ;
  assign n47501 = n4495 ^ n3007 ^ n607 ;
  assign n47502 = ( n4314 & ~n17005 ) | ( n4314 & n37186 ) | ( ~n17005 & n37186 ) ;
  assign n47503 = n7058 | n43866 ;
  assign n47504 = n19212 | n47503 ;
  assign n47505 = ( n2700 & ~n43883 ) | ( n2700 & n47504 ) | ( ~n43883 & n47504 ) ;
  assign n47506 = n11465 ^ n5615 ^ 1'b0 ;
  assign n47507 = n11587 ^ n9340 ^ 1'b0 ;
  assign n47508 = ~n47506 & n47507 ;
  assign n47509 = n18810 | n39585 ;
  assign n47510 = n47509 ^ n39702 ^ 1'b0 ;
  assign n47511 = n2195 & n39892 ;
  assign n47512 = ( n6242 & n10959 ) | ( n6242 & n31622 ) | ( n10959 & n31622 ) ;
  assign n47513 = ( n1661 & n19173 ) | ( n1661 & n20725 ) | ( n19173 & n20725 ) ;
  assign n47514 = n16819 ^ n8078 ^ n5853 ;
  assign n47515 = n15161 ^ n4231 ^ 1'b0 ;
  assign n47516 = n14604 ^ n9630 ^ n6471 ;
  assign n47517 = ( n7612 & n18796 ) | ( n7612 & ~n47516 ) | ( n18796 & ~n47516 ) ;
  assign n47518 = n47517 ^ n31619 ^ n25803 ;
  assign n47519 = ( n12535 & n17739 ) | ( n12535 & ~n32388 ) | ( n17739 & ~n32388 ) ;
  assign n47520 = ( n6760 & ~n32572 ) | ( n6760 & n47519 ) | ( ~n32572 & n47519 ) ;
  assign n47521 = ( n11788 & n17554 ) | ( n11788 & n31243 ) | ( n17554 & n31243 ) ;
  assign n47522 = n47521 ^ n24109 ^ n15990 ;
  assign n47523 = n24311 ^ n18721 ^ n10506 ;
  assign n47524 = ( n13619 & n14492 ) | ( n13619 & ~n47523 ) | ( n14492 & ~n47523 ) ;
  assign n47525 = n47524 ^ n18996 ^ n3989 ;
  assign n47526 = n19147 ^ n15101 ^ n1710 ;
  assign n47527 = n19193 | n30510 ;
  assign n47528 = n47526 | n47527 ;
  assign n47529 = ~n24995 & n40835 ;
  assign n47530 = n29382 & n47529 ;
  assign n47531 = n47530 ^ n27459 ^ n17776 ;
  assign n47532 = ( n16609 & ~n28018 ) | ( n16609 & n34040 ) | ( ~n28018 & n34040 ) ;
  assign n47539 = ( ~n675 & n2549 ) | ( ~n675 & n16236 ) | ( n2549 & n16236 ) ;
  assign n47535 = n10280 | n11698 ;
  assign n47536 = n3665 & ~n47535 ;
  assign n47537 = n47536 ^ n23823 ^ 1'b0 ;
  assign n47533 = n566 | n9853 ;
  assign n47534 = n21694 & ~n47533 ;
  assign n47538 = n47537 ^ n47534 ^ n17468 ;
  assign n47540 = n47539 ^ n47538 ^ n3650 ;
  assign n47541 = ( n20194 & ~n24126 ) | ( n20194 & n46891 ) | ( ~n24126 & n46891 ) ;
  assign n47542 = ( n38578 & n39191 ) | ( n38578 & n47541 ) | ( n39191 & n47541 ) ;
  assign n47543 = n30203 & n39289 ;
  assign n47544 = ( ~n25320 & n47542 ) | ( ~n25320 & n47543 ) | ( n47542 & n47543 ) ;
  assign n47545 = n20092 ^ n10814 ^ n10058 ;
  assign n47546 = n37751 ^ n24950 ^ n5194 ;
  assign n47547 = n47546 ^ n22205 ^ n16462 ;
  assign n47548 = ( n41637 & n41805 ) | ( n41637 & n47547 ) | ( n41805 & n47547 ) ;
  assign n47549 = ( n3240 & n12795 ) | ( n3240 & ~n18159 ) | ( n12795 & ~n18159 ) ;
  assign n47550 = n47549 ^ n35137 ^ 1'b0 ;
  assign n47551 = ( ~n524 & n15677 ) | ( ~n524 & n17624 ) | ( n15677 & n17624 ) ;
  assign n47552 = n47551 ^ n6812 ^ 1'b0 ;
  assign n47553 = ~n18493 & n47552 ;
  assign n47554 = ( n17016 & n40177 ) | ( n17016 & ~n47553 ) | ( n40177 & ~n47553 ) ;
  assign n47555 = n16746 ^ n12357 ^ n7921 ;
  assign n47556 = n45178 ^ n34504 ^ n6780 ;
  assign n47557 = n38518 ^ n20817 ^ n859 ;
  assign n47558 = ( ~n47555 & n47556 ) | ( ~n47555 & n47557 ) | ( n47556 & n47557 ) ;
  assign n47559 = n44327 ^ n29852 ^ n17746 ;
  assign n47560 = ( n19373 & n19415 ) | ( n19373 & ~n47559 ) | ( n19415 & ~n47559 ) ;
  assign n47561 = ( ~n12178 & n28722 ) | ( ~n12178 & n47243 ) | ( n28722 & n47243 ) ;
  assign n47562 = n47561 ^ n29285 ^ n12356 ;
  assign n47563 = n16819 ^ n14106 ^ 1'b0 ;
  assign n47564 = n6068 | n11920 ;
  assign n47565 = n13244 & ~n47564 ;
  assign n47566 = ( n42245 & n47563 ) | ( n42245 & n47565 ) | ( n47563 & n47565 ) ;
  assign n47571 = ( ~n1626 & n4523 ) | ( ~n1626 & n10635 ) | ( n4523 & n10635 ) ;
  assign n47568 = n21551 ^ n15157 ^ 1'b0 ;
  assign n47569 = ~n14277 & n47568 ;
  assign n47570 = n47569 ^ n40214 ^ 1'b0 ;
  assign n47567 = n42376 ^ n38011 ^ n17862 ;
  assign n47572 = n47571 ^ n47570 ^ n47567 ;
  assign n47573 = n10517 ^ n1095 ^ 1'b0 ;
  assign n47574 = n17159 | n47573 ;
  assign n47575 = ~n16419 & n30923 ;
  assign n47576 = n47575 ^ n30820 ^ 1'b0 ;
  assign n47577 = ~n27681 & n31581 ;
  assign n47578 = n15232 ^ n9143 ^ n4295 ;
  assign n47579 = n37899 ^ n34523 ^ n33088 ;
  assign n47580 = n37293 ^ n18280 ^ n9055 ;
  assign n47581 = ( ~n6880 & n33250 ) | ( ~n6880 & n47580 ) | ( n33250 & n47580 ) ;
  assign n47582 = n41980 ^ n23022 ^ n7352 ;
  assign n47583 = n44882 ^ n33704 ^ n33066 ;
  assign n47584 = ( n2908 & n29470 ) | ( n2908 & n47583 ) | ( n29470 & n47583 ) ;
  assign n47585 = n36275 ^ n16051 ^ 1'b0 ;
  assign n47586 = ( n15011 & ~n37940 ) | ( n15011 & n39847 ) | ( ~n37940 & n39847 ) ;
  assign n47587 = ( n1256 & ~n2322 ) | ( n1256 & n11249 ) | ( ~n2322 & n11249 ) ;
  assign n47588 = ( n661 & n1708 ) | ( n661 & ~n3419 ) | ( n1708 & ~n3419 ) ;
  assign n47589 = n47588 ^ n28464 ^ n12775 ;
  assign n47590 = n19982 ^ n10404 ^ 1'b0 ;
  assign n47591 = ( ~n22769 & n27558 ) | ( ~n22769 & n47590 ) | ( n27558 & n47590 ) ;
  assign n47592 = ( n29045 & n30459 ) | ( n29045 & n36632 ) | ( n30459 & n36632 ) ;
  assign n47593 = n47592 ^ n12706 ^ n974 ;
  assign n47594 = n13561 ^ n4785 ^ 1'b0 ;
  assign n47595 = n42420 & n47594 ;
  assign n47596 = n47595 ^ n24185 ^ n2978 ;
  assign n47602 = ( ~n21765 & n26455 ) | ( ~n21765 & n28615 ) | ( n26455 & n28615 ) ;
  assign n47600 = ( n7590 & n11751 ) | ( n7590 & ~n12109 ) | ( n11751 & ~n12109 ) ;
  assign n47601 = n47600 ^ n19000 ^ n8392 ;
  assign n47598 = n264 & ~n10379 ;
  assign n47597 = n26265 ^ n19231 ^ n6774 ;
  assign n47599 = n47598 ^ n47597 ^ n6554 ;
  assign n47603 = n47602 ^ n47601 ^ n47599 ;
  assign n47604 = n47032 ^ n20851 ^ n6341 ;
  assign n47605 = n47604 ^ n25982 ^ 1'b0 ;
  assign n47606 = n47605 ^ n44097 ^ n1036 ;
  assign n47607 = ( ~n816 & n21179 ) | ( ~n816 & n37357 ) | ( n21179 & n37357 ) ;
  assign n47608 = n13114 ^ n3911 ^ 1'b0 ;
  assign n47609 = n17357 ^ n7835 ^ n2320 ;
  assign n47610 = ( n3666 & n47608 ) | ( n3666 & ~n47609 ) | ( n47608 & ~n47609 ) ;
  assign n47611 = n18417 & n47610 ;
  assign n47612 = n47611 ^ n40997 ^ 1'b0 ;
  assign n47613 = n37706 ^ n20724 ^ 1'b0 ;
  assign n47614 = n26400 & ~n47613 ;
  assign n47615 = ( ~n21645 & n36995 ) | ( ~n21645 & n37662 ) | ( n36995 & n37662 ) ;
  assign n47617 = n14283 | n18663 ;
  assign n47618 = n34641 | n47617 ;
  assign n47616 = ( n2237 & n5721 ) | ( n2237 & ~n12441 ) | ( n5721 & ~n12441 ) ;
  assign n47619 = n47618 ^ n47616 ^ n3935 ;
  assign n47627 = n24110 ^ n18118 ^ n7127 ;
  assign n47628 = n47627 ^ n13054 ^ n320 ;
  assign n47621 = n28574 ^ n16508 ^ n7565 ;
  assign n47622 = n47621 ^ n19129 ^ n15819 ;
  assign n47623 = ( ~n4707 & n31273 ) | ( ~n4707 & n47622 ) | ( n31273 & n47622 ) ;
  assign n47620 = ( ~n2546 & n5066 ) | ( ~n2546 & n21262 ) | ( n5066 & n21262 ) ;
  assign n47624 = n47623 ^ n47620 ^ n19211 ;
  assign n47625 = ( n3314 & ~n30063 ) | ( n3314 & n40127 ) | ( ~n30063 & n40127 ) ;
  assign n47626 = ( n26906 & n47624 ) | ( n26906 & n47625 ) | ( n47624 & n47625 ) ;
  assign n47629 = n47628 ^ n47626 ^ n2840 ;
  assign n47630 = n32576 ^ n14231 ^ n3176 ;
  assign n47631 = n24579 ^ n19120 ^ 1'b0 ;
  assign n47632 = n9609 ^ n6424 ^ 1'b0 ;
  assign n47633 = n36904 ^ n30824 ^ n1301 ;
  assign n47634 = ( ~n10969 & n33197 ) | ( ~n10969 & n47633 ) | ( n33197 & n47633 ) ;
  assign n47635 = n47634 ^ n38363 ^ n11661 ;
  assign n47636 = n47635 ^ n37825 ^ n32009 ;
  assign n47637 = ( n10884 & n19189 ) | ( n10884 & ~n34230 ) | ( n19189 & ~n34230 ) ;
  assign n47638 = ( n1725 & n24934 ) | ( n1725 & n47637 ) | ( n24934 & n47637 ) ;
  assign n47639 = n47638 ^ n38670 ^ n13749 ;
  assign n47640 = ( ~n21711 & n47636 ) | ( ~n21711 & n47639 ) | ( n47636 & n47639 ) ;
  assign n47641 = n16536 ^ n15411 ^ n6057 ;
  assign n47642 = ( n1814 & ~n2894 ) | ( n1814 & n13127 ) | ( ~n2894 & n13127 ) ;
  assign n47643 = n25722 ^ n9757 ^ 1'b0 ;
  assign n47644 = n47642 | n47643 ;
  assign n47645 = ( n34760 & ~n47641 ) | ( n34760 & n47644 ) | ( ~n47641 & n47644 ) ;
  assign n47646 = ( n30178 & ~n40384 ) | ( n30178 & n42282 ) | ( ~n40384 & n42282 ) ;
  assign n47647 = ~n1341 & n36690 ;
  assign n47648 = n27393 & n47647 ;
  assign n47649 = n45197 ^ n39958 ^ n10567 ;
  assign n47650 = n47649 ^ n30582 ^ n11222 ;
  assign n47651 = n38181 ^ n28423 ^ n11076 ;
  assign n47652 = ( ~n13838 & n18045 ) | ( ~n13838 & n38408 ) | ( n18045 & n38408 ) ;
  assign n47653 = n38443 ^ n6139 ^ n4739 ;
  assign n47654 = n47653 ^ n24301 ^ n1629 ;
  assign n47655 = n10355 ^ n7443 ^ n1774 ;
  assign n47656 = n47655 ^ n27529 ^ n23285 ;
  assign n47663 = n18427 & n33924 ;
  assign n47657 = ( n13087 & ~n16059 ) | ( n13087 & n17000 ) | ( ~n16059 & n17000 ) ;
  assign n47658 = ~n16669 & n24519 ;
  assign n47659 = ( n38386 & ~n47657 ) | ( n38386 & n47658 ) | ( ~n47657 & n47658 ) ;
  assign n47660 = ( n4355 & n11003 ) | ( n4355 & n13114 ) | ( n11003 & n13114 ) ;
  assign n47661 = n47660 ^ n39708 ^ 1'b0 ;
  assign n47662 = n47659 | n47661 ;
  assign n47664 = n47663 ^ n47662 ^ n26601 ;
  assign n47667 = n7411 | n24516 ;
  assign n47668 = n1597 & ~n47667 ;
  assign n47665 = ( n17015 & n24826 ) | ( n17015 & ~n34462 ) | ( n24826 & ~n34462 ) ;
  assign n47666 = n9481 & ~n47665 ;
  assign n47669 = n47668 ^ n47666 ^ 1'b0 ;
  assign n47670 = ~n31253 & n46131 ;
  assign n47671 = ~n27360 & n47670 ;
  assign n47672 = n36589 ^ n16930 ^ n1952 ;
  assign n47673 = ( ~n3986 & n22723 ) | ( ~n3986 & n47672 ) | ( n22723 & n47672 ) ;
  assign n47674 = n40119 ^ n26265 ^ n4783 ;
  assign n47675 = ( n2856 & n40331 ) | ( n2856 & n47674 ) | ( n40331 & n47674 ) ;
  assign n47676 = n47675 ^ n31604 ^ n29199 ;
  assign n47677 = n22494 ^ n12580 ^ 1'b0 ;
  assign n47678 = ( ~n5600 & n21193 ) | ( ~n5600 & n27419 ) | ( n21193 & n27419 ) ;
  assign n47679 = ( ~n7089 & n21309 ) | ( ~n7089 & n22539 ) | ( n21309 & n22539 ) ;
  assign n47680 = ( ~n3296 & n21390 ) | ( ~n3296 & n44967 ) | ( n21390 & n44967 ) ;
  assign n47681 = ( n6477 & n25629 ) | ( n6477 & ~n47680 ) | ( n25629 & ~n47680 ) ;
  assign n47682 = n47681 ^ n13893 ^ 1'b0 ;
  assign n47683 = n16483 | n31487 ;
  assign n47684 = ( n4349 & n4726 ) | ( n4349 & ~n11323 ) | ( n4726 & ~n11323 ) ;
  assign n47685 = n40540 ^ n12291 ^ 1'b0 ;
  assign n47686 = ~n21724 & n47685 ;
  assign n47687 = n47684 & n47686 ;
  assign n47688 = n47687 ^ n21619 ^ 1'b0 ;
  assign n47693 = ( x2 & n30915 ) | ( x2 & ~n32837 ) | ( n30915 & ~n32837 ) ;
  assign n47689 = ( ~n3244 & n4654 ) | ( ~n3244 & n13019 ) | ( n4654 & n13019 ) ;
  assign n47690 = ( ~n9654 & n18239 ) | ( ~n9654 & n24125 ) | ( n18239 & n24125 ) ;
  assign n47691 = ( n43318 & n47689 ) | ( n43318 & ~n47690 ) | ( n47689 & ~n47690 ) ;
  assign n47692 = n8812 | n47691 ;
  assign n47694 = n47693 ^ n47692 ^ 1'b0 ;
  assign n47701 = n35104 ^ n26326 ^ n17042 ;
  assign n47698 = ( n3746 & ~n4197 ) | ( n3746 & n24200 ) | ( ~n4197 & n24200 ) ;
  assign n47699 = ( n3369 & n18059 ) | ( n3369 & n47698 ) | ( n18059 & n47698 ) ;
  assign n47695 = n19989 & n31335 ;
  assign n47696 = n47695 ^ n38910 ^ 1'b0 ;
  assign n47697 = ( ~n13992 & n47163 ) | ( ~n13992 & n47696 ) | ( n47163 & n47696 ) ;
  assign n47700 = n47699 ^ n47697 ^ 1'b0 ;
  assign n47702 = n47701 ^ n47700 ^ n17540 ;
  assign n47703 = n42974 ^ n39392 ^ n16362 ;
  assign n47704 = ( n3577 & n18646 ) | ( n3577 & ~n19914 ) | ( n18646 & ~n19914 ) ;
  assign n47705 = n7548 ^ n5218 ^ n3395 ;
  assign n47706 = n31757 ^ n7476 ^ n1573 ;
  assign n47707 = ( n10305 & n14679 ) | ( n10305 & n19267 ) | ( n14679 & n19267 ) ;
  assign n47708 = n43470 | n47707 ;
  assign n47709 = ~n11718 & n31236 ;
  assign n47711 = n16607 ^ n16035 ^ n1136 ;
  assign n47712 = n32794 ^ n14380 ^ 1'b0 ;
  assign n47713 = ~n47711 & n47712 ;
  assign n47714 = n47713 ^ n9521 ^ n6985 ;
  assign n47710 = n10053 & ~n32694 ;
  assign n47715 = n47714 ^ n47710 ^ 1'b0 ;
  assign n47716 = ( n7699 & ~n8126 ) | ( n7699 & n34776 ) | ( ~n8126 & n34776 ) ;
  assign n47717 = ( ~n3786 & n12828 ) | ( ~n3786 & n38067 ) | ( n12828 & n38067 ) ;
  assign n47718 = ( n13666 & n25432 ) | ( n13666 & ~n33619 ) | ( n25432 & ~n33619 ) ;
  assign n47719 = n25905 ^ n9934 ^ n399 ;
  assign n47720 = ( ~x192 & n9489 ) | ( ~x192 & n47719 ) | ( n9489 & n47719 ) ;
  assign n47721 = ( n22525 & n41188 ) | ( n22525 & ~n47720 ) | ( n41188 & ~n47720 ) ;
  assign n47722 = n34941 ^ n30853 ^ 1'b0 ;
  assign n47723 = n18410 ^ n12061 ^ n5659 ;
  assign n47724 = ( n9941 & ~n40278 ) | ( n9941 & n47723 ) | ( ~n40278 & n47723 ) ;
  assign n47725 = ( n47721 & ~n47722 ) | ( n47721 & n47724 ) | ( ~n47722 & n47724 ) ;
  assign n47726 = n33894 ^ n32483 ^ n7354 ;
  assign n47727 = n47726 ^ n46392 ^ n38096 ;
  assign n47728 = n21391 & n39598 ;
  assign n47729 = n47728 ^ n14256 ^ 1'b0 ;
  assign n47730 = n9926 ^ n3483 ^ n3110 ;
  assign n47731 = n46857 ^ n10555 ^ n3382 ;
  assign n47732 = ( n27380 & n47730 ) | ( n27380 & ~n47731 ) | ( n47730 & ~n47731 ) ;
  assign n47733 = n13225 & ~n17126 ;
  assign n47734 = n47733 ^ n20813 ^ 1'b0 ;
  assign n47735 = n47734 ^ n6193 ^ n1133 ;
  assign n47736 = n31107 ^ n30913 ^ n14107 ;
  assign n47737 = ( n8981 & n47735 ) | ( n8981 & n47736 ) | ( n47735 & n47736 ) ;
  assign n47738 = ( n4826 & n8013 ) | ( n4826 & n25351 ) | ( n8013 & n25351 ) ;
  assign n47740 = ( n2172 & ~n12395 ) | ( n2172 & n16969 ) | ( ~n12395 & n16969 ) ;
  assign n47739 = ( n3482 & n15150 ) | ( n3482 & n15356 ) | ( n15150 & n15356 ) ;
  assign n47741 = n47740 ^ n47739 ^ n606 ;
  assign n47742 = n47741 ^ n8828 ^ x61 ;
  assign n47743 = n4721 & n47742 ;
  assign n47744 = ~n47738 & n47743 ;
  assign n47745 = ( n1758 & n40487 ) | ( n1758 & n47744 ) | ( n40487 & n47744 ) ;
  assign n47746 = n22074 ^ n19843 ^ x128 ;
  assign n47747 = ( n13782 & ~n38198 ) | ( n13782 & n38207 ) | ( ~n38198 & n38207 ) ;
  assign n47748 = n47747 ^ n16841 ^ n8702 ;
  assign n47749 = n16048 ^ n6525 ^ n3780 ;
  assign n47750 = n34712 ^ n31508 ^ 1'b0 ;
  assign n47751 = ( n25942 & n26088 ) | ( n25942 & ~n47750 ) | ( n26088 & ~n47750 ) ;
  assign n47752 = n47751 ^ n41754 ^ 1'b0 ;
  assign n47753 = n2240 & ~n47752 ;
  assign n47754 = ~n21400 & n37721 ;
  assign n47755 = ~n20913 & n47754 ;
  assign n47756 = ( n5586 & n25343 ) | ( n5586 & n32884 ) | ( n25343 & n32884 ) ;
  assign n47759 = n36372 ^ n14829 ^ 1'b0 ;
  assign n47760 = ( n15570 & ~n47444 ) | ( n15570 & n47759 ) | ( ~n47444 & n47759 ) ;
  assign n47757 = n30023 ^ n18883 ^ n4359 ;
  assign n47758 = n47757 ^ n45752 ^ n1300 ;
  assign n47761 = n47760 ^ n47758 ^ n5871 ;
  assign n47762 = ( n46278 & n47756 ) | ( n46278 & ~n47761 ) | ( n47756 & ~n47761 ) ;
  assign n47763 = n40131 ^ n33647 ^ n23921 ;
  assign n47764 = ( ~n733 & n26677 ) | ( ~n733 & n43616 ) | ( n26677 & n43616 ) ;
  assign n47765 = ( n19085 & n21961 ) | ( n19085 & ~n36338 ) | ( n21961 & ~n36338 ) ;
  assign n47766 = n47765 ^ n37886 ^ n13486 ;
  assign n47767 = ~n29595 & n33732 ;
  assign n47768 = n47767 ^ n11645 ^ 1'b0 ;
  assign n47769 = n47768 ^ n16066 ^ n15062 ;
  assign n47770 = n44135 ^ n6326 ^ n3139 ;
  assign n47771 = n24004 ^ n21660 ^ n6336 ;
  assign n47772 = n44960 | n47771 ;
  assign n47773 = ( n3242 & n38873 ) | ( n3242 & n47772 ) | ( n38873 & n47772 ) ;
  assign n47774 = ( n28905 & ~n30853 ) | ( n28905 & n43534 ) | ( ~n30853 & n43534 ) ;
  assign n47775 = n1212 ^ n953 ^ 1'b0 ;
  assign n47776 = n23060 & n47775 ;
  assign n47777 = n20794 ^ n18031 ^ n6038 ;
  assign n47778 = n40780 ^ n32307 ^ 1'b0 ;
  assign n47779 = n36224 & n47778 ;
  assign n47780 = ( n41301 & ~n47777 ) | ( n41301 & n47779 ) | ( ~n47777 & n47779 ) ;
  assign n47781 = n45433 ^ n3446 ^ x101 ;
  assign n47782 = n46591 ^ n7125 ^ n6600 ;
  assign n47783 = n47782 ^ n2689 ^ 1'b0 ;
  assign n47784 = n15485 ^ n12697 ^ 1'b0 ;
  assign n47785 = n32684 ^ n20851 ^ n15262 ;
  assign n47786 = ( n25776 & n47784 ) | ( n25776 & ~n47785 ) | ( n47784 & ~n47785 ) ;
  assign n47787 = n38007 ^ n22710 ^ n275 ;
  assign n47788 = ( ~n10106 & n19406 ) | ( ~n10106 & n47787 ) | ( n19406 & n47787 ) ;
  assign n47789 = ( ~n2557 & n9183 ) | ( ~n2557 & n47788 ) | ( n9183 & n47788 ) ;
  assign n47790 = ( n25735 & n29183 ) | ( n25735 & n32500 ) | ( n29183 & n32500 ) ;
  assign n47791 = ( x176 & n10437 ) | ( x176 & ~n22045 ) | ( n10437 & ~n22045 ) ;
  assign n47792 = ( n38950 & n47790 ) | ( n38950 & n47791 ) | ( n47790 & n47791 ) ;
  assign n47793 = ( x28 & ~n5181 ) | ( x28 & n28148 ) | ( ~n5181 & n28148 ) ;
  assign n47794 = ( n1478 & n44846 ) | ( n1478 & n47793 ) | ( n44846 & n47793 ) ;
  assign n47795 = n44936 ^ n31557 ^ n26674 ;
  assign n47797 = ( ~n19467 & n27991 ) | ( ~n19467 & n34427 ) | ( n27991 & n34427 ) ;
  assign n47796 = n44510 ^ n30636 ^ n1188 ;
  assign n47798 = n47797 ^ n47796 ^ n38494 ;
  assign n47799 = ( ~n25824 & n31495 ) | ( ~n25824 & n36318 ) | ( n31495 & n36318 ) ;
  assign n47800 = n37025 ^ n17337 ^ 1'b0 ;
  assign n47801 = n33604 & ~n47800 ;
  assign n47802 = n47801 ^ n29498 ^ n12767 ;
  assign n47803 = n37993 ^ n23240 ^ n7748 ;
  assign n47804 = n13523 ^ n1186 ^ n372 ;
  assign n47805 = n47804 ^ n22038 ^ n1549 ;
  assign n47806 = ( ~n3219 & n5870 ) | ( ~n3219 & n47805 ) | ( n5870 & n47805 ) ;
  assign n47807 = n34749 ^ n19615 ^ n16135 ;
  assign n47808 = n47807 ^ n11389 ^ n8071 ;
  assign n47809 = ( n8256 & n35538 ) | ( n8256 & n44954 ) | ( n35538 & n44954 ) ;
  assign n47810 = n19493 ^ n5845 ^ n2492 ;
  assign n47811 = n11081 & n40835 ;
  assign n47812 = n18351 & n47811 ;
  assign n47813 = n45811 & n47812 ;
  assign n47814 = n17337 ^ n2225 ^ 1'b0 ;
  assign n47815 = ( n7287 & n28431 ) | ( n7287 & ~n47814 ) | ( n28431 & ~n47814 ) ;
  assign n47816 = n20111 ^ n14130 ^ n8279 ;
  assign n47817 = n47816 ^ n40558 ^ n26813 ;
  assign n47818 = n20602 ^ n16198 ^ n10562 ;
  assign n47819 = ( n1426 & n4459 ) | ( n1426 & n18251 ) | ( n4459 & n18251 ) ;
  assign n47820 = n47819 ^ n38350 ^ n603 ;
  assign n47821 = n47820 ^ n22511 ^ n19977 ;
  assign n47822 = n24802 ^ n11408 ^ 1'b0 ;
  assign n47823 = n25298 | n47822 ;
  assign n47824 = n39725 ^ n12337 ^ 1'b0 ;
  assign n47825 = n33728 ^ n19261 ^ n5104 ;
  assign n47826 = n47825 ^ n29739 ^ n8905 ;
  assign n47827 = ( n47823 & n47824 ) | ( n47823 & ~n47826 ) | ( n47824 & ~n47826 ) ;
  assign n47828 = ( n18434 & n35666 ) | ( n18434 & ~n45669 ) | ( n35666 & ~n45669 ) ;
  assign n47829 = n26140 & ~n41218 ;
  assign n47830 = n47829 ^ n7829 ^ 1'b0 ;
  assign n47831 = ( ~n3415 & n9795 ) | ( ~n3415 & n11523 ) | ( n9795 & n11523 ) ;
  assign n47832 = n47831 ^ n23282 ^ n3809 ;
  assign n47833 = n47832 ^ n36175 ^ n15170 ;
  assign n47834 = n47833 ^ n14358 ^ n14215 ;
  assign n47835 = n43534 ^ n15764 ^ n7126 ;
  assign n47836 = n33315 ^ n18298 ^ 1'b0 ;
  assign n47837 = n8667 & n9392 ;
  assign n47838 = n26262 ^ n15269 ^ n3221 ;
  assign n47839 = ( n5548 & n25207 ) | ( n5548 & ~n36597 ) | ( n25207 & ~n36597 ) ;
  assign n47840 = ( n11877 & n13364 ) | ( n11877 & ~n15426 ) | ( n13364 & ~n15426 ) ;
  assign n47841 = n47840 ^ n16037 ^ n713 ;
  assign n47842 = ( n12312 & n19898 ) | ( n12312 & ~n46465 ) | ( n19898 & ~n46465 ) ;
  assign n47843 = ( n17791 & n47841 ) | ( n17791 & ~n47842 ) | ( n47841 & ~n47842 ) ;
  assign n47844 = n4805 & ~n5470 ;
  assign n47845 = n45066 ^ n38440 ^ n6497 ;
  assign n47846 = ( n12192 & n45598 ) | ( n12192 & ~n47845 ) | ( n45598 & ~n47845 ) ;
  assign n47847 = n47846 ^ n29883 ^ n7558 ;
  assign n47848 = ( n7217 & n14477 ) | ( n7217 & n47847 ) | ( n14477 & n47847 ) ;
  assign n47849 = ( n3159 & n21551 ) | ( n3159 & ~n38546 ) | ( n21551 & ~n38546 ) ;
  assign n47850 = n47849 ^ n9607 ^ n4728 ;
  assign n47851 = ( ~n1948 & n5219 ) | ( ~n1948 & n17708 ) | ( n5219 & n17708 ) ;
  assign n47852 = ~n2172 & n43138 ;
  assign n47853 = n47851 & n47852 ;
  assign n47854 = n47853 ^ n31699 ^ n23160 ;
  assign n47855 = ( n7111 & ~n8433 ) | ( n7111 & n35888 ) | ( ~n8433 & n35888 ) ;
  assign n47856 = n47855 ^ n33720 ^ n25004 ;
  assign n47857 = n6444 & n26280 ;
  assign n47858 = n17125 & n47857 ;
  assign n47859 = ( ~n13985 & n45387 ) | ( ~n13985 & n45887 ) | ( n45387 & n45887 ) ;
  assign n47860 = n26666 ^ x21 ^ 1'b0 ;
  assign n47861 = n47860 ^ n14993 ^ n3988 ;
  assign n47862 = ( n4806 & n47088 ) | ( n4806 & ~n47861 ) | ( n47088 & ~n47861 ) ;
  assign n47863 = ~n41285 & n44072 ;
  assign n47866 = ( n6297 & ~n15079 ) | ( n6297 & n18645 ) | ( ~n15079 & n18645 ) ;
  assign n47867 = n47866 ^ n31987 ^ n25777 ;
  assign n47864 = n22198 ^ n10368 ^ n7972 ;
  assign n47865 = ( n6689 & n13169 ) | ( n6689 & ~n47864 ) | ( n13169 & ~n47864 ) ;
  assign n47868 = n47867 ^ n47865 ^ n4071 ;
  assign n47869 = n47791 ^ n21215 ^ n11181 ;
  assign n47870 = ( n9359 & n39814 ) | ( n9359 & ~n47869 ) | ( n39814 & ~n47869 ) ;
  assign n47871 = n32527 & n47870 ;
  assign n47872 = n42717 ^ n36547 ^ n17797 ;
  assign n47873 = n333 | n38686 ;
  assign n47874 = n32113 | n47873 ;
  assign n47875 = n47874 ^ n35303 ^ n28783 ;
  assign n47876 = n30368 ^ n24404 ^ n12041 ;
  assign n47877 = n47876 ^ n39454 ^ n31507 ;
  assign n47878 = n47877 ^ n42441 ^ n15260 ;
  assign n47879 = n31367 ^ n19111 ^ n2181 ;
  assign n47880 = n478 & n47879 ;
  assign n47881 = n47880 ^ n16246 ^ 1'b0 ;
  assign n47884 = n4588 | n15862 ;
  assign n47885 = n47884 ^ n29525 ^ 1'b0 ;
  assign n47882 = n24191 & n39478 ;
  assign n47883 = n47882 ^ n15493 ^ 1'b0 ;
  assign n47886 = n47885 ^ n47883 ^ n2517 ;
  assign n47890 = n3349 & ~n40613 ;
  assign n47891 = ~n5759 & n47890 ;
  assign n47887 = ( n15776 & n22956 ) | ( n15776 & ~n33022 ) | ( n22956 & ~n33022 ) ;
  assign n47888 = n26937 & ~n27560 ;
  assign n47889 = ( n37338 & n47887 ) | ( n37338 & ~n47888 ) | ( n47887 & ~n47888 ) ;
  assign n47892 = n47891 ^ n47889 ^ n27346 ;
  assign n47893 = ( n2122 & n3168 ) | ( n2122 & n23258 ) | ( n3168 & n23258 ) ;
  assign n47894 = n34278 ^ n22109 ^ n3091 ;
  assign n47895 = ( ~n3530 & n3588 ) | ( ~n3530 & n37847 ) | ( n3588 & n37847 ) ;
  assign n47896 = n37555 ^ n34377 ^ n19544 ;
  assign n47897 = ( n31639 & n47895 ) | ( n31639 & ~n47896 ) | ( n47895 & ~n47896 ) ;
  assign n47898 = n47894 & n47897 ;
  assign n47899 = n8527 ^ n421 ^ 1'b0 ;
  assign n47900 = n9365 & ~n47899 ;
  assign n47901 = ( ~n1497 & n27046 ) | ( ~n1497 & n47900 ) | ( n27046 & n47900 ) ;
  assign n47902 = n45077 ^ n21207 ^ n6993 ;
  assign n47903 = n47902 ^ n25618 ^ 1'b0 ;
  assign n47904 = n10380 ^ n7989 ^ n888 ;
  assign n47905 = n47904 ^ n40264 ^ n10209 ;
  assign n47906 = ( n15698 & n40616 ) | ( n15698 & ~n47905 ) | ( n40616 & ~n47905 ) ;
  assign n47907 = n44896 ^ n6962 ^ n6618 ;
  assign n47908 = n30792 ^ n14332 ^ n1674 ;
  assign n47909 = n47908 ^ n28851 ^ n17767 ;
  assign n47910 = ( n12222 & n14196 ) | ( n12222 & n24665 ) | ( n14196 & n24665 ) ;
  assign n47911 = ( ~n37249 & n41954 ) | ( ~n37249 & n47910 ) | ( n41954 & n47910 ) ;
  assign n47912 = n42078 ^ n33175 ^ n32489 ;
  assign n47913 = ( n10616 & n10839 ) | ( n10616 & n31569 ) | ( n10839 & n31569 ) ;
  assign n47914 = ( n26967 & ~n35070 ) | ( n26967 & n47913 ) | ( ~n35070 & n47913 ) ;
  assign n47923 = n31672 ^ n7043 ^ n1853 ;
  assign n47924 = n47923 ^ n43427 ^ n386 ;
  assign n47916 = x146 & n6021 ;
  assign n47917 = n47916 ^ n4184 ^ 1'b0 ;
  assign n47915 = n5869 & ~n20268 ;
  assign n47918 = n47917 ^ n47915 ^ 1'b0 ;
  assign n47919 = n47918 ^ n35880 ^ n1696 ;
  assign n47920 = ( n1777 & ~n15145 ) | ( n1777 & n16010 ) | ( ~n15145 & n16010 ) ;
  assign n47921 = n47920 ^ n37086 ^ n14866 ;
  assign n47922 = ( n28375 & n47919 ) | ( n28375 & ~n47921 ) | ( n47919 & ~n47921 ) ;
  assign n47925 = n47924 ^ n47922 ^ n6352 ;
  assign n47926 = n47925 ^ n14996 ^ 1'b0 ;
  assign n47927 = n32525 | n47926 ;
  assign n47928 = n1741 & n2685 ;
  assign n47929 = n7152 & n47928 ;
  assign n47930 = n47929 ^ n6620 ^ 1'b0 ;
  assign n47931 = n7907 ^ n7572 ^ n4375 ;
  assign n47932 = ( ~n2532 & n37797 ) | ( ~n2532 & n47931 ) | ( n37797 & n47931 ) ;
  assign n47933 = ( n11835 & ~n17553 ) | ( n11835 & n26248 ) | ( ~n17553 & n26248 ) ;
  assign n47934 = ( ~n26122 & n47932 ) | ( ~n26122 & n47933 ) | ( n47932 & n47933 ) ;
  assign n47935 = ( n15614 & ~n27443 ) | ( n15614 & n33557 ) | ( ~n27443 & n33557 ) ;
  assign n47936 = ( n9547 & ~n14352 ) | ( n9547 & n47935 ) | ( ~n14352 & n47935 ) ;
  assign n47937 = n46060 ^ n33254 ^ n30152 ;
  assign n47938 = ( n6293 & ~n13020 ) | ( n6293 & n47937 ) | ( ~n13020 & n47937 ) ;
  assign n47942 = ( n13825 & n38740 ) | ( n13825 & ~n44269 ) | ( n38740 & ~n44269 ) ;
  assign n47939 = ( n5368 & n6523 ) | ( n5368 & ~n21226 ) | ( n6523 & ~n21226 ) ;
  assign n47940 = ~n43382 & n47939 ;
  assign n47941 = n47940 ^ n9605 ^ 1'b0 ;
  assign n47943 = n47942 ^ n47941 ^ n11796 ;
  assign n47944 = n4807 | n6760 ;
  assign n47945 = n2530 & ~n47944 ;
  assign n47946 = ( n1555 & n2838 ) | ( n1555 & n14069 ) | ( n2838 & n14069 ) ;
  assign n47947 = ( n7313 & n16168 ) | ( n7313 & ~n47946 ) | ( n16168 & ~n47946 ) ;
  assign n47948 = n28089 ^ n12238 ^ 1'b0 ;
  assign n47949 = ~n9942 & n47948 ;
  assign n47950 = ( n47945 & ~n47947 ) | ( n47945 & n47949 ) | ( ~n47947 & n47949 ) ;
  assign n47951 = ( n3097 & n33137 ) | ( n3097 & ~n34063 ) | ( n33137 & ~n34063 ) ;
  assign n47952 = n45969 ^ n27850 ^ n9484 ;
  assign n47953 = ( n19676 & n32609 ) | ( n19676 & n47952 ) | ( n32609 & n47952 ) ;
  assign n47954 = n10252 | n12213 ;
  assign n47955 = n3298 & ~n22265 ;
  assign n47956 = n47955 ^ n43104 ^ 1'b0 ;
  assign n47957 = ( n5630 & n11008 ) | ( n5630 & n45674 ) | ( n11008 & n45674 ) ;
  assign n47958 = n29817 ^ n20663 ^ n4894 ;
  assign n47959 = ( n10338 & n10814 ) | ( n10338 & ~n47958 ) | ( n10814 & ~n47958 ) ;
  assign n47960 = n29927 ^ n18326 ^ n11307 ;
  assign n47961 = ( ~n17602 & n36528 ) | ( ~n17602 & n47960 ) | ( n36528 & n47960 ) ;
  assign n47962 = n47961 ^ n18557 ^ n17425 ;
  assign n47966 = n30993 ^ n9074 ^ 1'b0 ;
  assign n47967 = n41021 | n47966 ;
  assign n47965 = n25199 ^ n5160 ^ n3089 ;
  assign n47963 = n44859 ^ n20097 ^ n12815 ;
  assign n47964 = ( n21823 & ~n25179 ) | ( n21823 & n47963 ) | ( ~n25179 & n47963 ) ;
  assign n47968 = n47967 ^ n47965 ^ n47964 ;
  assign n47969 = ( ~n5145 & n20419 ) | ( ~n5145 & n39601 ) | ( n20419 & n39601 ) ;
  assign n47970 = n27615 ^ n18696 ^ n1767 ;
  assign n47971 = ( n25131 & ~n47969 ) | ( n25131 & n47970 ) | ( ~n47969 & n47970 ) ;
  assign n47972 = n47971 ^ n43198 ^ 1'b0 ;
  assign n47974 = n3596 ^ n1048 ^ 1'b0 ;
  assign n47973 = n18185 & ~n30860 ;
  assign n47975 = n47974 ^ n47973 ^ 1'b0 ;
  assign n47976 = ( ~n26186 & n47410 ) | ( ~n26186 & n47975 ) | ( n47410 & n47975 ) ;
  assign n47977 = n47788 ^ n22033 ^ 1'b0 ;
  assign n47978 = ( n862 & n20037 ) | ( n862 & ~n20834 ) | ( n20037 & ~n20834 ) ;
  assign n47979 = ( n17025 & ~n41354 ) | ( n17025 & n47978 ) | ( ~n41354 & n47978 ) ;
  assign n47980 = n8288 ^ n5901 ^ 1'b0 ;
  assign n47981 = n19025 & ~n47980 ;
  assign n47984 = ( ~n5521 & n16492 ) | ( ~n5521 & n21325 ) | ( n16492 & n21325 ) ;
  assign n47985 = ( ~n10937 & n22678 ) | ( ~n10937 & n47984 ) | ( n22678 & n47984 ) ;
  assign n47982 = n39317 ^ n20673 ^ n839 ;
  assign n47983 = n33030 & n47982 ;
  assign n47986 = n47985 ^ n47983 ^ 1'b0 ;
  assign n47987 = n27749 ^ n3374 ^ 1'b0 ;
  assign n47988 = n47987 ^ n41290 ^ n15326 ;
  assign n47989 = n43374 ^ n41782 ^ n21717 ;
  assign n47990 = n47988 & ~n47989 ;
  assign n47991 = ( n902 & ~n1071 ) | ( n902 & n7941 ) | ( ~n1071 & n7941 ) ;
  assign n47992 = n47991 ^ n15102 ^ n4306 ;
  assign n47993 = ( n1549 & ~n17069 ) | ( n1549 & n46914 ) | ( ~n17069 & n46914 ) ;
  assign n47994 = ( n42394 & n47992 ) | ( n42394 & ~n47993 ) | ( n47992 & ~n47993 ) ;
  assign n47995 = ( n12797 & ~n36120 ) | ( n12797 & n36481 ) | ( ~n36120 & n36481 ) ;
  assign n47996 = n47995 ^ n24932 ^ 1'b0 ;
  assign n47997 = n28505 ^ n22469 ^ n16737 ;
  assign n47998 = ( ~n11953 & n21025 ) | ( ~n11953 & n47997 ) | ( n21025 & n47997 ) ;
  assign n47999 = n20940 ^ n14520 ^ 1'b0 ;
  assign n48000 = n8916 & ~n47999 ;
  assign n48001 = ( n5206 & n16305 ) | ( n5206 & n34497 ) | ( n16305 & n34497 ) ;
  assign n48002 = ( ~n39264 & n48000 ) | ( ~n39264 & n48001 ) | ( n48000 & n48001 ) ;
  assign n48003 = ( n16967 & n18042 ) | ( n16967 & n48002 ) | ( n18042 & n48002 ) ;
  assign n48004 = n36286 ^ n24343 ^ n15400 ;
  assign n48005 = n37028 ^ n27853 ^ n3112 ;
  assign n48006 = n48005 ^ n9039 ^ 1'b0 ;
  assign n48007 = n10896 & ~n48006 ;
  assign n48008 = n16425 ^ n11420 ^ x140 ;
  assign n48009 = ( n21709 & n34347 ) | ( n21709 & ~n48008 ) | ( n34347 & ~n48008 ) ;
  assign n48010 = n5632 ^ n3368 ^ 1'b0 ;
  assign n48011 = n48009 & n48010 ;
  assign n48012 = n3112 ^ x27 ^ 1'b0 ;
  assign n48013 = n48012 ^ n35236 ^ n30548 ;
  assign n48014 = n25502 ^ n21937 ^ n5229 ;
  assign n48015 = ( n32550 & n35026 ) | ( n32550 & ~n48014 ) | ( n35026 & ~n48014 ) ;
  assign n48016 = ( n22038 & n48013 ) | ( n22038 & n48015 ) | ( n48013 & n48015 ) ;
  assign n48017 = n48016 ^ n20839 ^ n20339 ;
  assign n48022 = n16290 ^ n7414 ^ n7165 ;
  assign n48023 = n18543 | n48022 ;
  assign n48020 = n19984 ^ n16346 ^ n15326 ;
  assign n48018 = n19363 & ~n43010 ;
  assign n48019 = n3619 | n48018 ;
  assign n48021 = n48020 ^ n48019 ^ 1'b0 ;
  assign n48024 = n48023 ^ n48021 ^ n8429 ;
  assign n48025 = ~n781 & n10238 ;
  assign n48026 = n48025 ^ n15304 ^ 1'b0 ;
  assign n48027 = n48026 ^ n37524 ^ n22938 ;
  assign n48028 = n30025 ^ n22411 ^ 1'b0 ;
  assign n48029 = n13040 ^ n4814 ^ n789 ;
  assign n48030 = ( n11754 & n23857 ) | ( n11754 & n24525 ) | ( n23857 & n24525 ) ;
  assign n48031 = n48030 ^ n36368 ^ 1'b0 ;
  assign n48032 = ( n34578 & n48029 ) | ( n34578 & ~n48031 ) | ( n48029 & ~n48031 ) ;
  assign n48033 = ~n43202 & n48032 ;
  assign n48034 = n18432 ^ n10832 ^ n3907 ;
  assign n48035 = ( n2515 & n15116 ) | ( n2515 & n48034 ) | ( n15116 & n48034 ) ;
  assign n48036 = ( n18722 & n40381 ) | ( n18722 & n48035 ) | ( n40381 & n48035 ) ;
  assign n48037 = ~n12997 & n39688 ;
  assign n48038 = n35306 & n48037 ;
  assign n48039 = n48038 ^ n26022 ^ n14568 ;
  assign n48045 = n36904 ^ n21554 ^ n2205 ;
  assign n48043 = n9462 ^ n6471 ^ n5743 ;
  assign n48042 = ( n19910 & ~n24370 ) | ( n19910 & n27052 ) | ( ~n24370 & n27052 ) ;
  assign n48044 = n48043 ^ n48042 ^ x228 ;
  assign n48040 = n40207 ^ n20802 ^ n17691 ;
  assign n48041 = ( ~n30840 & n35660 ) | ( ~n30840 & n48040 ) | ( n35660 & n48040 ) ;
  assign n48046 = n48045 ^ n48044 ^ n48041 ;
  assign n48047 = n19924 | n37013 ;
  assign n48048 = n39268 | n48047 ;
  assign n48049 = ( n7737 & ~n9781 ) | ( n7737 & n12978 ) | ( ~n9781 & n12978 ) ;
  assign n48050 = ( n499 & n27214 ) | ( n499 & ~n48049 ) | ( n27214 & ~n48049 ) ;
  assign n48051 = n39430 & n48050 ;
  assign n48052 = ( n752 & ~n6509 ) | ( n752 & n30957 ) | ( ~n6509 & n30957 ) ;
  assign n48053 = n18781 & n48052 ;
  assign n48054 = ( n4623 & ~n34343 ) | ( n4623 & n48053 ) | ( ~n34343 & n48053 ) ;
  assign n48055 = ( n24191 & ~n27491 ) | ( n24191 & n47623 ) | ( ~n27491 & n47623 ) ;
  assign n48056 = n48055 ^ n12275 ^ x55 ;
  assign n48057 = n48056 ^ n33873 ^ n31869 ;
  assign n48058 = ( n27684 & n27868 ) | ( n27684 & n48057 ) | ( n27868 & n48057 ) ;
  assign n48059 = n17184 ^ n14487 ^ n4849 ;
  assign n48060 = ( ~n3294 & n26997 ) | ( ~n3294 & n48059 ) | ( n26997 & n48059 ) ;
  assign n48061 = n48060 ^ n34669 ^ n12969 ;
  assign n48062 = n9997 ^ n4475 ^ n1308 ;
  assign n48063 = n28584 ^ n3924 ^ n2273 ;
  assign n48064 = n48063 ^ n19017 ^ n1076 ;
  assign n48065 = n44654 ^ n7905 ^ n2277 ;
  assign n48066 = n48065 ^ n22867 ^ 1'b0 ;
  assign n48067 = n13615 ^ n5023 ^ n3376 ;
  assign n48068 = n48067 ^ n28170 ^ n23832 ;
  assign n48069 = n27434 ^ n11225 ^ n9658 ;
  assign n48070 = n48069 ^ n44691 ^ n23570 ;
  assign n48071 = ( ~n23291 & n25050 ) | ( ~n23291 & n48070 ) | ( n25050 & n48070 ) ;
  assign n48072 = ( n22308 & n23527 ) | ( n22308 & n36368 ) | ( n23527 & n36368 ) ;
  assign n48073 = n33486 ^ n16063 ^ n5207 ;
  assign n48074 = n48073 ^ n16382 ^ n6299 ;
  assign n48075 = n48074 ^ n35397 ^ n13095 ;
  assign n48076 = ( n17818 & ~n25895 ) | ( n17818 & n36657 ) | ( ~n25895 & n36657 ) ;
  assign n48077 = n22930 ^ n14161 ^ 1'b0 ;
  assign n48078 = n13814 & n20396 ;
  assign n48079 = n48078 ^ n29176 ^ 1'b0 ;
  assign n48080 = n48079 ^ n20071 ^ 1'b0 ;
  assign n48082 = ( n13980 & n24171 ) | ( n13980 & n33892 ) | ( n24171 & n33892 ) ;
  assign n48081 = n16448 ^ n15268 ^ n2677 ;
  assign n48083 = n48082 ^ n48081 ^ n6513 ;
  assign n48084 = n13293 ^ n4364 ^ n2912 ;
  assign n48085 = n3101 & ~n48084 ;
  assign n48086 = n48085 ^ n33248 ^ n21938 ;
  assign n48087 = ( ~n6606 & n21666 ) | ( ~n6606 & n43037 ) | ( n21666 & n43037 ) ;
  assign n48090 = n41426 ^ n21633 ^ n11708 ;
  assign n48088 = ( n3653 & ~n7353 ) | ( n3653 & n27897 ) | ( ~n7353 & n27897 ) ;
  assign n48089 = n48088 ^ n13342 ^ n11564 ;
  assign n48091 = n48090 ^ n48089 ^ n6100 ;
  assign n48095 = n22847 & ~n41968 ;
  assign n48096 = n48095 ^ n9961 ^ 1'b0 ;
  assign n48092 = n26699 ^ n21846 ^ n2206 ;
  assign n48093 = n48092 ^ n46333 ^ n34645 ;
  assign n48094 = ~n9240 & n48093 ;
  assign n48097 = n48096 ^ n48094 ^ 1'b0 ;
  assign n48098 = n21207 ^ n5576 ^ 1'b0 ;
  assign n48099 = n25590 & ~n48098 ;
  assign n48100 = n17768 | n28604 ;
  assign n48101 = n48099 | n48100 ;
  assign n48102 = n4644 & n9433 ;
  assign n48103 = n43079 | n48102 ;
  assign n48104 = n48101 | n48103 ;
  assign n48105 = ( n6596 & n7619 ) | ( n6596 & ~n9882 ) | ( n7619 & ~n9882 ) ;
  assign n48106 = n48105 ^ n32963 ^ n32663 ;
  assign n48107 = ( ~n38833 & n47002 ) | ( ~n38833 & n48106 ) | ( n47002 & n48106 ) ;
  assign n48109 = n34081 ^ n1181 ^ 1'b0 ;
  assign n48108 = ( ~n11647 & n15473 ) | ( ~n11647 & n37652 ) | ( n15473 & n37652 ) ;
  assign n48110 = n48109 ^ n48108 ^ n41423 ;
  assign n48111 = ( ~n5007 & n45560 ) | ( ~n5007 & n48110 ) | ( n45560 & n48110 ) ;
  assign n48112 = ( n16976 & n22568 ) | ( n16976 & n29616 ) | ( n22568 & n29616 ) ;
  assign n48113 = n3114 & n4414 ;
  assign n48114 = n48113 ^ n38643 ^ 1'b0 ;
  assign n48115 = n48112 | n48114 ;
  assign n48116 = ( n24635 & n28000 ) | ( n24635 & n40781 ) | ( n28000 & n40781 ) ;
  assign n48117 = n3804 | n30651 ;
  assign n48118 = ( n16024 & n22885 ) | ( n16024 & n25552 ) | ( n22885 & n25552 ) ;
  assign n48119 = ~n285 & n34604 ;
  assign n48120 = n28696 & n48119 ;
  assign n48121 = n13403 ^ n1897 ^ n1333 ;
  assign n48122 = n3391 | n29715 ;
  assign n48123 = ~n12702 & n48122 ;
  assign n48124 = ( n23778 & n40436 ) | ( n23778 & ~n48123 ) | ( n40436 & ~n48123 ) ;
  assign n48125 = n48124 ^ n12733 ^ n5024 ;
  assign n48126 = ( ~n47660 & n48121 ) | ( ~n47660 & n48125 ) | ( n48121 & n48125 ) ;
  assign n48127 = ( n2429 & ~n7584 ) | ( n2429 & n9433 ) | ( ~n7584 & n9433 ) ;
  assign n48128 = n48127 ^ n29541 ^ n4514 ;
  assign n48129 = ( n26080 & ~n41432 ) | ( n26080 & n48128 ) | ( ~n41432 & n48128 ) ;
  assign n48130 = ( ~n4630 & n39015 ) | ( ~n4630 & n44192 ) | ( n39015 & n44192 ) ;
  assign n48131 = ( n4995 & n33041 ) | ( n4995 & n39035 ) | ( n33041 & n39035 ) ;
  assign n48132 = ( n21576 & ~n29336 ) | ( n21576 & n36709 ) | ( ~n29336 & n36709 ) ;
  assign n48133 = n3495 & n48132 ;
  assign n48134 = n48133 ^ n8082 ^ 1'b0 ;
  assign n48135 = n48134 ^ n31858 ^ n8895 ;
  assign n48136 = ( n5238 & n15577 ) | ( n5238 & ~n31864 ) | ( n15577 & ~n31864 ) ;
  assign n48137 = ( n801 & n1458 ) | ( n801 & n48136 ) | ( n1458 & n48136 ) ;
  assign n48138 = n48137 ^ n28632 ^ n13672 ;
  assign n48139 = ( ~n8475 & n8731 ) | ( ~n8475 & n10107 ) | ( n8731 & n10107 ) ;
  assign n48140 = n48139 ^ n11622 ^ n11605 ;
  assign n48141 = n48140 ^ n31428 ^ n6911 ;
  assign n48144 = ( n11650 & ~n18527 ) | ( n11650 & n25664 ) | ( ~n18527 & n25664 ) ;
  assign n48145 = ( n10795 & n41629 ) | ( n10795 & n48144 ) | ( n41629 & n48144 ) ;
  assign n48142 = n8426 & ~n28111 ;
  assign n48143 = ( n28008 & n28617 ) | ( n28008 & n48142 ) | ( n28617 & n48142 ) ;
  assign n48146 = n48145 ^ n48143 ^ n34261 ;
  assign n48147 = n41024 ^ n38962 ^ 1'b0 ;
  assign n48148 = n33691 ^ n28704 ^ n4098 ;
  assign n48149 = ( n4412 & ~n31022 ) | ( n4412 & n32435 ) | ( ~n31022 & n32435 ) ;
  assign n48150 = ( n29276 & ~n48148 ) | ( n29276 & n48149 ) | ( ~n48148 & n48149 ) ;
  assign n48151 = n48150 ^ n20302 ^ n14171 ;
  assign n48152 = ( n5107 & n17567 ) | ( n5107 & ~n48151 ) | ( n17567 & ~n48151 ) ;
  assign n48153 = ( ~n2861 & n45631 ) | ( ~n2861 & n48152 ) | ( n45631 & n48152 ) ;
  assign n48154 = n1558 & n2015 ;
  assign n48155 = n48154 ^ n18001 ^ 1'b0 ;
  assign n48156 = ( ~n4468 & n34589 ) | ( ~n4468 & n48155 ) | ( n34589 & n48155 ) ;
  assign n48157 = ~n21478 & n30886 ;
  assign n48158 = ~n15589 & n48157 ;
  assign n48159 = ( ~n9440 & n11216 ) | ( ~n9440 & n12653 ) | ( n11216 & n12653 ) ;
  assign n48160 = ( n15793 & n48158 ) | ( n15793 & n48159 ) | ( n48158 & n48159 ) ;
  assign n48161 = ( ~n1156 & n19166 ) | ( ~n1156 & n24156 ) | ( n19166 & n24156 ) ;
  assign n48162 = n31562 | n35054 ;
  assign n48163 = n48162 ^ x80 ^ 1'b0 ;
  assign n48164 = ( ~n7265 & n19585 ) | ( ~n7265 & n48163 ) | ( n19585 & n48163 ) ;
  assign n48165 = ( ~n3443 & n5099 ) | ( ~n3443 & n13390 ) | ( n5099 & n13390 ) ;
  assign n48166 = ( ~n487 & n33342 ) | ( ~n487 & n48165 ) | ( n33342 & n48165 ) ;
  assign n48167 = n48166 ^ n46227 ^ n10211 ;
  assign n48168 = n48167 ^ n18277 ^ 1'b0 ;
  assign n48169 = n13571 | n48145 ;
  assign n48170 = n19294 & ~n48169 ;
  assign n48171 = n48170 ^ n44189 ^ n3236 ;
  assign n48172 = ( n3019 & ~n4955 ) | ( n3019 & n48171 ) | ( ~n4955 & n48171 ) ;
  assign n48173 = n7598 ^ n4064 ^ n2438 ;
  assign n48174 = ( n3168 & n11831 ) | ( n3168 & ~n48173 ) | ( n11831 & ~n48173 ) ;
  assign n48175 = n39231 ^ n6252 ^ n4967 ;
  assign n48176 = n9807 | n12701 ;
  assign n48177 = ~n48175 & n48176 ;
  assign n48178 = n48177 ^ n9434 ^ 1'b0 ;
  assign n48179 = n44921 ^ n37584 ^ n13983 ;
  assign n48180 = n23771 & n36760 ;
  assign n48181 = n40651 ^ n23383 ^ n20557 ;
  assign n48182 = ( n571 & n44479 ) | ( n571 & ~n48181 ) | ( n44479 & ~n48181 ) ;
  assign n48183 = ( ~n23265 & n29086 ) | ( ~n23265 & n43075 ) | ( n29086 & n43075 ) ;
  assign n48184 = n31205 ^ n29995 ^ 1'b0 ;
  assign n48185 = n22037 ^ n18199 ^ 1'b0 ;
  assign n48186 = n9748 ^ n4736 ^ 1'b0 ;
  assign n48187 = ~n14613 & n48186 ;
  assign n48188 = ( n8431 & ~n22236 ) | ( n8431 & n48187 ) | ( ~n22236 & n48187 ) ;
  assign n48189 = ( n8380 & n16545 ) | ( n8380 & n21351 ) | ( n16545 & n21351 ) ;
  assign n48190 = n48189 ^ n35509 ^ n1719 ;
  assign n48191 = n7282 & n35397 ;
  assign n48192 = n18133 & n48191 ;
  assign n48193 = n8611 | n33948 ;
  assign n48194 = n48193 ^ n41164 ^ 1'b0 ;
  assign n48195 = n34962 ^ n18188 ^ n7696 ;
  assign n48196 = ( n7020 & ~n27424 ) | ( n7020 & n48195 ) | ( ~n27424 & n48195 ) ;
  assign n48197 = ( ~n2959 & n8694 ) | ( ~n2959 & n11443 ) | ( n8694 & n11443 ) ;
  assign n48198 = n48197 ^ n15630 ^ n9907 ;
  assign n48199 = n20914 ^ n13996 ^ n7786 ;
  assign n48200 = n26553 ^ n18149 ^ n12250 ;
  assign n48201 = n40877 & n45604 ;
  assign n48202 = n5957 & n48201 ;
  assign n48203 = n12191 | n48202 ;
  assign n48205 = n35786 ^ n29308 ^ n9415 ;
  assign n48206 = ( n3496 & ~n12836 ) | ( n3496 & n48205 ) | ( ~n12836 & n48205 ) ;
  assign n48204 = ( n7721 & ~n14041 ) | ( n7721 & n38224 ) | ( ~n14041 & n38224 ) ;
  assign n48207 = n48206 ^ n48204 ^ n46554 ;
  assign n48209 = n1705 | n17158 ;
  assign n48210 = ( n8990 & n43546 ) | ( n8990 & ~n48209 ) | ( n43546 & ~n48209 ) ;
  assign n48208 = ( n13162 & n29956 ) | ( n13162 & ~n48038 ) | ( n29956 & ~n48038 ) ;
  assign n48211 = n48210 ^ n48208 ^ n1072 ;
  assign n48213 = ( n1637 & n13727 ) | ( n1637 & ~n23168 ) | ( n13727 & ~n23168 ) ;
  assign n48214 = n48213 ^ n19623 ^ 1'b0 ;
  assign n48215 = n15069 | n48214 ;
  assign n48212 = n45285 ^ n8909 ^ n2303 ;
  assign n48216 = n48215 ^ n48212 ^ n20059 ;
  assign n48219 = n2014 & ~n13329 ;
  assign n48217 = ( n722 & n4920 ) | ( n722 & ~n33507 ) | ( n4920 & ~n33507 ) ;
  assign n48218 = n48217 ^ n37676 ^ n418 ;
  assign n48220 = n48219 ^ n48218 ^ n29829 ;
  assign n48221 = ( x161 & n7744 ) | ( x161 & n19388 ) | ( n7744 & n19388 ) ;
  assign n48222 = n7219 ^ n2421 ^ 1'b0 ;
  assign n48223 = n2084 & ~n48222 ;
  assign n48224 = n48223 ^ n38534 ^ n15311 ;
  assign n48225 = ( n1725 & n48221 ) | ( n1725 & n48224 ) | ( n48221 & n48224 ) ;
  assign n48226 = ( ~n2371 & n17073 ) | ( ~n2371 & n43495 ) | ( n17073 & n43495 ) ;
  assign n48229 = ( n6508 & n17331 ) | ( n6508 & ~n36246 ) | ( n17331 & ~n36246 ) ;
  assign n48227 = n32228 ^ n29752 ^ 1'b0 ;
  assign n48228 = n30983 & ~n48227 ;
  assign n48230 = n48229 ^ n48228 ^ n35059 ;
  assign n48231 = n47410 ^ n35154 ^ 1'b0 ;
  assign n48232 = n41034 & ~n48231 ;
  assign n48233 = n48232 ^ n13183 ^ 1'b0 ;
  assign n48234 = ~n5911 & n48233 ;
  assign n48235 = n48234 ^ n43403 ^ n706 ;
  assign n48236 = ~n13486 & n20412 ;
  assign n48237 = ( ~n6539 & n13171 ) | ( ~n6539 & n15219 ) | ( n13171 & n15219 ) ;
  assign n48238 = n41662 & n48237 ;
  assign n48239 = n48238 ^ n12947 ^ 1'b0 ;
  assign n48240 = n37683 ^ n10016 ^ 1'b0 ;
  assign n48241 = n48240 ^ n21445 ^ n6581 ;
  assign n48242 = n48241 ^ n10454 ^ n9191 ;
  assign n48243 = ( n42719 & n48239 ) | ( n42719 & n48242 ) | ( n48239 & n48242 ) ;
  assign n48244 = ( n22244 & n28240 ) | ( n22244 & n39470 ) | ( n28240 & n39470 ) ;
  assign n48245 = n11717 ^ n4485 ^ n2898 ;
  assign n48246 = n48245 ^ n35368 ^ n15455 ;
  assign n48247 = n38538 ^ n35688 ^ n26031 ;
  assign n48252 = ( ~n14000 & n30690 ) | ( ~n14000 & n36937 ) | ( n30690 & n36937 ) ;
  assign n48250 = ( ~n2044 & n12527 ) | ( ~n2044 & n12555 ) | ( n12527 & n12555 ) ;
  assign n48251 = n48250 ^ n28097 ^ n17423 ;
  assign n48248 = ~n7506 & n19554 ;
  assign n48249 = n24715 & n48248 ;
  assign n48253 = n48252 ^ n48251 ^ n48249 ;
  assign n48254 = ( n16724 & n21209 ) | ( n16724 & ~n39842 ) | ( n21209 & ~n39842 ) ;
  assign n48255 = n48254 ^ n43880 ^ n21921 ;
  assign n48256 = ( n11566 & ~n12159 ) | ( n11566 & n35021 ) | ( ~n12159 & n35021 ) ;
  assign n48257 = n40892 ^ n28908 ^ n27117 ;
  assign n48258 = ( n7348 & ~n16827 ) | ( n7348 & n48257 ) | ( ~n16827 & n48257 ) ;
  assign n48259 = ( ~n9258 & n30535 ) | ( ~n9258 & n32429 ) | ( n30535 & n32429 ) ;
  assign n48260 = n48259 ^ n7222 ^ 1'b0 ;
  assign n48261 = n8601 ^ n5268 ^ 1'b0 ;
  assign n48262 = n31958 & n48261 ;
  assign n48263 = n48262 ^ n18869 ^ n1367 ;
  assign n48264 = ( n6675 & n15111 ) | ( n6675 & ~n48263 ) | ( n15111 & ~n48263 ) ;
  assign n48265 = n22024 ^ n12447 ^ n8279 ;
  assign n48266 = n36909 ^ n31062 ^ n13345 ;
  assign n48271 = n20176 ^ n5432 ^ n3597 ;
  assign n48268 = n21311 ^ n1075 ^ 1'b0 ;
  assign n48269 = n23232 & n48268 ;
  assign n48267 = n4863 | n44415 ;
  assign n48270 = n48269 ^ n48267 ^ 1'b0 ;
  assign n48272 = n48271 ^ n48270 ^ n7895 ;
  assign n48273 = n35524 ^ n34720 ^ n27916 ;
  assign n48274 = ( n625 & n26753 ) | ( n625 & n38844 ) | ( n26753 & n38844 ) ;
  assign n48275 = n5358 & ~n9923 ;
  assign n48276 = n40703 ^ n3628 ^ n2890 ;
  assign n48277 = ( n727 & ~n16567 ) | ( n727 & n18507 ) | ( ~n16567 & n18507 ) ;
  assign n48278 = n48277 ^ n32771 ^ n14483 ;
  assign n48279 = n40520 & n48278 ;
  assign n48283 = ( n5169 & n18487 ) | ( n5169 & n25333 ) | ( n18487 & n25333 ) ;
  assign n48280 = n16662 ^ n3206 ^ 1'b0 ;
  assign n48281 = n32875 | n48280 ;
  assign n48282 = n46319 & ~n48281 ;
  assign n48284 = n48283 ^ n48282 ^ n17309 ;
  assign n48287 = ( n15092 & n18052 ) | ( n15092 & n18628 ) | ( n18052 & n18628 ) ;
  assign n48285 = n1705 & ~n12031 ;
  assign n48286 = n48285 ^ n32622 ^ 1'b0 ;
  assign n48288 = n48287 ^ n48286 ^ 1'b0 ;
  assign n48290 = ( n1388 & n18223 ) | ( n1388 & ~n42635 ) | ( n18223 & ~n42635 ) ;
  assign n48291 = n48290 ^ n31297 ^ 1'b0 ;
  assign n48292 = ~n5379 & n48291 ;
  assign n48289 = n22340 ^ n21222 ^ n7147 ;
  assign n48293 = n48292 ^ n48289 ^ n42427 ;
  assign n48294 = ( ~n4462 & n13281 ) | ( ~n4462 & n16761 ) | ( n13281 & n16761 ) ;
  assign n48295 = n9534 | n37306 ;
  assign n48296 = n48295 ^ n44544 ^ 1'b0 ;
  assign n48297 = n12855 ^ n9047 ^ 1'b0 ;
  assign n48298 = n41945 & n48297 ;
  assign n48299 = ( n16824 & n20538 ) | ( n16824 & ~n27341 ) | ( n20538 & ~n27341 ) ;
  assign n48300 = n48299 ^ n10445 ^ n10275 ;
  assign n48301 = ( n1624 & n17005 ) | ( n1624 & ~n27500 ) | ( n17005 & ~n27500 ) ;
  assign n48302 = n48301 ^ n24015 ^ n9757 ;
  assign n48303 = ( n10367 & n12512 ) | ( n10367 & ~n48302 ) | ( n12512 & ~n48302 ) ;
  assign n48304 = ( n30158 & ~n39447 ) | ( n30158 & n48303 ) | ( ~n39447 & n48303 ) ;
  assign n48305 = ( ~n6841 & n8579 ) | ( ~n6841 & n11946 ) | ( n8579 & n11946 ) ;
  assign n48306 = n48305 ^ n40783 ^ n8554 ;
  assign n48307 = n48306 ^ n8665 ^ 1'b0 ;
  assign n48308 = n26453 ^ n25772 ^ n8484 ;
  assign n48309 = n48308 ^ n20373 ^ n1662 ;
  assign n48310 = n31343 ^ n27368 ^ n9171 ;
  assign n48311 = ( n446 & ~n9754 ) | ( n446 & n35475 ) | ( ~n9754 & n35475 ) ;
  assign n48312 = n42537 ^ n27642 ^ 1'b0 ;
  assign n48313 = ( ~n19740 & n35231 ) | ( ~n19740 & n48312 ) | ( n35231 & n48312 ) ;
  assign n48314 = n6372 & ~n13419 ;
  assign n48315 = n48314 ^ n39970 ^ 1'b0 ;
  assign n48316 = n36956 ^ n1824 ^ 1'b0 ;
  assign n48317 = ~n12052 & n48316 ;
  assign n48318 = ( n8229 & n23635 ) | ( n8229 & ~n35235 ) | ( n23635 & ~n35235 ) ;
  assign n48319 = n48318 ^ n12297 ^ n4683 ;
  assign n48320 = n48319 ^ n45220 ^ n11473 ;
  assign n48321 = ~n7053 & n38338 ;
  assign n48322 = ~n36687 & n48321 ;
  assign n48323 = n40147 ^ n2791 ^ 1'b0 ;
  assign n48324 = n48322 | n48323 ;
  assign n48325 = n48324 ^ n46735 ^ n20818 ;
  assign n48326 = n24213 ^ n21702 ^ n20481 ;
  assign n48327 = n48326 ^ n27292 ^ 1'b0 ;
  assign n48328 = ( ~n31666 & n33806 ) | ( ~n31666 & n36544 ) | ( n33806 & n36544 ) ;
  assign n48332 = n18981 & ~n20917 ;
  assign n48333 = n48332 ^ n42219 ^ 1'b0 ;
  assign n48329 = n31251 ^ n8734 ^ n7933 ;
  assign n48330 = n48329 ^ n32615 ^ 1'b0 ;
  assign n48331 = n14628 & n48330 ;
  assign n48334 = n48333 ^ n48331 ^ n42685 ;
  assign n48335 = ~n22139 & n27316 ;
  assign n48336 = n48335 ^ n16763 ^ 1'b0 ;
  assign n48337 = ( n12411 & n27193 ) | ( n12411 & ~n48336 ) | ( n27193 & ~n48336 ) ;
  assign n48338 = n48337 ^ n15732 ^ n11535 ;
  assign n48339 = ( n30315 & ~n30995 ) | ( n30315 & n40766 ) | ( ~n30995 & n40766 ) ;
  assign n48340 = n34418 | n48339 ;
  assign n48341 = n15157 & ~n48340 ;
  assign n48342 = n46251 ^ n32003 ^ n17374 ;
  assign n48343 = ( n2744 & ~n13840 ) | ( n2744 & n48342 ) | ( ~n13840 & n48342 ) ;
  assign n48344 = ~n961 & n43547 ;
  assign n48345 = ~n48343 & n48344 ;
  assign n48346 = n43388 ^ n42169 ^ n31863 ;
  assign n48348 = ( n6397 & ~n11945 ) | ( n6397 & n28376 ) | ( ~n11945 & n28376 ) ;
  assign n48347 = n41648 & ~n43325 ;
  assign n48349 = n48348 ^ n48347 ^ 1'b0 ;
  assign n48350 = ( n33245 & n47042 ) | ( n33245 & ~n48349 ) | ( n47042 & ~n48349 ) ;
  assign n48351 = n45406 ^ n44859 ^ n8691 ;
  assign n48354 = ( n22512 & n40786 ) | ( n22512 & n40938 ) | ( n40786 & n40938 ) ;
  assign n48352 = n28740 ^ n7262 ^ n1208 ;
  assign n48353 = n48352 ^ n44083 ^ n5539 ;
  assign n48355 = n48354 ^ n48353 ^ n16020 ;
  assign n48356 = n17959 | n39320 ;
  assign n48357 = ~n1084 & n42358 ;
  assign n48363 = n20460 ^ n17357 ^ n12359 ;
  assign n48358 = ~n1757 & n11083 ;
  assign n48359 = n48358 ^ n12057 ^ 1'b0 ;
  assign n48360 = ( x120 & n13361 ) | ( x120 & n48359 ) | ( n13361 & n48359 ) ;
  assign n48361 = n48360 ^ n24082 ^ n15000 ;
  assign n48362 = n48361 ^ n47851 ^ n30716 ;
  assign n48364 = n48363 ^ n48362 ^ n29912 ;
  assign n48365 = n48364 ^ n27061 ^ n8676 ;
  assign n48366 = n18382 ^ n16969 ^ n3831 ;
  assign n48367 = ( ~n39871 & n44773 ) | ( ~n39871 & n48366 ) | ( n44773 & n48366 ) ;
  assign n48368 = n48367 ^ n25316 ^ n11117 ;
  assign n48369 = n36578 ^ n34726 ^ n12708 ;
  assign n48370 = ( n4473 & n7010 ) | ( n4473 & n13357 ) | ( n7010 & n13357 ) ;
  assign n48371 = ~n684 & n21822 ;
  assign n48372 = n48371 ^ n9937 ^ 1'b0 ;
  assign n48373 = n31292 & n48372 ;
  assign n48374 = ~n48370 & n48373 ;
  assign n48375 = n27553 ^ n511 ^ 1'b0 ;
  assign n48377 = ( n1957 & ~n5996 ) | ( n1957 & n9138 ) | ( ~n5996 & n9138 ) ;
  assign n48376 = n25131 ^ n4523 ^ n3744 ;
  assign n48378 = n48377 ^ n48376 ^ n19107 ;
  assign n48379 = ( n1921 & n10772 ) | ( n1921 & n30324 ) | ( n10772 & n30324 ) ;
  assign n48380 = n37709 ^ n7489 ^ n7057 ;
  assign n48381 = n44864 ^ n22165 ^ n2470 ;
  assign n48382 = n46558 ^ n43486 ^ n4028 ;
  assign n48383 = n32734 ^ n25494 ^ 1'b0 ;
  assign n48384 = ( n11734 & n13473 ) | ( n11734 & n16611 ) | ( n13473 & n16611 ) ;
  assign n48385 = ( ~n280 & n25963 ) | ( ~n280 & n48384 ) | ( n25963 & n48384 ) ;
  assign n48386 = n48385 ^ n35520 ^ n26122 ;
  assign n48387 = n39842 ^ n37671 ^ n28877 ;
  assign n48388 = n37606 ^ n909 ^ 1'b0 ;
  assign n48389 = ( n894 & n6775 ) | ( n894 & n48388 ) | ( n6775 & n48388 ) ;
  assign n48394 = ( n2919 & n3617 ) | ( n2919 & n17719 ) | ( n3617 & n17719 ) ;
  assign n48390 = n22118 ^ n1664 ^ n690 ;
  assign n48391 = ( n3199 & ~n9950 ) | ( n3199 & n19204 ) | ( ~n9950 & n19204 ) ;
  assign n48392 = n48391 ^ n17858 ^ n16389 ;
  assign n48393 = ( n35219 & n48390 ) | ( n35219 & ~n48392 ) | ( n48390 & ~n48392 ) ;
  assign n48395 = n48394 ^ n48393 ^ n43700 ;
  assign n48396 = n3651 & ~n3790 ;
  assign n48397 = n48395 & n48396 ;
  assign n48398 = n5067 | n24500 ;
  assign n48399 = n48398 ^ n1653 ^ 1'b0 ;
  assign n48400 = n48399 ^ n42556 ^ n10909 ;
  assign n48401 = n13769 ^ x145 ^ 1'b0 ;
  assign n48402 = n48401 ^ n47939 ^ n10380 ;
  assign n48403 = n48402 ^ n36974 ^ n36871 ;
  assign n48404 = n2933 & ~n48403 ;
  assign n48405 = ~n48400 & n48404 ;
  assign n48406 = n28980 ^ n24467 ^ n9329 ;
  assign n48408 = ( n3654 & n5024 ) | ( n3654 & ~n32629 ) | ( n5024 & ~n32629 ) ;
  assign n48407 = n18301 ^ n9961 ^ n4120 ;
  assign n48409 = n48408 ^ n48407 ^ n18656 ;
  assign n48410 = n4463 & ~n25530 ;
  assign n48411 = n48410 ^ n10105 ^ 1'b0 ;
  assign n48412 = ( n4317 & n14264 ) | ( n4317 & ~n48411 ) | ( n14264 & ~n48411 ) ;
  assign n48413 = ( n6183 & n27285 ) | ( n6183 & ~n30699 ) | ( n27285 & ~n30699 ) ;
  assign n48414 = n48413 ^ n42365 ^ n1018 ;
  assign n48415 = ( ~n1173 & n5204 ) | ( ~n1173 & n14520 ) | ( n5204 & n14520 ) ;
  assign n48416 = ( n23669 & ~n30694 ) | ( n23669 & n48415 ) | ( ~n30694 & n48415 ) ;
  assign n48417 = ( n12940 & ~n40074 ) | ( n12940 & n48416 ) | ( ~n40074 & n48416 ) ;
  assign n48418 = n17357 ^ n14926 ^ n1121 ;
  assign n48419 = n48418 ^ n38671 ^ n8890 ;
  assign n48420 = n28279 ^ n11070 ^ n1620 ;
  assign n48421 = n48420 ^ n14202 ^ n10579 ;
  assign n48422 = n5193 & ~n18082 ;
  assign n48423 = ~n9225 & n48422 ;
  assign n48424 = ( n2010 & ~n28418 ) | ( n2010 & n48423 ) | ( ~n28418 & n48423 ) ;
  assign n48425 = ( n9317 & ~n20330 ) | ( n9317 & n25371 ) | ( ~n20330 & n25371 ) ;
  assign n48426 = ( n2392 & n48424 ) | ( n2392 & n48425 ) | ( n48424 & n48425 ) ;
  assign n48427 = n48426 ^ n11679 ^ 1'b0 ;
  assign n48428 = n45438 | n48427 ;
  assign n48429 = ~n14176 & n28515 ;
  assign n48430 = ~n15713 & n48429 ;
  assign n48431 = n4498 & n29878 ;
  assign n48432 = n48430 & n48431 ;
  assign n48433 = ( x73 & ~n14930 ) | ( x73 & n30131 ) | ( ~n14930 & n30131 ) ;
  assign n48434 = n41957 ^ n14791 ^ n13436 ;
  assign n48435 = ( n14744 & n22630 ) | ( n14744 & n48434 ) | ( n22630 & n48434 ) ;
  assign n48436 = n18816 ^ n8115 ^ 1'b0 ;
  assign n48437 = n42948 | n48436 ;
  assign n48438 = ~n10206 & n14380 ;
  assign n48439 = n48438 ^ n6277 ^ 1'b0 ;
  assign n48440 = n48439 ^ n30349 ^ n17932 ;
  assign n48441 = ( n11370 & n32196 ) | ( n11370 & n48440 ) | ( n32196 & n48440 ) ;
  assign n48442 = n42218 ^ n26551 ^ n23087 ;
  assign n48443 = n48442 ^ n10135 ^ n8363 ;
  assign n48447 = n17634 ^ n7568 ^ n5757 ;
  assign n48444 = ( n3571 & ~n16481 ) | ( n3571 & n16822 ) | ( ~n16481 & n16822 ) ;
  assign n48445 = n7371 & ~n47146 ;
  assign n48446 = ~n48444 & n48445 ;
  assign n48448 = n48447 ^ n48446 ^ n23076 ;
  assign n48449 = n26133 ^ n3881 ^ n371 ;
  assign n48451 = ( n1657 & n3181 ) | ( n1657 & ~n13661 ) | ( n3181 & ~n13661 ) ;
  assign n48450 = n22380 ^ n10134 ^ n4458 ;
  assign n48452 = n48451 ^ n48450 ^ n10060 ;
  assign n48453 = n26594 ^ n17050 ^ n6389 ;
  assign n48457 = ( n421 & n12609 ) | ( n421 & n14384 ) | ( n12609 & n14384 ) ;
  assign n48458 = n48457 ^ n38324 ^ n12327 ;
  assign n48454 = ( ~n7654 & n27533 ) | ( ~n7654 & n27977 ) | ( n27533 & n27977 ) ;
  assign n48455 = n48454 ^ n7063 ^ n808 ;
  assign n48456 = ( ~n11457 & n21826 ) | ( ~n11457 & n48455 ) | ( n21826 & n48455 ) ;
  assign n48459 = n48458 ^ n48456 ^ n37786 ;
  assign n48460 = n42834 ^ n13574 ^ n11765 ;
  assign n48461 = ( n4090 & n12012 ) | ( n4090 & ~n36395 ) | ( n12012 & ~n36395 ) ;
  assign n48462 = n44864 ^ n17547 ^ n15341 ;
  assign n48463 = n29244 ^ n25387 ^ 1'b0 ;
  assign n48464 = n48463 ^ n32168 ^ n21731 ;
  assign n48465 = ( ~n29812 & n33955 ) | ( ~n29812 & n39929 ) | ( n33955 & n39929 ) ;
  assign n48466 = n10678 & n11803 ;
  assign n48467 = ~n437 & n39430 ;
  assign n48468 = ~n17376 & n48467 ;
  assign n48469 = ~n27819 & n46083 ;
  assign n48470 = n25416 ^ n9492 ^ 1'b0 ;
  assign n48471 = ( n23215 & ~n32794 ) | ( n23215 & n48470 ) | ( ~n32794 & n48470 ) ;
  assign n48472 = n13840 ^ n11210 ^ n1010 ;
  assign n48473 = n35847 & ~n48472 ;
  assign n48474 = ( ~n1624 & n12462 ) | ( ~n1624 & n39875 ) | ( n12462 & n39875 ) ;
  assign n48475 = n48474 ^ n11564 ^ n6308 ;
  assign n48476 = ( ~n8355 & n32379 ) | ( ~n8355 & n37970 ) | ( n32379 & n37970 ) ;
  assign n48477 = n48476 ^ n46355 ^ n8111 ;
  assign n48478 = ( n8704 & n34489 ) | ( n8704 & ~n48477 ) | ( n34489 & ~n48477 ) ;
  assign n48479 = n14511 | n24423 ;
  assign n48480 = n48479 ^ n8593 ^ 1'b0 ;
  assign n48481 = n48480 ^ n13992 ^ n2069 ;
  assign n48482 = ( ~n23206 & n24852 ) | ( ~n23206 & n30701 ) | ( n24852 & n30701 ) ;
  assign n48483 = ( ~n9516 & n18942 ) | ( ~n9516 & n33682 ) | ( n18942 & n33682 ) ;
  assign n48484 = n6164 | n48483 ;
  assign n48485 = n18582 ^ n12707 ^ n9438 ;
  assign n48486 = n16908 & ~n29523 ;
  assign n48487 = ( n18803 & ~n48485 ) | ( n18803 & n48486 ) | ( ~n48485 & n48486 ) ;
  assign n48488 = n8317 & ~n48487 ;
  assign n48489 = ~n37596 & n48488 ;
  assign n48490 = ( n2925 & n4204 ) | ( n2925 & n5603 ) | ( n4204 & n5603 ) ;
  assign n48492 = ( n1103 & n2049 ) | ( n1103 & n19383 ) | ( n2049 & n19383 ) ;
  assign n48491 = n11854 ^ n7896 ^ n2923 ;
  assign n48493 = n48492 ^ n48491 ^ n27445 ;
  assign n48494 = ( n9366 & ~n48490 ) | ( n9366 & n48493 ) | ( ~n48490 & n48493 ) ;
  assign n48495 = ( n6323 & n7278 ) | ( n6323 & n45431 ) | ( n7278 & n45431 ) ;
  assign n48496 = ( n823 & n6513 ) | ( n823 & n40804 ) | ( n6513 & n40804 ) ;
  assign n48497 = ( n8810 & n17305 ) | ( n8810 & n29418 ) | ( n17305 & n29418 ) ;
  assign n48498 = ( n2106 & n7328 ) | ( n2106 & ~n10525 ) | ( n7328 & ~n10525 ) ;
  assign n48499 = ( n31458 & ~n39995 ) | ( n31458 & n45357 ) | ( ~n39995 & n45357 ) ;
  assign n48500 = n9295 | n13189 ;
  assign n48501 = n2649 & n23780 ;
  assign n48502 = ( n11300 & n34484 ) | ( n11300 & ~n48501 ) | ( n34484 & ~n48501 ) ;
  assign n48503 = n48502 ^ n37532 ^ n36764 ;
  assign n48504 = n45013 ^ n37015 ^ 1'b0 ;
  assign n48505 = ( x27 & ~n16726 ) | ( x27 & n48504 ) | ( ~n16726 & n48504 ) ;
  assign n48506 = n11539 ^ n5170 ^ n2037 ;
  assign n48507 = n48506 ^ n17033 ^ n12335 ;
  assign n48508 = ( ~n3796 & n5447 ) | ( ~n3796 & n34040 ) | ( n5447 & n34040 ) ;
  assign n48509 = n6850 & n48508 ;
  assign n48510 = n38001 ^ n22504 ^ n14059 ;
  assign n48511 = n10269 ^ n5109 ^ 1'b0 ;
  assign n48512 = n4178 ^ n3608 ^ 1'b0 ;
  assign n48513 = ~n7756 & n48512 ;
  assign n48514 = n48513 ^ n22010 ^ n21754 ;
  assign n48517 = ( n1468 & ~n3646 ) | ( n1468 & n43202 ) | ( ~n3646 & n43202 ) ;
  assign n48515 = ( n1983 & n9291 ) | ( n1983 & n23663 ) | ( n9291 & n23663 ) ;
  assign n48516 = n48515 ^ n20246 ^ n11479 ;
  assign n48518 = n48517 ^ n48516 ^ n2359 ;
  assign n48519 = ( n6561 & n24712 ) | ( n6561 & ~n32876 ) | ( n24712 & ~n32876 ) ;
  assign n48520 = n43381 ^ n32917 ^ n29715 ;
  assign n48521 = ( n4177 & ~n9923 ) | ( n4177 & n48520 ) | ( ~n9923 & n48520 ) ;
  assign n48522 = ( n4770 & n13713 ) | ( n4770 & n17789 ) | ( n13713 & n17789 ) ;
  assign n48523 = ( ~n8374 & n9647 ) | ( ~n8374 & n48522 ) | ( n9647 & n48522 ) ;
  assign n48524 = n19873 ^ n9923 ^ 1'b0 ;
  assign n48525 = n48523 & n48524 ;
  assign n48526 = ( n692 & n27351 ) | ( n692 & n48525 ) | ( n27351 & n48525 ) ;
  assign n48527 = ( n48519 & n48521 ) | ( n48519 & ~n48526 ) | ( n48521 & ~n48526 ) ;
  assign n48528 = n48439 ^ n22837 ^ n3216 ;
  assign n48529 = n28672 & ~n30376 ;
  assign n48530 = n28002 ^ n10407 ^ n3799 ;
  assign n48531 = n8635 ^ n2390 ^ 1'b0 ;
  assign n48532 = ( n41188 & n48530 ) | ( n41188 & ~n48531 ) | ( n48530 & ~n48531 ) ;
  assign n48533 = n48532 ^ n14712 ^ n8092 ;
  assign n48534 = n48533 ^ n29255 ^ n4083 ;
  assign n48535 = ( n37950 & n41092 ) | ( n37950 & ~n48534 ) | ( n41092 & ~n48534 ) ;
  assign n48536 = n46524 ^ n31719 ^ n30772 ;
  assign n48537 = ( n14419 & n22814 ) | ( n14419 & ~n34168 ) | ( n22814 & ~n34168 ) ;
  assign n48538 = ( n26553 & n35533 ) | ( n26553 & n48537 ) | ( n35533 & n48537 ) ;
  assign n48539 = n48538 ^ n45140 ^ n9053 ;
  assign n48540 = n44562 ^ n15659 ^ 1'b0 ;
  assign n48541 = n24174 & n48540 ;
  assign n48542 = ( n7383 & n39631 ) | ( n7383 & n46404 ) | ( n39631 & n46404 ) ;
  assign n48543 = ( n3952 & ~n5964 ) | ( n3952 & n32154 ) | ( ~n5964 & n32154 ) ;
  assign n48544 = n48543 ^ n37555 ^ n23747 ;
  assign n48545 = ( n15601 & n30157 ) | ( n15601 & ~n48544 ) | ( n30157 & ~n48544 ) ;
  assign n48546 = ( n46243 & ~n48542 ) | ( n46243 & n48545 ) | ( ~n48542 & n48545 ) ;
  assign n48547 = n34035 ^ n16436 ^ n5155 ;
  assign n48548 = ( n475 & n25231 ) | ( n475 & n36741 ) | ( n25231 & n36741 ) ;
  assign n48549 = n42052 ^ n38231 ^ n19262 ;
  assign n48550 = ( n35957 & n36547 ) | ( n35957 & ~n39003 ) | ( n36547 & ~n39003 ) ;
  assign n48553 = n45120 ^ n26651 ^ n25626 ;
  assign n48554 = x163 | n48553 ;
  assign n48555 = n48554 ^ n46703 ^ n14280 ;
  assign n48551 = ( n2651 & n11430 ) | ( n2651 & n23456 ) | ( n11430 & n23456 ) ;
  assign n48552 = n48551 ^ n31258 ^ n4968 ;
  assign n48556 = n48555 ^ n48552 ^ n6194 ;
  assign n48557 = n22294 ^ n21497 ^ n21095 ;
  assign n48558 = ( n12633 & n25405 ) | ( n12633 & n42100 ) | ( n25405 & n42100 ) ;
  assign n48559 = ~n12605 & n17268 ;
  assign n48560 = n48559 ^ n1321 ^ 1'b0 ;
  assign n48561 = ( n666 & n7551 ) | ( n666 & n11675 ) | ( n7551 & n11675 ) ;
  assign n48562 = ( n12621 & n18471 ) | ( n12621 & ~n48561 ) | ( n18471 & ~n48561 ) ;
  assign n48563 = n48562 ^ n27528 ^ n14839 ;
  assign n48564 = ( ~n3210 & n38110 ) | ( ~n3210 & n48563 ) | ( n38110 & n48563 ) ;
  assign n48565 = ( ~n7649 & n10875 ) | ( ~n7649 & n16119 ) | ( n10875 & n16119 ) ;
  assign n48566 = n48565 ^ n31123 ^ n17732 ;
  assign n48567 = n38337 ^ n8524 ^ 1'b0 ;
  assign n48568 = ( n17056 & ~n30038 ) | ( n17056 & n48567 ) | ( ~n30038 & n48567 ) ;
  assign n48569 = n48568 ^ n44412 ^ n39969 ;
  assign n48570 = n12061 | n17539 ;
  assign n48575 = ~n2453 & n17211 ;
  assign n48576 = n48575 ^ n16974 ^ 1'b0 ;
  assign n48573 = n3587 | n9782 ;
  assign n48574 = n48573 ^ n33336 ^ 1'b0 ;
  assign n48577 = n48576 ^ n48574 ^ n8285 ;
  assign n48578 = ( ~n37860 & n44737 ) | ( ~n37860 & n48577 ) | ( n44737 & n48577 ) ;
  assign n48571 = n38028 ^ n24409 ^ n6732 ;
  assign n48572 = n48571 ^ n42714 ^ n4001 ;
  assign n48579 = n48578 ^ n48572 ^ n29677 ;
  assign n48580 = n7387 ^ n6826 ^ 1'b0 ;
  assign n48581 = n19471 & n48580 ;
  assign n48582 = ( n2478 & n41844 ) | ( n2478 & ~n48581 ) | ( n41844 & ~n48581 ) ;
  assign n48583 = n48582 ^ n14074 ^ n1733 ;
  assign n48584 = ( n10873 & n37189 ) | ( n10873 & ~n44786 ) | ( n37189 & ~n44786 ) ;
  assign n48586 = n26186 ^ n25820 ^ n23358 ;
  assign n48585 = n46953 ^ n16899 ^ n5370 ;
  assign n48587 = n48586 ^ n48585 ^ n23304 ;
  assign n48588 = n11311 | n27292 ;
  assign n48589 = n48588 ^ n13498 ^ 1'b0 ;
  assign n48590 = n48589 ^ n16340 ^ 1'b0 ;
  assign n48591 = n48587 & ~n48590 ;
  assign n48593 = n6332 | n31745 ;
  assign n48594 = n8986 & ~n48593 ;
  assign n48592 = n40134 ^ n36038 ^ n21894 ;
  assign n48595 = n48594 ^ n48592 ^ n3524 ;
  assign n48596 = ( n1836 & n26477 ) | ( n1836 & n41509 ) | ( n26477 & n41509 ) ;
  assign n48597 = ( ~n8721 & n32066 ) | ( ~n8721 & n44983 ) | ( n32066 & n44983 ) ;
  assign n48598 = ( n18235 & n48596 ) | ( n18235 & n48597 ) | ( n48596 & n48597 ) ;
  assign n48599 = n20724 ^ n11406 ^ 1'b0 ;
  assign n48600 = n47695 ^ n33329 ^ 1'b0 ;
  assign n48601 = ( ~n1595 & n15808 ) | ( ~n1595 & n24771 ) | ( n15808 & n24771 ) ;
  assign n48602 = n5340 ^ n1295 ^ n1218 ;
  assign n48603 = n32638 & ~n48602 ;
  assign n48604 = ~n5522 & n48603 ;
  assign n48605 = n48604 ^ n31650 ^ n3804 ;
  assign n48606 = n25320 ^ n16289 ^ n9925 ;
  assign n48607 = ( n6276 & ~n13322 ) | ( n6276 & n48606 ) | ( ~n13322 & n48606 ) ;
  assign n48608 = n45702 ^ n36687 ^ n17565 ;
  assign n48609 = n15837 ^ n6211 ^ 1'b0 ;
  assign n48610 = n11560 & ~n48609 ;
  assign n48611 = ( ~n3154 & n7395 ) | ( ~n3154 & n17000 ) | ( n7395 & n17000 ) ;
  assign n48612 = ( n6849 & n46219 ) | ( n6849 & n48611 ) | ( n46219 & n48611 ) ;
  assign n48613 = ( n23482 & ~n25110 ) | ( n23482 & n46316 ) | ( ~n25110 & n46316 ) ;
  assign n48614 = ( ~n9292 & n18642 ) | ( ~n9292 & n19300 ) | ( n18642 & n19300 ) ;
  assign n48615 = n48614 ^ n26742 ^ n26717 ;
  assign n48616 = ( n7059 & n9377 ) | ( n7059 & n13742 ) | ( n9377 & n13742 ) ;
  assign n48617 = n15906 ^ n15171 ^ n3932 ;
  assign n48618 = n6469 & n23030 ;
  assign n48619 = n48618 ^ n26827 ^ n10071 ;
  assign n48620 = n37523 ^ n27175 ^ n11679 ;
  assign n48621 = ( n2529 & ~n39541 ) | ( n2529 & n48620 ) | ( ~n39541 & n48620 ) ;
  assign n48622 = n2124 & ~n8793 ;
  assign n48623 = ( n14366 & n21828 ) | ( n14366 & ~n25532 ) | ( n21828 & ~n25532 ) ;
  assign n48624 = n48623 ^ n27463 ^ n19925 ;
  assign n48625 = ~n7020 & n10932 ;
  assign n48626 = n48625 ^ n38986 ^ n23899 ;
  assign n48627 = n14764 ^ n14519 ^ n753 ;
  assign n48628 = ( n1094 & n30406 ) | ( n1094 & n43657 ) | ( n30406 & n43657 ) ;
  assign n48629 = ( ~n31084 & n32978 ) | ( ~n31084 & n48628 ) | ( n32978 & n48628 ) ;
  assign n48630 = n42625 ^ n16802 ^ n14652 ;
  assign n48631 = x223 | n31378 ;
  assign n48632 = n48631 ^ n11556 ^ n504 ;
  assign n48633 = n23124 ^ n12483 ^ n1971 ;
  assign n48634 = n28953 ^ n19867 ^ n12446 ;
  assign n48635 = n48634 ^ n10784 ^ n5344 ;
  assign n48636 = ( ~n5178 & n23846 ) | ( ~n5178 & n40751 ) | ( n23846 & n40751 ) ;
  assign n48637 = ( n3221 & n48635 ) | ( n3221 & ~n48636 ) | ( n48635 & ~n48636 ) ;
  assign n48638 = ( n32571 & ~n48633 ) | ( n32571 & n48637 ) | ( ~n48633 & n48637 ) ;
  assign n48639 = n38771 ^ n11214 ^ n10718 ;
  assign n48640 = ( n14014 & ~n27679 ) | ( n14014 & n39215 ) | ( ~n27679 & n39215 ) ;
  assign n48641 = n48640 ^ n22433 ^ n15068 ;
  assign n48643 = ( n11835 & ~n12202 ) | ( n11835 & n18351 ) | ( ~n12202 & n18351 ) ;
  assign n48644 = n48643 ^ n40940 ^ n36831 ;
  assign n48642 = n46172 ^ n24082 ^ n9503 ;
  assign n48645 = n48644 ^ n48642 ^ n38275 ;
  assign n48646 = n41454 ^ n6912 ^ n3789 ;
  assign n48647 = n7449 | n33157 ;
  assign n48648 = n48647 ^ n23101 ^ n23010 ;
  assign n48649 = n18783 | n19238 ;
  assign n48650 = n10403 | n48649 ;
  assign n48651 = n48650 ^ n43712 ^ n41113 ;
  assign n48652 = n24951 ^ n9522 ^ n8191 ;
  assign n48653 = ( n6435 & n9175 ) | ( n6435 & n48652 ) | ( n9175 & n48652 ) ;
  assign n48654 = n42333 ^ n24694 ^ n13430 ;
  assign n48655 = n48654 ^ n2426 ^ 1'b0 ;
  assign n48656 = ( n19919 & n24050 ) | ( n19919 & n48655 ) | ( n24050 & n48655 ) ;
  assign n48657 = n38352 & n48656 ;
  assign n48658 = ~n43514 & n48657 ;
  assign n48659 = ( n818 & n4807 ) | ( n818 & ~n6560 ) | ( n4807 & ~n6560 ) ;
  assign n48660 = ( n9956 & n15064 ) | ( n9956 & ~n48659 ) | ( n15064 & ~n48659 ) ;
  assign n48661 = n16606 | n47872 ;
  assign n48662 = n48661 ^ n31120 ^ 1'b0 ;
  assign n48665 = n29434 ^ n3237 ^ 1'b0 ;
  assign n48663 = n38227 ^ n14843 ^ x129 ;
  assign n48664 = ( n11510 & n12064 ) | ( n11510 & ~n48663 ) | ( n12064 & ~n48663 ) ;
  assign n48666 = n48665 ^ n48664 ^ n25228 ;
  assign n48667 = n16103 ^ n7849 ^ n738 ;
  assign n48668 = n39418 ^ n18910 ^ n14365 ;
  assign n48669 = ( n16097 & n48667 ) | ( n16097 & n48668 ) | ( n48667 & n48668 ) ;
  assign n48670 = n48669 ^ n34075 ^ 1'b0 ;
  assign n48671 = n48666 | n48670 ;
  assign n48672 = n19086 ^ n5151 ^ 1'b0 ;
  assign n48673 = n5379 | n48672 ;
  assign n48674 = n46860 ^ n37342 ^ n30315 ;
  assign n48675 = ( n17498 & ~n48673 ) | ( n17498 & n48674 ) | ( ~n48673 & n48674 ) ;
  assign n48676 = n28176 ^ n12732 ^ n7767 ;
  assign n48677 = ( n18462 & n21341 ) | ( n18462 & ~n22324 ) | ( n21341 & ~n22324 ) ;
  assign n48678 = n48677 ^ n30001 ^ n4092 ;
  assign n48679 = n48678 ^ n19104 ^ n16043 ;
  assign n48680 = ( n1830 & n4647 ) | ( n1830 & n10917 ) | ( n4647 & n10917 ) ;
  assign n48681 = ( n15117 & n25696 ) | ( n15117 & n48680 ) | ( n25696 & n48680 ) ;
  assign n48682 = n8894 ^ n6710 ^ n498 ;
  assign n48683 = ( n10658 & n22992 ) | ( n10658 & ~n48682 ) | ( n22992 & ~n48682 ) ;
  assign n48684 = n48683 ^ n45664 ^ n42590 ;
  assign n48685 = n37293 | n40734 ;
  assign n48686 = n23395 | n48685 ;
  assign n48687 = ( n37780 & ~n39706 ) | ( n37780 & n48686 ) | ( ~n39706 & n48686 ) ;
  assign n48688 = n42258 ^ n13040 ^ n5556 ;
  assign n48689 = n48688 ^ n31872 ^ n25461 ;
  assign n48690 = n23226 & n35747 ;
  assign n48691 = ~n19487 & n48690 ;
  assign n48692 = n25672 ^ n21131 ^ 1'b0 ;
  assign n48693 = n48691 | n48692 ;
  assign n48694 = ( n1960 & n7839 ) | ( n1960 & n42717 ) | ( n7839 & n42717 ) ;
  assign n48695 = n3209 & ~n48694 ;
  assign n48696 = ~n2038 & n48695 ;
  assign n48697 = ( n4285 & n30378 ) | ( n4285 & n35454 ) | ( n30378 & n35454 ) ;
  assign n48701 = ( n4418 & n8667 ) | ( n4418 & ~n27592 ) | ( n8667 & ~n27592 ) ;
  assign n48700 = n3554 | n5680 ;
  assign n48698 = ~n4307 & n40002 ;
  assign n48699 = n48698 ^ n48520 ^ 1'b0 ;
  assign n48702 = n48701 ^ n48700 ^ n48699 ;
  assign n48703 = n33113 ^ n10892 ^ 1'b0 ;
  assign n48704 = n37671 ^ n29251 ^ n759 ;
  assign n48705 = ( n11982 & n43103 ) | ( n11982 & ~n48704 ) | ( n43103 & ~n48704 ) ;
  assign n48706 = n48705 ^ n16248 ^ 1'b0 ;
  assign n48707 = n27064 ^ n24860 ^ n7869 ;
  assign n48708 = n7786 ^ n7066 ^ n2528 ;
  assign n48709 = n48708 ^ n31085 ^ n1524 ;
  assign n48710 = n48709 ^ n45178 ^ n42920 ;
  assign n48711 = ( ~n21377 & n33967 ) | ( ~n21377 & n38853 ) | ( n33967 & n38853 ) ;
  assign n48712 = n8834 | n28318 ;
  assign n48713 = n48712 ^ n22712 ^ 1'b0 ;
  assign n48714 = n15700 & n48713 ;
  assign n48715 = n48714 ^ n16888 ^ n11606 ;
  assign n48716 = n20017 & ~n47643 ;
  assign n48717 = n48716 ^ n20437 ^ 1'b0 ;
  assign n48718 = ~n6273 & n17101 ;
  assign n48719 = n48718 ^ n32666 ^ 1'b0 ;
  assign n48720 = n7236 & ~n24536 ;
  assign n48721 = n48720 ^ n21411 ^ 1'b0 ;
  assign n48722 = n16884 ^ n11007 ^ 1'b0 ;
  assign n48723 = n48722 ^ n41822 ^ n30111 ;
  assign n48724 = ( n16522 & n48721 ) | ( n16522 & n48723 ) | ( n48721 & n48723 ) ;
  assign n48725 = ( n1763 & ~n9414 ) | ( n1763 & n48724 ) | ( ~n9414 & n48724 ) ;
  assign n48729 = ( ~n556 & n10615 ) | ( ~n556 & n13788 ) | ( n10615 & n13788 ) ;
  assign n48727 = ( ~n6017 & n11339 ) | ( ~n6017 & n20001 ) | ( n11339 & n20001 ) ;
  assign n48728 = n48727 ^ n23686 ^ n647 ;
  assign n48726 = n39426 ^ n28867 ^ n13559 ;
  assign n48730 = n48729 ^ n48728 ^ n48726 ;
  assign n48731 = n33341 ^ n29119 ^ n20013 ;
  assign n48732 = n27311 ^ n15927 ^ n9932 ;
  assign n48733 = n44101 ^ n30826 ^ n12682 ;
  assign n48734 = n48733 ^ n5464 ^ n4499 ;
  assign n48735 = n22233 ^ n20141 ^ n15265 ;
  assign n48737 = ( n2249 & n11063 ) | ( n2249 & ~n15723 ) | ( n11063 & ~n15723 ) ;
  assign n48736 = ( n2795 & ~n11499 ) | ( n2795 & n38460 ) | ( ~n11499 & n38460 ) ;
  assign n48738 = n48737 ^ n48736 ^ n3162 ;
  assign n48743 = n30158 ^ n23137 ^ n14919 ;
  assign n48739 = n28211 ^ n8058 ^ n7024 ;
  assign n48740 = ( ~n25457 & n29582 ) | ( ~n25457 & n48739 ) | ( n29582 & n48739 ) ;
  assign n48741 = n48740 ^ n42954 ^ n30699 ;
  assign n48742 = ( n1584 & ~n36917 ) | ( n1584 & n48741 ) | ( ~n36917 & n48741 ) ;
  assign n48744 = n48743 ^ n48742 ^ n10819 ;
  assign n48745 = n35868 | n36924 ;
  assign n48746 = ~n16672 & n40082 ;
  assign n48747 = ~n13750 & n48746 ;
  assign n48748 = n43198 ^ n28251 ^ n18952 ;
  assign n48749 = n12366 & ~n35010 ;
  assign n48750 = n16826 ^ n5865 ^ n1564 ;
  assign n48752 = ( ~n3927 & n12369 ) | ( ~n3927 & n13848 ) | ( n12369 & n13848 ) ;
  assign n48751 = n13607 ^ n7337 ^ n1656 ;
  assign n48753 = n48752 ^ n48751 ^ n9407 ;
  assign n48754 = ( n1549 & n48750 ) | ( n1549 & n48753 ) | ( n48750 & n48753 ) ;
  assign n48755 = n9329 ^ n8924 ^ n380 ;
  assign n48756 = n48755 ^ n4840 ^ n850 ;
  assign n48757 = n48756 ^ n27606 ^ n11043 ;
  assign n48758 = n32269 ^ n23840 ^ n16102 ;
  assign n48759 = ( n7893 & ~n46264 ) | ( n7893 & n48758 ) | ( ~n46264 & n48758 ) ;
  assign n48760 = n48759 ^ n48040 ^ n16732 ;
  assign n48761 = ~n39012 & n46659 ;
  assign n48762 = n48761 ^ n30810 ^ 1'b0 ;
  assign n48763 = n48762 ^ n39226 ^ n35906 ;
  assign n48764 = n33653 & n38966 ;
  assign n48765 = n19358 & n48764 ;
  assign n48766 = ( n7486 & n24276 ) | ( n7486 & n30327 ) | ( n24276 & n30327 ) ;
  assign n48767 = ( n8284 & n48413 ) | ( n8284 & ~n48766 ) | ( n48413 & ~n48766 ) ;
  assign n48768 = ( n550 & n2912 ) | ( n550 & n9088 ) | ( n2912 & n9088 ) ;
  assign n48769 = n48768 ^ n44786 ^ n8412 ;
  assign n48770 = ( n24955 & n26688 ) | ( n24955 & n30707 ) | ( n26688 & n30707 ) ;
  assign n48771 = ( n39169 & ~n48769 ) | ( n39169 & n48770 ) | ( ~n48769 & n48770 ) ;
  assign n48773 = n40358 ^ n19282 ^ n15521 ;
  assign n48774 = n48773 ^ n25232 ^ n22559 ;
  assign n48772 = n29866 ^ n21353 ^ n12969 ;
  assign n48775 = n48774 ^ n48772 ^ n10275 ;
  assign n48776 = n41204 ^ n27853 ^ n9915 ;
  assign n48777 = ( ~n2262 & n3061 ) | ( ~n2262 & n33502 ) | ( n3061 & n33502 ) ;
  assign n48778 = ~n18157 & n48777 ;
  assign n48779 = n40513 & n48778 ;
  assign n48780 = n30771 ^ n30678 ^ n15162 ;
  assign n48781 = ( n27470 & n48779 ) | ( n27470 & ~n48780 ) | ( n48779 & ~n48780 ) ;
  assign n48782 = ( ~n13972 & n42616 ) | ( ~n13972 & n48781 ) | ( n42616 & n48781 ) ;
  assign n48783 = ( n2991 & ~n12110 ) | ( n2991 & n23831 ) | ( ~n12110 & n23831 ) ;
  assign n48784 = n48783 ^ n27448 ^ n4939 ;
  assign n48785 = n42715 ^ n41276 ^ n37218 ;
  assign n48786 = ( ~n46261 & n48784 ) | ( ~n46261 & n48785 ) | ( n48784 & n48785 ) ;
  assign n48787 = n23933 ^ n22320 ^ n15295 ;
  assign n48788 = ( n3495 & n41507 ) | ( n3495 & n48787 ) | ( n41507 & n48787 ) ;
  assign n48789 = n48788 ^ n20148 ^ n12306 ;
  assign n48790 = n21220 ^ n20325 ^ n7321 ;
  assign n48791 = n48790 ^ n24323 ^ n20928 ;
  assign n48792 = ( n8434 & ~n14657 ) | ( n8434 & n37606 ) | ( ~n14657 & n37606 ) ;
  assign n48793 = n8256 | n43019 ;
  assign n48794 = n48793 ^ n13531 ^ 1'b0 ;
  assign n48795 = n10122 & ~n11254 ;
  assign n48796 = n43096 & n48795 ;
  assign n48799 = ( n1117 & n12091 ) | ( n1117 & n36959 ) | ( n12091 & n36959 ) ;
  assign n48797 = n3473 & ~n40218 ;
  assign n48798 = n48797 ^ n25233 ^ 1'b0 ;
  assign n48800 = n48799 ^ n48798 ^ n21777 ;
  assign n48801 = ( n12126 & n25223 ) | ( n12126 & ~n48030 ) | ( n25223 & ~n48030 ) ;
  assign n48802 = n32270 ^ n23355 ^ n14004 ;
  assign n48803 = n43900 ^ n29662 ^ n19119 ;
  assign n48805 = n34997 ^ n10679 ^ n4068 ;
  assign n48804 = n7649 ^ n602 ^ 1'b0 ;
  assign n48806 = n48805 ^ n48804 ^ n33761 ;
  assign n48807 = ( n2534 & n7944 ) | ( n2534 & n45941 ) | ( n7944 & n45941 ) ;
  assign n48809 = ( n7475 & n30597 ) | ( n7475 & ~n37475 ) | ( n30597 & ~n37475 ) ;
  assign n48808 = n42261 ^ n39703 ^ n27317 ;
  assign n48810 = n48809 ^ n48808 ^ n33795 ;
  assign n48811 = n46688 ^ n43014 ^ n3285 ;
  assign n48812 = ( n23279 & n33825 ) | ( n23279 & ~n40794 ) | ( n33825 & ~n40794 ) ;
  assign n48813 = n48812 ^ n27446 ^ 1'b0 ;
  assign n48814 = n4096 & ~n48813 ;
  assign n48815 = ( n20710 & n34421 ) | ( n20710 & ~n48814 ) | ( n34421 & ~n48814 ) ;
  assign n48816 = n23828 ^ n6440 ^ 1'b0 ;
  assign n48817 = n46642 | n48816 ;
  assign n48819 = n28718 ^ n11097 ^ n8107 ;
  assign n48818 = ~n5141 & n17748 ;
  assign n48820 = n48819 ^ n48818 ^ 1'b0 ;
  assign n48821 = n18801 ^ n10669 ^ n2424 ;
  assign n48823 = n45509 | n45877 ;
  assign n48822 = n27240 | n37352 ;
  assign n48824 = n48823 ^ n48822 ^ 1'b0 ;
  assign n48825 = n48821 | n48824 ;
  assign n48826 = n27357 ^ n14174 ^ n13093 ;
  assign n48827 = n34972 ^ n19919 ^ n10809 ;
  assign n48828 = n48827 ^ n42086 ^ n28323 ;
  assign n48829 = ( n5136 & n48826 ) | ( n5136 & n48828 ) | ( n48826 & n48828 ) ;
  assign n48830 = n28444 ^ n13813 ^ 1'b0 ;
  assign n48831 = n39109 & ~n48830 ;
  assign n48832 = n48831 ^ n14518 ^ n3976 ;
  assign n48833 = n20108 ^ n16937 ^ n12418 ;
  assign n48834 = ( n9928 & n16702 ) | ( n9928 & ~n48833 ) | ( n16702 & ~n48833 ) ;
  assign n48835 = n48834 ^ n30259 ^ n28315 ;
  assign n48836 = n29385 ^ n23418 ^ n13981 ;
  assign n48837 = n21548 ^ n8194 ^ n7672 ;
  assign n48838 = n43191 ^ n33873 ^ n21645 ;
  assign n48839 = ( ~n7443 & n48837 ) | ( ~n7443 & n48838 ) | ( n48837 & n48838 ) ;
  assign n48840 = n48839 ^ n16215 ^ n9560 ;
  assign n48841 = n9826 ^ n5303 ^ n4172 ;
  assign n48842 = n14257 ^ n13437 ^ n9503 ;
  assign n48843 = n12460 ^ n7363 ^ 1'b0 ;
  assign n48844 = n5384 | n48843 ;
  assign n48845 = n11291 ^ n10165 ^ n2246 ;
  assign n48846 = n30362 ^ n5319 ^ n3012 ;
  assign n48847 = n48846 ^ n34107 ^ n9106 ;
  assign n48848 = n48847 ^ n13251 ^ n1683 ;
  assign n48849 = n9815 ^ n6383 ^ n2458 ;
  assign n48850 = ( n3452 & ~n20308 ) | ( n3452 & n48849 ) | ( ~n20308 & n48849 ) ;
  assign n48851 = n48848 & n48850 ;
  assign n48852 = ( ~n23952 & n48845 ) | ( ~n23952 & n48851 ) | ( n48845 & n48851 ) ;
  assign n48853 = n48852 ^ n32271 ^ n4917 ;
  assign n48854 = ( n19546 & n23795 ) | ( n19546 & ~n45933 ) | ( n23795 & ~n45933 ) ;
  assign n48858 = n338 & n48122 ;
  assign n48859 = n48858 ^ n31466 ^ 1'b0 ;
  assign n48855 = n7193 ^ n4811 ^ 1'b0 ;
  assign n48856 = n48855 ^ n34896 ^ 1'b0 ;
  assign n48857 = n48856 ^ n42069 ^ n9907 ;
  assign n48860 = n48859 ^ n48857 ^ n32361 ;
  assign n48861 = ( n12548 & n16015 ) | ( n12548 & n45051 ) | ( n16015 & n45051 ) ;
  assign n48862 = ( n16736 & n35420 ) | ( n16736 & n39871 ) | ( n35420 & n39871 ) ;
  assign n48863 = n48862 ^ n9258 ^ 1'b0 ;
  assign n48864 = ( n7022 & n46451 ) | ( n7022 & n48863 ) | ( n46451 & n48863 ) ;
  assign n48865 = ( ~n4390 & n36829 ) | ( ~n4390 & n39075 ) | ( n36829 & n39075 ) ;
  assign n48866 = n48865 ^ n39829 ^ n30506 ;
  assign n48867 = ( ~n4013 & n23998 ) | ( ~n4013 & n30618 ) | ( n23998 & n30618 ) ;
  assign n48868 = ( ~x117 & n9392 ) | ( ~x117 & n27909 ) | ( n9392 & n27909 ) ;
  assign n48870 = ( n4941 & n7771 ) | ( n4941 & ~n22098 ) | ( n7771 & ~n22098 ) ;
  assign n48869 = n33987 ^ n31587 ^ n7540 ;
  assign n48871 = n48870 ^ n48869 ^ n46561 ;
  assign n48872 = n14507 ^ n12145 ^ 1'b0 ;
  assign n48873 = ~n48871 & n48872 ;
  assign n48874 = n3392 & ~n13715 ;
  assign n48875 = ~n29125 & n48874 ;
  assign n48876 = n48875 ^ n6643 ^ 1'b0 ;
  assign n48877 = ( n3927 & n5897 ) | ( n3927 & ~n24374 ) | ( n5897 & ~n24374 ) ;
  assign n48878 = ( n809 & n2063 ) | ( n809 & n40747 ) | ( n2063 & n40747 ) ;
  assign n48879 = n44457 ^ n27558 ^ n5007 ;
  assign n48880 = n41208 ^ n23226 ^ n3012 ;
  assign n48881 = n25512 ^ n3541 ^ 1'b0 ;
  assign n48882 = n20280 & ~n48881 ;
  assign n48883 = n48882 ^ n25410 ^ n12850 ;
  assign n48884 = ( n48879 & n48880 ) | ( n48879 & ~n48883 ) | ( n48880 & ~n48883 ) ;
  assign n48885 = n24540 ^ n11578 ^ n6847 ;
  assign n48886 = n48885 ^ n21261 ^ n14611 ;
  assign n48887 = n48886 ^ n21641 ^ n3205 ;
  assign n48888 = ( n3730 & ~n44962 ) | ( n3730 & n48887 ) | ( ~n44962 & n48887 ) ;
  assign n48889 = n11526 ^ n3229 ^ 1'b0 ;
  assign n48890 = n2084 & ~n48889 ;
  assign n48896 = n29221 ^ n12803 ^ n9510 ;
  assign n48894 = ( ~n9092 & n12210 ) | ( ~n9092 & n13390 ) | ( n12210 & n13390 ) ;
  assign n48892 = ( n3405 & n8826 ) | ( n3405 & ~n18307 ) | ( n8826 & ~n18307 ) ;
  assign n48891 = n27852 ^ n25161 ^ 1'b0 ;
  assign n48893 = n48892 ^ n48891 ^ n1599 ;
  assign n48895 = n48894 ^ n48893 ^ n9238 ;
  assign n48897 = n48896 ^ n48895 ^ n6320 ;
  assign n48898 = ( ~n23955 & n37175 ) | ( ~n23955 & n39306 ) | ( n37175 & n39306 ) ;
  assign n48899 = ( n11256 & n11358 ) | ( n11256 & ~n19007 ) | ( n11358 & ~n19007 ) ;
  assign n48900 = ( ~n842 & n22445 ) | ( ~n842 & n48899 ) | ( n22445 & n48899 ) ;
  assign n48901 = ( n5530 & n17724 ) | ( n5530 & n19100 ) | ( n17724 & n19100 ) ;
  assign n48902 = n48901 ^ n10461 ^ 1'b0 ;
  assign n48903 = n40795 & n48902 ;
  assign n48904 = n37246 ^ n16730 ^ n4242 ;
  assign n48905 = n48904 ^ n42312 ^ n933 ;
  assign n48906 = x210 & ~n18239 ;
  assign n48907 = ( ~n302 & n1223 ) | ( ~n302 & n16926 ) | ( n1223 & n16926 ) ;
  assign n48908 = n48907 ^ n41496 ^ n14579 ;
  assign n48909 = n48908 ^ n40384 ^ 1'b0 ;
  assign n48913 = n46743 ^ n7186 ^ n5219 ;
  assign n48914 = n48913 ^ n24119 ^ n7288 ;
  assign n48910 = ( ~n14068 & n16812 ) | ( ~n14068 & n31892 ) | ( n16812 & n31892 ) ;
  assign n48911 = ( n1402 & n20136 ) | ( n1402 & ~n48910 ) | ( n20136 & ~n48910 ) ;
  assign n48912 = ( ~n23449 & n23998 ) | ( ~n23449 & n48911 ) | ( n23998 & n48911 ) ;
  assign n48915 = n48914 ^ n48912 ^ n30475 ;
  assign n48916 = ( x17 & n35075 ) | ( x17 & n48915 ) | ( n35075 & n48915 ) ;
  assign n48917 = ( n2977 & n14931 ) | ( n2977 & ~n48916 ) | ( n14931 & ~n48916 ) ;
  assign n48918 = ( n2349 & n9324 ) | ( n2349 & n24030 ) | ( n9324 & n24030 ) ;
  assign n48919 = n4326 ^ x182 ^ 1'b0 ;
  assign n48920 = ~n48918 & n48919 ;
  assign n48921 = ( n4500 & ~n17209 ) | ( n4500 & n37431 ) | ( ~n17209 & n37431 ) ;
  assign n48922 = n26102 & n48921 ;
  assign n48923 = n2916 | n48922 ;
  assign n48924 = n48923 ^ n26880 ^ 1'b0 ;
  assign n48925 = ( n1292 & n1299 ) | ( n1292 & ~n24837 ) | ( n1299 & ~n24837 ) ;
  assign n48926 = ( n15334 & n37653 ) | ( n15334 & n48925 ) | ( n37653 & n48925 ) ;
  assign n48927 = n48926 ^ n19954 ^ n4863 ;
  assign n48928 = n33621 ^ n24647 ^ n4882 ;
  assign n48929 = ( n15195 & n16941 ) | ( n15195 & ~n36579 ) | ( n16941 & ~n36579 ) ;
  assign n48930 = n32240 ^ n26053 ^ n9183 ;
  assign n48931 = ( n1373 & ~n48929 ) | ( n1373 & n48930 ) | ( ~n48929 & n48930 ) ;
  assign n48932 = n41766 ^ n27679 ^ n19000 ;
  assign n48933 = n19265 ^ n17108 ^ n3293 ;
  assign n48934 = ( n10937 & n48932 ) | ( n10937 & ~n48933 ) | ( n48932 & ~n48933 ) ;
  assign n48935 = ( n2305 & ~n14374 ) | ( n2305 & n19525 ) | ( ~n14374 & n19525 ) ;
  assign n48936 = n48935 ^ n4191 ^ 1'b0 ;
  assign n48937 = n4801 & ~n42403 ;
  assign n48938 = n36896 ^ n26611 ^ n25277 ;
  assign n48939 = n9601 & ~n42590 ;
  assign n48940 = ~n10870 & n48939 ;
  assign n48941 = ( n25384 & n48938 ) | ( n25384 & n48940 ) | ( n48938 & n48940 ) ;
  assign n48942 = n38425 ^ n8892 ^ 1'b0 ;
  assign n48943 = n3785 | n30258 ;
  assign n48944 = ( n4943 & ~n9953 ) | ( n4943 & n48943 ) | ( ~n9953 & n48943 ) ;
  assign n48946 = n27492 ^ n19388 ^ n8817 ;
  assign n48945 = n4703 | n25205 ;
  assign n48947 = n48946 ^ n48945 ^ 1'b0 ;
  assign n48948 = ( n6009 & n23385 ) | ( n6009 & n33894 ) | ( n23385 & n33894 ) ;
  assign n48949 = ( n17123 & ~n20484 ) | ( n17123 & n48948 ) | ( ~n20484 & n48948 ) ;
  assign n48950 = n14288 ^ n7854 ^ n5098 ;
  assign n48951 = n12002 & ~n48950 ;
  assign n48952 = ~n20505 & n48951 ;
  assign n48953 = ( ~n6904 & n10473 ) | ( ~n6904 & n48952 ) | ( n10473 & n48952 ) ;
  assign n48954 = ( n16002 & ~n33698 ) | ( n16002 & n48953 ) | ( ~n33698 & n48953 ) ;
  assign n48955 = ( ~n14195 & n24651 ) | ( ~n14195 & n27713 ) | ( n24651 & n27713 ) ;
  assign n48956 = n48955 ^ n2781 ^ 1'b0 ;
  assign n48957 = ( ~n23291 & n40747 ) | ( ~n23291 & n48956 ) | ( n40747 & n48956 ) ;
  assign n48958 = ( n4154 & ~n26190 ) | ( n4154 & n48957 ) | ( ~n26190 & n48957 ) ;
  assign n48959 = ( n34768 & n45078 ) | ( n34768 & ~n48958 ) | ( n45078 & ~n48958 ) ;
  assign n48960 = ( n19757 & n30009 ) | ( n19757 & ~n37611 ) | ( n30009 & ~n37611 ) ;
  assign n48961 = n41211 ^ n20458 ^ n4876 ;
  assign n48962 = ( n27351 & ~n33626 ) | ( n27351 & n37135 ) | ( ~n33626 & n37135 ) ;
  assign n48963 = ( n5603 & n26881 ) | ( n5603 & n48962 ) | ( n26881 & n48962 ) ;
  assign n48964 = ~n2211 & n11217 ;
  assign n48965 = n48964 ^ n9479 ^ 1'b0 ;
  assign n48966 = ( ~n13587 & n14201 ) | ( ~n13587 & n48965 ) | ( n14201 & n48965 ) ;
  assign n48967 = n38686 ^ n15328 ^ n5066 ;
  assign n48968 = n39425 ^ n26536 ^ n16753 ;
  assign n48969 = n48968 ^ n20996 ^ x40 ;
  assign n48970 = n47032 ^ n9661 ^ 1'b0 ;
  assign n48971 = n2110 & n48970 ;
  assign n48972 = n35052 ^ n34745 ^ n16139 ;
  assign n48973 = n40384 ^ n18456 ^ n16801 ;
  assign n48974 = ( n23329 & n27861 ) | ( n23329 & n28808 ) | ( n27861 & n28808 ) ;
  assign n48975 = n48974 ^ n38927 ^ 1'b0 ;
  assign n48976 = ~n37087 & n48975 ;
  assign n48977 = n48976 ^ n1171 ^ 1'b0 ;
  assign n48979 = ( ~n3219 & n21432 ) | ( ~n3219 & n28490 ) | ( n21432 & n28490 ) ;
  assign n48978 = n19741 ^ n6078 ^ n4082 ;
  assign n48980 = n48979 ^ n48978 ^ n8934 ;
  assign n48981 = ( ~n13865 & n37560 ) | ( ~n13865 & n41577 ) | ( n37560 & n41577 ) ;
  assign n48982 = ( n30292 & n32722 ) | ( n30292 & n48981 ) | ( n32722 & n48981 ) ;
  assign n48983 = ( x248 & n9707 ) | ( x248 & n25611 ) | ( n9707 & n25611 ) ;
  assign n48984 = n11948 ^ n7544 ^ 1'b0 ;
  assign n48985 = ( n10617 & n14734 ) | ( n10617 & ~n48984 ) | ( n14734 & ~n48984 ) ;
  assign n48986 = n28201 ^ n22032 ^ n17678 ;
  assign n48987 = ( n48983 & ~n48985 ) | ( n48983 & n48986 ) | ( ~n48985 & n48986 ) ;
  assign n48988 = n5441 | n44691 ;
  assign n48989 = n48988 ^ n9521 ^ 1'b0 ;
  assign n48990 = ( n9496 & n18527 ) | ( n9496 & ~n35554 ) | ( n18527 & ~n35554 ) ;
  assign n48991 = n14428 ^ n1211 ^ 1'b0 ;
  assign n48992 = n39819 ^ n23882 ^ n4189 ;
  assign n48993 = n8124 & ~n9839 ;
  assign n48994 = ~n5675 & n48993 ;
  assign n48995 = ( n10341 & n26575 ) | ( n10341 & ~n48994 ) | ( n26575 & ~n48994 ) ;
  assign n48996 = ( n22876 & ~n48992 ) | ( n22876 & n48995 ) | ( ~n48992 & n48995 ) ;
  assign n48997 = ( n4611 & n35573 ) | ( n4611 & n36546 ) | ( n35573 & n36546 ) ;
  assign n48998 = ( n6018 & n11816 ) | ( n6018 & n15261 ) | ( n11816 & n15261 ) ;
  assign n48999 = n27904 ^ n23617 ^ n8908 ;
  assign n49000 = n6109 & ~n24682 ;
  assign n49001 = ~n48999 & n49000 ;
  assign n49002 = ( n11720 & n48998 ) | ( n11720 & n49001 ) | ( n48998 & n49001 ) ;
  assign n49003 = ( n3724 & ~n8386 ) | ( n3724 & n19700 ) | ( ~n8386 & n19700 ) ;
  assign n49004 = n49003 ^ n41164 ^ n24895 ;
  assign n49005 = n19982 ^ n5178 ^ x155 ;
  assign n49006 = ( ~n39717 & n44425 ) | ( ~n39717 & n49005 ) | ( n44425 & n49005 ) ;
  assign n49007 = n33334 ^ n20669 ^ 1'b0 ;
  assign n49008 = n22887 & ~n49007 ;
  assign n49009 = ( n5401 & n42799 ) | ( n5401 & ~n49008 ) | ( n42799 & ~n49008 ) ;
  assign n49010 = n4318 & ~n7714 ;
  assign n49011 = n49009 & n49010 ;
  assign n49012 = n25161 & n29543 ;
  assign n49013 = ( n3831 & ~n7892 ) | ( n3831 & n17167 ) | ( ~n7892 & n17167 ) ;
  assign n49014 = n7754 & n49013 ;
  assign n49015 = n49012 & n49014 ;
  assign n49016 = ( ~n1641 & n45312 ) | ( ~n1641 & n47608 ) | ( n45312 & n47608 ) ;
  assign n49017 = ( n37020 & n39786 ) | ( n37020 & ~n49016 ) | ( n39786 & ~n49016 ) ;
  assign n49018 = ( ~n2892 & n5713 ) | ( ~n2892 & n39756 ) | ( n5713 & n39756 ) ;
  assign n49019 = n16066 | n49018 ;
  assign n49020 = n49019 ^ n31318 ^ n20407 ;
  assign n49021 = ( n3126 & ~n35942 ) | ( n3126 & n45828 ) | ( ~n35942 & n45828 ) ;
  assign n49022 = n24744 ^ n22397 ^ n8510 ;
  assign n49023 = ( n4779 & n26025 ) | ( n4779 & n42145 ) | ( n26025 & n42145 ) ;
  assign n49024 = n38020 ^ n31787 ^ n15620 ;
  assign n49025 = ( ~n8072 & n49023 ) | ( ~n8072 & n49024 ) | ( n49023 & n49024 ) ;
  assign n49026 = ( ~n596 & n4995 ) | ( ~n596 & n22320 ) | ( n4995 & n22320 ) ;
  assign n49027 = n49026 ^ n1494 ^ 1'b0 ;
  assign n49028 = n7325 & n49027 ;
  assign n49029 = n49028 ^ n40394 ^ n8292 ;
  assign n49030 = n18851 ^ n2098 ^ n1301 ;
  assign n49031 = n49030 ^ n37473 ^ n7848 ;
  assign n49032 = n26134 ^ n13610 ^ 1'b0 ;
  assign n49033 = n15744 | n15968 ;
  assign n49034 = n49033 ^ n6168 ^ 1'b0 ;
  assign n49035 = n26034 ^ n20591 ^ 1'b0 ;
  assign n49036 = n21550 ^ n17429 ^ n4342 ;
  assign n49037 = n25893 ^ n17208 ^ n13386 ;
  assign n49038 = ( n42022 & n49036 ) | ( n42022 & n49037 ) | ( n49036 & n49037 ) ;
  assign n49039 = ( ~n36852 & n41937 ) | ( ~n36852 & n49038 ) | ( n41937 & n49038 ) ;
  assign n49040 = n29392 ^ n14670 ^ n14570 ;
  assign n49041 = n33218 ^ n26037 ^ 1'b0 ;
  assign n49042 = n11877 & ~n11982 ;
  assign n49043 = n49042 ^ n2288 ^ 1'b0 ;
  assign n49044 = n49043 ^ n22041 ^ 1'b0 ;
  assign n49045 = n49041 | n49044 ;
  assign n49046 = ( ~n11967 & n22847 ) | ( ~n11967 & n49045 ) | ( n22847 & n49045 ) ;
  assign n49047 = n41826 ^ n40639 ^ n2085 ;
  assign n49048 = ( n10695 & n29392 ) | ( n10695 & ~n49047 ) | ( n29392 & ~n49047 ) ;
  assign n49049 = n24257 ^ n9788 ^ n7239 ;
  assign n49050 = n49049 ^ n13019 ^ n11392 ;
  assign n49053 = n10834 | n11254 ;
  assign n49054 = n49053 ^ n30911 ^ 1'b0 ;
  assign n49051 = n31039 & ~n35800 ;
  assign n49052 = n49051 ^ n3578 ^ n1746 ;
  assign n49055 = n49054 ^ n49052 ^ n15830 ;
  assign n49056 = n40541 ^ n25596 ^ 1'b0 ;
  assign n49057 = n32583 | n49056 ;
  assign n49058 = n26503 | n49057 ;
  assign n49059 = n20880 | n25591 ;
  assign n49060 = ~n13326 & n49059 ;
  assign n49061 = n49060 ^ n12634 ^ 1'b0 ;
  assign n49062 = n44190 ^ n35458 ^ n32923 ;
  assign n49063 = ( n16636 & ~n41746 ) | ( n16636 & n49062 ) | ( ~n41746 & n49062 ) ;
  assign n49064 = ( n16531 & ~n19320 ) | ( n16531 & n49063 ) | ( ~n19320 & n49063 ) ;
  assign n49065 = n39755 ^ n29861 ^ n7723 ;
  assign n49066 = n49065 ^ n46847 ^ n30709 ;
  assign n49067 = n32705 ^ n10707 ^ n4518 ;
  assign n49068 = ( n21666 & n29338 ) | ( n21666 & n49067 ) | ( n29338 & n49067 ) ;
  assign n49069 = n47309 ^ n28984 ^ 1'b0 ;
  assign n49070 = ( ~n13664 & n18444 ) | ( ~n13664 & n18984 ) | ( n18444 & n18984 ) ;
  assign n49071 = ( ~n775 & n6940 ) | ( ~n775 & n39864 ) | ( n6940 & n39864 ) ;
  assign n49072 = ( n5892 & n49070 ) | ( n5892 & n49071 ) | ( n49070 & n49071 ) ;
  assign n49073 = n20771 ^ n16545 ^ n6061 ;
  assign n49076 = n33388 ^ n13429 ^ n7743 ;
  assign n49074 = n12560 ^ n11639 ^ n5578 ;
  assign n49075 = n38942 & n49074 ;
  assign n49077 = n49076 ^ n49075 ^ n46045 ;
  assign n49080 = ( n4887 & ~n22406 ) | ( n4887 & n26588 ) | ( ~n22406 & n26588 ) ;
  assign n49078 = ( n5269 & n7893 ) | ( n5269 & n9858 ) | ( n7893 & n9858 ) ;
  assign n49079 = ~n40195 & n49078 ;
  assign n49081 = n49080 ^ n49079 ^ 1'b0 ;
  assign n49088 = ( n535 & n22346 ) | ( n535 & ~n40247 ) | ( n22346 & ~n40247 ) ;
  assign n49084 = ( n12828 & n18988 ) | ( n12828 & n42630 ) | ( n18988 & n42630 ) ;
  assign n49085 = n34347 ^ n6082 ^ n5705 ;
  assign n49086 = ~n49084 & n49085 ;
  assign n49087 = n49086 ^ n41326 ^ n14811 ;
  assign n49082 = ( n3893 & n11283 ) | ( n3893 & ~n21284 ) | ( n11283 & ~n21284 ) ;
  assign n49083 = ( n5014 & n32443 ) | ( n5014 & ~n49082 ) | ( n32443 & ~n49082 ) ;
  assign n49089 = n49088 ^ n49087 ^ n49083 ;
  assign n49093 = ~n19561 & n26635 ;
  assign n49094 = n49093 ^ n677 ^ 1'b0 ;
  assign n49090 = ( n7584 & n10970 ) | ( n7584 & ~n29263 ) | ( n10970 & ~n29263 ) ;
  assign n49091 = n9971 | n30931 ;
  assign n49092 = n49090 | n49091 ;
  assign n49095 = n49094 ^ n49092 ^ n1178 ;
  assign n49096 = n4891 ^ n2785 ^ x64 ;
  assign n49097 = n31484 ^ n18313 ^ n522 ;
  assign n49098 = ( n21215 & n27582 ) | ( n21215 & n33774 ) | ( n27582 & n33774 ) ;
  assign n49099 = ( ~n4042 & n20461 ) | ( ~n4042 & n49098 ) | ( n20461 & n49098 ) ;
  assign n49100 = ( n49096 & ~n49097 ) | ( n49096 & n49099 ) | ( ~n49097 & n49099 ) ;
  assign n49101 = ( n15850 & n21449 ) | ( n15850 & ~n40838 ) | ( n21449 & ~n40838 ) ;
  assign n49102 = ( n2994 & n34807 ) | ( n2994 & ~n49101 ) | ( n34807 & ~n49101 ) ;
  assign n49110 = n2274 | n46391 ;
  assign n49104 = ( n632 & ~n2241 ) | ( n632 & n6148 ) | ( ~n2241 & n6148 ) ;
  assign n49103 = n3549 & ~n18503 ;
  assign n49105 = n49104 ^ n49103 ^ 1'b0 ;
  assign n49106 = n19700 ^ n5243 ^ n3445 ;
  assign n49107 = n49106 ^ n26661 ^ n5164 ;
  assign n49108 = n35031 ^ n15134 ^ 1'b0 ;
  assign n49109 = ( n49105 & n49107 ) | ( n49105 & ~n49108 ) | ( n49107 & ~n49108 ) ;
  assign n49111 = n49110 ^ n49109 ^ n24268 ;
  assign n49112 = ( n6493 & ~n19075 ) | ( n6493 & n34997 ) | ( ~n19075 & n34997 ) ;
  assign n49113 = n48663 ^ n31439 ^ n21789 ;
  assign n49114 = n49113 ^ n2063 ^ 1'b0 ;
  assign n49115 = ( n26528 & ~n49112 ) | ( n26528 & n49114 ) | ( ~n49112 & n49114 ) ;
  assign n49116 = n18549 ^ n11619 ^ n11053 ;
  assign n49117 = n49116 ^ n9600 ^ 1'b0 ;
  assign n49118 = ~n9204 & n49117 ;
  assign n49119 = n49118 ^ n16970 ^ n15199 ;
  assign n49120 = n49119 ^ n31261 ^ n10411 ;
  assign n49121 = ( n44572 & n48262 ) | ( n44572 & ~n49120 ) | ( n48262 & ~n49120 ) ;
  assign n49122 = n1630 & n25842 ;
  assign n49123 = n49122 ^ n11525 ^ 1'b0 ;
  assign n49124 = n17892 ^ n16832 ^ 1'b0 ;
  assign n49125 = n46071 & ~n49124 ;
  assign n49126 = n38976 ^ n21785 ^ n9589 ;
  assign n49127 = n49126 ^ n28763 ^ n22275 ;
  assign n49128 = ( n31460 & ~n45371 ) | ( n31460 & n49127 ) | ( ~n45371 & n49127 ) ;
  assign n49129 = ~n1912 & n8294 ;
  assign n49130 = n49129 ^ n11247 ^ 1'b0 ;
  assign n49131 = ( ~n22656 & n25629 ) | ( ~n22656 & n49130 ) | ( n25629 & n49130 ) ;
  assign n49139 = n25001 & n27393 ;
  assign n49140 = n49139 ^ n26208 ^ n2668 ;
  assign n49141 = n49140 ^ n35996 ^ n4455 ;
  assign n49134 = n6914 ^ n6360 ^ n2944 ;
  assign n49132 = n19107 ^ n8428 ^ n7995 ;
  assign n49133 = n49132 ^ n7978 ^ n5997 ;
  assign n49135 = n49134 ^ n49133 ^ n2094 ;
  assign n49136 = ( n12707 & n21845 ) | ( n12707 & n22800 ) | ( n21845 & n22800 ) ;
  assign n49137 = n49136 ^ n47377 ^ n14074 ;
  assign n49138 = ( n5608 & n49135 ) | ( n5608 & ~n49137 ) | ( n49135 & ~n49137 ) ;
  assign n49142 = n49141 ^ n49138 ^ 1'b0 ;
  assign n49143 = ( ~n13288 & n21133 ) | ( ~n13288 & n27590 ) | ( n21133 & n27590 ) ;
  assign n49144 = ( ~n10908 & n25129 ) | ( ~n10908 & n37004 ) | ( n25129 & n37004 ) ;
  assign n49145 = n5219 ^ n476 ^ 1'b0 ;
  assign n49146 = ( n4528 & n6498 ) | ( n4528 & ~n45864 ) | ( n6498 & ~n45864 ) ;
  assign n49147 = n49146 ^ n14251 ^ x88 ;
  assign n49151 = ( n7704 & ~n8983 ) | ( n7704 & n32211 ) | ( ~n8983 & n32211 ) ;
  assign n49148 = n9143 ^ n5088 ^ 1'b0 ;
  assign n49149 = n4657 & ~n49148 ;
  assign n49150 = n49149 ^ n26073 ^ n25692 ;
  assign n49152 = n49151 ^ n49150 ^ n19889 ;
  assign n49153 = n11465 ^ n5277 ^ 1'b0 ;
  assign n49154 = n7786 ^ n3009 ^ n2583 ;
  assign n49155 = ( n17888 & n49153 ) | ( n17888 & ~n49154 ) | ( n49153 & ~n49154 ) ;
  assign n49156 = n49155 ^ n26192 ^ x60 ;
  assign n49157 = ( n28098 & n34373 ) | ( n28098 & n49156 ) | ( n34373 & n49156 ) ;
  assign n49158 = n49157 ^ n40011 ^ n9932 ;
  assign n49159 = n30186 ^ n30013 ^ 1'b0 ;
  assign n49160 = ~n11256 & n49159 ;
  assign n49161 = n2902 ^ n2046 ^ n1866 ;
  assign n49162 = n49161 ^ n7351 ^ n1735 ;
  assign n49163 = n49162 ^ n43663 ^ 1'b0 ;
  assign n49164 = n26994 & ~n49163 ;
  assign n49165 = ( n15693 & n43269 ) | ( n15693 & ~n43905 ) | ( n43269 & ~n43905 ) ;
  assign n49166 = ( n2657 & ~n13893 ) | ( n2657 & n29435 ) | ( ~n13893 & n29435 ) ;
  assign n49167 = ( n9024 & n24487 ) | ( n9024 & ~n26590 ) | ( n24487 & ~n26590 ) ;
  assign n49168 = n38805 ^ n20614 ^ n6880 ;
  assign n49169 = n49168 ^ n48921 ^ n18519 ;
  assign n49170 = ( ~n1112 & n23207 ) | ( ~n1112 & n47033 ) | ( n23207 & n47033 ) ;
  assign n49171 = n49170 ^ n18610 ^ n13940 ;
  assign n49172 = ( ~n4101 & n16890 ) | ( ~n4101 & n26847 ) | ( n16890 & n26847 ) ;
  assign n49173 = n49172 ^ n36436 ^ n8714 ;
  assign n49174 = n3561 | n49173 ;
  assign n49175 = n33531 & ~n49174 ;
  assign n49176 = ( n829 & n46514 ) | ( n829 & ~n49175 ) | ( n46514 & ~n49175 ) ;
  assign n49177 = ( ~n17668 & n33478 ) | ( ~n17668 & n42942 ) | ( n33478 & n42942 ) ;
  assign n49178 = ( n1193 & ~n1811 ) | ( n1193 & n9746 ) | ( ~n1811 & n9746 ) ;
  assign n49179 = n49178 ^ n41060 ^ n15812 ;
  assign n49180 = n11970 ^ n7642 ^ n5539 ;
  assign n49181 = ( n19999 & n22042 ) | ( n19999 & ~n49180 ) | ( n22042 & ~n49180 ) ;
  assign n49182 = n33388 | n49181 ;
  assign n49183 = n49182 ^ n14791 ^ 1'b0 ;
  assign n49187 = n31822 | n36590 ;
  assign n49185 = ( x246 & n5310 ) | ( x246 & ~n12627 ) | ( n5310 & ~n12627 ) ;
  assign n49186 = ( n4075 & ~n18101 ) | ( n4075 & n49185 ) | ( ~n18101 & n49185 ) ;
  assign n49188 = n49187 ^ n49186 ^ n21105 ;
  assign n49189 = n41216 | n49188 ;
  assign n49184 = n35105 ^ n19685 ^ n8480 ;
  assign n49190 = n49189 ^ n49184 ^ n16614 ;
  assign n49191 = n41217 ^ n35982 ^ n9395 ;
  assign n49195 = n25521 ^ n16324 ^ 1'b0 ;
  assign n49192 = ( n5206 & ~n28851 ) | ( n5206 & n34050 ) | ( ~n28851 & n34050 ) ;
  assign n49193 = n26845 | n40131 ;
  assign n49194 = n49192 & ~n49193 ;
  assign n49196 = n49195 ^ n49194 ^ n27308 ;
  assign n49197 = n22931 ^ n6564 ^ 1'b0 ;
  assign n49198 = n31427 & n49197 ;
  assign n49199 = ( n1563 & n6819 ) | ( n1563 & ~n49198 ) | ( n6819 & ~n49198 ) ;
  assign n49200 = n13448 ^ n9789 ^ n2274 ;
  assign n49201 = n49200 ^ n44209 ^ n25414 ;
  assign n49202 = ( n19104 & n49199 ) | ( n19104 & n49201 ) | ( n49199 & n49201 ) ;
  assign n49205 = ( ~n3395 & n9433 ) | ( ~n3395 & n17363 ) | ( n9433 & n17363 ) ;
  assign n49206 = n19929 & n49205 ;
  assign n49203 = n1054 | n6903 ;
  assign n49204 = n49203 ^ n41502 ^ 1'b0 ;
  assign n49207 = n49206 ^ n49204 ^ n16104 ;
  assign n49208 = ~n7446 & n30706 ;
  assign n49209 = n36399 & n49208 ;
  assign n49210 = n49209 ^ n45473 ^ n4807 ;
  assign n49211 = n23556 ^ n12136 ^ 1'b0 ;
  assign n49212 = n44724 ^ n2838 ^ n2653 ;
  assign n49219 = n34916 ^ n23734 ^ n3491 ;
  assign n49216 = n31962 ^ n28798 ^ n18910 ;
  assign n49214 = n34175 ^ n29181 ^ n26865 ;
  assign n49213 = n784 & ~n36206 ;
  assign n49215 = n49214 ^ n49213 ^ 1'b0 ;
  assign n49217 = n49216 ^ n49215 ^ n26847 ;
  assign n49218 = ( n21640 & n43695 ) | ( n21640 & ~n49217 ) | ( n43695 & ~n49217 ) ;
  assign n49220 = n49219 ^ n49218 ^ n45037 ;
  assign n49221 = n37358 ^ n17483 ^ n14304 ;
  assign n49222 = n49221 ^ n34943 ^ n6040 ;
  assign n49223 = n24656 & ~n25008 ;
  assign n49224 = ( n32542 & ~n44718 ) | ( n32542 & n49223 ) | ( ~n44718 & n49223 ) ;
  assign n49225 = n49224 ^ n41463 ^ x60 ;
  assign n49228 = n32379 ^ n4118 ^ 1'b0 ;
  assign n49226 = ( ~n4202 & n11689 ) | ( ~n4202 & n11926 ) | ( n11689 & n11926 ) ;
  assign n49227 = ( ~n17228 & n23663 ) | ( ~n17228 & n49226 ) | ( n23663 & n49226 ) ;
  assign n49229 = n49228 ^ n49227 ^ n39095 ;
  assign n49230 = ( n6494 & n18468 ) | ( n6494 & ~n33204 ) | ( n18468 & ~n33204 ) ;
  assign n49231 = n36068 ^ n24189 ^ n9386 ;
  assign n49232 = ( n34173 & n45287 ) | ( n34173 & n49231 ) | ( n45287 & n49231 ) ;
  assign n49233 = ( ~n8014 & n8711 ) | ( ~n8014 & n36365 ) | ( n8711 & n36365 ) ;
  assign n49234 = ( n4405 & n5344 ) | ( n4405 & n15102 ) | ( n5344 & n15102 ) ;
  assign n49235 = n4389 ^ n1109 ^ 1'b0 ;
  assign n49236 = n47609 | n49235 ;
  assign n49238 = ( n5280 & n8433 ) | ( n5280 & n12822 ) | ( n8433 & n12822 ) ;
  assign n49239 = ( n16501 & n18069 ) | ( n16501 & n49238 ) | ( n18069 & n49238 ) ;
  assign n49237 = n32859 ^ n29448 ^ n25408 ;
  assign n49240 = n49239 ^ n49237 ^ n9357 ;
  assign n49241 = n48067 ^ n24581 ^ n8055 ;
  assign n49242 = n15647 ^ n6855 ^ x236 ;
  assign n49243 = ( ~n20579 & n38763 ) | ( ~n20579 & n49242 ) | ( n38763 & n49242 ) ;
  assign n49244 = n49243 ^ n45396 ^ n3140 ;
  assign n49245 = n49244 ^ n38943 ^ 1'b0 ;
  assign n49246 = n13554 ^ n10086 ^ n4198 ;
  assign n49247 = n49246 ^ n18598 ^ n11845 ;
  assign n49248 = n48410 ^ n24423 ^ n14791 ;
  assign n49249 = n49248 ^ n27000 ^ n6858 ;
  assign n49250 = n44571 ^ n13468 ^ n3112 ;
  assign n49251 = n49250 ^ n4308 ^ 1'b0 ;
  assign n49252 = ( ~n1259 & n13473 ) | ( ~n1259 & n49251 ) | ( n13473 & n49251 ) ;
  assign n49253 = ( ~n11945 & n12165 ) | ( ~n11945 & n31017 ) | ( n12165 & n31017 ) ;
  assign n49254 = ( ~n1236 & n2528 ) | ( ~n1236 & n49253 ) | ( n2528 & n49253 ) ;
  assign n49255 = n31783 ^ n21185 ^ n2766 ;
  assign n49256 = x37 & ~n46947 ;
  assign n49257 = ~n49255 & n49256 ;
  assign n49258 = n4414 & ~n12782 ;
  assign n49259 = n21379 & n49258 ;
  assign n49260 = ( n1761 & n36021 ) | ( n1761 & n46906 ) | ( n36021 & n46906 ) ;
  assign n49261 = n11877 & ~n22222 ;
  assign n49262 = ( n22494 & n36046 ) | ( n22494 & n44216 ) | ( n36046 & n44216 ) ;
  assign n49263 = ( ~n8256 & n8385 ) | ( ~n8256 & n13059 ) | ( n8385 & n13059 ) ;
  assign n49264 = ( n13615 & n13726 ) | ( n13615 & n49263 ) | ( n13726 & n49263 ) ;
  assign n49265 = ( n31491 & n41149 ) | ( n31491 & ~n49264 ) | ( n41149 & ~n49264 ) ;
  assign n49266 = n49265 ^ n28419 ^ n21234 ;
  assign n49267 = ( n33721 & ~n37262 ) | ( n33721 & n49266 ) | ( ~n37262 & n49266 ) ;
  assign n49268 = n14332 ^ n13218 ^ n3054 ;
  assign n49269 = n23156 & ~n49268 ;
  assign n49270 = n10215 ^ n8456 ^ n1131 ;
  assign n49271 = n49270 ^ n33104 ^ n23447 ;
  assign n49272 = n25322 ^ n24312 ^ n19094 ;
  assign n49273 = n49272 ^ n36872 ^ n13420 ;
  assign n49275 = ( n16771 & n17147 ) | ( n16771 & n23360 ) | ( n17147 & n23360 ) ;
  assign n49274 = x47 & n48756 ;
  assign n49276 = n49275 ^ n49274 ^ n35034 ;
  assign n49277 = n1925 & n9829 ;
  assign n49278 = n49277 ^ n9640 ^ 1'b0 ;
  assign n49279 = n7904 & n49278 ;
  assign n49280 = n20943 & n49279 ;
  assign n49281 = n43738 ^ n3087 ^ 1'b0 ;
  assign n49282 = n10308 & n49281 ;
  assign n49283 = n24958 ^ n19774 ^ n9201 ;
  assign n49284 = n16950 ^ n14405 ^ n4099 ;
  assign n49285 = ( ~n792 & n39238 ) | ( ~n792 & n49284 ) | ( n39238 & n49284 ) ;
  assign n49286 = n14725 ^ n13347 ^ n1841 ;
  assign n49287 = n49286 ^ n20880 ^ n2793 ;
  assign n49288 = n6351 & n28271 ;
  assign n49289 = ~n49287 & n49288 ;
  assign n49290 = ( n22004 & ~n49285 ) | ( n22004 & n49289 ) | ( ~n49285 & n49289 ) ;
  assign n49291 = ( n37892 & n49283 ) | ( n37892 & ~n49290 ) | ( n49283 & ~n49290 ) ;
  assign n49292 = n20708 ^ n20128 ^ 1'b0 ;
  assign n49293 = ( n12799 & n29737 ) | ( n12799 & ~n33852 ) | ( n29737 & ~n33852 ) ;
  assign n49294 = n38240 ^ n33848 ^ 1'b0 ;
  assign n49295 = ( n2984 & ~n7399 ) | ( n2984 & n13405 ) | ( ~n7399 & n13405 ) ;
  assign n49296 = ( x147 & n3514 ) | ( x147 & ~n49295 ) | ( n3514 & ~n49295 ) ;
  assign n49297 = n49296 ^ n31557 ^ n28232 ;
  assign n49298 = n40731 ^ n18740 ^ 1'b0 ;
  assign n49299 = ( ~n1415 & n14349 ) | ( ~n1415 & n42858 ) | ( n14349 & n42858 ) ;
  assign n49300 = ( n13153 & ~n26631 ) | ( n13153 & n27400 ) | ( ~n26631 & n27400 ) ;
  assign n49301 = n49300 ^ n9895 ^ n3494 ;
  assign n49302 = n20459 & n36807 ;
  assign n49303 = n7783 ^ n2716 ^ n1100 ;
  assign n49304 = n49303 ^ n20640 ^ n12519 ;
  assign n49305 = n29683 ^ n16885 ^ n2438 ;
  assign n49306 = n49305 ^ n39496 ^ 1'b0 ;
  assign n49307 = n44954 ^ n13846 ^ n12701 ;
  assign n49308 = ( n11718 & n20039 ) | ( n11718 & ~n29649 ) | ( n20039 & ~n29649 ) ;
  assign n49309 = ( ~n45847 & n49307 ) | ( ~n45847 & n49308 ) | ( n49307 & n49308 ) ;
  assign n49310 = ( n13282 & n20843 ) | ( n13282 & n27398 ) | ( n20843 & n27398 ) ;
  assign n49311 = ( n5327 & n22964 ) | ( n5327 & ~n49310 ) | ( n22964 & ~n49310 ) ;
  assign n49312 = n4429 ^ n1044 ^ n782 ;
  assign n49313 = n41328 ^ n24190 ^ n4195 ;
  assign n49314 = n49313 ^ n440 ^ x226 ;
  assign n49315 = ( n11681 & ~n16334 ) | ( n11681 & n40273 ) | ( ~n16334 & n40273 ) ;
  assign n49316 = n43055 ^ n24539 ^ n13494 ;
  assign n49317 = ( n1551 & n20092 ) | ( n1551 & n23807 ) | ( n20092 & n23807 ) ;
  assign n49318 = ( ~n10396 & n49316 ) | ( ~n10396 & n49317 ) | ( n49316 & n49317 ) ;
  assign n49319 = ( ~n4988 & n49315 ) | ( ~n4988 & n49318 ) | ( n49315 & n49318 ) ;
  assign n49320 = n47034 ^ n35522 ^ n20834 ;
  assign n49321 = n11065 & ~n15189 ;
  assign n49322 = n28983 ^ n27811 ^ n2159 ;
  assign n49324 = ( n2058 & n32622 ) | ( n2058 & ~n44425 ) | ( n32622 & ~n44425 ) ;
  assign n49323 = ~n37733 & n47735 ;
  assign n49325 = n49324 ^ n49323 ^ 1'b0 ;
  assign n49326 = n49325 ^ n39602 ^ n10458 ;
  assign n49327 = n49326 ^ n44510 ^ n31568 ;
  assign n49328 = n34816 ^ n16948 ^ n8340 ;
  assign n49329 = n49328 ^ n36846 ^ n17745 ;
  assign n49333 = n12588 ^ n5078 ^ n998 ;
  assign n49334 = ( n6439 & ~n29526 ) | ( n6439 & n49333 ) | ( ~n29526 & n49333 ) ;
  assign n49330 = n1929 & n22723 ;
  assign n49331 = ~n44023 & n49330 ;
  assign n49332 = n49331 ^ n39015 ^ n30823 ;
  assign n49335 = n49334 ^ n49332 ^ n21246 ;
  assign n49336 = ( n31649 & ~n32360 ) | ( n31649 & n42929 ) | ( ~n32360 & n42929 ) ;
  assign n49337 = n21932 | n41888 ;
  assign n49338 = n49337 ^ n23647 ^ 1'b0 ;
  assign n49339 = n49338 ^ n16861 ^ n11645 ;
  assign n49340 = ~n39098 & n43876 ;
  assign n49341 = n43426 & n49340 ;
  assign n49342 = n49341 ^ n45767 ^ n2340 ;
  assign n49344 = ~n28492 & n36533 ;
  assign n49345 = n41813 & n49344 ;
  assign n49343 = n812 | n30368 ;
  assign n49346 = n49345 ^ n49343 ^ 1'b0 ;
  assign n49347 = n23084 & ~n28638 ;
  assign n49348 = ( n4615 & ~n10843 ) | ( n4615 & n49347 ) | ( ~n10843 & n49347 ) ;
  assign n49349 = n49348 ^ n29221 ^ n3256 ;
  assign n49350 = n47672 ^ n20586 ^ n11465 ;
  assign n49351 = n49350 ^ n3840 ^ n2727 ;
  assign n49352 = n33135 ^ n15696 ^ 1'b0 ;
  assign n49353 = ( x96 & n17067 ) | ( x96 & ~n20278 ) | ( n17067 & ~n20278 ) ;
  assign n49354 = ~n31415 & n49353 ;
  assign n49355 = n49354 ^ n40952 ^ n29450 ;
  assign n49357 = ( n17163 & n31210 ) | ( n17163 & n39076 ) | ( n31210 & n39076 ) ;
  assign n49356 = n3304 | n33204 ;
  assign n49358 = n49357 ^ n49356 ^ 1'b0 ;
  assign n49359 = ( ~n27161 & n27184 ) | ( ~n27161 & n49358 ) | ( n27184 & n49358 ) ;
  assign n49362 = n33076 ^ n11154 ^ 1'b0 ;
  assign n49363 = ~n30493 & n49362 ;
  assign n49360 = n21096 ^ n14140 ^ 1'b0 ;
  assign n49361 = n49360 ^ n3483 ^ x100 ;
  assign n49364 = n49363 ^ n49361 ^ n14826 ;
  assign n49365 = ~n48551 & n49364 ;
  assign n49366 = ( n10803 & n49359 ) | ( n10803 & ~n49365 ) | ( n49359 & ~n49365 ) ;
  assign n49367 = ( ~n3238 & n26757 ) | ( ~n3238 & n39271 ) | ( n26757 & n39271 ) ;
  assign n49368 = n49367 ^ n21632 ^ n4999 ;
  assign n49369 = n49067 ^ n15790 ^ n6354 ;
  assign n49370 = n6262 ^ n4085 ^ n951 ;
  assign n49371 = ( n275 & ~n23383 ) | ( n275 & n49370 ) | ( ~n23383 & n49370 ) ;
  assign n49372 = n49371 ^ n16480 ^ n9382 ;
  assign n49373 = n37610 ^ n7192 ^ n6399 ;
  assign n49374 = ( n3639 & n7819 ) | ( n3639 & ~n15158 ) | ( n7819 & ~n15158 ) ;
  assign n49375 = ( n5405 & n48333 ) | ( n5405 & n49374 ) | ( n48333 & n49374 ) ;
  assign n49376 = n2417 & ~n2943 ;
  assign n49377 = ( ~n1532 & n4798 ) | ( ~n1532 & n16563 ) | ( n4798 & n16563 ) ;
  assign n49378 = ( n17214 & n49376 ) | ( n17214 & ~n49377 ) | ( n49376 & ~n49377 ) ;
  assign n49381 = n1471 ^ n1052 ^ x5 ;
  assign n49382 = ( n17874 & n20541 ) | ( n17874 & ~n49381 ) | ( n20541 & ~n49381 ) ;
  assign n49383 = n49382 ^ n44960 ^ n12280 ;
  assign n49379 = ( n15575 & ~n18188 ) | ( n15575 & n25864 ) | ( ~n18188 & n25864 ) ;
  assign n49380 = n49379 ^ n26472 ^ n20395 ;
  assign n49384 = n49383 ^ n49380 ^ n36096 ;
  assign n49385 = n49384 ^ n30881 ^ x192 ;
  assign n49386 = ( n46548 & n49378 ) | ( n46548 & ~n49385 ) | ( n49378 & ~n49385 ) ;
  assign n49387 = n10005 ^ n9712 ^ n1197 ;
  assign n49388 = n42846 ^ n13271 ^ n3813 ;
  assign n49389 = n44107 ^ n43418 ^ n36757 ;
  assign n49395 = ( n18332 & n27581 ) | ( n18332 & n39302 ) | ( n27581 & n39302 ) ;
  assign n49394 = n22052 ^ n5767 ^ x137 ;
  assign n49390 = ( ~n17844 & n23916 ) | ( ~n17844 & n37909 ) | ( n23916 & n37909 ) ;
  assign n49391 = ( ~n10420 & n21428 ) | ( ~n10420 & n49390 ) | ( n21428 & n49390 ) ;
  assign n49392 = ( n18643 & ~n31712 ) | ( n18643 & n32808 ) | ( ~n31712 & n32808 ) ;
  assign n49393 = ( n4998 & ~n49391 ) | ( n4998 & n49392 ) | ( ~n49391 & n49392 ) ;
  assign n49396 = n49395 ^ n49394 ^ n49393 ;
  assign n49400 = n5399 ^ n3056 ^ 1'b0 ;
  assign n49401 = n21388 | n49400 ;
  assign n49398 = ( n14017 & n18333 ) | ( n14017 & n29494 ) | ( n18333 & n29494 ) ;
  assign n49399 = n49398 ^ n36150 ^ n34428 ;
  assign n49397 = n20640 ^ n3588 ^ n1194 ;
  assign n49402 = n49401 ^ n49399 ^ n49397 ;
  assign n49403 = ( ~n11290 & n32495 ) | ( ~n11290 & n43006 ) | ( n32495 & n43006 ) ;
  assign n49404 = n49403 ^ n27840 ^ 1'b0 ;
  assign n49405 = ~n17468 & n49404 ;
  assign n49406 = n37836 ^ n10439 ^ n3746 ;
  assign n49407 = ( n11775 & ~n12011 ) | ( n11775 & n40666 ) | ( ~n12011 & n40666 ) ;
  assign n49408 = ( x169 & ~n49406 ) | ( x169 & n49407 ) | ( ~n49406 & n49407 ) ;
  assign n49409 = ( n12646 & ~n16959 ) | ( n12646 & n22701 ) | ( ~n16959 & n22701 ) ;
  assign n49410 = n8576 & ~n14859 ;
  assign n49411 = ( n18163 & ~n49409 ) | ( n18163 & n49410 ) | ( ~n49409 & n49410 ) ;
  assign n49412 = n11886 ^ n11198 ^ n5534 ;
  assign n49413 = ( n4413 & n40877 ) | ( n4413 & n49412 ) | ( n40877 & n49412 ) ;
  assign n49418 = ( n15520 & ~n37825 ) | ( n15520 & n43977 ) | ( ~n37825 & n43977 ) ;
  assign n49414 = n12839 ^ n12126 ^ n1398 ;
  assign n49415 = n49414 ^ n14524 ^ n12583 ;
  assign n49416 = n49415 ^ n41386 ^ n2864 ;
  assign n49417 = ( n5414 & ~n25832 ) | ( n5414 & n49416 ) | ( ~n25832 & n49416 ) ;
  assign n49419 = n49418 ^ n49417 ^ n2028 ;
  assign n49420 = n39698 ^ n1443 ^ 1'b0 ;
  assign n49421 = n6351 ^ n3052 ^ n529 ;
  assign n49422 = n49421 ^ n46110 ^ n24985 ;
  assign n49423 = n42050 ^ n39340 ^ n14163 ;
  assign n49424 = n33892 ^ n11990 ^ n1553 ;
  assign n49425 = ( n406 & n6201 ) | ( n406 & ~n6714 ) | ( n6201 & ~n6714 ) ;
  assign n49426 = n49425 ^ n14972 ^ n8052 ;
  assign n49427 = ( n20676 & n40044 ) | ( n20676 & n49426 ) | ( n40044 & n49426 ) ;
  assign n49428 = n18555 & ~n38528 ;
  assign n49429 = n49428 ^ n21591 ^ 1'b0 ;
  assign n49430 = ( n8706 & n27772 ) | ( n8706 & ~n28548 ) | ( n27772 & ~n28548 ) ;
  assign n49431 = n49430 ^ n41468 ^ n31799 ;
  assign n49432 = ( ~n1406 & n12027 ) | ( ~n1406 & n28653 ) | ( n12027 & n28653 ) ;
  assign n49433 = n49432 ^ n21231 ^ n19812 ;
  assign n49434 = ~n3150 & n49433 ;
  assign n49435 = ~n23783 & n49434 ;
  assign n49436 = ( n7557 & n47601 ) | ( n7557 & n49435 ) | ( n47601 & n49435 ) ;
  assign n49437 = n18500 ^ n6506 ^ n1112 ;
  assign n49438 = ( n10741 & ~n19186 ) | ( n10741 & n49437 ) | ( ~n19186 & n49437 ) ;
  assign n49439 = n19211 ^ n11817 ^ n8333 ;
  assign n49440 = ( n34775 & n49438 ) | ( n34775 & ~n49439 ) | ( n49438 & ~n49439 ) ;
  assign n49441 = ( n22377 & n33875 ) | ( n22377 & ~n49347 ) | ( n33875 & ~n49347 ) ;
  assign n49442 = ( n8903 & n19815 ) | ( n8903 & n24804 ) | ( n19815 & n24804 ) ;
  assign n49443 = ( ~n4742 & n26006 ) | ( ~n4742 & n40809 ) | ( n26006 & n40809 ) ;
  assign n49444 = n40412 ^ n37425 ^ n10150 ;
  assign n49445 = n22820 & ~n49444 ;
  assign n49446 = ~n16428 & n49445 ;
  assign n49447 = ~n26184 & n43235 ;
  assign n49448 = n49447 ^ n23659 ^ 1'b0 ;
  assign n49449 = ( n27648 & n30973 ) | ( n27648 & n49448 ) | ( n30973 & n49448 ) ;
  assign n49450 = n49449 ^ n32887 ^ n32227 ;
  assign n49451 = n49450 ^ n2664 ^ 1'b0 ;
  assign n49452 = n23065 & n49451 ;
  assign n49453 = ( n3403 & n25968 ) | ( n3403 & n26069 ) | ( n25968 & n26069 ) ;
  assign n49454 = ( n14235 & n16956 ) | ( n14235 & ~n49453 ) | ( n16956 & ~n49453 ) ;
  assign n49455 = ( ~n21029 & n29608 ) | ( ~n21029 & n44596 ) | ( n29608 & n44596 ) ;
  assign n49456 = n20104 & ~n45866 ;
  assign n49457 = n19357 & ~n36307 ;
  assign n49458 = ( n3372 & n13935 ) | ( n3372 & n18889 ) | ( n13935 & n18889 ) ;
  assign n49459 = n49458 ^ n32973 ^ n9785 ;
  assign n49460 = n39443 ^ n27995 ^ 1'b0 ;
  assign n49461 = ( n2165 & ~n5729 ) | ( n2165 & n12220 ) | ( ~n5729 & n12220 ) ;
  assign n49462 = n49461 ^ n20098 ^ n6932 ;
  assign n49463 = n23755 & ~n38602 ;
  assign n49464 = n49463 ^ n27524 ^ 1'b0 ;
  assign n49465 = ( n37067 & n43895 ) | ( n37067 & ~n49464 ) | ( n43895 & ~n49464 ) ;
  assign n49466 = ( n1732 & n48401 ) | ( n1732 & ~n49465 ) | ( n48401 & ~n49465 ) ;
  assign n49467 = n47396 ^ n27533 ^ n10993 ;
  assign n49468 = ( n9021 & n15773 ) | ( n9021 & ~n44510 ) | ( n15773 & ~n44510 ) ;
  assign n49469 = ~n15757 & n49468 ;
  assign n49470 = n27894 | n49469 ;
  assign n49471 = ( n1757 & n16578 ) | ( n1757 & ~n49470 ) | ( n16578 & ~n49470 ) ;
  assign n49472 = ( n7795 & n8424 ) | ( n7795 & n20086 ) | ( n8424 & n20086 ) ;
  assign n49473 = n49472 ^ n35826 ^ n4915 ;
  assign n49474 = n47850 | n49473 ;
  assign n49475 = n49471 & ~n49474 ;
  assign n49476 = n22388 ^ n13874 ^ n4018 ;
  assign n49477 = n49476 ^ n18505 ^ n1651 ;
  assign n49478 = n49477 ^ n40602 ^ n15478 ;
  assign n49479 = n11663 & ~n37491 ;
  assign n49480 = n49479 ^ n19050 ^ 1'b0 ;
  assign n49481 = n49480 ^ n1734 ^ 1'b0 ;
  assign n49482 = n49478 & ~n49481 ;
  assign n49484 = n27589 ^ n15128 ^ n14788 ;
  assign n49485 = ( n14980 & ~n27668 ) | ( n14980 & n49484 ) | ( ~n27668 & n49484 ) ;
  assign n49486 = ( n8567 & ~n11153 ) | ( n8567 & n49485 ) | ( ~n11153 & n49485 ) ;
  assign n49487 = n49486 ^ n15017 ^ n7096 ;
  assign n49483 = n33943 ^ n31851 ^ n20816 ;
  assign n49488 = n49487 ^ n49483 ^ n7472 ;
  assign n49489 = n39343 ^ n32233 ^ n3948 ;
  assign n49490 = n49489 ^ n4387 ^ n2640 ;
  assign n49491 = n44910 ^ n12519 ^ n8991 ;
  assign n49492 = ~n5597 & n23156 ;
  assign n49493 = n7343 | n49492 ;
  assign n49494 = n35771 ^ n27924 ^ n9692 ;
  assign n49495 = ( ~n8269 & n13632 ) | ( ~n8269 & n49494 ) | ( n13632 & n49494 ) ;
  assign n49496 = ( ~n1647 & n4267 ) | ( ~n1647 & n42566 ) | ( n4267 & n42566 ) ;
  assign n49497 = n49496 ^ n39612 ^ n37553 ;
  assign n49498 = n6021 ^ n5159 ^ n4817 ;
  assign n49499 = ( n364 & n8159 ) | ( n364 & ~n49498 ) | ( n8159 & ~n49498 ) ;
  assign n49500 = n49499 ^ n24033 ^ n22092 ;
  assign n49501 = n12031 ^ n5429 ^ n1662 ;
  assign n49502 = n44115 ^ x193 ^ 1'b0 ;
  assign n49503 = n36881 & n49502 ;
  assign n49504 = ( ~n6737 & n16672 ) | ( ~n6737 & n26503 ) | ( n16672 & n26503 ) ;
  assign n49505 = n49504 ^ n41204 ^ 1'b0 ;
  assign n49506 = n34228 & n49505 ;
  assign n49507 = n44889 ^ n42484 ^ n17046 ;
  assign n49508 = ( n31748 & ~n38095 ) | ( n31748 & n49507 ) | ( ~n38095 & n49507 ) ;
  assign n49509 = n42221 ^ n29208 ^ n17123 ;
  assign n49515 = n610 & ~n26310 ;
  assign n49516 = n49515 ^ n15500 ^ 1'b0 ;
  assign n49517 = ( n35211 & n44602 ) | ( n35211 & ~n49516 ) | ( n44602 & ~n49516 ) ;
  assign n49513 = ( n1691 & n9175 ) | ( n1691 & n39231 ) | ( n9175 & n39231 ) ;
  assign n49514 = ( n8499 & n8603 ) | ( n8499 & ~n49513 ) | ( n8603 & ~n49513 ) ;
  assign n49510 = n1993 & ~n12800 ;
  assign n49511 = n5775 & n49510 ;
  assign n49512 = ( n10113 & n12381 ) | ( n10113 & n49511 ) | ( n12381 & n49511 ) ;
  assign n49518 = n49517 ^ n49514 ^ n49512 ;
  assign n49519 = ( ~n11098 & n14802 ) | ( ~n11098 & n39893 ) | ( n14802 & n39893 ) ;
  assign n49520 = n25815 ^ n22574 ^ n7825 ;
  assign n49521 = ( n10949 & n12869 ) | ( n10949 & ~n27606 ) | ( n12869 & ~n27606 ) ;
  assign n49522 = ( n8925 & n31165 ) | ( n8925 & ~n49521 ) | ( n31165 & ~n49521 ) ;
  assign n49523 = n17747 ^ n680 ^ 1'b0 ;
  assign n49524 = n48176 ^ n29928 ^ n21253 ;
  assign n49525 = ~n20212 & n24447 ;
  assign n49526 = n26035 ^ n19294 ^ x242 ;
  assign n49527 = n22369 ^ n12506 ^ n8531 ;
  assign n49528 = ( n24261 & n27650 ) | ( n24261 & ~n49527 ) | ( n27650 & ~n49527 ) ;
  assign n49529 = ( n5445 & ~n37882 ) | ( n5445 & n38242 ) | ( ~n37882 & n38242 ) ;
  assign n49530 = ( n4100 & n13868 ) | ( n4100 & ~n49529 ) | ( n13868 & ~n49529 ) ;
  assign n49531 = n18171 ^ n10824 ^ n1500 ;
  assign n49532 = n27533 ^ n5168 ^ x22 ;
  assign n49533 = ( n11215 & n34901 ) | ( n11215 & n49532 ) | ( n34901 & n49532 ) ;
  assign n49534 = ( n5376 & n14728 ) | ( n5376 & ~n41192 ) | ( n14728 & ~n41192 ) ;
  assign n49535 = n2043 | n38897 ;
  assign n49536 = ( n23144 & n34258 ) | ( n23144 & n49535 ) | ( n34258 & n49535 ) ;
  assign n49537 = ( n17005 & n22756 ) | ( n17005 & n49092 ) | ( n22756 & n49092 ) ;
  assign n49538 = n13812 & ~n24295 ;
  assign n49539 = n7224 & n49538 ;
  assign n49540 = n1449 & ~n49539 ;
  assign n49541 = n44935 & n49540 ;
  assign n49542 = ~n7742 & n39805 ;
  assign n49543 = n24592 & n49542 ;
  assign n49544 = n27907 ^ n17578 ^ n13835 ;
  assign n49545 = ( n3488 & ~n8604 ) | ( n3488 & n9541 ) | ( ~n8604 & n9541 ) ;
  assign n49546 = n36712 ^ n17503 ^ 1'b0 ;
  assign n49547 = ( n5395 & n49545 ) | ( n5395 & n49546 ) | ( n49545 & n49546 ) ;
  assign n49548 = n49547 ^ n47308 ^ n40394 ;
  assign n49549 = n45026 ^ n42796 ^ n27828 ;
  assign n49550 = n9472 & n35551 ;
  assign n49551 = ( n11582 & ~n40982 ) | ( n11582 & n49550 ) | ( ~n40982 & n49550 ) ;
  assign n49552 = ( n3814 & n11160 ) | ( n3814 & ~n11736 ) | ( n11160 & ~n11736 ) ;
  assign n49553 = ( n15170 & n23931 ) | ( n15170 & ~n49552 ) | ( n23931 & ~n49552 ) ;
  assign n49554 = n18908 ^ n16252 ^ n7809 ;
  assign n49555 = ( n13816 & n15374 ) | ( n13816 & ~n49554 ) | ( n15374 & ~n49554 ) ;
  assign n49556 = n31325 ^ n13487 ^ n11136 ;
  assign n49557 = n19663 ^ n10046 ^ n7967 ;
  assign n49558 = n4832 & ~n39195 ;
  assign n49559 = n49558 ^ n30072 ^ n16965 ;
  assign n49560 = n20549 | n27643 ;
  assign n49561 = n49560 ^ n29672 ^ 1'b0 ;
  assign n49562 = ( n12990 & n14209 ) | ( n12990 & ~n14665 ) | ( n14209 & ~n14665 ) ;
  assign n49563 = n14852 & ~n46169 ;
  assign n49564 = n49563 ^ n8894 ^ 1'b0 ;
  assign n49565 = ( x97 & ~n23743 ) | ( x97 & n49564 ) | ( ~n23743 & n49564 ) ;
  assign n49566 = n49565 ^ n42290 ^ n28191 ;
  assign n49567 = ( n26374 & n36662 ) | ( n26374 & n49566 ) | ( n36662 & n49566 ) ;
  assign n49570 = n1348 & ~n21889 ;
  assign n49571 = n4771 & n49570 ;
  assign n49572 = n49571 ^ n17140 ^ n9290 ;
  assign n49568 = n16762 & ~n38199 ;
  assign n49569 = ~n1667 & n49568 ;
  assign n49573 = n49572 ^ n49569 ^ n6074 ;
  assign n49574 = n12978 ^ n970 ^ 1'b0 ;
  assign n49575 = n49574 ^ n26335 ^ n1659 ;
  assign n49576 = n49575 ^ n41922 ^ n10081 ;
  assign n49577 = ( ~n1673 & n26434 ) | ( ~n1673 & n45060 ) | ( n26434 & n45060 ) ;
  assign n49578 = ( n2378 & n5352 ) | ( n2378 & n9395 ) | ( n5352 & n9395 ) ;
  assign n49581 = n8291 ^ n5086 ^ 1'b0 ;
  assign n49579 = n38610 ^ n28042 ^ n24475 ;
  assign n49580 = n49579 ^ n25380 ^ n4376 ;
  assign n49582 = n49581 ^ n49580 ^ n31067 ;
  assign n49583 = n39062 ^ n26343 ^ n14774 ;
  assign n49584 = ( n9148 & n14104 ) | ( n9148 & ~n49583 ) | ( n14104 & ~n49583 ) ;
  assign n49585 = ( n10181 & ~n14061 ) | ( n10181 & n20051 ) | ( ~n14061 & n20051 ) ;
  assign n49586 = n49585 ^ n32517 ^ n32079 ;
  assign n49587 = n40346 & n49586 ;
  assign n49588 = n49587 ^ n23084 ^ 1'b0 ;
  assign n49589 = ~n3759 & n13729 ;
  assign n49590 = n49589 ^ n32018 ^ 1'b0 ;
  assign n49591 = n49590 ^ n14357 ^ n8228 ;
  assign n49592 = n8986 ^ n2385 ^ 1'b0 ;
  assign n49593 = ~n18732 & n43618 ;
  assign n49594 = n49593 ^ n42936 ^ 1'b0 ;
  assign n49595 = ( n7875 & ~n30335 ) | ( n7875 & n49594 ) | ( ~n30335 & n49594 ) ;
  assign n49596 = n49595 ^ n38778 ^ n1763 ;
  assign n49597 = ( n5105 & n34323 ) | ( n5105 & n45369 ) | ( n34323 & n45369 ) ;
  assign n49598 = ( n1015 & ~n19598 ) | ( n1015 & n49597 ) | ( ~n19598 & n49597 ) ;
  assign n49599 = n31250 ^ n7598 ^ n1712 ;
  assign n49600 = ( n12919 & n17780 ) | ( n12919 & n49599 ) | ( n17780 & n49599 ) ;
  assign n49601 = n41327 ^ n29954 ^ n20412 ;
  assign n49602 = n49601 ^ n40787 ^ n19459 ;
  assign n49603 = n2626 ^ n2036 ^ 1'b0 ;
  assign n49604 = ( n3695 & n44669 ) | ( n3695 & ~n45190 ) | ( n44669 & ~n45190 ) ;
  assign n49605 = ( n33890 & ~n49603 ) | ( n33890 & n49604 ) | ( ~n49603 & n49604 ) ;
  assign n49606 = n34453 ^ n5022 ^ n4045 ;
  assign n49607 = ( n10418 & n24550 ) | ( n10418 & n38227 ) | ( n24550 & n38227 ) ;
  assign n49608 = ( ~n33484 & n49606 ) | ( ~n33484 & n49607 ) | ( n49606 & n49607 ) ;
  assign n49609 = ( n2492 & n10248 ) | ( n2492 & ~n10869 ) | ( n10248 & ~n10869 ) ;
  assign n49610 = n49223 ^ n15993 ^ 1'b0 ;
  assign n49611 = n4064 & n49610 ;
  assign n49614 = n18603 ^ n1866 ^ 1'b0 ;
  assign n49615 = n49614 ^ n22472 ^ n16695 ;
  assign n49612 = ( n11781 & n18216 ) | ( n11781 & n39605 ) | ( n18216 & n39605 ) ;
  assign n49613 = ~n9965 & n49612 ;
  assign n49616 = n49615 ^ n49613 ^ 1'b0 ;
  assign n49617 = ( ~n3965 & n11210 ) | ( ~n3965 & n29978 ) | ( n11210 & n29978 ) ;
  assign n49618 = ( ~n6122 & n43464 ) | ( ~n6122 & n49617 ) | ( n43464 & n49617 ) ;
  assign n49619 = ( ~n7112 & n12421 ) | ( ~n7112 & n34078 ) | ( n12421 & n34078 ) ;
  assign n49620 = n19274 & n49619 ;
  assign n49621 = n13589 ^ n3512 ^ n1610 ;
  assign n49622 = ( n1358 & n19495 ) | ( n1358 & n28413 ) | ( n19495 & n28413 ) ;
  assign n49623 = n8482 ^ n2700 ^ 1'b0 ;
  assign n49624 = n49623 ^ n33460 ^ n18436 ;
  assign n49625 = ~n1547 & n7995 ;
  assign n49626 = ( n1494 & ~n42410 ) | ( n1494 & n49625 ) | ( ~n42410 & n49625 ) ;
  assign n49627 = n3528 & n43383 ;
  assign n49628 = n4368 & n49627 ;
  assign n49629 = ( n5703 & n9322 ) | ( n5703 & n49628 ) | ( n9322 & n49628 ) ;
  assign n49630 = n28268 ^ n17051 ^ 1'b0 ;
  assign n49631 = n49630 ^ n45019 ^ n29134 ;
  assign n49632 = ( n9435 & ~n12218 ) | ( n9435 & n15269 ) | ( ~n12218 & n15269 ) ;
  assign n49633 = ~n37798 & n49632 ;
  assign n49634 = ~n47649 & n49633 ;
  assign n49636 = n29850 ^ n26699 ^ n350 ;
  assign n49635 = n37203 & ~n49494 ;
  assign n49637 = n49636 ^ n49635 ^ 1'b0 ;
  assign n49638 = n49637 ^ n40250 ^ n1690 ;
  assign n49639 = ( n11795 & ~n14966 ) | ( n11795 & n23249 ) | ( ~n14966 & n23249 ) ;
  assign n49640 = n6177 & ~n35428 ;
  assign n49641 = n49640 ^ n33728 ^ 1'b0 ;
  assign n49642 = n49641 ^ n30570 ^ n19425 ;
  assign n49643 = ( ~n6655 & n17347 ) | ( ~n6655 & n19251 ) | ( n17347 & n19251 ) ;
  assign n49644 = ( n1574 & n49642 ) | ( n1574 & ~n49643 ) | ( n49642 & ~n49643 ) ;
  assign n49646 = ( n26585 & ~n37111 ) | ( n26585 & n43380 ) | ( ~n37111 & n43380 ) ;
  assign n49645 = ( n7030 & n24781 ) | ( n7030 & n30498 ) | ( n24781 & n30498 ) ;
  assign n49647 = n49646 ^ n49645 ^ n16351 ;
  assign n49648 = ( n19013 & n49644 ) | ( n19013 & n49647 ) | ( n49644 & n49647 ) ;
  assign n49649 = n16263 & ~n19484 ;
  assign n49650 = ( ~n33907 & n35249 ) | ( ~n33907 & n49649 ) | ( n35249 & n49649 ) ;
  assign n49651 = ( ~n10939 & n11560 ) | ( ~n10939 & n49650 ) | ( n11560 & n49650 ) ;
  assign n49653 = n7841 ^ n7605 ^ n2164 ;
  assign n49654 = n49653 ^ n24035 ^ n22666 ;
  assign n49652 = ( n3074 & n19184 ) | ( n3074 & n36497 ) | ( n19184 & n36497 ) ;
  assign n49655 = n49654 ^ n49652 ^ n18356 ;
  assign n49656 = n18432 ^ n15070 ^ n5583 ;
  assign n49657 = n47083 ^ n30527 ^ n4892 ;
  assign n49661 = n2400 & n3458 ;
  assign n49662 = ( n4472 & n27637 ) | ( n4472 & n49661 ) | ( n27637 & n49661 ) ;
  assign n49659 = n19754 ^ n4848 ^ n4147 ;
  assign n49660 = n35112 | n49659 ;
  assign n49658 = n13513 | n44684 ;
  assign n49663 = n49662 ^ n49660 ^ n49658 ;
  assign n49664 = n10068 ^ n7352 ^ 1'b0 ;
  assign n49665 = n2575 | n49664 ;
  assign n49666 = n28473 ^ n26949 ^ n19525 ;
  assign n49667 = ( n6875 & n35797 ) | ( n6875 & ~n49173 ) | ( n35797 & ~n49173 ) ;
  assign n49668 = ( n22861 & ~n37342 ) | ( n22861 & n49667 ) | ( ~n37342 & n49667 ) ;
  assign n49670 = n37610 ^ n21793 ^ n20314 ;
  assign n49669 = ( n13793 & n28582 ) | ( n13793 & n37729 ) | ( n28582 & n37729 ) ;
  assign n49671 = n49670 ^ n49669 ^ n7521 ;
  assign n49672 = ( ~n13487 & n15411 ) | ( ~n13487 & n27309 ) | ( n15411 & n27309 ) ;
  assign n49673 = ( n23644 & ~n26025 ) | ( n23644 & n27469 ) | ( ~n26025 & n27469 ) ;
  assign n49674 = n49673 ^ n47689 ^ n42995 ;
  assign n49675 = ( n8484 & n13897 ) | ( n8484 & ~n14451 ) | ( n13897 & ~n14451 ) ;
  assign n49676 = n40750 ^ n967 ^ x140 ;
  assign n49677 = ( ~n27974 & n49675 ) | ( ~n27974 & n49676 ) | ( n49675 & n49676 ) ;
  assign n49678 = n35447 ^ n15479 ^ n14381 ;
  assign n49679 = ( n3670 & ~n24756 ) | ( n3670 & n49678 ) | ( ~n24756 & n49678 ) ;
  assign n49680 = ( n7021 & n14837 ) | ( n7021 & n49679 ) | ( n14837 & n49679 ) ;
  assign n49681 = n28899 ^ n13036 ^ n1557 ;
  assign n49682 = n20447 | n27473 ;
  assign n49683 = n26369 | n49682 ;
  assign n49684 = n8420 | n9700 ;
  assign n49685 = n49684 ^ n35946 ^ 1'b0 ;
  assign n49686 = n25460 ^ n8829 ^ n8657 ;
  assign n49687 = ( x168 & n9171 ) | ( x168 & n10040 ) | ( n9171 & n10040 ) ;
  assign n49688 = n23529 ^ n4202 ^ 1'b0 ;
  assign n49689 = n49688 ^ n46749 ^ 1'b0 ;
  assign n49690 = n49687 & n49689 ;
  assign n49691 = n3588 | n4410 ;
  assign n49692 = ( n13155 & n41202 ) | ( n13155 & n42274 ) | ( n41202 & n42274 ) ;
  assign n49693 = ( ~n4293 & n44104 ) | ( ~n4293 & n49692 ) | ( n44104 & n49692 ) ;
  assign n49696 = ( n427 & n8166 ) | ( n427 & n19332 ) | ( n8166 & n19332 ) ;
  assign n49697 = ( ~n22490 & n22799 ) | ( ~n22490 & n49696 ) | ( n22799 & n49696 ) ;
  assign n49694 = ( n1586 & ~n1748 ) | ( n1586 & n6400 ) | ( ~n1748 & n6400 ) ;
  assign n49695 = n49694 ^ n15369 ^ n11682 ;
  assign n49698 = n49697 ^ n49695 ^ n1627 ;
  assign n49699 = ( ~n912 & n7542 ) | ( ~n912 & n44892 ) | ( n7542 & n44892 ) ;
  assign n49703 = n10779 & n19985 ;
  assign n49704 = n45410 & n49703 ;
  assign n49700 = n29701 ^ n19686 ^ n12537 ;
  assign n49701 = n49700 ^ n43666 ^ 1'b0 ;
  assign n49702 = n49701 ^ n36061 ^ n1822 ;
  assign n49705 = n49704 ^ n49702 ^ n24980 ;
  assign n49706 = n49705 ^ n1733 ^ n1622 ;
  assign n49708 = ( n4623 & n9233 ) | ( n4623 & n49704 ) | ( n9233 & n49704 ) ;
  assign n49709 = ( ~n1535 & n19586 ) | ( ~n1535 & n49708 ) | ( n19586 & n49708 ) ;
  assign n49707 = n22806 ^ n8879 ^ n2336 ;
  assign n49710 = n49709 ^ n49707 ^ n8597 ;
  assign n49711 = n17990 ^ n15394 ^ n10794 ;
  assign n49712 = n49711 ^ n20002 ^ n11704 ;
  assign n49713 = n4203 & ~n39006 ;
  assign n49714 = ~n49712 & n49713 ;
  assign n49715 = ( n21215 & ~n27915 ) | ( n21215 & n30523 ) | ( ~n27915 & n30523 ) ;
  assign n49716 = ( ~n10893 & n16855 ) | ( ~n10893 & n33056 ) | ( n16855 & n33056 ) ;
  assign n49717 = n49716 ^ n23722 ^ n3957 ;
  assign n49718 = n49717 ^ n7754 ^ 1'b0 ;
  assign n49719 = n26589 ^ n4436 ^ n2046 ;
  assign n49720 = n49719 ^ n26349 ^ n299 ;
  assign n49721 = ( n9351 & ~n17101 ) | ( n9351 & n40115 ) | ( ~n17101 & n40115 ) ;
  assign n49722 = ( n15586 & n18127 ) | ( n15586 & ~n24098 ) | ( n18127 & ~n24098 ) ;
  assign n49723 = n49722 ^ n13183 ^ n6780 ;
  assign n49724 = n49723 ^ n4205 ^ n2469 ;
  assign n49725 = n49724 ^ n27307 ^ n20192 ;
  assign n49726 = ~n9633 & n41521 ;
  assign n49727 = ( n2861 & n17062 ) | ( n2861 & ~n35358 ) | ( n17062 & ~n35358 ) ;
  assign n49728 = ( n10097 & n46407 ) | ( n10097 & ~n49727 ) | ( n46407 & ~n49727 ) ;
  assign n49729 = n10743 ^ x108 ^ 1'b0 ;
  assign n49730 = n13530 & n49729 ;
  assign n49731 = n49730 ^ n37818 ^ n4863 ;
  assign n49732 = ( n12315 & n12702 ) | ( n12315 & ~n29127 ) | ( n12702 & ~n29127 ) ;
  assign n49733 = n49732 ^ n22802 ^ x79 ;
  assign n49736 = ( n16629 & n34153 ) | ( n16629 & n38278 ) | ( n34153 & n38278 ) ;
  assign n49734 = n9873 ^ n6487 ^ n1722 ;
  assign n49735 = ~n1633 & n49734 ;
  assign n49737 = n49736 ^ n49735 ^ 1'b0 ;
  assign n49738 = n13460 & ~n41077 ;
  assign n49739 = n20461 ^ n16633 ^ 1'b0 ;
  assign n49740 = ( n2959 & n9717 ) | ( n2959 & n42896 ) | ( n9717 & n42896 ) ;
  assign n49741 = ( n29511 & n49739 ) | ( n29511 & n49740 ) | ( n49739 & n49740 ) ;
  assign n49742 = n49741 ^ n48030 ^ n1693 ;
  assign n49743 = n17683 ^ n9174 ^ n4390 ;
  assign n49744 = ( ~n2834 & n7000 ) | ( ~n2834 & n10485 ) | ( n7000 & n10485 ) ;
  assign n49745 = ( n992 & ~n49743 ) | ( n992 & n49744 ) | ( ~n49743 & n49744 ) ;
  assign n49746 = ( n21050 & ~n36450 ) | ( n21050 & n37610 ) | ( ~n36450 & n37610 ) ;
  assign n49747 = n49746 ^ n30535 ^ n9557 ;
  assign n49748 = ( n20875 & n29770 ) | ( n20875 & ~n33927 ) | ( n29770 & ~n33927 ) ;
  assign n49749 = ( n21013 & n49747 ) | ( n21013 & n49748 ) | ( n49747 & n49748 ) ;
  assign n49750 = n49749 ^ n43029 ^ n29489 ;
  assign n49751 = n39481 ^ n30699 ^ n13317 ;
  assign n49752 = ( n7152 & n22604 ) | ( n7152 & n36446 ) | ( n22604 & n36446 ) ;
  assign n49753 = ( n42941 & n47005 ) | ( n42941 & ~n49752 ) | ( n47005 & ~n49752 ) ;
  assign n49754 = n29786 ^ n26899 ^ n21700 ;
  assign n49755 = ( n508 & n15137 ) | ( n508 & ~n38952 ) | ( n15137 & ~n38952 ) ;
  assign n49756 = ~n12052 & n49755 ;
  assign n49757 = n29995 & n49756 ;
  assign n49758 = ~n46824 & n49757 ;
  assign n49760 = n49507 ^ n9372 ^ x116 ;
  assign n49759 = n12646 & n19590 ;
  assign n49761 = n49760 ^ n49759 ^ 1'b0 ;
  assign n49762 = ( n3019 & ~n4159 ) | ( n3019 & n19107 ) | ( ~n4159 & n19107 ) ;
  assign n49763 = ( ~n1596 & n11898 ) | ( ~n1596 & n15810 ) | ( n11898 & n15810 ) ;
  assign n49764 = n32565 ^ n25848 ^ n25277 ;
  assign n49765 = n29666 ^ n17125 ^ n7711 ;
  assign n49766 = ( ~n18123 & n44165 ) | ( ~n18123 & n49765 ) | ( n44165 & n49765 ) ;
  assign n49767 = ( n7877 & ~n10714 ) | ( n7877 & n30998 ) | ( ~n10714 & n30998 ) ;
  assign n49768 = ( n16746 & n26523 ) | ( n16746 & ~n31301 ) | ( n26523 & ~n31301 ) ;
  assign n49769 = ( ~n2218 & n21951 ) | ( ~n2218 & n33459 ) | ( n21951 & n33459 ) ;
  assign n49770 = ( n8161 & n24094 ) | ( n8161 & n37513 ) | ( n24094 & n37513 ) ;
  assign n49771 = n34541 ^ n13529 ^ n909 ;
  assign n49772 = n35165 & ~n39552 ;
  assign n49773 = n49772 ^ n12533 ^ 1'b0 ;
  assign n49774 = ( n5272 & ~n36067 ) | ( n5272 & n38326 ) | ( ~n36067 & n38326 ) ;
  assign n49775 = ( n14242 & n16495 ) | ( n14242 & ~n31640 ) | ( n16495 & ~n31640 ) ;
  assign n49776 = n49775 ^ n13007 ^ 1'b0 ;
  assign n49777 = ( n22827 & n25038 ) | ( n22827 & ~n49776 ) | ( n25038 & ~n49776 ) ;
  assign n49778 = n45751 ^ n40452 ^ n25574 ;
  assign n49779 = n49778 ^ n30509 ^ n8370 ;
  assign n49780 = n22395 & n25018 ;
  assign n49781 = n37683 & n49780 ;
  assign n49782 = ( n28984 & n43564 ) | ( n28984 & ~n49781 ) | ( n43564 & ~n49781 ) ;
  assign n49783 = n11135 & ~n33254 ;
  assign n49784 = ( ~n2617 & n39425 ) | ( ~n2617 & n49783 ) | ( n39425 & n49783 ) ;
  assign n49785 = n16106 ^ n5998 ^ n5298 ;
  assign n49786 = n49785 ^ n35711 ^ n3097 ;
  assign n49787 = ( n10969 & n11359 ) | ( n10969 & ~n38088 ) | ( n11359 & ~n38088 ) ;
  assign n49788 = n49787 ^ n18216 ^ n17857 ;
  assign n49789 = ( n14317 & ~n33127 ) | ( n14317 & n49788 ) | ( ~n33127 & n49788 ) ;
  assign n49790 = n28273 ^ n18925 ^ n18430 ;
  assign n49791 = n49790 ^ n25896 ^ n18129 ;
  assign n49792 = ( n12546 & n22002 ) | ( n12546 & ~n49791 ) | ( n22002 & ~n49791 ) ;
  assign n49793 = n24287 & n41327 ;
  assign n49794 = n19538 ^ n18972 ^ 1'b0 ;
  assign n49795 = ~n20528 & n49794 ;
  assign n49796 = n31068 ^ n7479 ^ 1'b0 ;
  assign n49797 = n49795 & ~n49796 ;
  assign n49798 = n40131 ^ n39706 ^ n9100 ;
  assign n49799 = ( n4579 & n6696 ) | ( n4579 & ~n49798 ) | ( n6696 & ~n49798 ) ;
  assign n49800 = ~n22932 & n44541 ;
  assign n49801 = ( n6128 & n13398 ) | ( n6128 & n41474 ) | ( n13398 & n41474 ) ;
  assign n49802 = n8830 & ~n10775 ;
  assign n49803 = n39216 & n49802 ;
  assign n49804 = n49803 ^ n22457 ^ n19475 ;
  assign n49805 = n49804 ^ n20800 ^ n4671 ;
  assign n49806 = n17761 & n29850 ;
  assign n49807 = ( n7959 & n12111 ) | ( n7959 & ~n16658 ) | ( n12111 & ~n16658 ) ;
  assign n49808 = n49807 ^ n45035 ^ n6807 ;
  assign n49809 = ( n9156 & ~n43464 ) | ( n9156 & n47313 ) | ( ~n43464 & n47313 ) ;
  assign n49811 = ( ~n5105 & n13630 ) | ( ~n5105 & n23385 ) | ( n13630 & n23385 ) ;
  assign n49812 = n49811 ^ n5411 ^ 1'b0 ;
  assign n49810 = ( n7823 & ~n10740 ) | ( n7823 & n46076 ) | ( ~n10740 & n46076 ) ;
  assign n49813 = n49812 ^ n49810 ^ n25030 ;
  assign n49814 = n49813 ^ n28696 ^ n26230 ;
  assign n49815 = ( n9411 & n20143 ) | ( n9411 & ~n32789 ) | ( n20143 & ~n32789 ) ;
  assign n49816 = n10933 & ~n31092 ;
  assign n49817 = ~n49815 & n49816 ;
  assign n49818 = n23943 ^ n3895 ^ 1'b0 ;
  assign n49819 = n13266 & ~n49818 ;
  assign n49820 = n26698 ^ n2972 ^ 1'b0 ;
  assign n49821 = n7645 | n49820 ;
  assign n49822 = n6825 & ~n49821 ;
  assign n49823 = n49822 ^ n25298 ^ 1'b0 ;
  assign n49824 = ( ~n28326 & n34631 ) | ( ~n28326 & n49823 ) | ( n34631 & n49823 ) ;
  assign n49825 = n34465 ^ n23066 ^ 1'b0 ;
  assign n49826 = n6978 & n49825 ;
  assign n49827 = ( n30113 & ~n42261 ) | ( n30113 & n49826 ) | ( ~n42261 & n49826 ) ;
  assign n49829 = ( n6964 & n13252 ) | ( n6964 & n29845 ) | ( n13252 & n29845 ) ;
  assign n49828 = n12288 & n42864 ;
  assign n49830 = n49829 ^ n49828 ^ 1'b0 ;
  assign n49831 = n49830 ^ n29813 ^ 1'b0 ;
  assign n49832 = ( ~n9831 & n18941 ) | ( ~n9831 & n49831 ) | ( n18941 & n49831 ) ;
  assign n49833 = n18101 & ~n19570 ;
  assign n49834 = n49833 ^ n40653 ^ n27981 ;
  assign n49835 = ( n1149 & n33446 ) | ( n1149 & ~n42759 ) | ( n33446 & ~n42759 ) ;
  assign n49836 = n49835 ^ n49702 ^ n10177 ;
  assign n49837 = n13147 & ~n25539 ;
  assign n49838 = n49837 ^ n32486 ^ n18309 ;
  assign n49839 = n13186 | n49838 ;
  assign n49840 = n33852 ^ n8014 ^ 1'b0 ;
  assign n49841 = n49840 ^ n47958 ^ n15488 ;
  assign n49842 = ( n28628 & ~n49839 ) | ( n28628 & n49841 ) | ( ~n49839 & n49841 ) ;
  assign n49843 = n41031 ^ n21996 ^ n20035 ;
  assign n49844 = n13435 & n26772 ;
  assign n49845 = n49469 ^ n45477 ^ n8027 ;
  assign n49846 = n21818 ^ n1384 ^ 1'b0 ;
  assign n49847 = n36771 ^ n22017 ^ n13819 ;
  assign n49848 = ( ~n21953 & n49846 ) | ( ~n21953 & n49847 ) | ( n49846 & n49847 ) ;
  assign n49849 = ~n1410 & n9303 ;
  assign n49850 = n49849 ^ n32808 ^ n23190 ;
  assign n49851 = ( ~n28745 & n44569 ) | ( ~n28745 & n49850 ) | ( n44569 & n49850 ) ;
  assign n49852 = n37495 ^ n23452 ^ n3972 ;
  assign n49853 = ( n1795 & n11520 ) | ( n1795 & ~n40108 ) | ( n11520 & ~n40108 ) ;
  assign n49854 = n9673 & n49853 ;
  assign n49855 = n45870 ^ n35261 ^ 1'b0 ;
  assign n49856 = ( n1707 & n4694 ) | ( n1707 & ~n41193 ) | ( n4694 & ~n41193 ) ;
  assign n49857 = ( n1540 & n3387 ) | ( n1540 & n13762 ) | ( n3387 & n13762 ) ;
  assign n49858 = ( n11177 & n14195 ) | ( n11177 & ~n49857 ) | ( n14195 & ~n49857 ) ;
  assign n49859 = n40705 ^ n8563 ^ n3780 ;
  assign n49860 = n34362 ^ n27928 ^ 1'b0 ;
  assign n49861 = n49860 ^ n43880 ^ n17726 ;
  assign n49862 = ( n6530 & n15189 ) | ( n6530 & n25678 ) | ( n15189 & n25678 ) ;
  assign n49863 = ( n32923 & ~n38577 ) | ( n32923 & n49862 ) | ( ~n38577 & n49862 ) ;
  assign n49864 = ( n388 & ~n2349 ) | ( n388 & n4965 ) | ( ~n2349 & n4965 ) ;
  assign n49865 = n18626 | n29488 ;
  assign n49866 = n22011 | n49865 ;
  assign n49867 = ( n15569 & n24501 ) | ( n15569 & n49866 ) | ( n24501 & n49866 ) ;
  assign n49868 = ( ~n12056 & n33238 ) | ( ~n12056 & n42846 ) | ( n33238 & n42846 ) ;
  assign n49869 = ( n16505 & n49867 ) | ( n16505 & ~n49868 ) | ( n49867 & ~n49868 ) ;
  assign n49870 = ( ~n15934 & n49864 ) | ( ~n15934 & n49869 ) | ( n49864 & n49869 ) ;
  assign n49871 = n49870 ^ n10178 ^ n6085 ;
  assign n49872 = n45724 ^ n37551 ^ n23419 ;
  assign n49873 = n38218 ^ n11530 ^ n2654 ;
  assign n49874 = ( n28546 & ~n29099 ) | ( n28546 & n44521 ) | ( ~n29099 & n44521 ) ;
  assign n49875 = n36713 ^ n21008 ^ n5749 ;
  assign n49876 = n49875 ^ n8080 ^ n2341 ;
  assign n49877 = ( n4157 & n9229 ) | ( n4157 & n40492 ) | ( n9229 & n40492 ) ;
  assign n49878 = n49877 ^ n10549 ^ n4640 ;
  assign n49879 = ( ~n43203 & n45569 ) | ( ~n43203 & n49878 ) | ( n45569 & n49878 ) ;
  assign n49880 = ( n16293 & ~n16991 ) | ( n16293 & n27570 ) | ( ~n16991 & n27570 ) ;
  assign n49881 = n49880 ^ n7461 ^ 1'b0 ;
  assign n49882 = n6567 & ~n49881 ;
  assign n49883 = n24092 ^ n18038 ^ 1'b0 ;
  assign n49884 = n4241 & n49883 ;
  assign n49885 = n49884 ^ n5759 ^ n2528 ;
  assign n49886 = n782 & ~n4562 ;
  assign n49887 = n49886 ^ n3739 ^ n343 ;
  assign n49888 = n31211 ^ n17963 ^ n7904 ;
  assign n49889 = n46171 ^ n17597 ^ n16732 ;
  assign n49890 = ( n9128 & n49888 ) | ( n9128 & ~n49889 ) | ( n49888 & ~n49889 ) ;
  assign n49891 = n26039 ^ n5274 ^ n3487 ;
  assign n49892 = n49891 ^ n36609 ^ 1'b0 ;
  assign n49893 = ( n10903 & n42868 ) | ( n10903 & ~n45049 ) | ( n42868 & ~n45049 ) ;
  assign n49895 = ( ~n8434 & n9832 ) | ( ~n8434 & n35410 ) | ( n9832 & n35410 ) ;
  assign n49896 = ( n11875 & n48483 ) | ( n11875 & n49895 ) | ( n48483 & n49895 ) ;
  assign n49897 = n49896 ^ n15974 ^ n13782 ;
  assign n49894 = n23348 | n48823 ;
  assign n49898 = n49897 ^ n49894 ^ n7088 ;
  assign n49899 = n45820 ^ n14357 ^ n4393 ;
  assign n49900 = ( ~n4449 & n8869 ) | ( ~n4449 & n49899 ) | ( n8869 & n49899 ) ;
  assign n49901 = ( n2598 & n38071 ) | ( n2598 & ~n49900 ) | ( n38071 & ~n49900 ) ;
  assign n49902 = n23182 ^ n11186 ^ n7244 ;
  assign n49909 = ( n903 & ~n5117 ) | ( n903 & n15845 ) | ( ~n5117 & n15845 ) ;
  assign n49910 = ( n13477 & n35955 ) | ( n13477 & n49909 ) | ( n35955 & n49909 ) ;
  assign n49912 = n28192 ^ n24403 ^ n2341 ;
  assign n49911 = ( n10307 & n12451 ) | ( n10307 & ~n22238 ) | ( n12451 & ~n22238 ) ;
  assign n49913 = n49912 ^ n49911 ^ n8658 ;
  assign n49914 = n49910 & ~n49913 ;
  assign n49903 = n32232 ^ n21341 ^ 1'b0 ;
  assign n49904 = n7694 & ~n49903 ;
  assign n49905 = ( ~n9932 & n31282 ) | ( ~n9932 & n49904 ) | ( n31282 & n49904 ) ;
  assign n49906 = n49905 ^ n9690 ^ n3110 ;
  assign n49907 = n39237 & n49906 ;
  assign n49908 = ~n10929 & n49907 ;
  assign n49915 = n49914 ^ n49908 ^ 1'b0 ;
  assign n49916 = n3050 & ~n21442 ;
  assign n49917 = n49916 ^ n2233 ^ 1'b0 ;
  assign n49918 = n40019 ^ n17479 ^ n17374 ;
  assign n49919 = ( n3819 & ~n42847 ) | ( n3819 & n49918 ) | ( ~n42847 & n49918 ) ;
  assign n49920 = n6563 & n49919 ;
  assign n49921 = n49920 ^ n35956 ^ n11441 ;
  assign n49922 = n49921 ^ n34080 ^ n32774 ;
  assign n49923 = n41501 ^ n1080 ^ n887 ;
  assign n49924 = n41967 ^ n14617 ^ n6650 ;
  assign n49925 = ( n8928 & n29778 ) | ( n8928 & ~n44048 ) | ( n29778 & ~n44048 ) ;
  assign n49926 = ( ~n16944 & n49924 ) | ( ~n16944 & n49925 ) | ( n49924 & n49925 ) ;
  assign n49927 = ~n4531 & n20451 ;
  assign n49928 = n49927 ^ n4113 ^ 1'b0 ;
  assign n49929 = ( n15810 & n37599 ) | ( n15810 & n49928 ) | ( n37599 & n49928 ) ;
  assign n49930 = n2774 & ~n8233 ;
  assign n49931 = ( n4774 & n6435 ) | ( n4774 & ~n9159 ) | ( n6435 & ~n9159 ) ;
  assign n49932 = ( n11932 & ~n15895 ) | ( n11932 & n21842 ) | ( ~n15895 & n21842 ) ;
  assign n49933 = ( n46902 & n49931 ) | ( n46902 & n49932 ) | ( n49931 & n49932 ) ;
  assign n49934 = n906 & ~n17075 ;
  assign n49935 = n49933 & n49934 ;
  assign n49936 = ( ~n3655 & n27130 ) | ( ~n3655 & n49935 ) | ( n27130 & n49935 ) ;
  assign n49938 = n15926 ^ n6528 ^ 1'b0 ;
  assign n49939 = n22482 & n49938 ;
  assign n49937 = n19513 ^ n17475 ^ n14401 ;
  assign n49940 = n49939 ^ n49937 ^ n23722 ;
  assign n49941 = ( n9318 & n12695 ) | ( n9318 & ~n17188 ) | ( n12695 & ~n17188 ) ;
  assign n49942 = ( n23231 & n42387 ) | ( n23231 & ~n49941 ) | ( n42387 & ~n49941 ) ;
  assign n49943 = n17348 ^ n16818 ^ n11661 ;
  assign n49944 = ( n327 & n10306 ) | ( n327 & ~n49943 ) | ( n10306 & ~n49943 ) ;
  assign n49945 = ~n3281 & n46566 ;
  assign n49946 = n49944 & n49945 ;
  assign n49947 = n15177 & ~n34642 ;
  assign n49948 = n49947 ^ n35303 ^ 1'b0 ;
  assign n49949 = n42883 ^ n9958 ^ 1'b0 ;
  assign n49950 = n2184 | n5648 ;
  assign n49951 = n38113 ^ n26701 ^ n9985 ;
  assign n49952 = n21323 | n47112 ;
  assign n49953 = n49952 ^ n4620 ^ 1'b0 ;
  assign n49954 = n49953 ^ n23052 ^ n7875 ;
  assign n49955 = n31868 ^ n26164 ^ n18706 ;
  assign n49956 = ( n2978 & n11714 ) | ( n2978 & ~n48926 ) | ( n11714 & ~n48926 ) ;
  assign n49957 = ( n10776 & n27307 ) | ( n10776 & ~n33064 ) | ( n27307 & ~n33064 ) ;
  assign n49958 = ( n7785 & n11745 ) | ( n7785 & ~n49957 ) | ( n11745 & ~n49957 ) ;
  assign n49959 = n41398 ^ n41104 ^ n7352 ;
  assign n49960 = n49331 ^ n33731 ^ n3474 ;
  assign n49961 = ( ~n19677 & n31299 ) | ( ~n19677 & n49960 ) | ( n31299 & n49960 ) ;
  assign n49962 = n38529 ^ n21602 ^ n2335 ;
  assign n49963 = ( n1762 & n49961 ) | ( n1762 & n49962 ) | ( n49961 & n49962 ) ;
  assign n49964 = n20952 ^ n5532 ^ n1309 ;
  assign n49965 = ( n1206 & n4426 ) | ( n1206 & ~n8601 ) | ( n4426 & ~n8601 ) ;
  assign n49966 = n49965 ^ n48322 ^ 1'b0 ;
  assign n49967 = n49964 & n49966 ;
  assign n49968 = n17359 ^ n11230 ^ n2840 ;
  assign n49969 = n49968 ^ n21166 ^ n12881 ;
  assign n49970 = n48407 ^ n47396 ^ n34283 ;
  assign n49971 = ( n6359 & n12513 ) | ( n6359 & ~n23178 ) | ( n12513 & ~n23178 ) ;
  assign n49972 = ( ~n14046 & n24067 ) | ( ~n14046 & n49971 ) | ( n24067 & n49971 ) ;
  assign n49973 = n38929 ^ n34771 ^ n4806 ;
  assign n49974 = ( n5179 & ~n17974 ) | ( n5179 & n47388 ) | ( ~n17974 & n47388 ) ;
  assign n49975 = n19974 ^ n12695 ^ 1'b0 ;
  assign n49976 = n49975 ^ n7495 ^ n3027 ;
  assign n49977 = n33542 ^ n21227 ^ n12162 ;
  assign n49978 = ( n1275 & n7452 ) | ( n1275 & ~n49977 ) | ( n7452 & ~n49977 ) ;
  assign n49979 = ( ~n18592 & n23065 ) | ( ~n18592 & n34153 ) | ( n23065 & n34153 ) ;
  assign n49980 = n49979 ^ n4876 ^ 1'b0 ;
  assign n49981 = n18450 | n49980 ;
  assign n49982 = n49981 ^ n39811 ^ n20326 ;
  assign n49983 = ( ~n13134 & n29711 ) | ( ~n13134 & n49982 ) | ( n29711 & n49982 ) ;
  assign n49984 = ( n20214 & ~n49978 ) | ( n20214 & n49983 ) | ( ~n49978 & n49983 ) ;
  assign n49985 = n45740 ^ n17091 ^ 1'b0 ;
  assign n49986 = n7896 & ~n49985 ;
  assign n49987 = n34962 ^ n8294 ^ n4091 ;
  assign n49988 = ( n2167 & ~n3082 ) | ( n2167 & n49987 ) | ( ~n3082 & n49987 ) ;
  assign n49989 = n49988 ^ n8162 ^ n1914 ;
  assign n49990 = n14808 ^ n9416 ^ n6904 ;
  assign n49991 = n49990 ^ n40724 ^ n15576 ;
  assign n49992 = ( n1320 & ~n10571 ) | ( n1320 & n32922 ) | ( ~n10571 & n32922 ) ;
  assign n49993 = ( n5794 & n23469 ) | ( n5794 & ~n33535 ) | ( n23469 & ~n33535 ) ;
  assign n49994 = ( n27491 & n30066 ) | ( n27491 & ~n49993 ) | ( n30066 & ~n49993 ) ;
  assign n49995 = n22739 ^ n21974 ^ 1'b0 ;
  assign n49996 = n49994 & ~n49995 ;
  assign n49997 = n49996 ^ n34223 ^ n3572 ;
  assign n49998 = ( n7543 & ~n49992 ) | ( n7543 & n49997 ) | ( ~n49992 & n49997 ) ;
  assign n49999 = ( n11568 & n30096 ) | ( n11568 & ~n38404 ) | ( n30096 & ~n38404 ) ;
  assign n50000 = ( n1265 & ~n43652 ) | ( n1265 & n47442 ) | ( ~n43652 & n47442 ) ;
  assign n50001 = n22106 ^ n18996 ^ n17461 ;
  assign n50002 = ( n6919 & ~n7443 ) | ( n6919 & n9650 ) | ( ~n7443 & n9650 ) ;
  assign n50003 = n50002 ^ n48485 ^ n31303 ;
  assign n50004 = n44311 ^ n17348 ^ n13541 ;
  assign n50005 = n50004 ^ n27046 ^ n4793 ;
  assign n50006 = n39169 ^ n29115 ^ 1'b0 ;
  assign n50007 = ~n1772 & n3146 ;
  assign n50008 = n50007 ^ n48108 ^ 1'b0 ;
  assign n50009 = n22871 ^ n21251 ^ n18889 ;
  assign n50010 = n5991 ^ n1377 ^ n1276 ;
  assign n50011 = n50010 ^ n35309 ^ n17888 ;
  assign n50012 = n33834 ^ n5957 ^ 1'b0 ;
  assign n50013 = ~n50011 & n50012 ;
  assign n50014 = n50013 ^ n21077 ^ n590 ;
  assign n50015 = ( ~n8912 & n50009 ) | ( ~n8912 & n50014 ) | ( n50009 & n50014 ) ;
  assign n50016 = ( n7720 & n36441 ) | ( n7720 & n49833 ) | ( n36441 & n49833 ) ;
  assign n50017 = ( ~n1291 & n6494 ) | ( ~n1291 & n22307 ) | ( n6494 & n22307 ) ;
  assign n50018 = n50017 ^ n37664 ^ n16704 ;
  assign n50019 = n44083 ^ n13526 ^ n8985 ;
  assign n50020 = n50019 ^ n44455 ^ 1'b0 ;
  assign n50025 = ~n4647 & n19158 ;
  assign n50026 = n50025 ^ n4704 ^ 1'b0 ;
  assign n50024 = ~n11557 & n13616 ;
  assign n50027 = n50026 ^ n50024 ^ n16966 ;
  assign n50021 = n22012 ^ n20651 ^ n19976 ;
  assign n50022 = n50021 ^ n38074 ^ n7442 ;
  assign n50023 = n50022 ^ n21985 ^ n14671 ;
  assign n50028 = n50027 ^ n50023 ^ n16524 ;
  assign n50032 = n17108 ^ n10661 ^ 1'b0 ;
  assign n50033 = n5571 | n50032 ;
  assign n50029 = ( n9251 & n31027 ) | ( n9251 & ~n39130 ) | ( n31027 & ~n39130 ) ;
  assign n50030 = ( n6695 & n12098 ) | ( n6695 & ~n50029 ) | ( n12098 & ~n50029 ) ;
  assign n50031 = n50030 ^ n11228 ^ n5550 ;
  assign n50034 = n50033 ^ n50031 ^ n31327 ;
  assign n50035 = n9819 & n47213 ;
  assign n50036 = ( n5966 & n19319 ) | ( n5966 & ~n50035 ) | ( n19319 & ~n50035 ) ;
  assign n50037 = n28588 ^ n27097 ^ n20048 ;
  assign n50038 = n50037 ^ n33150 ^ n1137 ;
  assign n50039 = ~n34118 & n47489 ;
  assign n50040 = n29956 & n50039 ;
  assign n50042 = n27863 & ~n30047 ;
  assign n50041 = ( n6193 & n32380 ) | ( n6193 & n33025 ) | ( n32380 & n33025 ) ;
  assign n50043 = n50042 ^ n50041 ^ n1408 ;
  assign n50044 = n13995 ^ n10820 ^ 1'b0 ;
  assign n50045 = ( ~n2441 & n43190 ) | ( ~n2441 & n50044 ) | ( n43190 & n50044 ) ;
  assign n50046 = ( n6010 & ~n8358 ) | ( n6010 & n18690 ) | ( ~n8358 & n18690 ) ;
  assign n50047 = n46202 ^ n37202 ^ n13927 ;
  assign n50048 = n11815 & n33040 ;
  assign n50049 = ~n8515 & n50048 ;
  assign n50050 = ( ~n35077 & n36559 ) | ( ~n35077 & n50049 ) | ( n36559 & n50049 ) ;
  assign n50051 = n50050 ^ n949 ^ 1'b0 ;
  assign n50052 = ( ~n14829 & n28447 ) | ( ~n14829 & n31086 ) | ( n28447 & n31086 ) ;
  assign n50053 = ( n8785 & ~n19267 ) | ( n8785 & n21856 ) | ( ~n19267 & n21856 ) ;
  assign n50054 = n33732 ^ n18088 ^ n8807 ;
  assign n50055 = ( n10595 & ~n50053 ) | ( n10595 & n50054 ) | ( ~n50053 & n50054 ) ;
  assign n50056 = n41419 ^ n24555 ^ n10202 ;
  assign n50057 = n50056 ^ n40380 ^ n22318 ;
  assign n50059 = n39737 ^ n9786 ^ n7825 ;
  assign n50058 = n17858 & n24191 ;
  assign n50060 = n50059 ^ n50058 ^ 1'b0 ;
  assign n50061 = n24566 ^ n7918 ^ n7624 ;
  assign n50062 = n50061 ^ n30848 ^ n29288 ;
  assign n50063 = n33875 ^ n13556 ^ 1'b0 ;
  assign n50064 = n14659 | n50063 ;
  assign n50065 = ( n10621 & n27462 ) | ( n10621 & ~n50064 ) | ( n27462 & ~n50064 ) ;
  assign n50066 = ( n20986 & ~n39419 ) | ( n20986 & n45750 ) | ( ~n39419 & n45750 ) ;
  assign n50067 = n42917 ^ n13567 ^ n9480 ;
  assign n50068 = ( n3559 & n20154 ) | ( n3559 & ~n45081 ) | ( n20154 & ~n45081 ) ;
  assign n50069 = ( n2376 & n43025 ) | ( n2376 & ~n50068 ) | ( n43025 & ~n50068 ) ;
  assign n50070 = ( n48568 & n50067 ) | ( n48568 & ~n50069 ) | ( n50067 & ~n50069 ) ;
  assign n50071 = n40996 ^ n26035 ^ 1'b0 ;
  assign n50072 = n35337 ^ n20716 ^ n14920 ;
  assign n50073 = n50072 ^ n21992 ^ n12098 ;
  assign n50077 = n13750 ^ n10199 ^ n9625 ;
  assign n50074 = ( ~n7815 & n17199 ) | ( ~n7815 & n22429 ) | ( n17199 & n22429 ) ;
  assign n50075 = n31989 ^ n18325 ^ n16095 ;
  assign n50076 = ( ~n15141 & n50074 ) | ( ~n15141 & n50075 ) | ( n50074 & n50075 ) ;
  assign n50078 = n50077 ^ n50076 ^ n27690 ;
  assign n50080 = n32584 ^ n20186 ^ n16329 ;
  assign n50079 = n38364 ^ n17205 ^ 1'b0 ;
  assign n50081 = n50080 ^ n50079 ^ n19918 ;
  assign n50082 = n5813 & n11208 ;
  assign n50083 = ~n16463 & n43820 ;
  assign n50084 = n50083 ^ n13133 ^ 1'b0 ;
  assign n50085 = n18444 & ~n39762 ;
  assign n50086 = n50085 ^ n33732 ^ 1'b0 ;
  assign n50087 = ~n29028 & n41463 ;
  assign n50088 = ( n12628 & n28583 ) | ( n12628 & ~n46170 ) | ( n28583 & ~n46170 ) ;
  assign n50089 = n46501 | n48839 ;
  assign n50094 = ( n22978 & n34988 ) | ( n22978 & ~n38932 ) | ( n34988 & ~n38932 ) ;
  assign n50090 = n3954 & ~n28434 ;
  assign n50091 = n50090 ^ n31653 ^ 1'b0 ;
  assign n50092 = n50091 ^ n6595 ^ n3621 ;
  assign n50093 = ( n1333 & n12639 ) | ( n1333 & ~n50092 ) | ( n12639 & ~n50092 ) ;
  assign n50095 = n50094 ^ n50093 ^ n15237 ;
  assign n50096 = ( ~n25062 & n32803 ) | ( ~n25062 & n41240 ) | ( n32803 & n41240 ) ;
  assign n50097 = n50096 ^ n47521 ^ n14403 ;
  assign n50098 = ( n13064 & n30508 ) | ( n13064 & ~n35835 ) | ( n30508 & ~n35835 ) ;
  assign n50099 = ( n17480 & n30134 ) | ( n17480 & ~n50098 ) | ( n30134 & ~n50098 ) ;
  assign n50100 = n1537 & ~n11649 ;
  assign n50101 = ~n11291 & n39747 ;
  assign n50102 = n35947 & n50101 ;
  assign n50103 = ( n10902 & n13387 ) | ( n10902 & ~n30436 ) | ( n13387 & ~n30436 ) ;
  assign n50104 = ( ~n1802 & n2045 ) | ( ~n1802 & n11204 ) | ( n2045 & n11204 ) ;
  assign n50105 = ( n7466 & n19790 ) | ( n7466 & n50104 ) | ( n19790 & n50104 ) ;
  assign n50106 = n31489 & n50105 ;
  assign n50107 = n2609 | n50106 ;
  assign n50108 = n50103 | n50107 ;
  assign n50109 = n22312 ^ n11354 ^ 1'b0 ;
  assign n50110 = n50109 ^ n49621 ^ 1'b0 ;
  assign n50112 = ( n6966 & ~n12415 ) | ( n6966 & n19329 ) | ( ~n12415 & n19329 ) ;
  assign n50113 = n29960 ^ n14387 ^ n10005 ;
  assign n50114 = n24004 ^ n22545 ^ n11477 ;
  assign n50115 = n50114 ^ n40163 ^ n38059 ;
  assign n50116 = ( n50112 & n50113 ) | ( n50112 & n50115 ) | ( n50113 & n50115 ) ;
  assign n50111 = ( n24291 & n29367 ) | ( n24291 & n33545 ) | ( n29367 & n33545 ) ;
  assign n50117 = n50116 ^ n50111 ^ 1'b0 ;
  assign n50118 = ( n5546 & n9021 ) | ( n5546 & ~n20699 ) | ( n9021 & ~n20699 ) ;
  assign n50119 = ( n6029 & n16762 ) | ( n6029 & ~n50118 ) | ( n16762 & ~n50118 ) ;
  assign n50120 = n43861 ^ n2744 ^ n1584 ;
  assign n50121 = n25630 ^ n1430 ^ n1348 ;
  assign n50122 = ( n8286 & n10598 ) | ( n8286 & n38332 ) | ( n10598 & n38332 ) ;
  assign n50123 = n31270 ^ n17983 ^ n17245 ;
  assign n50124 = n33583 ^ n30281 ^ n24150 ;
  assign n50125 = ( n642 & n11907 ) | ( n642 & ~n43880 ) | ( n11907 & ~n43880 ) ;
  assign n50126 = ( ~n19100 & n50124 ) | ( ~n19100 & n50125 ) | ( n50124 & n50125 ) ;
  assign n50127 = ( n3404 & n16131 ) | ( n3404 & n34063 ) | ( n16131 & n34063 ) ;
  assign n50128 = ( n2824 & n11095 ) | ( n2824 & ~n50127 ) | ( n11095 & ~n50127 ) ;
  assign n50129 = ( x104 & n40874 ) | ( x104 & n50128 ) | ( n40874 & n50128 ) ;
  assign n50130 = n44755 ^ n15401 ^ n7371 ;
  assign n50131 = n29385 & ~n50130 ;
  assign n50132 = n50131 ^ n11139 ^ 1'b0 ;
  assign n50133 = n48935 ^ n43065 ^ n25724 ;
  assign n50134 = n14632 ^ n2935 ^ 1'b0 ;
  assign n50135 = n4549 & ~n50134 ;
  assign n50136 = ( n4648 & n13434 ) | ( n4648 & n50135 ) | ( n13434 & n50135 ) ;
  assign n50137 = ( n26217 & n41979 ) | ( n26217 & ~n44919 ) | ( n41979 & ~n44919 ) ;
  assign n50138 = n20782 ^ n4224 ^ n2478 ;
  assign n50139 = n11347 ^ n8149 ^ n1881 ;
  assign n50140 = n50139 ^ n13816 ^ n3123 ;
  assign n50141 = n50140 ^ n21696 ^ n8489 ;
  assign n50142 = n50141 ^ n2264 ^ 1'b0 ;
  assign n50143 = n50138 & n50142 ;
  assign n50144 = ( n3645 & n33485 ) | ( n3645 & n50143 ) | ( n33485 & n50143 ) ;
  assign n50145 = n2598 & n6248 ;
  assign n50146 = n29231 & n50145 ;
  assign n50147 = n50146 ^ n32095 ^ n15051 ;
  assign n50148 = ( n15103 & ~n21789 ) | ( n15103 & n50147 ) | ( ~n21789 & n50147 ) ;
  assign n50149 = n5134 | n23654 ;
  assign n50150 = n50149 ^ n20593 ^ 1'b0 ;
  assign n50151 = n50150 ^ n46038 ^ n19942 ;
  assign n50157 = n37606 ^ n20608 ^ 1'b0 ;
  assign n50152 = ~n15921 & n23506 ;
  assign n50153 = n28250 ^ n26306 ^ n8923 ;
  assign n50154 = ( n17519 & n50152 ) | ( n17519 & n50153 ) | ( n50152 & n50153 ) ;
  assign n50155 = n5557 & ~n50154 ;
  assign n50156 = n44746 & n50155 ;
  assign n50158 = n50157 ^ n50156 ^ n9021 ;
  assign n50159 = n13561 & n16156 ;
  assign n50160 = n11074 & n50159 ;
  assign n50161 = ( x138 & ~n22244 ) | ( x138 & n42406 ) | ( ~n22244 & n42406 ) ;
  assign n50162 = ( n7717 & n19341 ) | ( n7717 & n42781 ) | ( n19341 & n42781 ) ;
  assign n50163 = n50162 ^ n34736 ^ n384 ;
  assign n50164 = ( n27861 & n30860 ) | ( n27861 & ~n48773 ) | ( n30860 & ~n48773 ) ;
  assign n50165 = n30700 ^ n17653 ^ n16225 ;
  assign n50166 = ( ~n9594 & n22928 ) | ( ~n9594 & n50165 ) | ( n22928 & n50165 ) ;
  assign n50167 = n47714 ^ n38028 ^ n18784 ;
  assign n50168 = n50167 ^ n47601 ^ 1'b0 ;
  assign n50169 = n23182 ^ n6243 ^ 1'b0 ;
  assign n50170 = ~n21458 & n50169 ;
  assign n50171 = n50170 ^ n26453 ^ n19353 ;
  assign n50172 = n50171 ^ n8004 ^ 1'b0 ;
  assign n50173 = n17237 ^ n8467 ^ 1'b0 ;
  assign n50174 = ~n1354 & n50173 ;
  assign n50175 = n50174 ^ n21399 ^ n20073 ;
  assign n50176 = ( n10953 & ~n49833 ) | ( n10953 & n50175 ) | ( ~n49833 & n50175 ) ;
  assign n50177 = n48089 ^ n31825 ^ n1523 ;
  assign n50178 = n43113 ^ n35433 ^ n1662 ;
  assign n50179 = n50178 ^ n29978 ^ 1'b0 ;
  assign n50180 = ( n5949 & ~n45007 ) | ( n5949 & n50179 ) | ( ~n45007 & n50179 ) ;
  assign n50181 = n32474 & n50180 ;
  assign n50182 = ~n19450 & n50181 ;
  assign n50183 = n23643 ^ n22681 ^ n6092 ;
  assign n50184 = ~n5412 & n28495 ;
  assign n50185 = ~n10464 & n50184 ;
  assign n50186 = n11923 ^ n6289 ^ 1'b0 ;
  assign n50187 = n12256 ^ n12078 ^ 1'b0 ;
  assign n50188 = ( ~n50185 & n50186 ) | ( ~n50185 & n50187 ) | ( n50186 & n50187 ) ;
  assign n50189 = ( ~n4058 & n18981 ) | ( ~n4058 & n24018 ) | ( n18981 & n24018 ) ;
  assign n50190 = n50189 ^ n32875 ^ n19408 ;
  assign n50191 = ( n33664 & ~n37051 ) | ( n33664 & n43235 ) | ( ~n37051 & n43235 ) ;
  assign n50192 = ( n513 & ~n46046 ) | ( n513 & n50191 ) | ( ~n46046 & n50191 ) ;
  assign n50193 = n47333 ^ n24277 ^ n1261 ;
  assign n50194 = n40215 ^ n18686 ^ n17486 ;
  assign n50195 = n31395 ^ n7734 ^ n4342 ;
  assign n50196 = ( n21635 & n30483 ) | ( n21635 & n50195 ) | ( n30483 & n50195 ) ;
  assign n50197 = ( n2832 & ~n22142 ) | ( n2832 & n50196 ) | ( ~n22142 & n50196 ) ;
  assign n50199 = n16170 ^ n14794 ^ n2219 ;
  assign n50200 = ( n6287 & ~n17201 ) | ( n6287 & n50199 ) | ( ~n17201 & n50199 ) ;
  assign n50201 = n50200 ^ n33926 ^ 1'b0 ;
  assign n50198 = n17869 | n30383 ;
  assign n50202 = n50201 ^ n50198 ^ 1'b0 ;
  assign n50203 = ( n1204 & ~n7658 ) | ( n1204 & n15137 ) | ( ~n7658 & n15137 ) ;
  assign n50204 = n39697 ^ n23924 ^ n20236 ;
  assign n50205 = ( n806 & n32577 ) | ( n806 & ~n44107 ) | ( n32577 & ~n44107 ) ;
  assign n50206 = n10810 | n22791 ;
  assign n50207 = n50206 ^ n37623 ^ n865 ;
  assign n50208 = n35420 ^ x25 ^ 1'b0 ;
  assign n50209 = ( ~n11959 & n18023 ) | ( ~n11959 & n37818 ) | ( n18023 & n37818 ) ;
  assign n50210 = n6188 ^ n1324 ^ 1'b0 ;
  assign n50211 = n30750 ^ n27104 ^ n14183 ;
  assign n50212 = ( n3114 & ~n27085 ) | ( n3114 & n50211 ) | ( ~n27085 & n50211 ) ;
  assign n50213 = n50212 ^ n49834 ^ 1'b0 ;
  assign n50214 = n6546 & n50213 ;
  assign n50215 = n17624 ^ n14562 ^ 1'b0 ;
  assign n50216 = n18537 & ~n50215 ;
  assign n50217 = n24721 | n25074 ;
  assign n50218 = n50216 | n50217 ;
  assign n50219 = ( ~n23145 & n30957 ) | ( ~n23145 & n33065 ) | ( n30957 & n33065 ) ;
  assign n50220 = ( n6866 & n16977 ) | ( n6866 & ~n35846 ) | ( n16977 & ~n35846 ) ;
  assign n50221 = n598 & ~n23143 ;
  assign n50222 = ( n4724 & ~n35264 ) | ( n4724 & n50221 ) | ( ~n35264 & n50221 ) ;
  assign n50223 = ( n26682 & n50220 ) | ( n26682 & ~n50222 ) | ( n50220 & ~n50222 ) ;
  assign n50224 = ( ~n8356 & n19537 ) | ( ~n8356 & n43691 ) | ( n19537 & n43691 ) ;
  assign n50225 = ~n39320 & n44534 ;
  assign n50226 = n10770 & n50225 ;
  assign n50227 = n50226 ^ n47865 ^ n31998 ;
  assign n50228 = ( n5330 & n50224 ) | ( n5330 & ~n50227 ) | ( n50224 & ~n50227 ) ;
  assign n50229 = n24473 ^ n4366 ^ 1'b0 ;
  assign n50230 = n27195 | n50229 ;
  assign n50231 = ( n7395 & n42729 ) | ( n7395 & ~n50230 ) | ( n42729 & ~n50230 ) ;
  assign n50232 = ( n18086 & ~n19356 ) | ( n18086 & n47816 ) | ( ~n19356 & n47816 ) ;
  assign n50233 = ( ~n11817 & n35726 ) | ( ~n11817 & n50232 ) | ( n35726 & n50232 ) ;
  assign n50234 = n11449 & n14907 ;
  assign n50235 = n50234 ^ n25257 ^ 1'b0 ;
  assign n50236 = n16468 ^ n7434 ^ n713 ;
  assign n50237 = n46744 & n50236 ;
  assign n50238 = ( n17480 & n50235 ) | ( n17480 & ~n50237 ) | ( n50235 & ~n50237 ) ;
  assign n50239 = n16607 ^ n14689 ^ n9494 ;
  assign n50240 = n37385 ^ n8940 ^ n4629 ;
  assign n50241 = ( n8849 & n38800 ) | ( n8849 & ~n50240 ) | ( n38800 & ~n50240 ) ;
  assign n50242 = n4274 & n4835 ;
  assign n50243 = ( n15293 & ~n25704 ) | ( n15293 & n50242 ) | ( ~n25704 & n50242 ) ;
  assign n50244 = ( n24897 & ~n28226 ) | ( n24897 & n50243 ) | ( ~n28226 & n50243 ) ;
  assign n50245 = n16115 ^ n8910 ^ 1'b0 ;
  assign n50246 = n50244 & n50245 ;
  assign n50247 = n4551 & n18529 ;
  assign n50248 = ( n7388 & ~n19721 ) | ( n7388 & n21101 ) | ( ~n19721 & n21101 ) ;
  assign n50249 = ( n5432 & n50247 ) | ( n5432 & ~n50248 ) | ( n50247 & ~n50248 ) ;
  assign n50250 = n30199 ^ n13063 ^ n3511 ;
  assign n50251 = ( n10551 & n20892 ) | ( n10551 & n36906 ) | ( n20892 & n36906 ) ;
  assign n50252 = n28764 & ~n42333 ;
  assign n50253 = ~n36605 & n50252 ;
  assign n50254 = n50253 ^ n39679 ^ n22936 ;
  assign n50255 = n8673 | n35732 ;
  assign n50256 = n50255 ^ n30006 ^ 1'b0 ;
  assign n50257 = ( n1611 & ~n21337 ) | ( n1611 & n39765 ) | ( ~n21337 & n39765 ) ;
  assign n50258 = n31296 & n50257 ;
  assign n50259 = n25609 | n50258 ;
  assign n50260 = n50259 ^ n19316 ^ 1'b0 ;
  assign n50261 = n50256 | n50260 ;
  assign n50262 = n31779 ^ n4748 ^ 1'b0 ;
  assign n50264 = n2980 ^ n2840 ^ n1175 ;
  assign n50265 = ( n8686 & n11482 ) | ( n8686 & ~n50264 ) | ( n11482 & ~n50264 ) ;
  assign n50263 = n44838 ^ n35764 ^ n11283 ;
  assign n50266 = n50265 ^ n50263 ^ n48880 ;
  assign n50267 = n22861 ^ n14483 ^ 1'b0 ;
  assign n50268 = n23174 ^ n14868 ^ n4605 ;
  assign n50269 = n8433 & n50268 ;
  assign n50270 = ( n3878 & ~n24807 ) | ( n3878 & n25871 ) | ( ~n24807 & n25871 ) ;
  assign n50271 = n50270 ^ n38305 ^ n19509 ;
  assign n50272 = n25129 ^ n17147 ^ n14355 ;
  assign n50273 = ( n17953 & n46506 ) | ( n17953 & ~n50272 ) | ( n46506 & ~n50272 ) ;
  assign n50274 = n14261 ^ n12397 ^ 1'b0 ;
  assign n50275 = ( n3000 & n22319 ) | ( n3000 & ~n41067 ) | ( n22319 & ~n41067 ) ;
  assign n50276 = n45917 ^ n42640 ^ n36152 ;
  assign n50278 = ( ~n9265 & n17199 ) | ( ~n9265 & n35329 ) | ( n17199 & n35329 ) ;
  assign n50277 = n43780 ^ n9263 ^ n6747 ;
  assign n50279 = n50278 ^ n50277 ^ n28328 ;
  assign n50280 = ( ~n29424 & n41057 ) | ( ~n29424 & n50279 ) | ( n41057 & n50279 ) ;
  assign n50281 = n28250 ^ n12326 ^ n3181 ;
  assign n50282 = n50281 ^ n25458 ^ 1'b0 ;
  assign n50283 = n33782 ^ n30897 ^ 1'b0 ;
  assign n50284 = ( n47757 & n50282 ) | ( n47757 & n50283 ) | ( n50282 & n50283 ) ;
  assign n50285 = n30554 ^ n28997 ^ n294 ;
  assign n50286 = n50285 ^ n49354 ^ n19425 ;
  assign n50287 = n37746 ^ n33021 ^ n14381 ;
  assign n50288 = n50287 ^ n31676 ^ n16840 ;
  assign n50289 = n50288 ^ n38095 ^ n28361 ;
  assign n50290 = ( x165 & ~n5290 ) | ( x165 & n28929 ) | ( ~n5290 & n28929 ) ;
  assign n50291 = ( n2515 & ~n3878 ) | ( n2515 & n10843 ) | ( ~n3878 & n10843 ) ;
  assign n50293 = ( ~n2515 & n13718 ) | ( ~n2515 & n43029 ) | ( n13718 & n43029 ) ;
  assign n50294 = ( ~n378 & n31979 ) | ( ~n378 & n50293 ) | ( n31979 & n50293 ) ;
  assign n50292 = ( n1712 & n4447 ) | ( n1712 & n47523 ) | ( n4447 & n47523 ) ;
  assign n50295 = n50294 ^ n50292 ^ n39447 ;
  assign n50296 = n47396 ^ n3594 ^ 1'b0 ;
  assign n50297 = ( n25941 & ~n40194 ) | ( n25941 & n47735 ) | ( ~n40194 & n47735 ) ;
  assign n50298 = ( n6250 & ~n33647 ) | ( n6250 & n36100 ) | ( ~n33647 & n36100 ) ;
  assign n50299 = ( n7696 & n19220 ) | ( n7696 & n50298 ) | ( n19220 & n50298 ) ;
  assign n50300 = n14450 & n19792 ;
  assign n50301 = ~n5255 & n50300 ;
  assign n50302 = n38235 ^ n17053 ^ n5159 ;
  assign n50303 = ( n13589 & ~n21413 ) | ( n13589 & n44686 ) | ( ~n21413 & n44686 ) ;
  assign n50304 = n6886 | n20235 ;
  assign n50305 = ( n13391 & ~n13999 ) | ( n13391 & n50304 ) | ( ~n13999 & n50304 ) ;
  assign n50308 = ~n21950 & n26378 ;
  assign n50309 = n50308 ^ n28043 ^ 1'b0 ;
  assign n50306 = n32837 ^ n19491 ^ n14094 ;
  assign n50307 = ( n7011 & n26717 ) | ( n7011 & ~n50306 ) | ( n26717 & ~n50306 ) ;
  assign n50310 = n50309 ^ n50307 ^ 1'b0 ;
  assign n50311 = n34171 ^ n14758 ^ n12936 ;
  assign n50312 = ( n1256 & ~n6926 ) | ( n1256 & n14178 ) | ( ~n6926 & n14178 ) ;
  assign n50313 = n50312 ^ n46033 ^ n3268 ;
  assign n50314 = n15212 ^ n5766 ^ n3621 ;
  assign n50315 = n16808 ^ n16104 ^ n12037 ;
  assign n50316 = n37342 ^ n24746 ^ n18041 ;
  assign n50317 = ( n14017 & n50315 ) | ( n14017 & n50316 ) | ( n50315 & n50316 ) ;
  assign n50318 = ( x114 & n10519 ) | ( x114 & n25656 ) | ( n10519 & n25656 ) ;
  assign n50319 = ~n2712 & n14362 ;
  assign n50320 = n50319 ^ n4115 ^ 1'b0 ;
  assign n50321 = n936 & ~n24611 ;
  assign n50322 = n39925 & n50321 ;
  assign n50323 = n50322 ^ n19238 ^ 1'b0 ;
  assign n50324 = n41856 ^ n30881 ^ n30221 ;
  assign n50325 = n9404 ^ n5818 ^ n1365 ;
  assign n50326 = ( n7794 & n13726 ) | ( n7794 & ~n18390 ) | ( n13726 & ~n18390 ) ;
  assign n50327 = n50326 ^ n22844 ^ n15889 ;
  assign n50328 = ( ~n31607 & n50325 ) | ( ~n31607 & n50327 ) | ( n50325 & n50327 ) ;
  assign n50329 = n38005 ^ n29370 ^ n3815 ;
  assign n50330 = n50329 ^ n3116 ^ x230 ;
  assign n50331 = n16702 ^ n4694 ^ 1'b0 ;
  assign n50332 = ( n3045 & n12797 ) | ( n3045 & n23741 ) | ( n12797 & n23741 ) ;
  assign n50333 = n50332 ^ n35587 ^ n14214 ;
  assign n50334 = ( n32507 & n43875 ) | ( n32507 & n50333 ) | ( n43875 & n50333 ) ;
  assign n50335 = n50334 ^ n12977 ^ 1'b0 ;
  assign n50336 = n6921 ^ n5737 ^ n1701 ;
  assign n50337 = ( n8982 & n12888 ) | ( n8982 & ~n50336 ) | ( n12888 & ~n50336 ) ;
  assign n50338 = n46716 ^ n25856 ^ n16687 ;
  assign n50339 = ( ~n11806 & n13736 ) | ( ~n11806 & n50338 ) | ( n13736 & n50338 ) ;
  assign n50340 = ( ~n2703 & n6413 ) | ( ~n2703 & n12587 ) | ( n6413 & n12587 ) ;
  assign n50341 = n20787 & n50340 ;
  assign n50342 = ( n2927 & n4359 ) | ( n2927 & ~n5220 ) | ( n4359 & ~n5220 ) ;
  assign n50343 = n14509 ^ n1636 ^ 1'b0 ;
  assign n50344 = n50342 & n50343 ;
  assign n50345 = n48043 ^ n41574 ^ n12541 ;
  assign n50346 = n50345 ^ n36005 ^ n21958 ;
  assign n50347 = ( n18052 & n18294 ) | ( n18052 & n22618 ) | ( n18294 & n22618 ) ;
  assign n50348 = ( n3731 & n4041 ) | ( n3731 & ~n14012 ) | ( n4041 & ~n14012 ) ;
  assign n50349 = n22042 ^ n9665 ^ n8330 ;
  assign n50350 = ( x43 & n13360 ) | ( x43 & ~n22820 ) | ( n13360 & ~n22820 ) ;
  assign n50351 = ( n25540 & n50349 ) | ( n25540 & ~n50350 ) | ( n50349 & ~n50350 ) ;
  assign n50352 = n46828 ^ n8286 ^ 1'b0 ;
  assign n50353 = ( ~n5074 & n25007 ) | ( ~n5074 & n50352 ) | ( n25007 & n50352 ) ;
  assign n50354 = n19295 ^ n12403 ^ n7736 ;
  assign n50355 = n50354 ^ n14507 ^ n11092 ;
  assign n50356 = n24643 ^ n18116 ^ n13040 ;
  assign n50357 = ( ~n15007 & n16417 ) | ( ~n15007 & n50356 ) | ( n16417 & n50356 ) ;
  assign n50358 = ( ~n20140 & n50355 ) | ( ~n20140 & n50357 ) | ( n50355 & n50357 ) ;
  assign n50359 = n17889 & ~n19347 ;
  assign n50360 = n50359 ^ n7500 ^ n1711 ;
  assign n50361 = n19806 ^ n679 ^ 1'b0 ;
  assign n50362 = ~n34428 & n50361 ;
  assign n50363 = n44028 ^ n16250 ^ n1877 ;
  assign n50364 = n50363 ^ n36759 ^ n6520 ;
  assign n50365 = n28418 ^ n22669 ^ n7459 ;
  assign n50366 = ( n10675 & n12744 ) | ( n10675 & ~n32837 ) | ( n12744 & ~n32837 ) ;
  assign n50367 = n50366 ^ n39500 ^ n29694 ;
  assign n50368 = n42045 ^ n23280 ^ 1'b0 ;
  assign n50369 = ( x212 & n9535 ) | ( x212 & ~n33559 ) | ( n9535 & ~n33559 ) ;
  assign n50370 = n44759 ^ n23974 ^ n20532 ;
  assign n50371 = n50370 ^ n18218 ^ n2239 ;
  assign n50372 = n50371 ^ n12755 ^ x106 ;
  assign n50373 = ( ~n7328 & n12146 ) | ( ~n7328 & n13664 ) | ( n12146 & n13664 ) ;
  assign n50374 = n50373 ^ n29466 ^ n5736 ;
  assign n50375 = n50374 ^ n43352 ^ n10420 ;
  assign n50376 = ~n10108 & n48292 ;
  assign n50377 = n50376 ^ n1084 ^ 1'b0 ;
  assign n50379 = n6615 & n20886 ;
  assign n50378 = ~n5975 & n31243 ;
  assign n50380 = n50379 ^ n50378 ^ 1'b0 ;
  assign n50381 = ( n4060 & n6724 ) | ( n4060 & n7563 ) | ( n6724 & n7563 ) ;
  assign n50382 = n27253 ^ n7475 ^ n2652 ;
  assign n50383 = ( n11970 & n20632 ) | ( n11970 & n22531 ) | ( n20632 & n22531 ) ;
  assign n50384 = ( n27904 & n50382 ) | ( n27904 & n50383 ) | ( n50382 & n50383 ) ;
  assign n50385 = n10014 | n21114 ;
  assign n50386 = n50385 ^ n48292 ^ n19386 ;
  assign n50388 = n22907 ^ n21195 ^ n13517 ;
  assign n50387 = n7751 & ~n33303 ;
  assign n50389 = n50388 ^ n50387 ^ 1'b0 ;
  assign n50390 = ( n7635 & ~n27034 ) | ( n7635 & n50389 ) | ( ~n27034 & n50389 ) ;
  assign n50391 = n15583 ^ n4018 ^ 1'b0 ;
  assign n50392 = n39805 & n50391 ;
  assign n50393 = ~n14540 & n34001 ;
  assign n50394 = ( ~n7597 & n35609 ) | ( ~n7597 & n36761 ) | ( n35609 & n36761 ) ;
  assign n50395 = n21302 & ~n33323 ;
  assign n50396 = ~n31753 & n50395 ;
  assign n50397 = n40002 ^ n14222 ^ n5209 ;
  assign n50398 = n50397 ^ n48787 ^ n9471 ;
  assign n50399 = n17710 ^ n15960 ^ n8042 ;
  assign n50400 = n29090 ^ n19747 ^ n10498 ;
  assign n50401 = ( n10956 & ~n34241 ) | ( n10956 & n50400 ) | ( ~n34241 & n50400 ) ;
  assign n50402 = ( n6778 & n50399 ) | ( n6778 & ~n50401 ) | ( n50399 & ~n50401 ) ;
  assign n50403 = ( n12201 & n19545 ) | ( n12201 & n23597 ) | ( n19545 & n23597 ) ;
  assign n50404 = n50403 ^ n47913 ^ n47571 ;
  assign n50405 = x132 ^ x31 ^ 1'b0 ;
  assign n50406 = ( n15388 & n37994 ) | ( n15388 & ~n48568 ) | ( n37994 & ~n48568 ) ;
  assign n50407 = ( n47831 & n50405 ) | ( n47831 & n50406 ) | ( n50405 & n50406 ) ;
  assign n50408 = n41999 ^ n32614 ^ n20091 ;
  assign n50409 = ( n11347 & ~n11792 ) | ( n11347 & n25690 ) | ( ~n11792 & n25690 ) ;
  assign n50410 = n50409 ^ n14242 ^ n11948 ;
  assign n50411 = n18363 ^ n9618 ^ n8298 ;
  assign n50412 = ( n30604 & n44016 ) | ( n30604 & n50411 ) | ( n44016 & n50411 ) ;
  assign n50413 = ( n1902 & ~n10643 ) | ( n1902 & n50412 ) | ( ~n10643 & n50412 ) ;
  assign n50414 = n28930 & n49525 ;
  assign n50415 = n50414 ^ n37085 ^ 1'b0 ;
  assign n50419 = ( n6261 & n7156 ) | ( n6261 & ~n29680 ) | ( n7156 & ~n29680 ) ;
  assign n50418 = n7266 ^ n4476 ^ n1850 ;
  assign n50420 = n50419 ^ n50418 ^ n6522 ;
  assign n50421 = n50420 ^ n31905 ^ n10304 ;
  assign n50416 = n19591 ^ n18892 ^ n13790 ;
  assign n50417 = n50416 ^ n39007 ^ n21069 ;
  assign n50422 = n50421 ^ n50417 ^ n43739 ;
  assign n50423 = ( n12755 & ~n37825 ) | ( n12755 & n45679 ) | ( ~n37825 & n45679 ) ;
  assign n50424 = ( ~n7923 & n20344 ) | ( ~n7923 & n23615 ) | ( n20344 & n23615 ) ;
  assign n50425 = ( n452 & n26072 ) | ( n452 & ~n39178 ) | ( n26072 & ~n39178 ) ;
  assign n50426 = ( n11238 & n33573 ) | ( n11238 & ~n35691 ) | ( n33573 & ~n35691 ) ;
  assign n50427 = ( n1292 & n14632 ) | ( n1292 & ~n26699 ) | ( n14632 & ~n26699 ) ;
  assign n50428 = n34655 ^ n27727 ^ 1'b0 ;
  assign n50429 = n9084 | n50428 ;
  assign n50430 = ( ~n44487 & n50427 ) | ( ~n44487 & n50429 ) | ( n50427 & n50429 ) ;
  assign n50431 = n1244 & ~n7346 ;
  assign n50432 = n9395 & n50431 ;
  assign n50433 = ( n7603 & ~n12962 ) | ( n7603 & n50432 ) | ( ~n12962 & n50432 ) ;
  assign n50434 = n50433 ^ n24179 ^ n4163 ;
  assign n50435 = n28033 & n50434 ;
  assign n50439 = ( n11101 & ~n29430 ) | ( n11101 & n50094 ) | ( ~n29430 & n50094 ) ;
  assign n50436 = n25212 ^ n1786 ^ n724 ;
  assign n50437 = ( n5445 & n42857 ) | ( n5445 & n50436 ) | ( n42857 & n50436 ) ;
  assign n50438 = ( ~n4090 & n29282 ) | ( ~n4090 & n50437 ) | ( n29282 & n50437 ) ;
  assign n50440 = n50439 ^ n50438 ^ n13799 ;
  assign n50441 = n3495 & n10168 ;
  assign n50442 = ~n19535 & n50441 ;
  assign n50443 = n24327 ^ n17000 ^ n2420 ;
  assign n50444 = n3572 & ~n17666 ;
  assign n50445 = n50444 ^ n5757 ^ 1'b0 ;
  assign n50446 = ( n23045 & n50443 ) | ( n23045 & n50445 ) | ( n50443 & n50445 ) ;
  assign n50447 = n50446 ^ n14464 ^ n7746 ;
  assign n50448 = ( n8152 & n50442 ) | ( n8152 & n50447 ) | ( n50442 & n50447 ) ;
  assign n50449 = ( n1264 & ~n22887 ) | ( n1264 & n50448 ) | ( ~n22887 & n50448 ) ;
  assign n50450 = n47744 ^ n47698 ^ n30638 ;
  assign n50451 = n13321 | n50450 ;
  assign n50452 = n41719 & ~n42999 ;
  assign n50453 = n5005 & n50452 ;
  assign n50454 = n40351 ^ n34740 ^ n26763 ;
  assign n50455 = ( ~n581 & n21334 ) | ( ~n581 & n50454 ) | ( n21334 & n50454 ) ;
  assign n50456 = n37697 ^ n29516 ^ n8938 ;
  assign n50457 = n14618 ^ n12242 ^ n5781 ;
  assign n50458 = n50457 ^ n26610 ^ 1'b0 ;
  assign n50459 = ( n15960 & n17220 ) | ( n15960 & ~n32401 ) | ( n17220 & ~n32401 ) ;
  assign n50460 = n50459 ^ n50113 ^ n5047 ;
  assign n50461 = ( n889 & ~n39876 ) | ( n889 & n50460 ) | ( ~n39876 & n50460 ) ;
  assign n50462 = ( x5 & n7264 ) | ( x5 & ~n15759 ) | ( n7264 & ~n15759 ) ;
  assign n50463 = n30103 ^ n16528 ^ n2609 ;
  assign n50464 = n50463 ^ n44848 ^ n11750 ;
  assign n50465 = n46216 ^ n10144 ^ 1'b0 ;
  assign n50466 = ( n26781 & ~n33400 ) | ( n26781 & n37068 ) | ( ~n33400 & n37068 ) ;
  assign n50467 = ( ~n6279 & n12706 ) | ( ~n6279 & n41432 ) | ( n12706 & n41432 ) ;
  assign n50468 = ( ~n18767 & n42593 ) | ( ~n18767 & n50467 ) | ( n42593 & n50467 ) ;
  assign n50469 = ( n21336 & ~n33745 ) | ( n21336 & n45989 ) | ( ~n33745 & n45989 ) ;
  assign n50470 = ( n10743 & ~n18842 ) | ( n10743 & n37609 ) | ( ~n18842 & n37609 ) ;
  assign n50471 = ( ~n31947 & n38725 ) | ( ~n31947 & n47642 ) | ( n38725 & n47642 ) ;
  assign n50472 = ( ~x190 & n10218 ) | ( ~x190 & n26960 ) | ( n10218 & n26960 ) ;
  assign n50474 = n4771 | n22950 ;
  assign n50475 = n7480 & ~n50474 ;
  assign n50473 = n15892 ^ n15334 ^ n5111 ;
  assign n50476 = n50475 ^ n50473 ^ n33695 ;
  assign n50477 = ( n2003 & n7583 ) | ( n2003 & n39226 ) | ( n7583 & n39226 ) ;
  assign n50478 = n50477 ^ n12275 ^ n10925 ;
  assign n50479 = ( n481 & ~n2309 ) | ( n481 & n37928 ) | ( ~n2309 & n37928 ) ;
  assign n50480 = ~n6317 & n47038 ;
  assign n50481 = n4113 & n50480 ;
  assign n50482 = n11701 & ~n19948 ;
  assign n50483 = ( n7424 & n8133 ) | ( n7424 & n50482 ) | ( n8133 & n50482 ) ;
  assign n50484 = n50483 ^ n18922 ^ 1'b0 ;
  assign n50485 = n4448 & ~n50484 ;
  assign n50486 = n43259 ^ n31046 ^ n938 ;
  assign n50487 = n50486 ^ n22043 ^ n1467 ;
  assign n50488 = ( ~n15082 & n38824 ) | ( ~n15082 & n50268 ) | ( n38824 & n50268 ) ;
  assign n50489 = n48602 ^ n22653 ^ n19829 ;
  assign n50490 = n19457 & n33256 ;
  assign n50491 = ( n11924 & n50489 ) | ( n11924 & ~n50490 ) | ( n50489 & ~n50490 ) ;
  assign n50492 = ( n4315 & n6437 ) | ( n4315 & n13527 ) | ( n6437 & n13527 ) ;
  assign n50494 = n16425 ^ n12496 ^ n5802 ;
  assign n50493 = ( n6734 & n6770 ) | ( n6734 & n33118 ) | ( n6770 & n33118 ) ;
  assign n50495 = n50494 ^ n50493 ^ n29511 ;
  assign n50496 = ( ~x89 & n50492 ) | ( ~x89 & n50495 ) | ( n50492 & n50495 ) ;
  assign n50497 = ( ~n6819 & n20114 ) | ( ~n6819 & n35245 ) | ( n20114 & n35245 ) ;
  assign n50498 = ( ~n3028 & n3539 ) | ( ~n3028 & n34402 ) | ( n3539 & n34402 ) ;
  assign n50499 = ( n14975 & n31907 ) | ( n14975 & n50498 ) | ( n31907 & n50498 ) ;
  assign n50500 = n4377 & ~n50499 ;
  assign n50501 = ( n2922 & n12462 ) | ( n2922 & n16934 ) | ( n12462 & n16934 ) ;
  assign n50502 = ( n15546 & ~n34046 ) | ( n15546 & n50501 ) | ( ~n34046 & n50501 ) ;
  assign n50503 = n4499 & ~n34366 ;
  assign n50504 = n7539 & n50503 ;
  assign n50505 = n13215 ^ n3749 ^ n3689 ;
  assign n50506 = ( n29596 & n36908 ) | ( n29596 & ~n50505 ) | ( n36908 & ~n50505 ) ;
  assign n50507 = n47191 ^ n35445 ^ n4370 ;
  assign n50508 = n26386 ^ n25892 ^ n24550 ;
  assign n50509 = ( n7361 & n48144 ) | ( n7361 & n50508 ) | ( n48144 & n50508 ) ;
  assign n50510 = n27738 ^ n26064 ^ n17364 ;
  assign n50511 = n50510 ^ n13896 ^ n4772 ;
  assign n50512 = n47198 ^ n27770 ^ n24459 ;
  assign n50513 = n50512 ^ n29379 ^ n4844 ;
  assign n50514 = n37456 ^ n31495 ^ n10430 ;
  assign n50515 = n28483 ^ n16318 ^ 1'b0 ;
  assign n50516 = n50515 ^ n26829 ^ n10326 ;
  assign n50517 = n31844 ^ n24193 ^ n7089 ;
  assign n50525 = n6831 & n10828 ;
  assign n50526 = n50525 ^ n10357 ^ 1'b0 ;
  assign n50527 = n50526 ^ n33903 ^ n8189 ;
  assign n50528 = ( n9197 & ~n15600 ) | ( n9197 & n50527 ) | ( ~n15600 & n50527 ) ;
  assign n50529 = ( n12156 & ~n23659 ) | ( n12156 & n50528 ) | ( ~n23659 & n50528 ) ;
  assign n50518 = ( n2064 & n13714 ) | ( n2064 & ~n38976 ) | ( n13714 & ~n38976 ) ;
  assign n50520 = n24350 ^ n14209 ^ x185 ;
  assign n50521 = n23743 & n50520 ;
  assign n50522 = n50521 ^ n9786 ^ 1'b0 ;
  assign n50519 = n41921 ^ n14431 ^ n10096 ;
  assign n50523 = n50522 ^ n50519 ^ n23284 ;
  assign n50524 = ( ~n33628 & n50518 ) | ( ~n33628 & n50523 ) | ( n50518 & n50523 ) ;
  assign n50530 = n50529 ^ n50524 ^ n7899 ;
  assign n50531 = n8614 & ~n26185 ;
  assign n50532 = n3285 & ~n31048 ;
  assign n50533 = n39929 ^ n16018 ^ n13631 ;
  assign n50534 = ( n4393 & n23772 ) | ( n4393 & ~n50533 ) | ( n23772 & ~n50533 ) ;
  assign n50535 = n50532 & n50534 ;
  assign n50536 = ~n50531 & n50535 ;
  assign n50537 = ~n8035 & n25576 ;
  assign n50538 = n50537 ^ n6300 ^ 1'b0 ;
  assign n50540 = ( n3047 & n13005 ) | ( n3047 & n24921 ) | ( n13005 & n24921 ) ;
  assign n50541 = n50540 ^ n20238 ^ n19666 ;
  assign n50539 = n15324 ^ n12843 ^ n7206 ;
  assign n50542 = n50541 ^ n50539 ^ n12530 ;
  assign n50543 = n26614 ^ n25748 ^ 1'b0 ;
  assign n50544 = ( n18576 & n37285 ) | ( n18576 & n47185 ) | ( n37285 & n47185 ) ;
  assign n50545 = ( n13634 & n28286 ) | ( n13634 & n48642 ) | ( n28286 & n48642 ) ;
  assign n50546 = n30875 & ~n33724 ;
  assign n50547 = n35874 ^ n33976 ^ 1'b0 ;
  assign n50548 = n26068 ^ n3218 ^ n372 ;
  assign n50549 = n50548 ^ n19522 ^ 1'b0 ;
  assign n50550 = n42169 ^ n20099 ^ n12674 ;
  assign n50551 = n40903 ^ n18004 ^ 1'b0 ;
  assign n50552 = n50551 ^ n26832 ^ n13589 ;
  assign n50553 = n50552 ^ n7396 ^ n7112 ;
  assign n50554 = n4619 & ~n33021 ;
  assign n50555 = n41112 ^ n23963 ^ 1'b0 ;
  assign n50556 = n50554 | n50555 ;
  assign n50557 = n24369 ^ n23340 ^ n15196 ;
  assign n50558 = n50557 ^ n40853 ^ n10651 ;
  assign n50559 = n50558 ^ n18988 ^ n14450 ;
  assign n50560 = ( n4474 & ~n10901 ) | ( n4474 & n20275 ) | ( ~n10901 & n20275 ) ;
  assign n50561 = n50560 ^ n40367 ^ n1711 ;
  assign n50562 = n46589 ^ n29282 ^ n15487 ;
  assign n50563 = n8334 & n50562 ;
  assign n50564 = n45699 & n50563 ;
  assign n50565 = ( n50559 & n50561 ) | ( n50559 & n50564 ) | ( n50561 & n50564 ) ;
  assign n50566 = n43700 ^ n10773 ^ n2268 ;
  assign n50567 = n50566 ^ n19762 ^ n17810 ;
  assign n50568 = n22260 ^ n14365 ^ n1766 ;
  assign n50569 = ( n11197 & n17065 ) | ( n11197 & ~n32860 ) | ( n17065 & ~n32860 ) ;
  assign n50570 = n50569 ^ n16429 ^ n15915 ;
  assign n50571 = n18500 ^ n17446 ^ n1919 ;
  assign n50572 = ( ~n8584 & n20288 ) | ( ~n8584 & n24742 ) | ( n20288 & n24742 ) ;
  assign n50573 = ( n14428 & n24367 ) | ( n14428 & ~n24640 ) | ( n24367 & ~n24640 ) ;
  assign n50574 = ( n6741 & n17475 ) | ( n6741 & n28377 ) | ( n17475 & n28377 ) ;
  assign n50575 = n50574 ^ n3559 ^ n1133 ;
  assign n50576 = ( n4905 & n18325 ) | ( n4905 & ~n29699 ) | ( n18325 & ~n29699 ) ;
  assign n50579 = n32628 ^ n26050 ^ n10948 ;
  assign n50577 = n11808 ^ n3270 ^ n804 ;
  assign n50578 = ( n26003 & ~n27346 ) | ( n26003 & n50577 ) | ( ~n27346 & n50577 ) ;
  assign n50580 = n50579 ^ n50578 ^ n8392 ;
  assign n50581 = ( n545 & ~n15775 ) | ( n545 & n17287 ) | ( ~n15775 & n17287 ) ;
  assign n50582 = ( n33478 & ~n36175 ) | ( n33478 & n45237 ) | ( ~n36175 & n45237 ) ;
  assign n50583 = ( n22074 & ~n50581 ) | ( n22074 & n50582 ) | ( ~n50581 & n50582 ) ;
  assign n50586 = ( ~n3958 & n4493 ) | ( ~n3958 & n8301 ) | ( n4493 & n8301 ) ;
  assign n50587 = n50586 ^ n20021 ^ n13364 ;
  assign n50584 = n11616 ^ n7128 ^ 1'b0 ;
  assign n50585 = ~n35945 & n50584 ;
  assign n50588 = n50587 ^ n50585 ^ n45283 ;
  assign n50589 = ( n19623 & ~n22302 ) | ( n19623 & n31589 ) | ( ~n22302 & n31589 ) ;
  assign n50590 = n47255 ^ n38975 ^ n33292 ;
  assign n50591 = n50590 ^ n38427 ^ n23615 ;
  assign n50592 = n46653 ^ n26930 ^ n2910 ;
  assign n50593 = ( n14132 & n25219 ) | ( n14132 & ~n29897 ) | ( n25219 & ~n29897 ) ;
  assign n50594 = ( n14949 & n27218 ) | ( n14949 & n50593 ) | ( n27218 & n50593 ) ;
  assign n50595 = ( n22210 & n50592 ) | ( n22210 & ~n50594 ) | ( n50592 & ~n50594 ) ;
  assign n50596 = n48489 ^ n44097 ^ 1'b0 ;
  assign n50597 = n43996 & n50596 ;
  assign n50598 = ~n7084 & n43987 ;
  assign n50599 = n50598 ^ n3822 ^ 1'b0 ;
  assign n50600 = ( n25505 & ~n28030 ) | ( n25505 & n34054 ) | ( ~n28030 & n34054 ) ;
  assign n50601 = n17147 ^ n4312 ^ 1'b0 ;
  assign n50602 = ( n445 & n13085 ) | ( n445 & ~n50601 ) | ( n13085 & ~n50601 ) ;
  assign n50603 = n35715 ^ n4979 ^ n3627 ;
  assign n50604 = n33937 ^ n3658 ^ 1'b0 ;
  assign n50605 = n31079 ^ n25638 ^ n8633 ;
  assign n50606 = n27644 ^ n6686 ^ n2626 ;
  assign n50607 = ( n6414 & n34210 ) | ( n6414 & ~n50606 ) | ( n34210 & ~n50606 ) ;
  assign n50608 = n50607 ^ n17174 ^ n12238 ;
  assign n50609 = ~n50605 & n50608 ;
  assign n50610 = ( n13393 & n14751 ) | ( n13393 & ~n44465 ) | ( n14751 & ~n44465 ) ;
  assign n50611 = n50610 ^ n24642 ^ 1'b0 ;
  assign n50612 = n7667 & n31243 ;
  assign n50613 = n50612 ^ n10520 ^ 1'b0 ;
  assign n50614 = ( n12736 & n13266 ) | ( n12736 & n50613 ) | ( n13266 & n50613 ) ;
  assign n50615 = n20999 ^ n7383 ^ n2768 ;
  assign n50616 = ( n8267 & n37850 ) | ( n8267 & ~n38459 ) | ( n37850 & ~n38459 ) ;
  assign n50617 = n50616 ^ n39878 ^ n37073 ;
  assign n50618 = ~n7385 & n42751 ;
  assign n50619 = n50618 ^ n1005 ^ 1'b0 ;
  assign n50620 = n17684 ^ n15767 ^ 1'b0 ;
  assign n50621 = n5665 & ~n11145 ;
  assign n50622 = n9278 & n50621 ;
  assign n50623 = ( n7918 & n16034 ) | ( n7918 & ~n50622 ) | ( n16034 & ~n50622 ) ;
  assign n50624 = n13661 & n16488 ;
  assign n50625 = n50624 ^ n4953 ^ 1'b0 ;
  assign n50626 = n50625 ^ n4454 ^ n1899 ;
  assign n50627 = ( n9623 & ~n48423 ) | ( n9623 & n50626 ) | ( ~n48423 & n50626 ) ;
  assign n50631 = n42919 ^ n29308 ^ n10185 ;
  assign n50628 = ( n25498 & n26284 ) | ( n25498 & n26446 ) | ( n26284 & n26446 ) ;
  assign n50629 = ( n12200 & n37926 ) | ( n12200 & ~n50628 ) | ( n37926 & ~n50628 ) ;
  assign n50630 = ( n9210 & n14873 ) | ( n9210 & n50629 ) | ( n14873 & n50629 ) ;
  assign n50632 = n50631 ^ n50630 ^ n21641 ;
  assign n50633 = ( n15329 & n33978 ) | ( n15329 & n50632 ) | ( n33978 & n50632 ) ;
  assign n50634 = n8310 | n19067 ;
  assign n50635 = n50634 ^ n49318 ^ n8668 ;
  assign n50636 = n27945 ^ n18782 ^ n16694 ;
  assign n50637 = n28281 ^ n2600 ^ n1729 ;
  assign n50638 = ( n7028 & n11326 ) | ( n7028 & ~n50637 ) | ( n11326 & ~n50637 ) ;
  assign n50639 = n6000 | n17949 ;
  assign n50640 = n50639 ^ n8314 ^ 1'b0 ;
  assign n50641 = ~n29549 & n39495 ;
  assign n50642 = n50640 & n50641 ;
  assign n50643 = ~n5299 & n16544 ;
  assign n50647 = n36039 ^ n13773 ^ n11214 ;
  assign n50644 = n16895 ^ n12465 ^ n6328 ;
  assign n50645 = n50644 ^ n33531 ^ n14590 ;
  assign n50646 = ( ~n20184 & n26337 ) | ( ~n20184 & n50645 ) | ( n26337 & n50645 ) ;
  assign n50648 = n50647 ^ n50646 ^ n4580 ;
  assign n50649 = n6706 & n34444 ;
  assign n50650 = n50649 ^ n5746 ^ 1'b0 ;
  assign n50651 = n31364 ^ n17768 ^ n9719 ;
  assign n50654 = n7020 | n31390 ;
  assign n50655 = n50654 ^ n1301 ^ 1'b0 ;
  assign n50652 = n3121 & ~n3883 ;
  assign n50653 = n50652 ^ n45199 ^ 1'b0 ;
  assign n50656 = n50655 ^ n50653 ^ n11074 ;
  assign n50657 = ( n50650 & n50651 ) | ( n50650 & ~n50656 ) | ( n50651 & ~n50656 ) ;
  assign n50658 = n49332 ^ n43668 ^ n14462 ;
  assign n50659 = n34874 ^ n20750 ^ n15241 ;
  assign n50660 = x230 & ~n36582 ;
  assign n50661 = ~n44532 & n50660 ;
  assign n50662 = ( n12400 & n33267 ) | ( n12400 & ~n50661 ) | ( n33267 & ~n50661 ) ;
  assign n50663 = n50662 ^ n28472 ^ n25409 ;
  assign n50664 = n41291 ^ n17599 ^ n2630 ;
  assign n50665 = ( n12458 & ~n13223 ) | ( n12458 & n50664 ) | ( ~n13223 & n50664 ) ;
  assign n50666 = n50665 ^ n16676 ^ n4045 ;
  assign n50667 = ( n3150 & n13057 ) | ( n3150 & ~n34253 ) | ( n13057 & ~n34253 ) ;
  assign n50668 = n50667 ^ n808 ^ 1'b0 ;
  assign n50669 = ~n30515 & n50668 ;
  assign n50670 = n6452 | n14218 ;
  assign n50673 = n28802 ^ n11007 ^ 1'b0 ;
  assign n50671 = ( ~n1992 & n3472 ) | ( ~n1992 & n15374 ) | ( n3472 & n15374 ) ;
  assign n50672 = x184 & ~n50671 ;
  assign n50674 = n50673 ^ n50672 ^ n2745 ;
  assign n50675 = ( n8803 & ~n39470 ) | ( n8803 & n50674 ) | ( ~n39470 & n50674 ) ;
  assign n50676 = n21234 ^ n16881 ^ 1'b0 ;
  assign n50677 = n50676 ^ n33035 ^ n32918 ;
  assign n50678 = n833 | n4424 ;
  assign n50679 = ~n988 & n18296 ;
  assign n50680 = ( n16202 & ~n50678 ) | ( n16202 & n50679 ) | ( ~n50678 & n50679 ) ;
  assign n50681 = n50680 ^ n13962 ^ n2719 ;
  assign n50682 = ( n5036 & n40093 ) | ( n5036 & ~n48060 ) | ( n40093 & ~n48060 ) ;
  assign n50683 = n43959 ^ n30756 ^ n1597 ;
  assign n50684 = n8934 & n36783 ;
  assign n50685 = ~n3463 & n50684 ;
  assign n50686 = ( ~n3561 & n18577 ) | ( ~n3561 & n27773 ) | ( n18577 & n27773 ) ;
  assign n50688 = n32781 & n44298 ;
  assign n50689 = n50688 ^ n44816 ^ 1'b0 ;
  assign n50687 = n33221 ^ n26007 ^ n269 ;
  assign n50690 = n50689 ^ n50687 ^ n14042 ;
  assign n50691 = ( ~n4718 & n50686 ) | ( ~n4718 & n50690 ) | ( n50686 & n50690 ) ;
  assign n50692 = n11204 ^ n7914 ^ n2431 ;
  assign n50696 = ( n8171 & ~n10684 ) | ( n8171 & n28328 ) | ( ~n10684 & n28328 ) ;
  assign n50694 = n16701 | n45969 ;
  assign n50695 = n50694 ^ n36418 ^ n23004 ;
  assign n50693 = n37126 ^ n36150 ^ n11269 ;
  assign n50697 = n50696 ^ n50695 ^ n50693 ;
  assign n50698 = n29947 ^ n16283 ^ n13953 ;
  assign n50699 = ( ~n11064 & n30315 ) | ( ~n11064 & n48783 ) | ( n30315 & n48783 ) ;
  assign n50700 = ( n11505 & n18450 ) | ( n11505 & ~n50699 ) | ( n18450 & ~n50699 ) ;
  assign n50701 = n49866 ^ n38981 ^ n33875 ;
  assign n50702 = n50701 ^ n45925 ^ n18791 ;
  assign n50703 = n16925 & ~n50702 ;
  assign n50704 = n50703 ^ n37650 ^ n28233 ;
  assign n50705 = n35549 ^ n9952 ^ n747 ;
  assign n50708 = n334 & ~n1324 ;
  assign n50709 = n50708 ^ n42603 ^ 1'b0 ;
  assign n50706 = ( ~n466 & n7072 ) | ( ~n466 & n34505 ) | ( n7072 & n34505 ) ;
  assign n50707 = ~n19126 & n50706 ;
  assign n50710 = n50709 ^ n50707 ^ 1'b0 ;
  assign n50711 = n29711 | n50710 ;
  assign n50712 = n26158 & ~n50711 ;
  assign n50713 = ( n20914 & ~n41422 ) | ( n20914 & n46844 ) | ( ~n41422 & n46844 ) ;
  assign n50714 = n38881 ^ n28417 ^ n13864 ;
  assign n50717 = n6887 ^ n6335 ^ 1'b0 ;
  assign n50718 = n50717 ^ n42022 ^ 1'b0 ;
  assign n50719 = ( n11991 & ~n38041 ) | ( n11991 & n50718 ) | ( ~n38041 & n50718 ) ;
  assign n50715 = n45750 ^ n27137 ^ n18184 ;
  assign n50716 = ( ~n18601 & n29997 ) | ( ~n18601 & n50715 ) | ( n29997 & n50715 ) ;
  assign n50720 = n50719 ^ n50716 ^ n14156 ;
  assign n50721 = n8555 | n12601 ;
  assign n50722 = n50721 ^ n11454 ^ n11068 ;
  assign n50725 = ( n4445 & n21828 ) | ( n4445 & n26384 ) | ( n21828 & n26384 ) ;
  assign n50723 = ( ~n5479 & n19141 ) | ( ~n5479 & n47443 ) | ( n19141 & n47443 ) ;
  assign n50724 = ( n7616 & n18988 ) | ( n7616 & n50723 ) | ( n18988 & n50723 ) ;
  assign n50726 = n50725 ^ n50724 ^ n27646 ;
  assign n50727 = n40116 ^ n38113 ^ n24850 ;
  assign n50728 = n24383 ^ n15237 ^ n4563 ;
  assign n50729 = n1583 | n17916 ;
  assign n50730 = ( n4926 & n12436 ) | ( n4926 & ~n13586 ) | ( n12436 & ~n13586 ) ;
  assign n50731 = n21312 | n50730 ;
  assign n50732 = n50731 ^ n24359 ^ 1'b0 ;
  assign n50733 = ( n9934 & ~n32864 ) | ( n9934 & n50732 ) | ( ~n32864 & n50732 ) ;
  assign n50734 = ( n1512 & n46402 ) | ( n1512 & n50733 ) | ( n46402 & n50733 ) ;
  assign n50735 = ~n27072 & n36597 ;
  assign n50736 = n9097 ^ n4197 ^ 1'b0 ;
  assign n50737 = ( n10223 & n37629 ) | ( n10223 & n50736 ) | ( n37629 & n50736 ) ;
  assign n50738 = n15293 & n23004 ;
  assign n50739 = ~n13720 & n50738 ;
  assign n50740 = ( n7094 & n35620 ) | ( n7094 & n50739 ) | ( n35620 & n50739 ) ;
  assign n50741 = ( n21422 & ~n24829 ) | ( n21422 & n31173 ) | ( ~n24829 & n31173 ) ;
  assign n50742 = n50741 ^ n44467 ^ n22512 ;
  assign n50743 = n49821 ^ n29142 ^ 1'b0 ;
  assign n50744 = n22514 ^ n5717 ^ 1'b0 ;
  assign n50745 = n20507 | n50744 ;
  assign n50746 = ( n10778 & n33621 ) | ( n10778 & n50745 ) | ( n33621 & n50745 ) ;
  assign n50747 = n24830 ^ n13301 ^ n6570 ;
  assign n50748 = n50747 ^ n39873 ^ n16025 ;
  assign n50751 = ( n18179 & n18492 ) | ( n18179 & n45502 ) | ( n18492 & n45502 ) ;
  assign n50749 = ( ~n6430 & n11676 ) | ( ~n6430 & n37165 ) | ( n11676 & n37165 ) ;
  assign n50750 = n50749 ^ n32833 ^ n10949 ;
  assign n50752 = n50751 ^ n50750 ^ n6200 ;
  assign n50753 = ( ~n15793 & n18639 ) | ( ~n15793 & n50752 ) | ( n18639 & n50752 ) ;
  assign n50754 = n10163 ^ n5918 ^ n2634 ;
  assign n50755 = n37518 ^ n12008 ^ n6828 ;
  assign n50756 = n50755 ^ n27938 ^ n25303 ;
  assign n50757 = ( n31152 & n50754 ) | ( n31152 & n50756 ) | ( n50754 & n50756 ) ;
  assign n50758 = n28951 | n41088 ;
  assign n50759 = ( n3016 & n16179 ) | ( n3016 & ~n22559 ) | ( n16179 & ~n22559 ) ;
  assign n50760 = ( ~n2929 & n6482 ) | ( ~n2929 & n7107 ) | ( n6482 & n7107 ) ;
  assign n50761 = ( n9855 & n29511 ) | ( n9855 & ~n50760 ) | ( n29511 & ~n50760 ) ;
  assign n50762 = n2061 & n17272 ;
  assign n50763 = n50762 ^ n43213 ^ 1'b0 ;
  assign n50764 = ( n35929 & n48933 ) | ( n35929 & ~n50763 ) | ( n48933 & ~n50763 ) ;
  assign n50765 = ( n1893 & n8624 ) | ( n1893 & ~n50764 ) | ( n8624 & ~n50764 ) ;
  assign n50766 = ( n3152 & n25541 ) | ( n3152 & ~n50765 ) | ( n25541 & ~n50765 ) ;
  assign n50767 = ( n9406 & n41533 ) | ( n9406 & n48370 ) | ( n41533 & n48370 ) ;
  assign n50768 = n36179 ^ n851 ^ 1'b0 ;
  assign n50769 = n12547 | n50768 ;
  assign n50770 = n26867 ^ n7432 ^ 1'b0 ;
  assign n50771 = n18181 | n50770 ;
  assign n50772 = ( ~n45761 & n50769 ) | ( ~n45761 & n50771 ) | ( n50769 & n50771 ) ;
  assign n50773 = n50772 ^ n45550 ^ n30579 ;
  assign n50774 = ( n21681 & ~n25192 ) | ( n21681 & n39585 ) | ( ~n25192 & n39585 ) ;
  assign n50775 = ( n17307 & ~n18660 ) | ( n17307 & n48513 ) | ( ~n18660 & n48513 ) ;
  assign n50776 = n50775 ^ n32792 ^ n6766 ;
  assign n50777 = n13282 ^ n7256 ^ 1'b0 ;
  assign n50778 = n43581 | n50777 ;
  assign n50779 = n50778 ^ n47735 ^ n36881 ;
  assign n50780 = ( n4525 & ~n50776 ) | ( n4525 & n50779 ) | ( ~n50776 & n50779 ) ;
  assign n50781 = n19353 ^ n15753 ^ 1'b0 ;
  assign n50782 = ( ~n9911 & n10190 ) | ( ~n9911 & n14032 ) | ( n10190 & n14032 ) ;
  assign n50783 = n7636 ^ n6902 ^ n664 ;
  assign n50784 = ~n44841 & n50783 ;
  assign n50785 = n50782 & n50784 ;
  assign n50786 = ( n21994 & ~n25083 ) | ( n21994 & n47739 ) | ( ~n25083 & n47739 ) ;
  assign n50787 = ( n11487 & n48721 ) | ( n11487 & ~n50786 ) | ( n48721 & ~n50786 ) ;
  assign n50788 = ( n1131 & ~n25049 ) | ( n1131 & n36224 ) | ( ~n25049 & n36224 ) ;
  assign n50789 = ( n18701 & ~n26733 ) | ( n18701 & n50788 ) | ( ~n26733 & n50788 ) ;
  assign n50790 = ( n417 & n34287 ) | ( n417 & n46824 ) | ( n34287 & n46824 ) ;
  assign n50791 = ( n464 & n1440 ) | ( n464 & ~n3828 ) | ( n1440 & ~n3828 ) ;
  assign n50792 = n50791 ^ n46593 ^ n29245 ;
  assign n50793 = ~n3741 & n11511 ;
  assign n50794 = n50793 ^ n48856 ^ 1'b0 ;
  assign n50795 = n50794 ^ n28364 ^ n4201 ;
  assign n50796 = ( n23469 & n25791 ) | ( n23469 & n50795 ) | ( n25791 & n50795 ) ;
  assign n50797 = n16632 ^ n10395 ^ 1'b0 ;
  assign n50798 = n32602 ^ n15909 ^ n2534 ;
  assign n50799 = ( n16562 & n50797 ) | ( n16562 & ~n50798 ) | ( n50797 & ~n50798 ) ;
  assign n50800 = ( n16206 & n25062 ) | ( n16206 & n50799 ) | ( n25062 & n50799 ) ;
  assign n50801 = ( n13532 & n15935 ) | ( n13532 & n26949 ) | ( n15935 & n26949 ) ;
  assign n50802 = n35760 ^ n27342 ^ n12077 ;
  assign n50803 = ( n2818 & ~n50801 ) | ( n2818 & n50802 ) | ( ~n50801 & n50802 ) ;
  assign n50804 = ~n6626 & n11385 ;
  assign n50805 = n3466 & n50804 ;
  assign n50806 = n24382 ^ n16935 ^ n3449 ;
  assign n50807 = ( ~n19429 & n50805 ) | ( ~n19429 & n50806 ) | ( n50805 & n50806 ) ;
  assign n50808 = ( n2795 & n8993 ) | ( n2795 & ~n26574 ) | ( n8993 & ~n26574 ) ;
  assign n50809 = n18010 & ~n36995 ;
  assign n50810 = n27943 & n50809 ;
  assign n50811 = n47331 & ~n50810 ;
  assign n50812 = ~n48537 & n50811 ;
  assign n50813 = n39392 ^ n3349 ^ 1'b0 ;
  assign n50814 = n17597 & ~n50813 ;
  assign n50815 = n12609 ^ n6467 ^ n2778 ;
  assign n50816 = n50815 ^ n38447 ^ 1'b0 ;
  assign n50817 = n40176 ^ n14094 ^ 1'b0 ;
  assign n50818 = n50817 ^ n37819 ^ n3943 ;
  assign n50819 = n14575 ^ n10062 ^ n593 ;
  assign n50820 = ( n32392 & n44694 ) | ( n32392 & n50819 ) | ( n44694 & n50819 ) ;
  assign n50821 = ( n8040 & n29950 ) | ( n8040 & n30255 ) | ( n29950 & n30255 ) ;
  assign n50822 = n50821 ^ n41048 ^ n5146 ;
  assign n50823 = n20559 | n38555 ;
  assign n50824 = n40459 ^ n6655 ^ n823 ;
  assign n50825 = ( n10096 & n25828 ) | ( n10096 & n33159 ) | ( n25828 & n33159 ) ;
  assign n50826 = ( n7525 & n20883 ) | ( n7525 & ~n50825 ) | ( n20883 & ~n50825 ) ;
  assign n50827 = ( n50823 & ~n50824 ) | ( n50823 & n50826 ) | ( ~n50824 & n50826 ) ;
  assign n50828 = ( n19868 & n27642 ) | ( n19868 & ~n42031 ) | ( n27642 & ~n42031 ) ;
  assign n50829 = n24335 ^ n10763 ^ n5974 ;
  assign n50830 = n9434 | n12029 ;
  assign n50831 = n12154 & ~n50830 ;
  assign n50832 = ( n5780 & ~n25038 ) | ( n5780 & n50831 ) | ( ~n25038 & n50831 ) ;
  assign n50833 = ( n34791 & n47600 ) | ( n34791 & n50832 ) | ( n47600 & n50832 ) ;
  assign n50834 = n45387 ^ n39525 ^ n16911 ;
  assign n50835 = n17328 & n35900 ;
  assign n50836 = ~n15557 & n50835 ;
  assign n50837 = ( n11988 & n26325 ) | ( n11988 & ~n32114 ) | ( n26325 & ~n32114 ) ;
  assign n50838 = n20341 & ~n37419 ;
  assign n50839 = ~n18185 & n18557 ;
  assign n50840 = n50839 ^ n7857 ^ n7478 ;
  assign n50841 = n50840 ^ n9021 ^ n4235 ;
  assign n50842 = ( n10094 & n26477 ) | ( n10094 & ~n38386 ) | ( n26477 & ~n38386 ) ;
  assign n50843 = ( n436 & n20472 ) | ( n436 & ~n39154 ) | ( n20472 & ~n39154 ) ;
  assign n50844 = n11481 ^ n5558 ^ n5104 ;
  assign n50845 = ( n2856 & n4700 ) | ( n2856 & n50844 ) | ( n4700 & n50844 ) ;
  assign n50846 = n47131 ^ n10493 ^ x233 ;
  assign n50847 = n33985 & n49366 ;
  assign n50848 = n25237 & n50847 ;
  assign n50849 = ( n9145 & n21811 ) | ( n9145 & n33347 ) | ( n21811 & n33347 ) ;
  assign n50850 = ~n14276 & n50849 ;
  assign n50851 = ( n1025 & ~n1127 ) | ( n1025 & n41332 ) | ( ~n1127 & n41332 ) ;
  assign n50854 = n10193 ^ n7038 ^ 1'b0 ;
  assign n50853 = n31787 ^ n21872 ^ n3191 ;
  assign n50852 = n24004 ^ n3798 ^ n3427 ;
  assign n50855 = n50854 ^ n50853 ^ n50852 ;
  assign n50856 = n50709 ^ n18695 ^ n8751 ;
  assign n50857 = n35957 ^ n33141 ^ 1'b0 ;
  assign n50858 = n13678 | n50857 ;
  assign n50859 = n50858 ^ n38902 ^ n19042 ;
  assign n50860 = n12812 ^ n11951 ^ n10960 ;
  assign n50861 = n45000 ^ n37874 ^ n13120 ;
  assign n50862 = n33362 ^ n13075 ^ n7061 ;
  assign n50863 = n50862 ^ n36857 ^ n2672 ;
  assign n50864 = n40434 ^ n9030 ^ 1'b0 ;
  assign n50865 = n50864 ^ n24150 ^ n19762 ;
  assign n50866 = n50865 ^ n12305 ^ n5856 ;
  assign n50867 = ( x41 & n37919 ) | ( x41 & n50866 ) | ( n37919 & n50866 ) ;
  assign n50868 = ~n9270 & n39141 ;
  assign n50869 = ( n2406 & ~n5004 ) | ( n2406 & n50868 ) | ( ~n5004 & n50868 ) ;
  assign n50870 = n45869 ^ n40002 ^ n5930 ;
  assign n50871 = ( ~n17267 & n50869 ) | ( ~n17267 & n50870 ) | ( n50869 & n50870 ) ;
  assign n50872 = ( x181 & n8451 ) | ( x181 & ~n39130 ) | ( n8451 & ~n39130 ) ;
  assign n50873 = n22173 ^ n9008 ^ n1349 ;
  assign n50874 = ( ~n36840 & n43477 ) | ( ~n36840 & n50873 ) | ( n43477 & n50873 ) ;
  assign n50875 = n10651 | n12725 ;
  assign n50876 = n26249 & ~n50875 ;
  assign n50877 = n50876 ^ n16210 ^ 1'b0 ;
  assign n50878 = n22578 | n50877 ;
  assign n50879 = n50878 ^ n30754 ^ n5852 ;
  assign n50880 = n36286 ^ n33805 ^ x13 ;
  assign n50881 = ( n15474 & n44832 ) | ( n15474 & n50880 ) | ( n44832 & n50880 ) ;
  assign n50882 = n38473 ^ n21972 ^ n1405 ;
  assign n50883 = ( ~n4460 & n19731 ) | ( ~n4460 & n50882 ) | ( n19731 & n50882 ) ;
  assign n50884 = n30552 ^ n28952 ^ 1'b0 ;
  assign n50885 = n22821 | n37315 ;
  assign n50886 = n50885 ^ n2825 ^ 1'b0 ;
  assign n50887 = n22326 ^ n1356 ^ 1'b0 ;
  assign n50888 = ( n2967 & n35485 ) | ( n2967 & ~n39890 ) | ( n35485 & ~n39890 ) ;
  assign n50889 = n15734 & n42161 ;
  assign n50890 = ( n760 & ~n2633 ) | ( n760 & n39788 ) | ( ~n2633 & n39788 ) ;
  assign n50891 = ( n4540 & n9760 ) | ( n4540 & ~n50890 ) | ( n9760 & ~n50890 ) ;
  assign n50892 = ( ~n21402 & n50889 ) | ( ~n21402 & n50891 ) | ( n50889 & n50891 ) ;
  assign n50893 = ( n24254 & ~n24338 ) | ( n24254 & n27287 ) | ( ~n24338 & n27287 ) ;
  assign n50894 = ( n20060 & ~n43358 ) | ( n20060 & n45752 ) | ( ~n43358 & n45752 ) ;
  assign n50899 = ~n11449 & n17343 ;
  assign n50900 = n50899 ^ n16028 ^ n8290 ;
  assign n50898 = n26241 ^ n17293 ^ n5902 ;
  assign n50895 = n25713 ^ n16311 ^ n3843 ;
  assign n50896 = n3904 & ~n50895 ;
  assign n50897 = n1038 & n50896 ;
  assign n50901 = n50900 ^ n50898 ^ n50897 ;
  assign n50902 = n32667 ^ n28354 ^ n14203 ;
  assign n50903 = n45083 ^ n33231 ^ n4886 ;
  assign n50904 = n50903 ^ n21195 ^ n20572 ;
  assign n50905 = n50904 ^ n39957 ^ 1'b0 ;
  assign n50906 = n3150 | n29976 ;
  assign n50907 = n50906 ^ n5350 ^ 1'b0 ;
  assign n50908 = n21937 & ~n50907 ;
  assign n50909 = n30116 ^ n28450 ^ n8141 ;
  assign n50910 = n50909 ^ n28586 ^ n22215 ;
  assign n50911 = n31771 ^ n21633 ^ n3130 ;
  assign n50912 = ( n35465 & n44832 ) | ( n35465 & ~n50911 ) | ( n44832 & ~n50911 ) ;
  assign n50913 = n50912 ^ n4515 ^ 1'b0 ;
  assign n50914 = n4144 & ~n50913 ;
  assign n50915 = n16835 | n42692 ;
  assign n50916 = n50915 ^ n22961 ^ 1'b0 ;
  assign n50917 = n15184 & n50916 ;
  assign n50918 = n13485 | n30635 ;
  assign n50919 = ( ~n8980 & n18321 ) | ( ~n8980 & n23790 ) | ( n18321 & n23790 ) ;
  assign n50920 = n50919 ^ n4123 ^ n2530 ;
  assign n50921 = n50920 ^ n45679 ^ n19242 ;
  assign n50922 = n30291 ^ n623 ^ 1'b0 ;
  assign n50923 = ~n18614 & n50922 ;
  assign n50924 = ( n12884 & n17590 ) | ( n12884 & n50923 ) | ( n17590 & n50923 ) ;
  assign n50925 = n29829 ^ n10878 ^ n4925 ;
  assign n50926 = ( n8870 & ~n11263 ) | ( n8870 & n14161 ) | ( ~n11263 & n14161 ) ;
  assign n50927 = ( n2783 & ~n43137 ) | ( n2783 & n43926 ) | ( ~n43137 & n43926 ) ;
  assign n50928 = ( n11081 & n50926 ) | ( n11081 & ~n50927 ) | ( n50926 & ~n50927 ) ;
  assign n50929 = ( x168 & n7759 ) | ( x168 & n27506 ) | ( n7759 & n27506 ) ;
  assign n50930 = n50929 ^ n33561 ^ n26962 ;
  assign n50931 = ( n356 & n12903 ) | ( n356 & ~n50930 ) | ( n12903 & ~n50930 ) ;
  assign n50932 = ( n5660 & n6782 ) | ( n5660 & ~n39468 ) | ( n6782 & ~n39468 ) ;
  assign n50933 = ( n10543 & n26345 ) | ( n10543 & ~n30409 ) | ( n26345 & ~n30409 ) ;
  assign n50934 = ( n16408 & n50932 ) | ( n16408 & ~n50933 ) | ( n50932 & ~n50933 ) ;
  assign n50935 = ( n20829 & n24557 ) | ( n20829 & ~n26248 ) | ( n24557 & ~n26248 ) ;
  assign n50936 = n37799 & ~n50935 ;
  assign n50937 = n50934 & n50936 ;
  assign n50938 = ( ~n1476 & n29941 ) | ( ~n1476 & n50268 ) | ( n29941 & n50268 ) ;
  assign n50939 = ( n4468 & n30127 ) | ( n4468 & ~n50938 ) | ( n30127 & ~n50938 ) ;
  assign n50940 = ( n6022 & n21302 ) | ( n6022 & ~n40957 ) | ( n21302 & ~n40957 ) ;
  assign n50941 = n50940 ^ n45196 ^ n42417 ;
  assign n50942 = n15388 & ~n33943 ;
  assign n50943 = n12256 & n18865 ;
  assign n50944 = n50943 ^ n6014 ^ 1'b0 ;
  assign n50945 = n50944 ^ n31432 ^ n15944 ;
  assign n50946 = n25041 ^ n24557 ^ n4984 ;
  assign n50947 = n50946 ^ n42261 ^ n14076 ;
  assign n50948 = ( ~n15020 & n30832 ) | ( ~n15020 & n39837 ) | ( n30832 & n39837 ) ;
  assign n50949 = ( n26542 & n50947 ) | ( n26542 & n50948 ) | ( n50947 & n50948 ) ;
  assign n50950 = n46514 ^ n10567 ^ n1555 ;
  assign n50951 = n25770 & n40512 ;
  assign n50952 = n34064 ^ n18440 ^ 1'b0 ;
  assign n50953 = n7000 | n50952 ;
  assign n50954 = n50953 ^ n27532 ^ n21127 ;
  assign n50955 = n35372 ^ n13096 ^ n7883 ;
  assign n50956 = ( n14630 & n15117 ) | ( n14630 & ~n43939 ) | ( n15117 & ~n43939 ) ;
  assign n50957 = ( n33408 & n41476 ) | ( n33408 & n50956 ) | ( n41476 & n50956 ) ;
  assign n50958 = ( n22838 & n50955 ) | ( n22838 & n50957 ) | ( n50955 & n50957 ) ;
  assign n50959 = n6927 & n24784 ;
  assign n50960 = n18821 & n50959 ;
  assign n50961 = n8374 | n50818 ;
  assign n50962 = n50412 | n50961 ;
  assign n50963 = n29190 ^ n21645 ^ n20946 ;
  assign n50964 = n50963 ^ n30707 ^ n10306 ;
  assign n50965 = n50964 ^ n30691 ^ n23060 ;
  assign n50967 = ( n9219 & n16411 ) | ( n9219 & ~n18589 ) | ( n16411 & ~n18589 ) ;
  assign n50966 = ( n4244 & n4739 ) | ( n4244 & ~n24469 ) | ( n4739 & ~n24469 ) ;
  assign n50968 = n50967 ^ n50966 ^ n38103 ;
  assign n50969 = n21206 & n39606 ;
  assign n50970 = n5368 | n5726 ;
  assign n50971 = n50970 ^ n25796 ^ n9299 ;
  assign n50972 = n18657 & ~n37989 ;
  assign n50973 = n1279 & n50972 ;
  assign n50975 = n24846 ^ n1796 ^ 1'b0 ;
  assign n50976 = ~n20964 & n50975 ;
  assign n50974 = ( ~n34710 & n35267 ) | ( ~n34710 & n50508 ) | ( n35267 & n50508 ) ;
  assign n50977 = n50976 ^ n50974 ^ n7171 ;
  assign n50978 = ( n21672 & n50973 ) | ( n21672 & n50977 ) | ( n50973 & n50977 ) ;
  assign n50979 = n14900 & ~n37143 ;
  assign n50980 = n1982 & ~n18832 ;
  assign n50981 = n22279 & n50980 ;
  assign n50982 = n6514 ^ n394 ^ 1'b0 ;
  assign n50983 = ( n7899 & n21239 ) | ( n7899 & n29183 ) | ( n21239 & n29183 ) ;
  assign n50984 = n42656 ^ n26806 ^ n16454 ;
  assign n50985 = ( n19359 & ~n50983 ) | ( n19359 & n50984 ) | ( ~n50983 & n50984 ) ;
  assign n50986 = ( n7444 & n10237 ) | ( n7444 & ~n45286 ) | ( n10237 & ~n45286 ) ;
  assign n50987 = n38358 ^ n13628 ^ n8536 ;
  assign n50988 = ( n12519 & n16934 ) | ( n12519 & ~n50987 ) | ( n16934 & ~n50987 ) ;
  assign n50989 = n50988 ^ n38446 ^ n30437 ;
  assign n50990 = ( ~n14704 & n14705 ) | ( ~n14704 & n50989 ) | ( n14705 & n50989 ) ;
  assign n50991 = ( ~n394 & n37518 ) | ( ~n394 & n43650 ) | ( n37518 & n43650 ) ;
  assign n50992 = n50991 ^ n24765 ^ n10174 ;
  assign n50993 = n50992 ^ n47129 ^ n9377 ;
  assign n50994 = n26234 ^ n8240 ^ n3596 ;
  assign n50995 = ( n13190 & ~n40370 ) | ( n13190 & n40603 ) | ( ~n40370 & n40603 ) ;
  assign n50996 = ( ~n2984 & n10295 ) | ( ~n2984 & n19987 ) | ( n10295 & n19987 ) ;
  assign n50997 = ( n30227 & n48750 ) | ( n30227 & n50996 ) | ( n48750 & n50996 ) ;
  assign n50998 = ( n10161 & ~n13496 ) | ( n10161 & n16072 ) | ( ~n13496 & n16072 ) ;
  assign n50999 = ( ~n14122 & n17181 ) | ( ~n14122 & n19608 ) | ( n17181 & n19608 ) ;
  assign n51000 = ( n29737 & n50998 ) | ( n29737 & n50999 ) | ( n50998 & n50999 ) ;
  assign n51001 = ( n6090 & ~n50997 ) | ( n6090 & n51000 ) | ( ~n50997 & n51000 ) ;
  assign n51002 = ( x108 & n5177 ) | ( x108 & n25782 ) | ( n5177 & n25782 ) ;
  assign n51003 = n15624 ^ n10421 ^ n1830 ;
  assign n51004 = n51003 ^ n7847 ^ 1'b0 ;
  assign n51005 = ( n15050 & n51002 ) | ( n15050 & n51004 ) | ( n51002 & n51004 ) ;
  assign n51006 = n13179 | n21654 ;
  assign n51007 = n51006 ^ n18688 ^ 1'b0 ;
  assign n51008 = ~n16748 & n43328 ;
  assign n51009 = ~n51007 & n51008 ;
  assign n51010 = n27901 ^ n20749 ^ n1396 ;
  assign n51011 = ~n14786 & n51010 ;
  assign n51012 = n51011 ^ n33001 ^ 1'b0 ;
  assign n51013 = ( ~n5536 & n9147 ) | ( ~n5536 & n44604 ) | ( n9147 & n44604 ) ;
  assign n51014 = ( n7700 & n30287 ) | ( n7700 & ~n51013 ) | ( n30287 & ~n51013 ) ;
  assign n51015 = n22817 ^ n17551 ^ n14077 ;
  assign n51016 = ( n37886 & ~n50653 ) | ( n37886 & n51015 ) | ( ~n50653 & n51015 ) ;
  assign n51017 = n41809 ^ n23670 ^ n16932 ;
  assign n51018 = n9853 ^ n7425 ^ n1621 ;
  assign n51019 = ( n4109 & ~n14183 ) | ( n4109 & n33385 ) | ( ~n14183 & n33385 ) ;
  assign n51020 = ( n9885 & n36426 ) | ( n9885 & ~n51019 ) | ( n36426 & ~n51019 ) ;
  assign n51021 = ( n12304 & n51018 ) | ( n12304 & n51020 ) | ( n51018 & n51020 ) ;
  assign n51022 = n23882 ^ n7707 ^ n5214 ;
  assign n51023 = n37425 ^ n13790 ^ n5301 ;
  assign n51024 = ( n2042 & ~n44985 ) | ( n2042 & n51023 ) | ( ~n44985 & n51023 ) ;
  assign n51025 = n12212 ^ n7800 ^ n5852 ;
  assign n51026 = ( n2748 & n33041 ) | ( n2748 & n51025 ) | ( n33041 & n51025 ) ;
  assign n51027 = n17077 ^ n10116 ^ n8773 ;
  assign n51028 = ( ~n3240 & n10050 ) | ( ~n3240 & n46094 ) | ( n10050 & n46094 ) ;
  assign n51029 = ( n48957 & n49382 ) | ( n48957 & ~n51028 ) | ( n49382 & ~n51028 ) ;
  assign n51030 = n30615 ^ n18994 ^ n8325 ;
  assign n51031 = ( n17667 & ~n18255 ) | ( n17667 & n51030 ) | ( ~n18255 & n51030 ) ;
  assign n51032 = n51031 ^ n11560 ^ 1'b0 ;
  assign n51033 = n25274 & ~n51032 ;
  assign n51034 = n4785 ^ n4088 ^ 1'b0 ;
  assign n51035 = n10118 & n51034 ;
  assign n51036 = ( ~n5698 & n9504 ) | ( ~n5698 & n11079 ) | ( n9504 & n11079 ) ;
  assign n51037 = ( n20243 & n25274 ) | ( n20243 & ~n28269 ) | ( n25274 & ~n28269 ) ;
  assign n51038 = n51037 ^ n39364 ^ n5836 ;
  assign n51039 = n25874 | n40259 ;
  assign n51040 = n51039 ^ n36315 ^ n11925 ;
  assign n51041 = n45597 ^ n23538 ^ 1'b0 ;
  assign n51042 = n5101 | n51041 ;
  assign n51043 = n38894 ^ n28664 ^ n9159 ;
  assign n51044 = ( n37218 & ~n45111 ) | ( n37218 & n51043 ) | ( ~n45111 & n51043 ) ;
  assign n51045 = ( n48594 & ~n51042 ) | ( n48594 & n51044 ) | ( ~n51042 & n51044 ) ;
  assign n51046 = ( n417 & ~n14360 ) | ( n417 & n27888 ) | ( ~n14360 & n27888 ) ;
  assign n51047 = ~n17244 & n45511 ;
  assign n51048 = ~n35290 & n51047 ;
  assign n51049 = ( n40444 & ~n51046 ) | ( n40444 & n51048 ) | ( ~n51046 & n51048 ) ;
  assign n51051 = ( n3951 & n5954 ) | ( n3951 & ~n42976 ) | ( n5954 & ~n42976 ) ;
  assign n51052 = n51051 ^ n49504 ^ n19449 ;
  assign n51050 = ( n7295 & ~n28741 ) | ( n7295 & n40292 ) | ( ~n28741 & n40292 ) ;
  assign n51053 = n51052 ^ n51050 ^ n49231 ;
  assign n51054 = n5060 & n6780 ;
  assign n51055 = ( n4967 & n44650 ) | ( n4967 & n51054 ) | ( n44650 & n51054 ) ;
  assign n51056 = ( n25921 & n33734 ) | ( n25921 & ~n51055 ) | ( n33734 & ~n51055 ) ;
  assign n51057 = n51056 ^ n46543 ^ n28484 ;
  assign n51058 = ( n12539 & n16520 ) | ( n12539 & ~n24478 ) | ( n16520 & ~n24478 ) ;
  assign n51059 = n7085 ^ n2643 ^ 1'b0 ;
  assign n51060 = n11706 & ~n51059 ;
  assign n51061 = ( n3497 & n20876 ) | ( n3497 & ~n51060 ) | ( n20876 & ~n51060 ) ;
  assign n51062 = n7894 & ~n45477 ;
  assign n51063 = ~n29009 & n51062 ;
  assign n51064 = ( n5592 & n6223 ) | ( n5592 & n15953 ) | ( n6223 & n15953 ) ;
  assign n51065 = n17867 | n25377 ;
  assign n51066 = n25377 & ~n51065 ;
  assign n51067 = ( n24922 & n32741 ) | ( n24922 & n51066 ) | ( n32741 & n51066 ) ;
  assign n51068 = n51067 ^ n25094 ^ n5324 ;
  assign n51069 = n51068 ^ n22701 ^ n20370 ;
  assign n51070 = n34220 & ~n51069 ;
  assign n51071 = ( n26488 & ~n31037 ) | ( n26488 & n44348 ) | ( ~n31037 & n44348 ) ;
  assign n51072 = n51071 ^ n13185 ^ n1887 ;
  assign n51073 = ( n6249 & ~n19736 ) | ( n6249 & n20031 ) | ( ~n19736 & n20031 ) ;
  assign n51074 = ( n9063 & ~n48008 ) | ( n9063 & n51073 ) | ( ~n48008 & n51073 ) ;
  assign n51077 = n16334 ^ n14457 ^ n8227 ;
  assign n51078 = ( n11237 & n11652 ) | ( n11237 & n51077 ) | ( n11652 & n51077 ) ;
  assign n51075 = ( ~n5004 & n10022 ) | ( ~n5004 & n11021 ) | ( n10022 & n11021 ) ;
  assign n51076 = n51075 ^ n13961 ^ n8103 ;
  assign n51079 = n51078 ^ n51076 ^ x152 ;
  assign n51080 = n26369 & n49907 ;
  assign n51081 = ~n28093 & n42880 ;
  assign n51082 = n18916 | n51081 ;
  assign n51083 = ( n22416 & ~n33088 ) | ( n22416 & n37726 ) | ( ~n33088 & n37726 ) ;
  assign n51084 = n51083 ^ n23028 ^ 1'b0 ;
  assign n51085 = n25477 ^ n14566 ^ n11051 ;
  assign n51086 = n51085 ^ n36657 ^ n24655 ;
  assign n51087 = n45750 ^ n22273 ^ 1'b0 ;
  assign n51088 = n31017 | n51087 ;
  assign n51089 = n14057 | n51088 ;
  assign n51090 = n51089 ^ n18561 ^ 1'b0 ;
  assign n51091 = x153 & ~n11705 ;
  assign n51092 = n51091 ^ n22587 ^ 1'b0 ;
  assign n51093 = ( n2787 & n25436 ) | ( n2787 & ~n38242 ) | ( n25436 & ~n38242 ) ;
  assign n51094 = ( n1533 & n21535 ) | ( n1533 & ~n51093 ) | ( n21535 & ~n51093 ) ;
  assign n51095 = n44543 ^ n40711 ^ n26671 ;
  assign n51096 = n34569 ^ n9333 ^ n2081 ;
  assign n51097 = n45150 ^ n37249 ^ n13711 ;
  assign n51098 = ( n14805 & ~n16220 ) | ( n14805 & n51097 ) | ( ~n16220 & n51097 ) ;
  assign n51099 = ~n12001 & n51098 ;
  assign n51100 = n51099 ^ n3409 ^ 1'b0 ;
  assign n51101 = n51100 ^ n34286 ^ n15205 ;
  assign n51102 = ( ~n8281 & n51096 ) | ( ~n8281 & n51101 ) | ( n51096 & n51101 ) ;
  assign n51103 = n26775 ^ n11922 ^ n3393 ;
  assign n51104 = ( n1766 & ~n5683 ) | ( n1766 & n47481 ) | ( ~n5683 & n47481 ) ;
  assign n51105 = n22583 ^ n12904 ^ n4653 ;
  assign n51106 = n51105 ^ n37778 ^ n27589 ;
  assign n51107 = ( n8957 & n12274 ) | ( n8957 & ~n33092 ) | ( n12274 & ~n33092 ) ;
  assign n51108 = ( n21115 & n28670 ) | ( n21115 & ~n51107 ) | ( n28670 & ~n51107 ) ;
  assign n51109 = n51108 ^ n48571 ^ n15735 ;
  assign n51110 = n28363 ^ n449 ^ 1'b0 ;
  assign n51111 = n7338 | n51110 ;
  assign n51112 = n15299 | n32671 ;
  assign n51113 = n2011 & ~n51112 ;
  assign n51114 = n36495 & n43786 ;
  assign n51115 = ( n7858 & n40273 ) | ( n7858 & ~n51114 ) | ( n40273 & ~n51114 ) ;
  assign n51116 = ( n40022 & ~n49285 ) | ( n40022 & n51115 ) | ( ~n49285 & n51115 ) ;
  assign n51117 = ( ~n5082 & n5808 ) | ( ~n5082 & n7592 ) | ( n5808 & n7592 ) ;
  assign n51118 = n51117 ^ n8465 ^ n6326 ;
  assign n51119 = ~n2014 & n8464 ;
  assign n51120 = n51119 ^ n14579 ^ 1'b0 ;
  assign n51121 = n51120 ^ n33531 ^ n19694 ;
  assign n51122 = ( n16867 & n51118 ) | ( n16867 & ~n51121 ) | ( n51118 & ~n51121 ) ;
  assign n51125 = ( n5983 & ~n7506 ) | ( n5983 & n13563 ) | ( ~n7506 & n13563 ) ;
  assign n51126 = ( ~n22615 & n43370 ) | ( ~n22615 & n51125 ) | ( n43370 & n51125 ) ;
  assign n51127 = n51126 ^ n31844 ^ 1'b0 ;
  assign n51124 = ( n1388 & n16105 ) | ( n1388 & n30428 ) | ( n16105 & n30428 ) ;
  assign n51128 = n51127 ^ n51124 ^ n606 ;
  assign n51123 = ( n14976 & n21961 ) | ( n14976 & n29558 ) | ( n21961 & n29558 ) ;
  assign n51129 = n51128 ^ n51123 ^ n45665 ;
  assign n51130 = ( n4210 & n11595 ) | ( n4210 & n35970 ) | ( n11595 & n35970 ) ;
  assign n51131 = n39525 ^ n27595 ^ n13867 ;
  assign n51132 = ( n6753 & ~n36974 ) | ( n6753 & n51131 ) | ( ~n36974 & n51131 ) ;
  assign n51133 = ( n18072 & n40885 ) | ( n18072 & n51132 ) | ( n40885 & n51132 ) ;
  assign n51134 = ( n13291 & ~n14427 ) | ( n13291 & n46278 ) | ( ~n14427 & n46278 ) ;
  assign n51135 = ( ~n14325 & n22883 ) | ( ~n14325 & n51134 ) | ( n22883 & n51134 ) ;
  assign n51136 = n51133 & n51135 ;
  assign n51137 = n28102 ^ n26658 ^ n17054 ;
  assign n51138 = n51137 ^ n18902 ^ n12264 ;
  assign n51139 = ( n6826 & n25683 ) | ( n6826 & ~n48377 ) | ( n25683 & ~n48377 ) ;
  assign n51140 = n51139 ^ n38021 ^ n27102 ;
  assign n51141 = n4377 & n19854 ;
  assign n51142 = ( n1626 & n7952 ) | ( n1626 & n34686 ) | ( n7952 & n34686 ) ;
  assign n51143 = n51142 ^ n20683 ^ n9895 ;
  assign n51144 = n23987 ^ n9496 ^ 1'b0 ;
  assign n51145 = ~n12611 & n51144 ;
  assign n51148 = n36450 ^ n24148 ^ n6023 ;
  assign n51149 = ( n5782 & n27125 ) | ( n5782 & ~n51148 ) | ( n27125 & ~n51148 ) ;
  assign n51147 = n12943 & n39090 ;
  assign n51150 = n51149 ^ n51147 ^ 1'b0 ;
  assign n51151 = n7763 & n51150 ;
  assign n51152 = n51151 ^ n37877 ^ 1'b0 ;
  assign n51146 = n41543 ^ n28136 ^ n18966 ;
  assign n51153 = n51152 ^ n51146 ^ n3005 ;
  assign n51154 = ( ~n2974 & n11341 ) | ( ~n2974 & n50221 ) | ( n11341 & n50221 ) ;
  assign n51155 = n51154 ^ n12545 ^ n2060 ;
  assign n51156 = n24059 ^ n11883 ^ n1649 ;
  assign n51160 = n23381 ^ n20923 ^ n3496 ;
  assign n51157 = ( n8283 & n19471 ) | ( n8283 & ~n32020 ) | ( n19471 & ~n32020 ) ;
  assign n51158 = n51157 ^ n10679 ^ n546 ;
  assign n51159 = ( n18642 & n49978 ) | ( n18642 & ~n51158 ) | ( n49978 & ~n51158 ) ;
  assign n51161 = n51160 ^ n51159 ^ n24743 ;
  assign n51162 = ( ~n11291 & n29721 ) | ( ~n11291 & n51161 ) | ( n29721 & n51161 ) ;
  assign n51164 = n10141 & n16228 ;
  assign n51165 = n51164 ^ n6748 ^ 1'b0 ;
  assign n51163 = n30993 ^ n21702 ^ n14332 ;
  assign n51166 = n51165 ^ n51163 ^ n32799 ;
  assign n51167 = n40286 ^ n16609 ^ n5477 ;
  assign n51168 = ( n24773 & ~n34052 ) | ( n24773 & n40761 ) | ( ~n34052 & n40761 ) ;
  assign n51169 = n11654 & n31284 ;
  assign n51170 = n33743 ^ n10885 ^ n10794 ;
  assign n51171 = n7487 & ~n37391 ;
  assign n51172 = n51171 ^ n18869 ^ 1'b0 ;
  assign n51173 = n30857 ^ n1206 ^ 1'b0 ;
  assign n51174 = n42848 | n51173 ;
  assign n51175 = n39340 ^ n38892 ^ n15193 ;
  assign n51176 = n48773 ^ n48055 ^ n36904 ;
  assign n51178 = ( n14791 & n20911 ) | ( n14791 & n27745 ) | ( n20911 & n27745 ) ;
  assign n51177 = n50817 ^ n45604 ^ n41411 ;
  assign n51179 = n51178 ^ n51177 ^ n27987 ;
  assign n51180 = ( n8284 & n32084 ) | ( n8284 & n51179 ) | ( n32084 & n51179 ) ;
  assign n51181 = n51180 ^ n42367 ^ n28220 ;
  assign n51182 = n51181 ^ n50272 ^ n13341 ;
  assign n51183 = n28136 ^ n12983 ^ n11485 ;
  assign n51184 = ( n23137 & ~n29357 ) | ( n23137 & n51183 ) | ( ~n29357 & n51183 ) ;
  assign n51185 = ( n8340 & n21850 ) | ( n8340 & ~n51184 ) | ( n21850 & ~n51184 ) ;
  assign n51186 = n42656 ^ n16189 ^ n11897 ;
  assign n51187 = ( n10340 & n20094 ) | ( n10340 & ~n51186 ) | ( n20094 & ~n51186 ) ;
  assign n51188 = ( n3030 & ~n3540 ) | ( n3030 & n10197 ) | ( ~n3540 & n10197 ) ;
  assign n51189 = n16071 | n27817 ;
  assign n51190 = n51189 ^ n8990 ^ 1'b0 ;
  assign n51191 = n51190 ^ n23220 ^ n10811 ;
  assign n51192 = ( n15401 & n51188 ) | ( n15401 & n51191 ) | ( n51188 & n51191 ) ;
  assign n51193 = n2502 & n43434 ;
  assign n51194 = n51193 ^ n25110 ^ 1'b0 ;
  assign n51195 = n51194 ^ n18402 ^ n16757 ;
  assign n51197 = n18603 ^ n9272 ^ n6874 ;
  assign n51196 = ( n5101 & n24653 ) | ( n5101 & n28972 ) | ( n24653 & n28972 ) ;
  assign n51198 = n51197 ^ n51196 ^ n24537 ;
  assign n51199 = ( n18583 & n29354 ) | ( n18583 & ~n43201 ) | ( n29354 & ~n43201 ) ;
  assign n51200 = n2518 & n51199 ;
  assign n51201 = ~n12275 & n51200 ;
  assign n51202 = n39368 ^ n28750 ^ n3488 ;
  assign n51203 = ( n3526 & n15102 ) | ( n3526 & ~n33536 ) | ( n15102 & ~n33536 ) ;
  assign n51204 = n22743 ^ n9996 ^ 1'b0 ;
  assign n51205 = n46699 ^ n38361 ^ n19802 ;
  assign n51206 = ( n9658 & ~n51204 ) | ( n9658 & n51205 ) | ( ~n51204 & n51205 ) ;
  assign n51207 = n31335 ^ n12228 ^ n5292 ;
  assign n51208 = ( ~n10278 & n31409 ) | ( ~n10278 & n34843 ) | ( n31409 & n34843 ) ;
  assign n51209 = ( ~n2916 & n32547 ) | ( ~n2916 & n51208 ) | ( n32547 & n51208 ) ;
  assign n51210 = n9879 & n51209 ;
  assign n51211 = ( n1344 & n12880 ) | ( n1344 & n20563 ) | ( n12880 & n20563 ) ;
  assign n51213 = ( n990 & n2374 ) | ( n990 & n4306 ) | ( n2374 & n4306 ) ;
  assign n51212 = ( n6559 & ~n24450 ) | ( n6559 & n50216 ) | ( ~n24450 & n50216 ) ;
  assign n51214 = n51213 ^ n51212 ^ n11677 ;
  assign n51215 = n38495 ^ n29765 ^ n21511 ;
  assign n51216 = n27974 ^ n10975 ^ n7597 ;
  assign n51217 = ( ~n31803 & n33022 ) | ( ~n31803 & n43278 ) | ( n33022 & n43278 ) ;
  assign n51218 = ( ~n29531 & n51216 ) | ( ~n29531 & n51217 ) | ( n51216 & n51217 ) ;
  assign n51219 = n15549 & n24018 ;
  assign n51220 = ( n4480 & n14012 ) | ( n4480 & n51219 ) | ( n14012 & n51219 ) ;
  assign n51221 = ~n26761 & n51220 ;
  assign n51222 = n23365 & n51221 ;
  assign n51225 = ( n767 & n2659 ) | ( n767 & n6045 ) | ( n2659 & n6045 ) ;
  assign n51223 = ( ~n8097 & n26508 ) | ( ~n8097 & n48043 ) | ( n26508 & n48043 ) ;
  assign n51224 = n51223 ^ n26968 ^ n10271 ;
  assign n51226 = n51225 ^ n51224 ^ n12064 ;
  assign n51227 = ( n8822 & ~n9741 ) | ( n8822 & n19978 ) | ( ~n9741 & n19978 ) ;
  assign n51228 = ( n34206 & n35929 ) | ( n34206 & n51227 ) | ( n35929 & n51227 ) ;
  assign n51229 = ( n1584 & n18636 ) | ( n1584 & ~n42770 ) | ( n18636 & ~n42770 ) ;
  assign n51230 = ( n2272 & n14828 ) | ( n2272 & n51229 ) | ( n14828 & n51229 ) ;
  assign n51231 = ( n3686 & n6340 ) | ( n3686 & ~n22125 ) | ( n6340 & ~n22125 ) ;
  assign n51232 = n34162 ^ n25521 ^ n19025 ;
  assign n51233 = n41337 ^ n35062 ^ n33193 ;
  assign n51234 = ( n10704 & ~n25164 ) | ( n10704 & n51233 ) | ( ~n25164 & n51233 ) ;
  assign n51235 = ( ~n26188 & n32329 ) | ( ~n26188 & n51234 ) | ( n32329 & n51234 ) ;
  assign n51236 = n48805 ^ n43319 ^ n26247 ;
  assign n51237 = ( ~n11585 & n11770 ) | ( ~n11585 & n27111 ) | ( n11770 & n27111 ) ;
  assign n51238 = n36741 ^ n13648 ^ n3995 ;
  assign n51239 = n42437 ^ n26479 ^ n20494 ;
  assign n51240 = n51239 ^ n12231 ^ n4383 ;
  assign n51241 = ( n3632 & ~n11934 ) | ( n3632 & n51240 ) | ( ~n11934 & n51240 ) ;
  assign n51242 = n33217 ^ n23759 ^ n20567 ;
  assign n51243 = n44670 ^ n7511 ^ x56 ;
  assign n51244 = ( ~n16820 & n26414 ) | ( ~n16820 & n51081 ) | ( n26414 & n51081 ) ;
  assign n51245 = n48657 ^ n14728 ^ 1'b0 ;
  assign n51246 = n38835 ^ n21377 ^ 1'b0 ;
  assign n51247 = ( n19851 & n47681 ) | ( n19851 & n51246 ) | ( n47681 & n51246 ) ;
  assign n51248 = ( n8960 & ~n50854 ) | ( n8960 & n51247 ) | ( ~n50854 & n51247 ) ;
  assign n51249 = n22902 ^ n7159 ^ 1'b0 ;
  assign n51250 = n2853 & n12274 ;
  assign n51251 = n51250 ^ n5085 ^ n4832 ;
  assign n51253 = n19736 ^ n5728 ^ n2292 ;
  assign n51252 = ( n20619 & ~n27817 ) | ( n20619 & n31544 ) | ( ~n27817 & n31544 ) ;
  assign n51254 = n51253 ^ n51252 ^ n16904 ;
  assign n51255 = n32741 ^ n30178 ^ 1'b0 ;
  assign n51256 = n20598 ^ n20468 ^ 1'b0 ;
  assign n51257 = n42855 ^ n12948 ^ 1'b0 ;
  assign n51258 = n31644 & ~n51257 ;
  assign n51259 = n20597 ^ n4178 ^ n2406 ;
  assign n51260 = n36307 ^ n16195 ^ 1'b0 ;
  assign n51261 = ( n16414 & n36691 ) | ( n16414 & n51260 ) | ( n36691 & n51260 ) ;
  assign n51262 = n41474 ^ n2761 ^ n473 ;
  assign n51263 = n2010 & ~n16796 ;
  assign n51264 = n51263 ^ n35780 ^ 1'b0 ;
  assign n51265 = n15624 ^ n7901 ^ 1'b0 ;
  assign n51266 = n34728 ^ n2637 ^ 1'b0 ;
  assign n51267 = ( ~n9038 & n9095 ) | ( ~n9038 & n51266 ) | ( n9095 & n51266 ) ;
  assign n51268 = ( ~n46240 & n51265 ) | ( ~n46240 & n51267 ) | ( n51265 & n51267 ) ;
  assign n51269 = ( n14234 & n40522 ) | ( n14234 & ~n44207 ) | ( n40522 & ~n44207 ) ;
  assign n51270 = ( n4394 & n5622 ) | ( n4394 & n19922 ) | ( n5622 & n19922 ) ;
  assign n51271 = n39055 & ~n51270 ;
  assign n51272 = n48360 ^ n20916 ^ n10652 ;
  assign n51275 = n4389 ^ n3094 ^ n632 ;
  assign n51276 = ( n7756 & n10261 ) | ( n7756 & ~n51275 ) | ( n10261 & ~n51275 ) ;
  assign n51277 = ( n1328 & n5470 ) | ( n1328 & ~n51276 ) | ( n5470 & ~n51276 ) ;
  assign n51273 = n25839 ^ n8354 ^ n1056 ;
  assign n51274 = n51273 ^ n6035 ^ 1'b0 ;
  assign n51278 = n51277 ^ n51274 ^ n35156 ;
  assign n51279 = n25360 ^ n567 ^ 1'b0 ;
  assign n51280 = n27299 ^ n16440 ^ n13459 ;
  assign n51281 = ( n6191 & n25220 ) | ( n6191 & ~n30502 ) | ( n25220 & ~n30502 ) ;
  assign n51282 = n51281 ^ n5327 ^ n2598 ;
  assign n51283 = n836 & n8004 ;
  assign n51284 = n51283 ^ n37739 ^ 1'b0 ;
  assign n51285 = n42100 & n51284 ;
  assign n51286 = ~n29124 & n51285 ;
  assign n51287 = ( n1208 & n15603 ) | ( n1208 & n33170 ) | ( n15603 & n33170 ) ;
  assign n51288 = n9241 & n49062 ;
  assign n51289 = n25208 & ~n40906 ;
  assign n51290 = n1824 & ~n34688 ;
  assign n51291 = ( n9421 & n23413 ) | ( n9421 & n51290 ) | ( n23413 & n51290 ) ;
  assign n51292 = ( n19861 & ~n36913 ) | ( n19861 & n40487 ) | ( ~n36913 & n40487 ) ;
  assign n51293 = ( ~n24957 & n37372 ) | ( ~n24957 & n38903 ) | ( n37372 & n38903 ) ;
  assign n51294 = ( n4020 & n6028 ) | ( n4020 & ~n13942 ) | ( n6028 & ~n13942 ) ;
  assign n51295 = ( ~n22669 & n44158 ) | ( ~n22669 & n51294 ) | ( n44158 & n51294 ) ;
  assign n51296 = n41383 ^ n11054 ^ 1'b0 ;
  assign n51297 = n2223 | n43636 ;
  assign n51298 = n28934 | n51297 ;
  assign n51299 = ( n7539 & n11258 ) | ( n7539 & ~n26368 ) | ( n11258 & ~n26368 ) ;
  assign n51300 = n38580 ^ n34885 ^ 1'b0 ;
  assign n51301 = n35438 ^ n12422 ^ n3391 ;
  assign n51302 = ( n22952 & n49875 ) | ( n22952 & n51301 ) | ( n49875 & n51301 ) ;
  assign n51303 = ( ~n2864 & n51300 ) | ( ~n2864 & n51302 ) | ( n51300 & n51302 ) ;
  assign n51304 = ( n7105 & n8838 ) | ( n7105 & n24043 ) | ( n8838 & n24043 ) ;
  assign n51305 = ( ~n15952 & n38270 ) | ( ~n15952 & n42218 ) | ( n38270 & n42218 ) ;
  assign n51312 = n25283 ^ n13527 ^ 1'b0 ;
  assign n51313 = n51312 ^ n16548 ^ n4644 ;
  assign n51314 = n51313 ^ n22406 ^ n3668 ;
  assign n51307 = ( n3342 & ~n3843 ) | ( n3342 & n19250 ) | ( ~n3843 & n19250 ) ;
  assign n51308 = n51307 ^ n7591 ^ n6097 ;
  assign n51309 = n51308 ^ n47526 ^ n6244 ;
  assign n51310 = n51309 ^ n20715 ^ n2507 ;
  assign n51306 = ( n4417 & n25259 ) | ( n4417 & ~n30222 ) | ( n25259 & ~n30222 ) ;
  assign n51311 = n51310 ^ n51306 ^ 1'b0 ;
  assign n51315 = n51314 ^ n51311 ^ n21896 ;
  assign n51316 = n36590 ^ n6964 ^ n6160 ;
  assign n51317 = n16043 & n51316 ;
  assign n51318 = ( n12192 & n29020 ) | ( n12192 & n41298 ) | ( n29020 & n41298 ) ;
  assign n51319 = n51318 ^ n20533 ^ n20425 ;
  assign n51320 = n22869 ^ n8099 ^ n6440 ;
  assign n51321 = n51320 ^ n20540 ^ n7962 ;
  assign n51322 = n51321 ^ n17366 ^ n14352 ;
  assign n51323 = n20782 | n24638 ;
  assign n51324 = n42953 ^ n23251 ^ n12125 ;
  assign n51325 = ( ~n4867 & n10638 ) | ( ~n4867 & n15576 ) | ( n10638 & n15576 ) ;
  assign n51326 = ( ~n262 & n14639 ) | ( ~n262 & n51325 ) | ( n14639 & n51325 ) ;
  assign n51327 = n51326 ^ n15570 ^ n14136 ;
  assign n51328 = ( n19905 & ~n33628 ) | ( n19905 & n51327 ) | ( ~n33628 & n51327 ) ;
  assign n51329 = ( n10624 & n12864 ) | ( n10624 & ~n51328 ) | ( n12864 & ~n51328 ) ;
  assign n51330 = ( n5024 & n5283 ) | ( n5024 & n15579 ) | ( n5283 & n15579 ) ;
  assign n51331 = n51330 ^ n22348 ^ n1293 ;
  assign n51332 = n51331 ^ n25135 ^ n19684 ;
  assign n51335 = n38318 ^ n27430 ^ n17770 ;
  assign n51336 = ( ~n733 & n33815 ) | ( ~n733 & n51335 ) | ( n33815 & n51335 ) ;
  assign n51333 = n45886 ^ n17069 ^ n2069 ;
  assign n51334 = n51333 ^ n31947 ^ n12674 ;
  assign n51337 = n51336 ^ n51334 ^ n1609 ;
  assign n51338 = ( n4642 & ~n14045 ) | ( n4642 & n22082 ) | ( ~n14045 & n22082 ) ;
  assign n51339 = n51338 ^ n14884 ^ n14653 ;
  assign n51340 = ~n7312 & n12955 ;
  assign n51341 = n51340 ^ n44446 ^ n17110 ;
  assign n51342 = n4212 & ~n16267 ;
  assign n51343 = n16932 & n51342 ;
  assign n51344 = n22218 ^ n20163 ^ n11060 ;
  assign n51345 = n45475 ^ n25896 ^ n23464 ;
  assign n51347 = n19623 ^ n14977 ^ n12886 ;
  assign n51348 = ( ~n34329 & n37158 ) | ( ~n34329 & n51347 ) | ( n37158 & n51347 ) ;
  assign n51346 = n27016 ^ n20249 ^ n15036 ;
  assign n51349 = n51348 ^ n51346 ^ n11948 ;
  assign n51350 = ( n28004 & n36758 ) | ( n28004 & n51349 ) | ( n36758 & n51349 ) ;
  assign n51352 = ( ~n4784 & n7522 ) | ( ~n4784 & n47311 ) | ( n7522 & n47311 ) ;
  assign n51351 = n40476 ^ n33100 ^ n28727 ;
  assign n51353 = n51352 ^ n51351 ^ n28659 ;
  assign n51354 = ( n8738 & ~n43162 ) | ( n8738 & n50401 ) | ( ~n43162 & n50401 ) ;
  assign n51355 = ( n6958 & ~n11389 ) | ( n6958 & n11722 ) | ( ~n11389 & n11722 ) ;
  assign n51356 = ( n23528 & ~n51354 ) | ( n23528 & n51355 ) | ( ~n51354 & n51355 ) ;
  assign n51357 = ( n14256 & n24009 ) | ( n14256 & ~n28822 ) | ( n24009 & ~n28822 ) ;
  assign n51358 = ( n6426 & n12454 ) | ( n6426 & ~n21249 ) | ( n12454 & ~n21249 ) ;
  assign n51359 = ( n16325 & ~n26908 ) | ( n16325 & n46459 ) | ( ~n26908 & n46459 ) ;
  assign n51360 = n13470 & ~n51359 ;
  assign n51361 = n51360 ^ n38822 ^ 1'b0 ;
  assign n51364 = n5122 ^ n1049 ^ 1'b0 ;
  assign n51365 = n49113 & n51364 ;
  assign n51363 = ( n8724 & ~n18817 ) | ( n8724 & n28220 ) | ( ~n18817 & n28220 ) ;
  assign n51362 = ( n20534 & n37970 ) | ( n20534 & ~n51227 ) | ( n37970 & ~n51227 ) ;
  assign n51366 = n51365 ^ n51363 ^ n51362 ;
  assign n51367 = ( x226 & ~n4238 ) | ( x226 & n37204 ) | ( ~n4238 & n37204 ) ;
  assign n51368 = n28329 ^ n22027 ^ n5414 ;
  assign n51369 = ( n5156 & ~n10634 ) | ( n5156 & n33494 ) | ( ~n10634 & n33494 ) ;
  assign n51370 = ( n29255 & n39309 ) | ( n29255 & ~n51369 ) | ( n39309 & ~n51369 ) ;
  assign n51371 = n40468 ^ n6351 ^ n3679 ;
  assign n51372 = ( n19615 & ~n30253 ) | ( n19615 & n51371 ) | ( ~n30253 & n51371 ) ;
  assign n51373 = n51372 ^ n27396 ^ n23760 ;
  assign n51374 = ( n1118 & ~n19370 ) | ( n1118 & n32487 ) | ( ~n19370 & n32487 ) ;
  assign n51375 = ( n2838 & n11329 ) | ( n2838 & n51374 ) | ( n11329 & n51374 ) ;
  assign n51376 = ( n21567 & n22028 ) | ( n21567 & n46434 ) | ( n22028 & n46434 ) ;
  assign n51377 = n33531 ^ n16253 ^ n16252 ;
  assign n51378 = ~n27530 & n51377 ;
  assign n51379 = ~n10050 & n51378 ;
  assign n51380 = n51379 ^ n30844 ^ 1'b0 ;
  assign n51381 = n33281 ^ n21878 ^ n16059 ;
  assign n51382 = n18581 ^ n16069 ^ n15501 ;
  assign n51383 = ( n11477 & n35744 ) | ( n11477 & n51382 ) | ( n35744 & n51382 ) ;
  assign n51384 = ( n32694 & n51381 ) | ( n32694 & n51383 ) | ( n51381 & n51383 ) ;
  assign n51385 = n25112 ^ n4298 ^ 1'b0 ;
  assign n51386 = n14989 & n51385 ;
  assign n51387 = n10279 | n27130 ;
  assign n51388 = n9601 | n51387 ;
  assign n51389 = n39936 ^ n14469 ^ 1'b0 ;
  assign n51390 = ~n26952 & n51389 ;
  assign n51391 = ( n13014 & n44784 ) | ( n13014 & n51390 ) | ( n44784 & n51390 ) ;
  assign n51392 = n43260 ^ n24203 ^ n14166 ;
  assign n51394 = ( n1801 & ~n4447 ) | ( n1801 & n11528 ) | ( ~n4447 & n11528 ) ;
  assign n51393 = n39470 ^ n39076 ^ n17407 ;
  assign n51395 = n51394 ^ n51393 ^ n4851 ;
  assign n51396 = ( n3891 & ~n19267 ) | ( n3891 & n50903 ) | ( ~n19267 & n50903 ) ;
  assign n51397 = ( n17583 & ~n41636 ) | ( n17583 & n44505 ) | ( ~n41636 & n44505 ) ;
  assign n51398 = ( n15643 & ~n22548 ) | ( n15643 & n37093 ) | ( ~n22548 & n37093 ) ;
  assign n51399 = n51398 ^ n39384 ^ 1'b0 ;
  assign n51400 = ( n8623 & n21994 ) | ( n8623 & n22831 ) | ( n21994 & n22831 ) ;
  assign n51401 = ( ~n21093 & n41268 ) | ( ~n21093 & n51400 ) | ( n41268 & n51400 ) ;
  assign n51403 = ( n2265 & n10776 ) | ( n2265 & ~n17951 ) | ( n10776 & ~n17951 ) ;
  assign n51402 = n33516 ^ n30209 ^ n21567 ;
  assign n51404 = n51403 ^ n51402 ^ n11775 ;
  assign n51405 = ( n5838 & ~n8208 ) | ( n5838 & n33317 ) | ( ~n8208 & n33317 ) ;
  assign n51406 = n51405 ^ n40483 ^ n7306 ;
  assign n51407 = n36900 ^ n12579 ^ 1'b0 ;
  assign n51408 = ( n5958 & n14662 ) | ( n5958 & n36152 ) | ( n14662 & n36152 ) ;
  assign n51409 = n51408 ^ n32969 ^ n5888 ;
  assign n51410 = n25703 & ~n51409 ;
  assign n51411 = ( n17542 & n18123 ) | ( n17542 & ~n24991 ) | ( n18123 & ~n24991 ) ;
  assign n51412 = ( n17704 & n30023 ) | ( n17704 & n51411 ) | ( n30023 & n51411 ) ;
  assign n51413 = n11611 ^ n6409 ^ n5193 ;
  assign n51414 = ( n1666 & n30931 ) | ( n1666 & ~n51413 ) | ( n30931 & ~n51413 ) ;
  assign n51415 = n51414 ^ n16681 ^ n3152 ;
  assign n51416 = ( ~n19466 & n50585 ) | ( ~n19466 & n51415 ) | ( n50585 & n51415 ) ;
  assign n51417 = ( n12915 & ~n27518 ) | ( n12915 & n28642 ) | ( ~n27518 & n28642 ) ;
  assign n51418 = n51417 ^ n3015 ^ n1452 ;
  assign n51419 = n39532 ^ n29526 ^ n7390 ;
  assign n51420 = ( n7706 & ~n9257 ) | ( n7706 & n31752 ) | ( ~n9257 & n31752 ) ;
  assign n51421 = n51420 ^ n10431 ^ n8226 ;
  assign n51422 = ( ~n7441 & n20597 ) | ( ~n7441 & n38736 ) | ( n20597 & n38736 ) ;
  assign n51423 = n41344 ^ n23604 ^ n4932 ;
  assign n51424 = ( ~n12936 & n48339 ) | ( ~n12936 & n51423 ) | ( n48339 & n51423 ) ;
  assign n51425 = ( x192 & n51422 ) | ( x192 & n51424 ) | ( n51422 & n51424 ) ;
  assign n51426 = n14231 & ~n41621 ;
  assign n51427 = n51426 ^ n10137 ^ 1'b0 ;
  assign n51428 = n13918 ^ n12636 ^ 1'b0 ;
  assign n51429 = n27189 | n51428 ;
  assign n51430 = n49383 ^ n48353 ^ n10808 ;
  assign n51431 = n8276 & ~n9026 ;
  assign n51432 = n51431 ^ n4739 ^ 1'b0 ;
  assign n51433 = ( n664 & ~n1403 ) | ( n664 & n51432 ) | ( ~n1403 & n51432 ) ;
  assign n51438 = ( ~n22810 & n23102 ) | ( ~n22810 & n47127 ) | ( n23102 & n47127 ) ;
  assign n51435 = ( n5649 & n16042 ) | ( n5649 & ~n28745 ) | ( n16042 & ~n28745 ) ;
  assign n51434 = n32710 ^ n31272 ^ n23020 ;
  assign n51436 = n51435 ^ n51434 ^ n9281 ;
  assign n51437 = n51436 ^ n35207 ^ n1724 ;
  assign n51439 = n51438 ^ n51437 ^ n39040 ;
  assign n51440 = ( ~n13349 & n15421 ) | ( ~n13349 & n35857 ) | ( n15421 & n35857 ) ;
  assign n51441 = ( n36058 & n43399 ) | ( n36058 & ~n49860 ) | ( n43399 & ~n49860 ) ;
  assign n51442 = ( n11216 & ~n20186 ) | ( n11216 & n21370 ) | ( ~n20186 & n21370 ) ;
  assign n51443 = n25318 ^ n4897 ^ n3654 ;
  assign n51444 = n51443 ^ n45663 ^ n6807 ;
  assign n51445 = n13354 ^ n5660 ^ n2159 ;
  assign n51446 = ( n20407 & n20743 ) | ( n20407 & ~n40957 ) | ( n20743 & ~n40957 ) ;
  assign n51447 = n51446 ^ n47711 ^ n28037 ;
  assign n51448 = ( n2249 & n3886 ) | ( n2249 & ~n51447 ) | ( n3886 & ~n51447 ) ;
  assign n51449 = ( ~n31550 & n51445 ) | ( ~n31550 & n51448 ) | ( n51445 & n51448 ) ;
  assign n51451 = n44967 ^ n43616 ^ n1665 ;
  assign n51450 = n31242 ^ n7698 ^ n7520 ;
  assign n51452 = n51451 ^ n51450 ^ n36384 ;
  assign n51453 = n45203 & ~n49089 ;
  assign n51454 = n51453 ^ n25498 ^ 1'b0 ;
  assign n51456 = n38299 ^ n21986 ^ n14794 ;
  assign n51455 = ~n40117 & n47548 ;
  assign n51457 = n51456 ^ n51455 ^ 1'b0 ;
  assign n51458 = ( ~n8108 & n26501 ) | ( ~n8108 & n27452 ) | ( n26501 & n27452 ) ;
  assign n51459 = ( ~n29243 & n45002 ) | ( ~n29243 & n51458 ) | ( n45002 & n51458 ) ;
  assign n51460 = ( n33963 & ~n48127 ) | ( n33963 & n49250 ) | ( ~n48127 & n49250 ) ;
  assign n51461 = n51460 ^ n40447 ^ n39876 ;
  assign n51462 = ( n9213 & ~n13361 ) | ( n9213 & n18888 ) | ( ~n13361 & n18888 ) ;
  assign n51463 = ( n8484 & ~n20922 ) | ( n8484 & n51462 ) | ( ~n20922 & n51462 ) ;
  assign n51464 = ( ~x132 & n28490 ) | ( ~x132 & n33944 ) | ( n28490 & n33944 ) ;
  assign n51465 = n44854 ^ n44844 ^ n22104 ;
  assign n51466 = ( n923 & n1310 ) | ( n923 & ~n21035 ) | ( n1310 & ~n21035 ) ;
  assign n51467 = ( n19786 & n40227 ) | ( n19786 & ~n46361 ) | ( n40227 & ~n46361 ) ;
  assign n51468 = n26721 | n29693 ;
  assign n51469 = n5749 | n51468 ;
  assign n51470 = n51469 ^ n51093 ^ n25265 ;
  assign n51471 = n38768 ^ n18998 ^ n2470 ;
  assign n51472 = n9788 & n20464 ;
  assign n51473 = n51472 ^ n44533 ^ 1'b0 ;
  assign n51475 = ( ~n2237 & n6525 ) | ( ~n2237 & n27199 ) | ( n6525 & n27199 ) ;
  assign n51474 = ( n4092 & ~n20689 ) | ( n4092 & n36347 ) | ( ~n20689 & n36347 ) ;
  assign n51476 = n51475 ^ n51474 ^ 1'b0 ;
  assign n51477 = ( n5651 & n13563 ) | ( n5651 & n18557 ) | ( n13563 & n18557 ) ;
  assign n51478 = n51477 ^ n37264 ^ n15346 ;
  assign n51479 = ( n1963 & ~n13623 ) | ( n1963 & n19084 ) | ( ~n13623 & n19084 ) ;
  assign n51480 = ( ~n2710 & n9815 ) | ( ~n2710 & n51479 ) | ( n9815 & n51479 ) ;
  assign n51481 = ( ~n16253 & n20363 ) | ( ~n16253 & n20865 ) | ( n20363 & n20865 ) ;
  assign n51482 = ( n30371 & ~n40807 ) | ( n30371 & n43048 ) | ( ~n40807 & n43048 ) ;
  assign n51483 = ( n3573 & ~n23963 ) | ( n3573 & n38221 ) | ( ~n23963 & n38221 ) ;
  assign n51484 = n51483 ^ n42972 ^ n1024 ;
  assign n51485 = n3703 | n9401 ;
  assign n51486 = n51485 ^ n7208 ^ 1'b0 ;
  assign n51487 = n50694 ^ n27241 ^ n25513 ;
  assign n51488 = ( n32059 & n50147 ) | ( n32059 & ~n51487 ) | ( n50147 & ~n51487 ) ;
  assign n51489 = n51488 ^ n18848 ^ 1'b0 ;
  assign n51490 = n29103 & n51489 ;
  assign n51491 = ( n689 & ~n2469 ) | ( n689 & n51490 ) | ( ~n2469 & n51490 ) ;
  assign n51492 = ~n1888 & n29060 ;
  assign n51493 = n51492 ^ n5063 ^ 1'b0 ;
  assign n51494 = n47238 ^ n25687 ^ n21160 ;
  assign n51495 = ( n7747 & n24114 ) | ( n7747 & ~n34554 ) | ( n24114 & ~n34554 ) ;
  assign n51496 = ( n26176 & n31664 ) | ( n26176 & n38567 ) | ( n31664 & n38567 ) ;
  assign n51497 = ( n356 & ~n730 ) | ( n356 & n5565 ) | ( ~n730 & n5565 ) ;
  assign n51498 = ~n19356 & n45180 ;
  assign n51499 = n24722 ^ n24561 ^ 1'b0 ;
  assign n51500 = ( n3607 & n19401 ) | ( n3607 & ~n51499 ) | ( n19401 & ~n51499 ) ;
  assign n51501 = n33156 ^ n8073 ^ 1'b0 ;
  assign n51502 = ( n51498 & n51500 ) | ( n51498 & n51501 ) | ( n51500 & n51501 ) ;
  assign n51503 = n48856 ^ n7206 ^ n3968 ;
  assign n51504 = n13466 & n35872 ;
  assign n51505 = n51504 ^ n13760 ^ n13459 ;
  assign n51506 = ( n11473 & ~n12021 ) | ( n11473 & n45074 ) | ( ~n12021 & n45074 ) ;
  assign n51507 = ( ~n11163 & n31840 ) | ( ~n11163 & n51506 ) | ( n31840 & n51506 ) ;
  assign n51508 = ~n15759 & n17705 ;
  assign n51509 = ~n38574 & n51508 ;
  assign n51510 = n3510 & n39767 ;
  assign n51511 = n51510 ^ n15024 ^ 1'b0 ;
  assign n51514 = ~n2889 & n30409 ;
  assign n51515 = n51514 ^ n26144 ^ n19663 ;
  assign n51513 = ( n6952 & n28657 ) | ( n6952 & n37877 ) | ( n28657 & n37877 ) ;
  assign n51512 = ( n6648 & ~n12881 ) | ( n6648 & n23718 ) | ( ~n12881 & n23718 ) ;
  assign n51516 = n51515 ^ n51513 ^ n51512 ;
  assign n51518 = n24460 ^ n12204 ^ n9114 ;
  assign n51517 = n10043 & ~n18810 ;
  assign n51519 = n51518 ^ n51517 ^ n32681 ;
  assign n51521 = n11788 | n32767 ;
  assign n51522 = n4075 & ~n51521 ;
  assign n51520 = ( n18815 & n30470 ) | ( n18815 & ~n39561 ) | ( n30470 & ~n39561 ) ;
  assign n51523 = n51522 ^ n51520 ^ n3692 ;
  assign n51524 = n51523 ^ n37436 ^ n17314 ;
  assign n51525 = ( n27213 & ~n33430 ) | ( n27213 & n38784 ) | ( ~n33430 & n38784 ) ;
  assign n51526 = ( n20419 & n46318 ) | ( n20419 & ~n51525 ) | ( n46318 & ~n51525 ) ;
  assign n51527 = n27593 ^ n13159 ^ n10828 ;
  assign n51528 = ( n1802 & n27110 ) | ( n1802 & n51527 ) | ( n27110 & n51527 ) ;
  assign n51529 = ( n5226 & n5956 ) | ( n5226 & n38137 ) | ( n5956 & n38137 ) ;
  assign n51533 = n22850 ^ n22799 ^ n20202 ;
  assign n51530 = n29201 ^ n26292 ^ 1'b0 ;
  assign n51531 = ~n17777 & n51530 ;
  assign n51532 = n51531 ^ n39879 ^ n1502 ;
  assign n51534 = n51533 ^ n51532 ^ n27544 ;
  assign n51535 = n36504 ^ n20060 ^ n3479 ;
  assign n51536 = n23627 | n26250 ;
  assign n51537 = ( n315 & n28872 ) | ( n315 & n36149 ) | ( n28872 & n36149 ) ;
  assign n51538 = n20376 | n51537 ;
  assign n51539 = ~n1809 & n51538 ;
  assign n51540 = n51539 ^ n5057 ^ 1'b0 ;
  assign n51541 = ( n44998 & n51536 ) | ( n44998 & n51540 ) | ( n51536 & n51540 ) ;
  assign n51542 = ( n2796 & ~n9628 ) | ( n2796 & n20875 ) | ( ~n9628 & n20875 ) ;
  assign n51543 = ( ~n21386 & n22205 ) | ( ~n21386 & n51542 ) | ( n22205 & n51542 ) ;
  assign n51544 = n1104 & ~n51543 ;
  assign n51545 = ~n1321 & n51544 ;
  assign n51546 = ( n20827 & n29134 ) | ( n20827 & n34113 ) | ( n29134 & n34113 ) ;
  assign n51547 = n37532 & ~n51546 ;
  assign n51548 = ~x53 & n51547 ;
  assign n51549 = n32525 ^ n22686 ^ n9088 ;
  assign n51550 = ( ~n30056 & n38642 ) | ( ~n30056 & n41565 ) | ( n38642 & n41565 ) ;
  assign n51551 = ( ~n19966 & n51549 ) | ( ~n19966 & n51550 ) | ( n51549 & n51550 ) ;
  assign n51552 = n38122 ^ n31409 ^ n25739 ;
  assign n51553 = n51537 ^ n19634 ^ 1'b0 ;
  assign n51554 = ( ~n29318 & n49209 ) | ( ~n29318 & n51553 ) | ( n49209 & n51553 ) ;
  assign n51564 = n10762 ^ n519 ^ 1'b0 ;
  assign n51565 = n15200 | n51564 ;
  assign n51559 = n32821 ^ n21613 ^ n21375 ;
  assign n51560 = n51559 ^ n34971 ^ n9087 ;
  assign n51561 = ( n5993 & n35290 ) | ( n5993 & ~n51560 ) | ( n35290 & ~n51560 ) ;
  assign n51562 = n28263 & ~n51561 ;
  assign n51555 = n13553 ^ n2376 ^ 1'b0 ;
  assign n51556 = ( n468 & n5312 ) | ( n468 & n51555 ) | ( n5312 & n51555 ) ;
  assign n51557 = n51556 ^ n26873 ^ n1735 ;
  assign n51558 = n13306 & n51557 ;
  assign n51563 = n51562 ^ n51558 ^ 1'b0 ;
  assign n51566 = n51565 ^ n51563 ^ n8804 ;
  assign n51567 = ( ~n1534 & n30732 ) | ( ~n1534 & n45688 ) | ( n30732 & n45688 ) ;
  assign n51570 = ( ~n21594 & n24253 ) | ( ~n21594 & n27650 ) | ( n24253 & n27650 ) ;
  assign n51568 = ( n3316 & ~n11765 ) | ( n3316 & n16443 ) | ( ~n11765 & n16443 ) ;
  assign n51569 = ( ~n1305 & n22472 ) | ( ~n1305 & n51568 ) | ( n22472 & n51568 ) ;
  assign n51571 = n51570 ^ n51569 ^ n5696 ;
  assign n51572 = ( n3740 & n5862 ) | ( n3740 & n8943 ) | ( n5862 & n8943 ) ;
  assign n51573 = ( ~n6718 & n48871 ) | ( ~n6718 & n51572 ) | ( n48871 & n51572 ) ;
  assign n51574 = n29055 ^ n28696 ^ n7724 ;
  assign n51576 = ~n3767 & n9616 ;
  assign n51575 = n27926 & ~n36894 ;
  assign n51577 = n51576 ^ n51575 ^ 1'b0 ;
  assign n51578 = n51577 ^ n554 ^ 1'b0 ;
  assign n51579 = n37641 & ~n51578 ;
  assign n51580 = n27330 ^ n3251 ^ 1'b0 ;
  assign n51581 = n15757 & n51580 ;
  assign n51582 = n34457 ^ n18221 ^ n14051 ;
  assign n51583 = ( n42269 & n51581 ) | ( n42269 & n51582 ) | ( n51581 & n51582 ) ;
  assign n51584 = n39377 ^ n13388 ^ 1'b0 ;
  assign n51585 = ( n25359 & ~n33783 ) | ( n25359 & n51584 ) | ( ~n33783 & n51584 ) ;
  assign n51586 = ( n5629 & ~n9766 ) | ( n5629 & n51585 ) | ( ~n9766 & n51585 ) ;
  assign n51587 = n16900 & ~n25838 ;
  assign n51588 = n51587 ^ n30422 ^ 1'b0 ;
  assign n51589 = n51588 ^ n35974 ^ n6286 ;
  assign n51590 = n22175 ^ n6668 ^ n4378 ;
  assign n51591 = ( n15468 & n32468 ) | ( n15468 & n34264 ) | ( n32468 & n34264 ) ;
  assign n51592 = n6665 & n36311 ;
  assign n51593 = ( n12315 & n43344 ) | ( n12315 & n44179 ) | ( n43344 & n44179 ) ;
  assign n51594 = ( n12536 & n24312 ) | ( n12536 & n51593 ) | ( n24312 & n51593 ) ;
  assign n51595 = n47516 ^ n30840 ^ n17044 ;
  assign n51596 = ( ~n1454 & n6188 ) | ( ~n1454 & n30965 ) | ( n6188 & n30965 ) ;
  assign n51597 = n51596 ^ n43468 ^ n35423 ;
  assign n51598 = ( n16756 & n51595 ) | ( n16756 & n51597 ) | ( n51595 & n51597 ) ;
  assign n51599 = n5763 & ~n18194 ;
  assign n51600 = n51599 ^ n23901 ^ 1'b0 ;
  assign n51601 = n4760 | n38198 ;
  assign n51602 = n13044 & ~n51601 ;
  assign n51603 = n9256 & n41782 ;
  assign n51604 = n51602 & n51603 ;
  assign n51612 = n43523 ^ n22213 ^ n826 ;
  assign n51613 = n51612 ^ n23596 ^ 1'b0 ;
  assign n51614 = n39481 & n51613 ;
  assign n51605 = ( n10470 & n12904 ) | ( n10470 & ~n16538 ) | ( n12904 & ~n16538 ) ;
  assign n51606 = n10690 & n50955 ;
  assign n51607 = ~n51605 & n51606 ;
  assign n51608 = n51607 ^ n11546 ^ 1'b0 ;
  assign n51609 = n51608 ^ n13432 ^ 1'b0 ;
  assign n51610 = n51609 ^ n11834 ^ 1'b0 ;
  assign n51611 = n12038 & n51610 ;
  assign n51615 = n51614 ^ n51611 ^ n5014 ;
  assign n51616 = n44957 ^ n36917 ^ n18223 ;
  assign n51617 = n45216 ^ n11392 ^ n7035 ;
  assign n51618 = ( n3339 & ~n26011 ) | ( n3339 & n51617 ) | ( ~n26011 & n51617 ) ;
  assign n51619 = ( n5271 & n24976 ) | ( n5271 & ~n29953 ) | ( n24976 & ~n29953 ) ;
  assign n51620 = ( n3465 & n26032 ) | ( n3465 & n51619 ) | ( n26032 & n51619 ) ;
  assign n51621 = n15439 & n51620 ;
  assign n51622 = n34052 ^ n20893 ^ n6233 ;
  assign n51623 = ( n3928 & n17157 ) | ( n3928 & ~n34869 ) | ( n17157 & ~n34869 ) ;
  assign n51624 = n13440 ^ n3275 ^ 1'b0 ;
  assign n51625 = n24139 ^ n8964 ^ 1'b0 ;
  assign n51626 = n45767 ^ n30686 ^ n26729 ;
  assign n51627 = ( n13065 & ~n46914 ) | ( n13065 & n51626 ) | ( ~n46914 & n51626 ) ;
  assign n51628 = ( ~n9848 & n44597 ) | ( ~n9848 & n51627 ) | ( n44597 & n51627 ) ;
  assign n51634 = n50196 ^ n31103 ^ n4010 ;
  assign n51631 = ( ~n472 & n1707 ) | ( ~n472 & n1845 ) | ( n1707 & n1845 ) ;
  assign n51629 = n32439 ^ n11795 ^ n8013 ;
  assign n51630 = ( n6648 & n17963 ) | ( n6648 & n51629 ) | ( n17963 & n51629 ) ;
  assign n51632 = n51631 ^ n51630 ^ n1238 ;
  assign n51633 = n2787 & ~n51632 ;
  assign n51635 = n51634 ^ n51633 ^ 1'b0 ;
  assign n51636 = ~n2557 & n34936 ;
  assign n51637 = n51636 ^ n4478 ^ 1'b0 ;
  assign n51638 = n13923 & n51637 ;
  assign n51639 = n43357 ^ n24865 ^ n19740 ;
  assign n51640 = ( n2953 & ~n28737 ) | ( n2953 & n51639 ) | ( ~n28737 & n51639 ) ;
  assign n51641 = n42090 ^ n15958 ^ n8925 ;
  assign n51642 = ( ~n18946 & n19572 ) | ( ~n18946 & n23226 ) | ( n19572 & n23226 ) ;
  assign n51643 = n17780 & ~n42119 ;
  assign n51644 = n35651 ^ n35130 ^ n29512 ;
  assign n51645 = ( n12673 & ~n21863 ) | ( n12673 & n40439 ) | ( ~n21863 & n40439 ) ;
  assign n51647 = ( n3076 & n12273 ) | ( n3076 & n26018 ) | ( n12273 & n26018 ) ;
  assign n51646 = n4533 ^ n3266 ^ n854 ;
  assign n51648 = n51647 ^ n51646 ^ n35738 ;
  assign n51649 = ( n9625 & n21725 ) | ( n9625 & n51648 ) | ( n21725 & n51648 ) ;
  assign n51650 = n38631 ^ n29221 ^ n19771 ;
  assign n51651 = n6351 & ~n21833 ;
  assign n51652 = n50631 & n51651 ;
  assign n51653 = n23475 ^ n16443 ^ n3674 ;
  assign n51654 = n51653 ^ n41677 ^ n22670 ;
  assign n51655 = ( n6636 & ~n9353 ) | ( n6636 & n15403 ) | ( ~n9353 & n15403 ) ;
  assign n51656 = ( n10506 & n16258 ) | ( n10506 & n51655 ) | ( n16258 & n51655 ) ;
  assign n51657 = ( n709 & n11136 ) | ( n709 & ~n14559 ) | ( n11136 & ~n14559 ) ;
  assign n51658 = n47488 ^ n40699 ^ n18418 ;
  assign n51659 = n51658 ^ n25025 ^ n9785 ;
  assign n51660 = ( n3718 & ~n8447 ) | ( n3718 & n21112 ) | ( ~n8447 & n21112 ) ;
  assign n51661 = ( n4484 & n7072 ) | ( n4484 & ~n51660 ) | ( n7072 & ~n51660 ) ;
  assign n51662 = n29122 ^ n1940 ^ n1465 ;
  assign n51663 = ( n1517 & ~n2803 ) | ( n1517 & n45618 ) | ( ~n2803 & n45618 ) ;
  assign n51664 = n34912 ^ n12116 ^ 1'b0 ;
  assign n51665 = n24038 & ~n51664 ;
  assign n51666 = ( n1137 & n5338 ) | ( n1137 & n51665 ) | ( n5338 & n51665 ) ;
  assign n51667 = n51666 ^ n26291 ^ n10129 ;
  assign n51669 = ( n1748 & n21375 ) | ( n1748 & ~n34156 ) | ( n21375 & ~n34156 ) ;
  assign n51668 = ~n4135 & n14228 ;
  assign n51670 = n51669 ^ n51668 ^ 1'b0 ;
  assign n51671 = n15870 & ~n23237 ;
  assign n51672 = ( ~n18184 & n26954 ) | ( ~n18184 & n37877 ) | ( n26954 & n37877 ) ;
  assign n51673 = n20106 ^ n11458 ^ n7565 ;
  assign n51674 = n32990 & ~n51673 ;
  assign n51675 = ( n31672 & n34234 ) | ( n31672 & n39075 ) | ( n34234 & n39075 ) ;
  assign n51676 = n51675 ^ n30411 ^ n10129 ;
  assign n51683 = ( n3947 & n15918 ) | ( n3947 & n45557 ) | ( n15918 & n45557 ) ;
  assign n51680 = n20412 ^ n7952 ^ n5872 ;
  assign n51677 = n14417 | n25136 ;
  assign n51678 = n20459 | n51677 ;
  assign n51679 = n51678 ^ n34168 ^ n5301 ;
  assign n51681 = n51680 ^ n51679 ^ n41894 ;
  assign n51682 = n51681 ^ n13292 ^ 1'b0 ;
  assign n51684 = n51683 ^ n51682 ^ n35551 ;
  assign n51685 = n41361 ^ n20931 ^ n7014 ;
  assign n51686 = n28290 ^ n25362 ^ 1'b0 ;
  assign n51687 = ( ~n3158 & n34158 ) | ( ~n3158 & n51686 ) | ( n34158 & n51686 ) ;
  assign n51688 = n51687 ^ n12985 ^ n4943 ;
  assign n51689 = ( n6455 & n14555 ) | ( n6455 & n19028 ) | ( n14555 & n19028 ) ;
  assign n51690 = ( ~n7667 & n12848 ) | ( ~n7667 & n51689 ) | ( n12848 & n51689 ) ;
  assign n51692 = ( x18 & ~n12530 ) | ( x18 & n41947 ) | ( ~n12530 & n41947 ) ;
  assign n51693 = n51692 ^ n24593 ^ n5167 ;
  assign n51691 = n4207 & n46251 ;
  assign n51694 = n51693 ^ n51691 ^ 1'b0 ;
  assign n51695 = ( n4289 & ~n13128 ) | ( n4289 & n51308 ) | ( ~n13128 & n51308 ) ;
  assign n51696 = ( ~n6656 & n10302 ) | ( ~n6656 & n50751 ) | ( n10302 & n50751 ) ;
  assign n51697 = ( n9972 & n11843 ) | ( n9972 & ~n28468 ) | ( n11843 & ~n28468 ) ;
  assign n51698 = ( n51695 & ~n51696 ) | ( n51695 & n51697 ) | ( ~n51696 & n51697 ) ;
  assign n51699 = n28550 ^ n4025 ^ n1881 ;
  assign n51701 = n43103 ^ n20666 ^ n1770 ;
  assign n51702 = n51701 ^ n20991 ^ n4285 ;
  assign n51700 = ( n26097 & ~n39168 ) | ( n26097 & n39432 ) | ( ~n39168 & n39432 ) ;
  assign n51703 = n51702 ^ n51700 ^ n36232 ;
  assign n51704 = n47034 ^ n6476 ^ n2209 ;
  assign n51705 = n41850 ^ n19572 ^ n4733 ;
  assign n51706 = ( n16189 & n20290 ) | ( n16189 & ~n45744 ) | ( n20290 & ~n45744 ) ;
  assign n51707 = n50272 ^ n15072 ^ n6296 ;
  assign n51708 = ( ~n1513 & n32196 ) | ( ~n1513 & n47234 ) | ( n32196 & n47234 ) ;
  assign n51709 = ( n7959 & n21382 ) | ( n7959 & ~n50416 ) | ( n21382 & ~n50416 ) ;
  assign n51710 = ( n1636 & n12102 ) | ( n1636 & n51709 ) | ( n12102 & n51709 ) ;
  assign n51711 = n45066 ^ n376 ^ 1'b0 ;
  assign n51712 = n51710 & n51711 ;
  assign n51713 = ~n3440 & n21679 ;
  assign n51714 = n51713 ^ n21585 ^ 1'b0 ;
  assign n51715 = n49357 ^ n45830 ^ 1'b0 ;
  assign n51716 = ~n14371 & n32026 ;
  assign n51717 = n50938 ^ n9498 ^ n7426 ;
  assign n51718 = ( n14978 & n46299 ) | ( n14978 & ~n51717 ) | ( n46299 & ~n51717 ) ;
  assign n51719 = ( n21408 & n26371 ) | ( n21408 & n30443 ) | ( n26371 & n30443 ) ;
  assign n51720 = n24426 ^ n7490 ^ n3124 ;
  assign n51721 = ( n32920 & ~n51719 ) | ( n32920 & n51720 ) | ( ~n51719 & n51720 ) ;
  assign n51722 = ( n1412 & n21286 ) | ( n1412 & ~n40002 ) | ( n21286 & ~n40002 ) ;
  assign n51723 = n40270 ^ n30848 ^ n4964 ;
  assign n51724 = ( n31572 & ~n51722 ) | ( n31572 & n51723 ) | ( ~n51722 & n51723 ) ;
  assign n51725 = ( n4248 & n19108 ) | ( n4248 & ~n24671 ) | ( n19108 & ~n24671 ) ;
  assign n51726 = ( ~n14235 & n14853 ) | ( ~n14235 & n17835 ) | ( n14853 & n17835 ) ;
  assign n51727 = n9056 & ~n51726 ;
  assign n51728 = ~n1452 & n51727 ;
  assign n51729 = ( n35069 & n51725 ) | ( n35069 & ~n51728 ) | ( n51725 & ~n51728 ) ;
  assign n51730 = ( n14380 & n30565 ) | ( n14380 & ~n38942 ) | ( n30565 & ~n38942 ) ;
  assign n51731 = n40379 ^ n25806 ^ n8913 ;
  assign n51732 = n51731 ^ n19520 ^ n19411 ;
  assign n51733 = n22098 ^ n20379 ^ n1411 ;
  assign n51734 = n47432 | n51733 ;
  assign n51735 = n11099 & ~n51734 ;
  assign n51736 = ( n261 & n12975 ) | ( n261 & n22911 ) | ( n12975 & n22911 ) ;
  assign n51737 = n32408 ^ n22772 ^ 1'b0 ;
  assign n51738 = n51736 & ~n51737 ;
  assign n51739 = n26684 ^ n21720 ^ n10505 ;
  assign n51740 = n51739 ^ n33094 ^ n1781 ;
  assign n51741 = n25240 ^ n1810 ^ 1'b0 ;
  assign n51742 = ~n1640 & n51741 ;
  assign n51743 = n51742 ^ n39938 ^ n3719 ;
  assign n51744 = n40654 | n51743 ;
  assign n51745 = ( n22503 & ~n50357 ) | ( n22503 & n51744 ) | ( ~n50357 & n51744 ) ;
  assign n51746 = ( ~n7324 & n17164 ) | ( ~n7324 & n51745 ) | ( n17164 & n51745 ) ;
  assign n51747 = n37710 ^ n3858 ^ 1'b0 ;
  assign n51748 = n15868 ^ n8058 ^ 1'b0 ;
  assign n51749 = n15373 ^ n4506 ^ 1'b0 ;
  assign n51750 = n51748 | n51749 ;
  assign n51751 = ( ~n516 & n16084 ) | ( ~n516 & n51750 ) | ( n16084 & n51750 ) ;
  assign n51752 = ( n4355 & n11887 ) | ( n4355 & n34343 ) | ( n11887 & n34343 ) ;
  assign n51755 = n33511 ^ n9555 ^ n5911 ;
  assign n51753 = n13260 ^ n11463 ^ 1'b0 ;
  assign n51754 = n19275 & n51753 ;
  assign n51756 = n51755 ^ n51754 ^ n45886 ;
  assign n51757 = n46039 ^ n6798 ^ n304 ;
  assign n51758 = n17723 & ~n38333 ;
  assign n51759 = n13934 & n51758 ;
  assign n51761 = ( ~n3587 & n12069 ) | ( ~n3587 & n24104 ) | ( n12069 & n24104 ) ;
  assign n51760 = n10103 ^ n3431 ^ x42 ;
  assign n51762 = n51761 ^ n51760 ^ n24659 ;
  assign n51763 = ( n6871 & ~n40311 ) | ( n6871 & n51762 ) | ( ~n40311 & n51762 ) ;
  assign n51764 = ( n19685 & n51759 ) | ( n19685 & n51763 ) | ( n51759 & n51763 ) ;
  assign n51767 = n21367 ^ n14663 ^ n7610 ;
  assign n51765 = n35485 ^ n9032 ^ n1427 ;
  assign n51766 = n51765 ^ n24448 ^ n6197 ;
  assign n51768 = n51767 ^ n51766 ^ n25274 ;
  assign n51769 = ( n6362 & ~n15897 ) | ( n6362 & n28671 ) | ( ~n15897 & n28671 ) ;
  assign n51770 = n29514 ^ n9374 ^ 1'b0 ;
  assign n51771 = n14612 & n51770 ;
  assign n51772 = n51771 ^ n19588 ^ n5267 ;
  assign n51773 = n26472 ^ n10636 ^ n5450 ;
  assign n51774 = n51773 ^ n27305 ^ 1'b0 ;
  assign n51775 = ~n18719 & n51774 ;
  assign n51776 = n51775 ^ n35595 ^ n2096 ;
  assign n51777 = n27959 ^ n6897 ^ 1'b0 ;
  assign n51778 = n31807 ^ n28689 ^ n27008 ;
  assign n51779 = n51778 ^ n37406 ^ n24990 ;
  assign n51780 = ( n18565 & n20735 ) | ( n18565 & n51779 ) | ( n20735 & n51779 ) ;
  assign n51781 = ( n13316 & ~n13441 ) | ( n13316 & n45588 ) | ( ~n13441 & n45588 ) ;
  assign n51782 = ( n6253 & ~n18330 ) | ( n6253 & n40700 ) | ( ~n18330 & n40700 ) ;
  assign n51783 = n51782 ^ n50109 ^ n38942 ;
  assign n51784 = n38760 | n43772 ;
  assign n51785 = n35093 ^ n26793 ^ n19610 ;
  assign n51786 = n51785 ^ n21033 ^ 1'b0 ;
  assign n51787 = n3470 & n51786 ;
  assign n51788 = n6639 ^ n1975 ^ 1'b0 ;
  assign n51789 = ( n13934 & n30291 ) | ( n13934 & ~n51788 ) | ( n30291 & ~n51788 ) ;
  assign n51790 = ( n2105 & ~n5834 ) | ( n2105 & n23624 ) | ( ~n5834 & n23624 ) ;
  assign n51791 = n51790 ^ n21937 ^ n16126 ;
  assign n51792 = n51791 ^ n49849 ^ 1'b0 ;
  assign n51793 = n18960 ^ n11717 ^ n10765 ;
  assign n51794 = n51793 ^ n30962 ^ n21082 ;
  assign n51795 = ( n24898 & n46104 ) | ( n24898 & ~n47941 ) | ( n46104 & ~n47941 ) ;
  assign n51796 = n30552 ^ n29186 ^ n13438 ;
  assign n51797 = ( n18430 & ~n37389 ) | ( n18430 & n39994 ) | ( ~n37389 & n39994 ) ;
  assign n51798 = n51797 ^ n37320 ^ n18608 ;
  assign n51799 = n9689 & n26368 ;
  assign n51800 = n11698 ^ n6147 ^ 1'b0 ;
  assign n51801 = ( n12204 & n51799 ) | ( n12204 & ~n51800 ) | ( n51799 & ~n51800 ) ;
  assign n51802 = n40144 ^ n27507 ^ n8047 ;
  assign n51803 = n39570 ^ n17958 ^ n2855 ;
  assign n51804 = ~n4968 & n51803 ;
  assign n51805 = ~n42654 & n51804 ;
  assign n51809 = n25409 & n45267 ;
  assign n51806 = ~n14652 & n16629 ;
  assign n51807 = n51806 ^ n15097 ^ 1'b0 ;
  assign n51808 = n51807 ^ n17932 ^ 1'b0 ;
  assign n51810 = n51809 ^ n51808 ^ n34858 ;
  assign n51811 = ~n11542 & n12809 ;
  assign n51812 = ( n24732 & n41898 ) | ( n24732 & n51811 ) | ( n41898 & n51811 ) ;
  assign n51813 = n51812 ^ n39820 ^ n18747 ;
  assign n51814 = ( n4342 & n4385 ) | ( n4342 & n11674 ) | ( n4385 & n11674 ) ;
  assign n51815 = ( n4310 & n12383 ) | ( n4310 & ~n51814 ) | ( n12383 & ~n51814 ) ;
  assign n51816 = ~n17389 & n43968 ;
  assign n51817 = n8483 | n13232 ;
  assign n51818 = n29095 & ~n51817 ;
  assign n51819 = ( n4913 & n47686 ) | ( n4913 & n51818 ) | ( n47686 & n51818 ) ;
  assign n51820 = n22406 ^ n14251 ^ x234 ;
  assign n51821 = n12182 ^ n10452 ^ n2003 ;
  assign n51822 = ( ~n32887 & n51820 ) | ( ~n32887 & n51821 ) | ( n51820 & n51821 ) ;
  assign n51823 = n51822 ^ n38279 ^ n17562 ;
  assign n51824 = ( n3634 & n34969 ) | ( n3634 & ~n37193 ) | ( n34969 & ~n37193 ) ;
  assign n51827 = n15129 ^ n13503 ^ n4318 ;
  assign n51828 = n51827 ^ n26148 ^ n2745 ;
  assign n51825 = n3920 & n4995 ;
  assign n51826 = n51825 ^ n31742 ^ n24017 ;
  assign n51829 = n51828 ^ n51826 ^ n28600 ;
  assign n51830 = n38291 ^ n32644 ^ n29301 ;
  assign n51831 = n26003 ^ n20041 ^ n7202 ;
  assign n51834 = n26925 ^ n9652 ^ n6974 ;
  assign n51835 = n36404 | n51834 ;
  assign n51836 = ~n45077 & n51835 ;
  assign n51837 = n11339 & n51836 ;
  assign n51832 = n1210 | n36302 ;
  assign n51833 = n24768 | n51832 ;
  assign n51838 = n51837 ^ n51833 ^ n30443 ;
  assign n51840 = ~n40917 & n43399 ;
  assign n51839 = n46039 ^ n36132 ^ n5090 ;
  assign n51841 = n51840 ^ n51839 ^ n12591 ;
  assign n51842 = ~n12250 & n24076 ;
  assign n51843 = n51842 ^ n24752 ^ 1'b0 ;
  assign n51844 = ( ~n1289 & n15724 ) | ( ~n1289 & n51843 ) | ( n15724 & n51843 ) ;
  assign n51845 = n35265 ^ n25267 ^ n4073 ;
  assign n51846 = n47201 ^ n40328 ^ n6567 ;
  assign n51847 = ( n2962 & n28304 ) | ( n2962 & n51846 ) | ( n28304 & n51846 ) ;
  assign n51848 = n44910 ^ n20689 ^ 1'b0 ;
  assign n51849 = ~n25968 & n51848 ;
  assign n51850 = n33342 ^ n19201 ^ 1'b0 ;
  assign n51851 = n39999 | n51850 ;
  assign n51852 = ( n22189 & ~n37179 ) | ( n22189 & n51851 ) | ( ~n37179 & n51851 ) ;
  assign n51853 = n38211 ^ n26738 ^ n21377 ;
  assign n51854 = n23186 ^ n21171 ^ n1662 ;
  assign n51855 = n51854 ^ n19019 ^ 1'b0 ;
  assign n51856 = n25405 & n35915 ;
  assign n51857 = n36458 ^ n6494 ^ n2915 ;
  assign n51858 = n44585 ^ n34329 ^ n13120 ;
  assign n51859 = ( n12489 & n19570 ) | ( n12489 & n51858 ) | ( n19570 & n51858 ) ;
  assign n51860 = n51859 ^ n41149 ^ n6837 ;
  assign n51861 = n51860 ^ n47016 ^ n7015 ;
  assign n51863 = ( n8552 & n32508 ) | ( n8552 & ~n45695 ) | ( n32508 & ~n45695 ) ;
  assign n51862 = n25729 ^ n16830 ^ 1'b0 ;
  assign n51864 = n51863 ^ n51862 ^ n11975 ;
  assign n51865 = n20991 ^ n14041 ^ n9380 ;
  assign n51866 = ( n3282 & ~n3986 ) | ( n3282 & n8945 ) | ( ~n3986 & n8945 ) ;
  assign n51867 = ( n32532 & n51865 ) | ( n32532 & n51866 ) | ( n51865 & n51866 ) ;
  assign n51868 = n50044 ^ n38477 ^ n17409 ;
  assign n51869 = n51868 ^ n24956 ^ n18558 ;
  assign n51870 = ( n274 & n5253 ) | ( n274 & ~n12294 ) | ( n5253 & ~n12294 ) ;
  assign n51871 = n51870 ^ n20448 ^ n7598 ;
  assign n51872 = n44367 ^ n9797 ^ n289 ;
  assign n51873 = ( n46935 & n51871 ) | ( n46935 & ~n51872 ) | ( n51871 & ~n51872 ) ;
  assign n51874 = n12093 & ~n43555 ;
  assign n51875 = n51874 ^ n3938 ^ 1'b0 ;
  assign n51876 = ( n5915 & n8833 ) | ( n5915 & ~n34211 ) | ( n8833 & ~n34211 ) ;
  assign n51877 = ( n3797 & n51875 ) | ( n3797 & n51876 ) | ( n51875 & n51876 ) ;
  assign n51878 = n34799 ^ n21579 ^ n1674 ;
  assign n51879 = n857 & n2524 ;
  assign n51880 = n9992 & n51879 ;
  assign n51881 = n51880 ^ n8287 ^ 1'b0 ;
  assign n51882 = ~n50832 & n51881 ;
  assign n51883 = n51878 & n51882 ;
  assign n51884 = n51883 ^ n24252 ^ x5 ;
  assign n51885 = ( n5794 & ~n27830 ) | ( n5794 & n38018 ) | ( ~n27830 & n38018 ) ;
  assign n51886 = n33132 ^ n3651 ^ n2284 ;
  assign n51887 = n462 & n8511 ;
  assign n51888 = n51887 ^ n18282 ^ 1'b0 ;
  assign n51889 = n44159 ^ n25230 ^ n8324 ;
  assign n51891 = x241 & ~n16638 ;
  assign n51892 = n51891 ^ n28176 ^ 1'b0 ;
  assign n51893 = n51892 ^ n39404 ^ n8974 ;
  assign n51894 = ( n8968 & n14506 ) | ( n8968 & n51893 ) | ( n14506 & n51893 ) ;
  assign n51890 = n29425 ^ n26108 ^ n12372 ;
  assign n51895 = n51894 ^ n51890 ^ n39999 ;
  assign n51896 = n51895 ^ n33120 ^ n2304 ;
  assign n51897 = ( n6496 & ~n20592 ) | ( n6496 & n29082 ) | ( ~n20592 & n29082 ) ;
  assign n51898 = n3317 | n8857 ;
  assign n51899 = n13763 & ~n51898 ;
  assign n51900 = ( n9754 & n13384 ) | ( n9754 & ~n51899 ) | ( n13384 & ~n51899 ) ;
  assign n51901 = n24317 | n43382 ;
  assign n51902 = n51901 ^ n50412 ^ 1'b0 ;
  assign n51903 = ( ~n12342 & n31080 ) | ( ~n12342 & n51902 ) | ( n31080 & n51902 ) ;
  assign n51904 = n30985 ^ n7279 ^ n6517 ;
  assign n51905 = ( n45440 & ~n46687 ) | ( n45440 & n51904 ) | ( ~n46687 & n51904 ) ;
  assign n51906 = ( n2478 & n3942 ) | ( n2478 & ~n29946 ) | ( n3942 & ~n29946 ) ;
  assign n51907 = ( n22120 & n31689 ) | ( n22120 & ~n51906 ) | ( n31689 & ~n51906 ) ;
  assign n51908 = ( n1244 & ~n3486 ) | ( n1244 & n40147 ) | ( ~n3486 & n40147 ) ;
  assign n51909 = ( n6538 & n17234 ) | ( n6538 & n26767 ) | ( n17234 & n26767 ) ;
  assign n51910 = ~n5417 & n33342 ;
  assign n51911 = ~n25431 & n51910 ;
  assign n51912 = n51909 & ~n51911 ;
  assign n51913 = n5765 | n37189 ;
  assign n51914 = n13942 | n51913 ;
  assign n51915 = ( n37019 & ~n51912 ) | ( n37019 & n51914 ) | ( ~n51912 & n51914 ) ;
  assign n51916 = n6471 & ~n13905 ;
  assign n51917 = n51916 ^ n28466 ^ 1'b0 ;
  assign n51918 = ( n15468 & ~n24269 ) | ( n15468 & n44883 ) | ( ~n24269 & n44883 ) ;
  assign n51920 = n1174 | n7906 ;
  assign n51919 = ( n8044 & n8259 ) | ( n8044 & ~n24596 ) | ( n8259 & ~n24596 ) ;
  assign n51921 = n51920 ^ n51919 ^ 1'b0 ;
  assign n51922 = n51921 ^ n28891 ^ n28057 ;
  assign n51923 = n49151 ^ n2180 ^ x103 ;
  assign n51924 = n51923 ^ n42587 ^ 1'b0 ;
  assign n51927 = ( n15444 & n21028 ) | ( n15444 & ~n49965 ) | ( n21028 & ~n49965 ) ;
  assign n51928 = n51927 ^ n28786 ^ n1197 ;
  assign n51929 = n51928 ^ n48034 ^ n4950 ;
  assign n51930 = ( n9858 & ~n14401 ) | ( n9858 & n51929 ) | ( ~n14401 & n51929 ) ;
  assign n51925 = n49076 ^ n37986 ^ n29683 ;
  assign n51926 = ( n2337 & ~n40412 ) | ( n2337 & n51925 ) | ( ~n40412 & n51925 ) ;
  assign n51931 = n51930 ^ n51926 ^ n26370 ;
  assign n51939 = ( n11410 & n18414 ) | ( n11410 & ~n18830 ) | ( n18414 & ~n18830 ) ;
  assign n51933 = ( n9219 & n14022 ) | ( n9219 & n42586 ) | ( n14022 & n42586 ) ;
  assign n51934 = n51933 ^ n39487 ^ n24943 ;
  assign n51935 = n14348 & n51934 ;
  assign n51936 = ~n44771 & n51935 ;
  assign n51932 = n1780 & n5471 ;
  assign n51937 = n51936 ^ n51932 ^ 1'b0 ;
  assign n51938 = n51937 ^ n32263 ^ n15840 ;
  assign n51940 = n51939 ^ n51938 ^ n27492 ;
  assign n51941 = n51940 ^ n33883 ^ n16053 ;
  assign n51942 = n21691 ^ n14072 ^ 1'b0 ;
  assign n51944 = n21079 ^ n17677 ^ n9289 ;
  assign n51945 = n51944 ^ n3669 ^ 1'b0 ;
  assign n51943 = ( n2452 & n6690 ) | ( n2452 & n50895 ) | ( n6690 & n50895 ) ;
  assign n51946 = n51945 ^ n51943 ^ n41509 ;
  assign n51947 = n46269 ^ n10759 ^ n5917 ;
  assign n51948 = n35364 & ~n36480 ;
  assign n51949 = ~n16853 & n51948 ;
  assign n51950 = n51895 ^ n11466 ^ 1'b0 ;
  assign n51951 = ~n51949 & n51950 ;
  assign n51952 = n41684 & ~n51260 ;
  assign n51955 = n11444 | n26514 ;
  assign n51953 = ( n1729 & n7272 ) | ( n1729 & n7446 ) | ( n7272 & n7446 ) ;
  assign n51954 = n51953 ^ n34889 ^ n22008 ;
  assign n51956 = n51955 ^ n51954 ^ n20290 ;
  assign n51957 = n51934 ^ n28078 ^ x212 ;
  assign n51958 = ( n7659 & n13175 ) | ( n7659 & ~n50363 ) | ( n13175 & ~n50363 ) ;
  assign n51959 = n51958 ^ n26297 ^ n23540 ;
  assign n51960 = ( n46397 & ~n50235 ) | ( n46397 & n51959 ) | ( ~n50235 & n51959 ) ;
  assign n51961 = n44278 ^ n23964 ^ n4836 ;
  assign n51962 = ( n10133 & n14671 ) | ( n10133 & n51181 ) | ( n14671 & n51181 ) ;
  assign n51965 = n31161 ^ n19140 ^ n12705 ;
  assign n51966 = ( n5101 & n20165 ) | ( n5101 & n51965 ) | ( n20165 & n51965 ) ;
  assign n51963 = n18254 & n30909 ;
  assign n51964 = n51963 ^ n26471 ^ 1'b0 ;
  assign n51967 = n51966 ^ n51964 ^ n49579 ;
  assign n51971 = ~n19198 & n22764 ;
  assign n51969 = n17902 ^ n8041 ^ 1'b0 ;
  assign n51968 = n15264 & n50399 ;
  assign n51970 = n51969 ^ n51968 ^ 1'b0 ;
  assign n51972 = n51971 ^ n51970 ^ 1'b0 ;
  assign n51973 = ( n10227 & n21030 ) | ( n10227 & n45937 ) | ( n21030 & n45937 ) ;
  assign n51974 = ( n12861 & n39073 ) | ( n12861 & ~n47627 ) | ( n39073 & ~n47627 ) ;
  assign n51975 = ( ~n691 & n5626 ) | ( ~n691 & n49432 ) | ( n5626 & n49432 ) ;
  assign n51976 = n51975 ^ n34664 ^ n8958 ;
  assign n51977 = ( n11379 & n51974 ) | ( n11379 & n51976 ) | ( n51974 & n51976 ) ;
  assign n51978 = n51977 ^ n46701 ^ n38662 ;
  assign n51979 = n29087 ^ n22921 ^ n16316 ;
  assign n51980 = n38768 ^ n26044 ^ n4386 ;
  assign n51981 = ( ~n23128 & n38916 ) | ( ~n23128 & n51980 ) | ( n38916 & n51980 ) ;
  assign n51982 = ( n39587 & ~n43019 ) | ( n39587 & n51981 ) | ( ~n43019 & n51981 ) ;
  assign n51983 = n39994 ^ n35168 ^ n617 ;
  assign n51984 = ( n27751 & n47320 ) | ( n27751 & n51983 ) | ( n47320 & n51983 ) ;
  assign n51985 = n39844 ^ n28551 ^ n5475 ;
  assign n51986 = n51985 ^ n35996 ^ n4710 ;
  assign n51987 = ( n22769 & n22985 ) | ( n22769 & n28628 ) | ( n22985 & n28628 ) ;
  assign n51988 = ( n13308 & n19478 ) | ( n13308 & ~n29126 ) | ( n19478 & ~n29126 ) ;
  assign n51989 = n33764 & n51988 ;
  assign n51990 = n15952 ^ n13662 ^ n7748 ;
  assign n51991 = n17440 & n51990 ;
  assign n51992 = ( n26496 & n29228 ) | ( n26496 & n51991 ) | ( n29228 & n51991 ) ;
  assign n51993 = ( n40794 & n51989 ) | ( n40794 & ~n51992 ) | ( n51989 & ~n51992 ) ;
  assign n51994 = ( n1298 & ~n13003 ) | ( n1298 & n31861 ) | ( ~n13003 & n31861 ) ;
  assign n51995 = ( n15174 & n21577 ) | ( n15174 & ~n51994 ) | ( n21577 & ~n51994 ) ;
  assign n51996 = n12484 & n21162 ;
  assign n51997 = n50501 ^ n39207 ^ n25192 ;
  assign n51998 = n15522 ^ n11270 ^ 1'b0 ;
  assign n51999 = ( n1062 & n31422 ) | ( n1062 & ~n51998 ) | ( n31422 & ~n51998 ) ;
  assign n52000 = n28131 ^ n12806 ^ n3196 ;
  assign n52001 = n39987 ^ n33777 ^ n6230 ;
  assign n52006 = ~n4033 & n10964 ;
  assign n52007 = ~n14291 & n52006 ;
  assign n52002 = ( n19493 & ~n20254 ) | ( n19493 & n25017 ) | ( ~n20254 & n25017 ) ;
  assign n52003 = n4157 | n12631 ;
  assign n52004 = n52003 ^ n10644 ^ 1'b0 ;
  assign n52005 = ( n42580 & n52002 ) | ( n42580 & n52004 ) | ( n52002 & n52004 ) ;
  assign n52008 = n52007 ^ n52005 ^ n12707 ;
  assign n52009 = ( n18625 & n36865 ) | ( n18625 & ~n52008 ) | ( n36865 & ~n52008 ) ;
  assign n52010 = n35664 ^ n26540 ^ 1'b0 ;
  assign n52012 = ( n1749 & n18870 ) | ( n1749 & n26979 ) | ( n18870 & n26979 ) ;
  assign n52011 = ( n4054 & n12502 ) | ( n4054 & n26337 ) | ( n12502 & n26337 ) ;
  assign n52013 = n52012 ^ n52011 ^ n5516 ;
  assign n52014 = n49788 ^ n33755 ^ n28585 ;
  assign n52015 = n4002 & n6368 ;
  assign n52016 = n26448 & n52015 ;
  assign n52017 = n22682 ^ n9057 ^ 1'b0 ;
  assign n52018 = n9850 & n52017 ;
  assign n52019 = n52018 ^ n32911 ^ n6791 ;
  assign n52020 = n48891 ^ n7004 ^ 1'b0 ;
  assign n52021 = ( ~n2706 & n4250 ) | ( ~n2706 & n4514 ) | ( n4250 & n4514 ) ;
  assign n52022 = ( x227 & n33057 ) | ( x227 & ~n52021 ) | ( n33057 & ~n52021 ) ;
  assign n52023 = n34794 ^ n1858 ^ n1282 ;
  assign n52025 = n40179 ^ n20254 ^ n3355 ;
  assign n52024 = n43830 ^ n25941 ^ n11095 ;
  assign n52026 = n52025 ^ n52024 ^ n6398 ;
  assign n52027 = ( n38948 & n52023 ) | ( n38948 & n52026 ) | ( n52023 & n52026 ) ;
  assign n52028 = ( n18238 & n27453 ) | ( n18238 & ~n48892 ) | ( n27453 & ~n48892 ) ;
  assign n52029 = ( n7866 & n30396 ) | ( n7866 & n43274 ) | ( n30396 & n43274 ) ;
  assign n52030 = n52029 ^ n26597 ^ n19812 ;
  assign n52031 = n47721 ^ n43970 ^ n502 ;
  assign n52032 = ( n51205 & n52030 ) | ( n51205 & ~n52031 ) | ( n52030 & ~n52031 ) ;
  assign n52033 = n27962 ^ n18275 ^ n16976 ;
  assign n52034 = ( ~n25455 & n37822 ) | ( ~n25455 & n52033 ) | ( n37822 & n52033 ) ;
  assign n52035 = ~n481 & n1799 ;
  assign n52036 = n52035 ^ n15289 ^ 1'b0 ;
  assign n52037 = n6535 & ~n31483 ;
  assign n52038 = ~n52036 & n52037 ;
  assign n52039 = n52038 ^ n32714 ^ n7072 ;
  assign n52040 = x223 & n1987 ;
  assign n52041 = n52040 ^ n5601 ^ 1'b0 ;
  assign n52042 = n41962 ^ n30646 ^ 1'b0 ;
  assign n52043 = n37456 ^ n21110 ^ n3796 ;
  assign n52044 = n52043 ^ n20185 ^ 1'b0 ;
  assign n52045 = n1014 & n52044 ;
  assign n52046 = n52045 ^ n44026 ^ n36195 ;
  assign n52047 = ( ~n21574 & n37438 ) | ( ~n21574 & n38056 ) | ( n37438 & n38056 ) ;
  assign n52048 = ( n19501 & n33966 ) | ( n19501 & ~n38894 ) | ( n33966 & ~n38894 ) ;
  assign n52049 = n49326 ^ n949 ^ n295 ;
  assign n52050 = n5037 ^ x120 ^ 1'b0 ;
  assign n52051 = ~n15205 & n52050 ;
  assign n52052 = ( n25179 & ~n49155 ) | ( n25179 & n52051 ) | ( ~n49155 & n52051 ) ;
  assign n52053 = n7707 & n12240 ;
  assign n52054 = n15256 & n52053 ;
  assign n52055 = n17718 & ~n46208 ;
  assign n52056 = ~n18260 & n52055 ;
  assign n52057 = ( ~n2239 & n11136 ) | ( ~n2239 & n39714 ) | ( n11136 & n39714 ) ;
  assign n52058 = ( ~n52054 & n52056 ) | ( ~n52054 & n52057 ) | ( n52056 & n52057 ) ;
  assign n52059 = n48819 ^ n46753 ^ n1563 ;
  assign n52060 = ( n3216 & n8760 ) | ( n3216 & ~n52059 ) | ( n8760 & ~n52059 ) ;
  assign n52061 = n52060 ^ n44040 ^ n19511 ;
  assign n52062 = n24093 & ~n25718 ;
  assign n52063 = n52062 ^ n4022 ^ 1'b0 ;
  assign n52064 = n39753 ^ n30225 ^ n19792 ;
  assign n52065 = n52064 ^ n6218 ^ n5757 ;
  assign n52066 = n5414 | n36756 ;
  assign n52067 = ( n13256 & ~n19270 ) | ( n13256 & n52066 ) | ( ~n19270 & n52066 ) ;
  assign n52068 = n50256 ^ n49265 ^ n39848 ;
  assign n52069 = n52067 & ~n52068 ;
  assign n52070 = n52065 & n52069 ;
  assign n52071 = n39595 ^ n19107 ^ n18767 ;
  assign n52072 = ( n7608 & n25667 ) | ( n7608 & n52071 ) | ( n25667 & n52071 ) ;
  assign n52073 = n25851 ^ n363 ^ 1'b0 ;
  assign n52074 = n51527 ^ n11934 ^ n6072 ;
  assign n52075 = ( n3237 & n19981 ) | ( n3237 & n26595 ) | ( n19981 & n26595 ) ;
  assign n52076 = ( n11124 & n13450 ) | ( n11124 & n29378 ) | ( n13450 & n29378 ) ;
  assign n52077 = n2129 & n44028 ;
  assign n52078 = ~n52076 & n52077 ;
  assign n52079 = ( n5302 & n52075 ) | ( n5302 & ~n52078 ) | ( n52075 & ~n52078 ) ;
  assign n52080 = ( n17406 & n25878 ) | ( n17406 & ~n44768 ) | ( n25878 & ~n44768 ) ;
  assign n52081 = ( n4178 & n19330 ) | ( n4178 & n52080 ) | ( n19330 & n52080 ) ;
  assign n52082 = n52081 ^ n44551 ^ n24701 ;
  assign n52083 = ( n6188 & n19175 ) | ( n6188 & n52082 ) | ( n19175 & n52082 ) ;
  assign n52084 = n29516 ^ n22429 ^ n14112 ;
  assign n52085 = ( n11559 & n13439 ) | ( n11559 & ~n52084 ) | ( n13439 & ~n52084 ) ;
  assign n52086 = ( n5876 & n21361 ) | ( n5876 & ~n27655 ) | ( n21361 & ~n27655 ) ;
  assign n52087 = ( n20054 & ~n21265 ) | ( n20054 & n52086 ) | ( ~n21265 & n52086 ) ;
  assign n52088 = n40613 ^ n31317 ^ n4184 ;
  assign n52089 = n26744 & ~n34208 ;
  assign n52090 = n22583 & n52089 ;
  assign n52091 = ~n15971 & n19898 ;
  assign n52092 = n52091 ^ n51098 ^ 1'b0 ;
  assign n52093 = n39656 ^ n31697 ^ 1'b0 ;
  assign n52094 = ( n18050 & ~n38351 ) | ( n18050 & n43126 ) | ( ~n38351 & n43126 ) ;
  assign n52095 = n30902 ^ n5944 ^ 1'b0 ;
  assign n52096 = ( ~n11276 & n52094 ) | ( ~n11276 & n52095 ) | ( n52094 & n52095 ) ;
  assign n52097 = ( n5829 & n6425 ) | ( n5829 & n18025 ) | ( n6425 & n18025 ) ;
  assign n52098 = n34568 ^ n25709 ^ n9193 ;
  assign n52099 = ( ~n30074 & n52097 ) | ( ~n30074 & n52098 ) | ( n52097 & n52098 ) ;
  assign n52100 = ( n1597 & n27485 ) | ( n1597 & ~n31437 ) | ( n27485 & ~n31437 ) ;
  assign n52101 = n50533 ^ n43756 ^ n14052 ;
  assign n52102 = ( n25384 & n44914 ) | ( n25384 & ~n46900 ) | ( n44914 & ~n46900 ) ;
  assign n52103 = ( n681 & ~n2835 ) | ( n681 & n24920 ) | ( ~n2835 & n24920 ) ;
  assign n52104 = ( n42027 & n49979 ) | ( n42027 & ~n52103 ) | ( n49979 & ~n52103 ) ;
  assign n52105 = ( n8767 & n34229 ) | ( n8767 & ~n52104 ) | ( n34229 & ~n52104 ) ;
  assign n52106 = n19915 ^ n11204 ^ 1'b0 ;
  assign n52107 = n38908 | n52106 ;
  assign n52108 = n26182 ^ n24290 ^ 1'b0 ;
  assign n52109 = n27669 & n52108 ;
  assign n52110 = ( n34117 & n52107 ) | ( n34117 & n52109 ) | ( n52107 & n52109 ) ;
  assign n52111 = ( n17881 & ~n20858 ) | ( n17881 & n36162 ) | ( ~n20858 & n36162 ) ;
  assign n52112 = ( ~n10720 & n20343 ) | ( ~n10720 & n27377 ) | ( n20343 & n27377 ) ;
  assign n52113 = ~n45508 & n52112 ;
  assign n52114 = ( ~n2958 & n24672 ) | ( ~n2958 & n52113 ) | ( n24672 & n52113 ) ;
  assign n52115 = n39035 ^ n30212 ^ n20341 ;
  assign n52116 = n25681 ^ n9989 ^ n1611 ;
  assign n52117 = ( n11286 & n41146 ) | ( n11286 & n52116 ) | ( n41146 & n52116 ) ;
  assign n52118 = n46838 ^ n31514 ^ n6458 ;
  assign n52119 = n22262 ^ n16477 ^ n8096 ;
  assign n52120 = ( ~n5339 & n42761 ) | ( ~n5339 & n52119 ) | ( n42761 & n52119 ) ;
  assign n52121 = ( ~n8578 & n11613 ) | ( ~n8578 & n21008 ) | ( n11613 & n21008 ) ;
  assign n52122 = n38799 ^ n10721 ^ n6977 ;
  assign n52123 = ( n10673 & ~n35623 ) | ( n10673 & n52122 ) | ( ~n35623 & n52122 ) ;
  assign n52124 = n44443 ^ n39647 ^ n15137 ;
  assign n52125 = ( ~n25825 & n27987 ) | ( ~n25825 & n41104 ) | ( n27987 & n41104 ) ;
  assign n52126 = ( n52123 & ~n52124 ) | ( n52123 & n52125 ) | ( ~n52124 & n52125 ) ;
  assign n52127 = ( n24454 & ~n37616 ) | ( n24454 & n52126 ) | ( ~n37616 & n52126 ) ;
  assign n52128 = n46179 ^ n14748 ^ n7332 ;
  assign n52129 = n50191 ^ n40270 ^ n2943 ;
  assign n52130 = ~n15494 & n41959 ;
  assign n52131 = n52130 ^ n3815 ^ 1'b0 ;
  assign n52132 = n11757 ^ n4425 ^ 1'b0 ;
  assign n52133 = ~n26773 & n52132 ;
  assign n52134 = n16488 ^ n6350 ^ n3428 ;
  assign n52135 = ( ~n6381 & n33053 ) | ( ~n6381 & n39601 ) | ( n33053 & n39601 ) ;
  assign n52136 = n22401 ^ n8010 ^ 1'b0 ;
  assign n52137 = n52136 ^ n23740 ^ n20015 ;
  assign n52138 = ( n5925 & n26460 ) | ( n5925 & n34156 ) | ( n26460 & n34156 ) ;
  assign n52139 = n37618 ^ n20660 ^ n2298 ;
  assign n52140 = ~n4465 & n32821 ;
  assign n52141 = n52140 ^ n43695 ^ n13547 ;
  assign n52142 = ( n49783 & n52139 ) | ( n49783 & ~n52141 ) | ( n52139 & ~n52141 ) ;
  assign n52143 = ( n30907 & n52138 ) | ( n30907 & n52142 ) | ( n52138 & n52142 ) ;
  assign n52144 = n42639 ^ n31184 ^ 1'b0 ;
  assign n52145 = n36723 ^ n35177 ^ 1'b0 ;
  assign n52146 = ( n3963 & ~n35721 ) | ( n3963 & n48394 ) | ( ~n35721 & n48394 ) ;
  assign n52147 = n42170 ^ n5005 ^ n2552 ;
  assign n52148 = n36294 ^ n13093 ^ 1'b0 ;
  assign n52149 = n52147 | n52148 ;
  assign n52150 = n19722 ^ n16146 ^ n9080 ;
  assign n52151 = n52150 ^ n26075 ^ n9934 ;
  assign n52152 = n13830 ^ n5852 ^ n3272 ;
  assign n52153 = ( n5091 & ~n18211 ) | ( n5091 & n52152 ) | ( ~n18211 & n52152 ) ;
  assign n52154 = ( n11814 & n34076 ) | ( n11814 & n36847 ) | ( n34076 & n36847 ) ;
  assign n52155 = n36959 ^ n8488 ^ 1'b0 ;
  assign n52156 = ( ~n3870 & n25888 ) | ( ~n3870 & n46893 ) | ( n25888 & n46893 ) ;
  assign n52157 = ( n18247 & ~n25710 ) | ( n18247 & n30647 ) | ( ~n25710 & n30647 ) ;
  assign n52158 = n52157 ^ n50671 ^ n17417 ;
  assign n52159 = n52158 ^ n36011 ^ n14588 ;
  assign n52160 = n27934 ^ n19876 ^ n17646 ;
  assign n52161 = n52160 ^ n27862 ^ n20908 ;
  assign n52162 = n18654 ^ n15517 ^ n14220 ;
  assign n52163 = ( n2627 & n36222 ) | ( n2627 & n40729 ) | ( n36222 & n40729 ) ;
  assign n52164 = ( n24119 & ~n27943 ) | ( n24119 & n28512 ) | ( ~n27943 & n28512 ) ;
  assign n52165 = n52164 ^ n10873 ^ 1'b0 ;
  assign n52166 = ~n5997 & n52165 ;
  assign n52167 = n37731 ^ n13246 ^ n9110 ;
  assign n52168 = n6126 ^ n1668 ^ 1'b0 ;
  assign n52169 = n52168 ^ n32684 ^ n7363 ;
  assign n52170 = ~n42882 & n52169 ;
  assign n52171 = ~n52167 & n52170 ;
  assign n52172 = ( n37032 & n41113 ) | ( n37032 & ~n52043 ) | ( n41113 & ~n52043 ) ;
  assign n52173 = n48799 ^ n1408 ^ 1'b0 ;
  assign n52174 = ~n13251 & n46995 ;
  assign n52175 = ( n5140 & ~n16211 ) | ( n5140 & n52174 ) | ( ~n16211 & n52174 ) ;
  assign n52176 = n8291 & ~n15881 ;
  assign n52177 = n52176 ^ n4234 ^ 1'b0 ;
  assign n52178 = ( n16888 & ~n52175 ) | ( n16888 & n52177 ) | ( ~n52175 & n52177 ) ;
  assign n52179 = n40110 & ~n52178 ;
  assign n52180 = n37856 ^ n34004 ^ n18597 ;
  assign n52181 = n52180 ^ n19323 ^ n2723 ;
  assign n52182 = n52181 ^ n50236 ^ n41583 ;
  assign n52183 = n27060 ^ n4462 ^ n1028 ;
  assign n52184 = ( n25510 & n26402 ) | ( n25510 & n52183 ) | ( n26402 & n52183 ) ;
  assign n52185 = ( n13341 & n39207 ) | ( n13341 & ~n52184 ) | ( n39207 & ~n52184 ) ;
  assign n52186 = ( n22835 & ~n25575 ) | ( n22835 & n29497 ) | ( ~n25575 & n29497 ) ;
  assign n52187 = ( n5098 & n7129 ) | ( n5098 & ~n19733 ) | ( n7129 & ~n19733 ) ;
  assign n52188 = n52187 ^ n12911 ^ n2968 ;
  assign n52189 = ( n1631 & ~n2780 ) | ( n1631 & n46127 ) | ( ~n2780 & n46127 ) ;
  assign n52190 = n51321 ^ n14285 ^ n9227 ;
  assign n52191 = n5069 & n52190 ;
  assign n52192 = ( ~n25900 & n50278 ) | ( ~n25900 & n52191 ) | ( n50278 & n52191 ) ;
  assign n52193 = ( ~n9711 & n18966 ) | ( ~n9711 & n38252 ) | ( n18966 & n38252 ) ;
  assign n52194 = ( n7324 & n50445 ) | ( n7324 & n52193 ) | ( n50445 & n52193 ) ;
  assign n52195 = n15149 | n52194 ;
  assign n52196 = ( n25786 & n29872 ) | ( n25786 & n52195 ) | ( n29872 & n52195 ) ;
  assign n52197 = n30379 | n52196 ;
  assign n52198 = n34066 & ~n52197 ;
  assign n52199 = ( n11319 & n21428 ) | ( n11319 & n29950 ) | ( n21428 & n29950 ) ;
  assign n52200 = ( n9659 & ~n21470 ) | ( n9659 & n44848 ) | ( ~n21470 & n44848 ) ;
  assign n52201 = ( n25195 & n31597 ) | ( n25195 & n52200 ) | ( n31597 & n52200 ) ;
  assign n52202 = n51028 ^ n2099 ^ 1'b0 ;
  assign n52203 = n52202 ^ n27650 ^ n9030 ;
  assign n52204 = n15404 ^ n10793 ^ 1'b0 ;
  assign n52205 = n9322 & n52204 ;
  assign n52206 = ( n25906 & n39864 ) | ( n25906 & n52205 ) | ( n39864 & n52205 ) ;
  assign n52207 = ( n3764 & n26742 ) | ( n3764 & ~n52206 ) | ( n26742 & ~n52206 ) ;
  assign n52212 = n12541 ^ n7615 ^ x2 ;
  assign n52208 = ( ~n609 & n5229 ) | ( ~n609 & n7015 ) | ( n5229 & n7015 ) ;
  assign n52209 = ( n25090 & ~n41288 ) | ( n25090 & n52208 ) | ( ~n41288 & n52208 ) ;
  assign n52210 = ( n9166 & n52195 ) | ( n9166 & ~n52209 ) | ( n52195 & ~n52209 ) ;
  assign n52211 = n52210 ^ n26770 ^ n20080 ;
  assign n52213 = n52212 ^ n52211 ^ n3222 ;
  assign n52214 = n24602 ^ n21707 ^ n5721 ;
  assign n52215 = ( ~n2733 & n32438 ) | ( ~n2733 & n52214 ) | ( n32438 & n52214 ) ;
  assign n52216 = n42305 ^ n39496 ^ n13179 ;
  assign n52217 = n52216 ^ n34360 ^ n7533 ;
  assign n52218 = ( n3303 & n6926 ) | ( n3303 & n9245 ) | ( n6926 & n9245 ) ;
  assign n52219 = n5901 & n7392 ;
  assign n52220 = ~x36 & n52219 ;
  assign n52221 = ( x235 & n3155 ) | ( x235 & n52220 ) | ( n3155 & n52220 ) ;
  assign n52222 = ( n11938 & n37436 ) | ( n11938 & n52221 ) | ( n37436 & n52221 ) ;
  assign n52223 = n17899 & n52222 ;
  assign n52224 = n52218 & n52223 ;
  assign n52225 = ( ~n17056 & n38455 ) | ( ~n17056 & n41130 ) | ( n38455 & n41130 ) ;
  assign n52226 = n52225 ^ n9926 ^ n5346 ;
  assign n52227 = n27464 ^ n17379 ^ n11771 ;
  assign n52228 = ( n11558 & n11919 ) | ( n11558 & n52227 ) | ( n11919 & n52227 ) ;
  assign n52229 = n22800 ^ n16116 ^ n1653 ;
  assign n52230 = n49630 ^ n31899 ^ n1132 ;
  assign n52231 = n26303 ^ n14169 ^ n7789 ;
  assign n52232 = n23785 ^ n18100 ^ n17442 ;
  assign n52233 = n12394 & ~n37907 ;
  assign n52234 = ~n15017 & n52233 ;
  assign n52235 = ( ~n43446 & n46733 ) | ( ~n43446 & n52234 ) | ( n46733 & n52234 ) ;
  assign n52236 = n52235 ^ n10629 ^ x37 ;
  assign n52237 = ( n15958 & n17475 ) | ( n15958 & ~n37020 ) | ( n17475 & ~n37020 ) ;
  assign n52240 = n49993 ^ n26493 ^ n6494 ;
  assign n52238 = ( n265 & n2483 ) | ( n265 & n8433 ) | ( n2483 & n8433 ) ;
  assign n52239 = n52238 ^ n19326 ^ n7502 ;
  assign n52241 = n52240 ^ n52239 ^ n22516 ;
  assign n52242 = ~n36430 & n44195 ;
  assign n52243 = ~n30700 & n52242 ;
  assign n52248 = ( n11364 & ~n33031 ) | ( n11364 & n34039 ) | ( ~n33031 & n34039 ) ;
  assign n52249 = ( ~n6717 & n21135 ) | ( ~n6717 & n52248 ) | ( n21135 & n52248 ) ;
  assign n52245 = n22721 ^ n13046 ^ n3294 ;
  assign n52244 = n4927 | n9165 ;
  assign n52246 = n52245 ^ n52244 ^ 1'b0 ;
  assign n52247 = n52246 ^ n19133 ^ n6281 ;
  assign n52250 = n52249 ^ n52247 ^ n23243 ;
  assign n52251 = n20364 ^ n5326 ^ 1'b0 ;
  assign n52252 = ( n43937 & n45583 ) | ( n43937 & n51134 ) | ( n45583 & n51134 ) ;
  assign n52253 = n52252 ^ n49514 ^ n11034 ;
  assign n52254 = ( n3119 & ~n52251 ) | ( n3119 & n52253 ) | ( ~n52251 & n52253 ) ;
  assign n52255 = ( n3435 & n30346 ) | ( n3435 & ~n35998 ) | ( n30346 & ~n35998 ) ;
  assign n52256 = n44073 ^ n4040 ^ 1'b0 ;
  assign n52257 = n52256 ^ n34879 ^ n32680 ;
  assign n52258 = n52257 ^ n18462 ^ n16335 ;
  assign n52259 = ( n2307 & ~n10550 ) | ( n2307 & n30458 ) | ( ~n10550 & n30458 ) ;
  assign n52260 = n52259 ^ n39967 ^ n10316 ;
  assign n52261 = ( n8318 & ~n29540 ) | ( n8318 & n30656 ) | ( ~n29540 & n30656 ) ;
  assign n52264 = ( ~n5148 & n7819 ) | ( ~n5148 & n41809 ) | ( n7819 & n41809 ) ;
  assign n52262 = n12565 ^ n4306 ^ 1'b0 ;
  assign n52263 = n38099 | n52262 ;
  assign n52265 = n52264 ^ n52263 ^ n6335 ;
  assign n52266 = n52265 ^ n28210 ^ n967 ;
  assign n52267 = ( n8092 & ~n30154 ) | ( n8092 & n52266 ) | ( ~n30154 & n52266 ) ;
  assign n52268 = ( n22222 & n52261 ) | ( n22222 & ~n52267 ) | ( n52261 & ~n52267 ) ;
  assign n52269 = ( n2011 & ~n3069 ) | ( n2011 & n8078 ) | ( ~n3069 & n8078 ) ;
  assign n52270 = ~n19519 & n29157 ;
  assign n52271 = ( n537 & n6180 ) | ( n537 & ~n52270 ) | ( n6180 & ~n52270 ) ;
  assign n52272 = ( ~n37729 & n52269 ) | ( ~n37729 & n52271 ) | ( n52269 & n52271 ) ;
  assign n52273 = ( n3217 & n20171 ) | ( n3217 & n38171 ) | ( n20171 & n38171 ) ;
  assign n52274 = ( n25977 & n42432 ) | ( n25977 & ~n52273 ) | ( n42432 & ~n52273 ) ;
  assign n52275 = n32147 | n46354 ;
  assign n52276 = n52275 ^ n20433 ^ n12378 ;
  assign n52277 = n5079 & ~n26952 ;
  assign n52278 = n31049 & n52277 ;
  assign n52279 = ( n14189 & n42761 ) | ( n14189 & ~n50974 ) | ( n42761 & ~n50974 ) ;
  assign n52280 = ( n3259 & n8315 ) | ( n3259 & n50844 ) | ( n8315 & n50844 ) ;
  assign n52281 = ( n20461 & ~n51835 ) | ( n20461 & n52280 ) | ( ~n51835 & n52280 ) ;
  assign n52282 = n9857 ^ n3455 ^ 1'b0 ;
  assign n52283 = n893 | n52282 ;
  assign n52284 = n52283 ^ n42310 ^ n29262 ;
  assign n52285 = ( n1204 & n3989 ) | ( n1204 & ~n23169 ) | ( n3989 & ~n23169 ) ;
  assign n52286 = n52285 ^ n22042 ^ 1'b0 ;
  assign n52287 = n38377 & n52286 ;
  assign n52288 = n8877 & n52287 ;
  assign n52289 = n50581 ^ n27256 ^ 1'b0 ;
  assign n52290 = n46546 ^ n36083 ^ n22445 ;
  assign n52291 = n45235 ^ n14785 ^ n1046 ;
  assign n52292 = ( ~n17834 & n25576 ) | ( ~n17834 & n52291 ) | ( n25576 & n52291 ) ;
  assign n52295 = ( x71 & n493 ) | ( x71 & ~n25810 ) | ( n493 & ~n25810 ) ;
  assign n52293 = n25624 ^ n9580 ^ 1'b0 ;
  assign n52294 = ( n18575 & n26654 ) | ( n18575 & n52293 ) | ( n26654 & n52293 ) ;
  assign n52296 = n52295 ^ n52294 ^ n6100 ;
  assign n52297 = n44421 | n52296 ;
  assign n52298 = n6989 & ~n52297 ;
  assign n52299 = n28948 ^ n27224 ^ 1'b0 ;
  assign n52300 = ( n9308 & ~n21108 ) | ( n9308 & n33460 ) | ( ~n21108 & n33460 ) ;
  assign n52301 = ( n49862 & n52299 ) | ( n49862 & ~n52300 ) | ( n52299 & ~n52300 ) ;
  assign n52302 = n25304 ^ n16820 ^ n2673 ;
  assign n52303 = n34362 & ~n52302 ;
  assign n52304 = n52301 & n52303 ;
  assign n52305 = ( n335 & ~n2183 ) | ( n335 & n4936 ) | ( ~n2183 & n4936 ) ;
  assign n52306 = n52305 ^ n22097 ^ n12188 ;
  assign n52307 = ( n24544 & n26298 ) | ( n24544 & n29210 ) | ( n26298 & n29210 ) ;
  assign n52309 = n32334 ^ n26536 ^ n257 ;
  assign n52310 = ( n5400 & n16213 ) | ( n5400 & n52309 ) | ( n16213 & n52309 ) ;
  assign n52311 = ( n5388 & n13294 ) | ( n5388 & ~n52310 ) | ( n13294 & ~n52310 ) ;
  assign n52308 = ( ~n1308 & n5275 ) | ( ~n1308 & n36271 ) | ( n5275 & n36271 ) ;
  assign n52312 = n52311 ^ n52308 ^ n13735 ;
  assign n52313 = n2412 & n20773 ;
  assign n52314 = n52313 ^ n17591 ^ 1'b0 ;
  assign n52315 = n52314 ^ n36238 ^ n16304 ;
  assign n52316 = ( n293 & ~n38987 ) | ( n293 & n40512 ) | ( ~n38987 & n40512 ) ;
  assign n52317 = n50146 ^ n16355 ^ n14732 ;
  assign n52318 = ( n9836 & ~n27686 ) | ( n9836 & n36764 ) | ( ~n27686 & n36764 ) ;
  assign n52319 = ( n8743 & ~n32979 ) | ( n8743 & n52318 ) | ( ~n32979 & n52318 ) ;
  assign n52320 = n44298 ^ n14591 ^ n8616 ;
  assign n52324 = n45569 ^ n37427 ^ 1'b0 ;
  assign n52325 = n40974 & ~n52324 ;
  assign n52323 = n25850 & ~n33546 ;
  assign n52326 = n52325 ^ n52323 ^ 1'b0 ;
  assign n52321 = n44572 ^ n34016 ^ n4911 ;
  assign n52322 = ~n44918 & n52321 ;
  assign n52327 = n52326 ^ n52322 ^ 1'b0 ;
  assign n52328 = n11604 & ~n40167 ;
  assign n52329 = ( n2942 & n12779 ) | ( n2942 & n52328 ) | ( n12779 & n52328 ) ;
  assign n52330 = ~n5837 & n35245 ;
  assign n52331 = ( n22830 & n25110 ) | ( n22830 & ~n52330 ) | ( n25110 & ~n52330 ) ;
  assign n52332 = ( ~n20229 & n46552 ) | ( ~n20229 & n50483 ) | ( n46552 & n50483 ) ;
  assign n52333 = n17611 ^ n8546 ^ n4980 ;
  assign n52334 = n52333 ^ n21595 ^ n5195 ;
  assign n52335 = ( ~n959 & n17965 ) | ( ~n959 & n34339 ) | ( n17965 & n34339 ) ;
  assign n52336 = ( n27419 & n45762 ) | ( n27419 & n52335 ) | ( n45762 & n52335 ) ;
  assign n52337 = n52336 ^ n21371 ^ n2268 ;
  assign n52338 = n17663 ^ n15296 ^ n10791 ;
  assign n52339 = ( n47073 & n48286 ) | ( n47073 & n52338 ) | ( n48286 & n52338 ) ;
  assign n52340 = ( n17374 & n27650 ) | ( n17374 & n52339 ) | ( n27650 & n52339 ) ;
  assign n52341 = n12938 | n22821 ;
  assign n52342 = ( n43799 & n43982 ) | ( n43799 & n52341 ) | ( n43982 & n52341 ) ;
  assign n52343 = ( n18575 & n29520 ) | ( n18575 & n47609 ) | ( n29520 & n47609 ) ;
  assign n52344 = n24611 ^ n23848 ^ 1'b0 ;
  assign n52345 = ( ~n2748 & n8238 ) | ( ~n2748 & n47218 ) | ( n8238 & n47218 ) ;
  assign n52346 = n45501 ^ n25933 ^ n1615 ;
  assign n52347 = ( n16072 & ~n38102 ) | ( n16072 & n52346 ) | ( ~n38102 & n52346 ) ;
  assign n52348 = ( n14542 & ~n14726 ) | ( n14542 & n45285 ) | ( ~n14726 & n45285 ) ;
  assign n52349 = n26003 ^ n21823 ^ 1'b0 ;
  assign n52350 = n52349 ^ n30916 ^ n6299 ;
  assign n52354 = n16441 & ~n28081 ;
  assign n52355 = n52354 ^ n37802 ^ 1'b0 ;
  assign n52351 = n45426 ^ n31778 ^ n1805 ;
  assign n52352 = ~n6042 & n42608 ;
  assign n52353 = ( n10925 & n52351 ) | ( n10925 & ~n52352 ) | ( n52351 & ~n52352 ) ;
  assign n52356 = n52355 ^ n52353 ^ n16967 ;
  assign n52357 = ( n8762 & n35047 ) | ( n8762 & ~n39923 ) | ( n35047 & ~n39923 ) ;
  assign n52358 = n52357 ^ n49829 ^ n23750 ;
  assign n52359 = n23825 ^ n22864 ^ n18296 ;
  assign n52360 = ( n13100 & n18077 ) | ( n13100 & n52359 ) | ( n18077 & n52359 ) ;
  assign n52361 = n17520 ^ n12280 ^ n10280 ;
  assign n52362 = ( n13722 & n16328 ) | ( n13722 & n24580 ) | ( n16328 & n24580 ) ;
  assign n52363 = ( n25059 & n37227 ) | ( n25059 & ~n42862 ) | ( n37227 & ~n42862 ) ;
  assign n52364 = ( ~n52361 & n52362 ) | ( ~n52361 & n52363 ) | ( n52362 & n52363 ) ;
  assign n52365 = ( ~n19052 & n52360 ) | ( ~n19052 & n52364 ) | ( n52360 & n52364 ) ;
  assign n52366 = n3219 & ~n20279 ;
  assign n52367 = n52366 ^ n28111 ^ 1'b0 ;
  assign n52368 = n12523 ^ n4574 ^ n3784 ;
  assign n52369 = n52368 ^ n28930 ^ n9667 ;
  assign n52370 = n21691 ^ n16803 ^ n579 ;
  assign n52371 = n52370 ^ n21502 ^ n19693 ;
  assign n52372 = ( n10953 & n21291 ) | ( n10953 & n52371 ) | ( n21291 & n52371 ) ;
  assign n52374 = n45368 ^ n30578 ^ n27462 ;
  assign n52373 = n13603 ^ n7130 ^ n5382 ;
  assign n52375 = n52374 ^ n52373 ^ n3779 ;
  assign n52376 = ( n5390 & n42624 ) | ( n5390 & ~n52375 ) | ( n42624 & ~n52375 ) ;
  assign n52377 = n16834 ^ n2190 ^ 1'b0 ;
  assign n52378 = ~n48910 & n52377 ;
  assign n52379 = n52378 ^ n33167 ^ n28976 ;
  assign n52380 = n42634 ^ n20640 ^ n9980 ;
  assign n52382 = n41883 ^ n20001 ^ n13974 ;
  assign n52383 = ( n12693 & n23449 ) | ( n12693 & n52382 ) | ( n23449 & n52382 ) ;
  assign n52381 = n18657 ^ n10490 ^ n6638 ;
  assign n52384 = n52383 ^ n52381 ^ n26630 ;
  assign n52385 = ( n1320 & n10849 ) | ( n1320 & n52384 ) | ( n10849 & n52384 ) ;
  assign n52386 = ( n1614 & ~n13940 ) | ( n1614 & n52385 ) | ( ~n13940 & n52385 ) ;
  assign n52387 = ( n696 & n18085 ) | ( n696 & ~n52386 ) | ( n18085 & ~n52386 ) ;
  assign n52388 = ( n11147 & n12983 ) | ( n11147 & n20549 ) | ( n12983 & n20549 ) ;
  assign n52389 = ( ~n340 & n21703 ) | ( ~n340 & n52388 ) | ( n21703 & n52388 ) ;
  assign n52390 = ( n2411 & n6410 ) | ( n2411 & n52389 ) | ( n6410 & n52389 ) ;
  assign n52391 = n52390 ^ n36260 ^ n35135 ;
  assign n52392 = ( n28328 & n32183 ) | ( n28328 & n52391 ) | ( n32183 & n52391 ) ;
  assign n52393 = ( n15438 & n35982 ) | ( n15438 & ~n45100 ) | ( n35982 & ~n45100 ) ;
  assign n52394 = n52393 ^ n34010 ^ n30967 ;
  assign n52395 = n30308 ^ n7636 ^ 1'b0 ;
  assign n52396 = n18842 & ~n52395 ;
  assign n52397 = n52396 ^ n52330 ^ 1'b0 ;
  assign n52398 = n52397 ^ n46698 ^ n26759 ;
  assign n52399 = n20924 ^ n20579 ^ 1'b0 ;
  assign n52400 = n52398 | n52399 ;
  assign n52401 = ( n5690 & n13044 ) | ( n5690 & n41148 ) | ( n13044 & n41148 ) ;
  assign n52402 = n52401 ^ n39974 ^ n16574 ;
  assign n52403 = n32295 ^ n29392 ^ n21042 ;
  assign n52404 = n858 & ~n6040 ;
  assign n52405 = ( n37281 & n44311 ) | ( n37281 & ~n52404 ) | ( n44311 & ~n52404 ) ;
  assign n52406 = n12898 & n27176 ;
  assign n52407 = n52406 ^ n21436 ^ 1'b0 ;
  assign n52408 = n52407 ^ n24355 ^ 1'b0 ;
  assign n52410 = n8524 ^ n530 ^ 1'b0 ;
  assign n52409 = n34552 ^ n20632 ^ n10145 ;
  assign n52411 = n52410 ^ n52409 ^ 1'b0 ;
  assign n52415 = ( ~n1108 & n7486 ) | ( ~n1108 & n13506 ) | ( n7486 & n13506 ) ;
  assign n52416 = ( n15058 & ~n19198 ) | ( n15058 & n52415 ) | ( ~n19198 & n52415 ) ;
  assign n52417 = n52416 ^ n30772 ^ n12782 ;
  assign n52413 = ( x113 & n3768 ) | ( x113 & ~n16604 ) | ( n3768 & ~n16604 ) ;
  assign n52414 = ( n11970 & n20084 ) | ( n11970 & ~n52413 ) | ( n20084 & ~n52413 ) ;
  assign n52418 = n52417 ^ n52414 ^ n8349 ;
  assign n52412 = n47090 ^ n36221 ^ n4364 ;
  assign n52419 = n52418 ^ n52412 ^ n14405 ;
  assign n52420 = n25257 ^ n4118 ^ n3659 ;
  assign n52421 = n52420 ^ n1593 ^ 1'b0 ;
  assign n52422 = n52421 ^ n47592 ^ 1'b0 ;
  assign n52423 = ~n3987 & n16970 ;
  assign n52424 = ~n4785 & n52423 ;
  assign n52425 = ( ~n19233 & n43959 ) | ( ~n19233 & n52424 ) | ( n43959 & n52424 ) ;
  assign n52426 = n52425 ^ n9412 ^ 1'b0 ;
  assign n52427 = n10969 ^ n7966 ^ 1'b0 ;
  assign n52428 = n464 & n52427 ;
  assign n52429 = ( n4930 & n16095 ) | ( n4930 & n52428 ) | ( n16095 & n52428 ) ;
  assign n52430 = n52429 ^ n20416 ^ 1'b0 ;
  assign n52431 = ~n39388 & n52430 ;
  assign n52432 = ~n17048 & n32052 ;
  assign n52433 = ( ~n8216 & n48470 ) | ( ~n8216 & n52432 ) | ( n48470 & n52432 ) ;
  assign n52434 = n29221 ^ n15349 ^ n13506 ;
  assign n52435 = n41167 ^ n34988 ^ n29190 ;
  assign n52436 = ( n12963 & n35991 ) | ( n12963 & n52435 ) | ( n35991 & n52435 ) ;
  assign n52437 = n32093 ^ n12300 ^ n7982 ;
  assign n52438 = ( n17867 & n36044 ) | ( n17867 & ~n52437 ) | ( n36044 & ~n52437 ) ;
  assign n52439 = ~n15702 & n39537 ;
  assign n52440 = ( n8763 & n9038 ) | ( n8763 & n11794 ) | ( n9038 & n11794 ) ;
  assign n52441 = n52440 ^ n7890 ^ n4403 ;
  assign n52442 = n19041 ^ n7232 ^ n6930 ;
  assign n52443 = ( n52439 & n52441 ) | ( n52439 & ~n52442 ) | ( n52441 & ~n52442 ) ;
  assign n52444 = n52443 ^ n17711 ^ n3067 ;
  assign n52446 = n21801 ^ n15279 ^ n7232 ;
  assign n52445 = n5386 & n19786 ;
  assign n52447 = n52446 ^ n52445 ^ 1'b0 ;
  assign n52448 = ( ~n19307 & n25851 ) | ( ~n19307 & n52447 ) | ( n25851 & n52447 ) ;
  assign n52449 = n17046 ^ n14225 ^ n10544 ;
  assign n52450 = ( n21442 & n52448 ) | ( n21442 & ~n52449 ) | ( n52448 & ~n52449 ) ;
  assign n52455 = n32486 ^ n14638 ^ 1'b0 ;
  assign n52451 = n5908 ^ n5536 ^ n1726 ;
  assign n52452 = ( n4668 & n23399 ) | ( n4668 & ~n52451 ) | ( n23399 & ~n52451 ) ;
  assign n52453 = n52452 ^ n48998 ^ n23081 ;
  assign n52454 = n52453 ^ n31989 ^ n15727 ;
  assign n52456 = n52455 ^ n52454 ^ n14702 ;
  assign n52457 = n52456 ^ n45145 ^ n561 ;
  assign n52458 = ( ~n2875 & n6950 ) | ( ~n2875 & n14109 ) | ( n6950 & n14109 ) ;
  assign n52459 = ( n16047 & ~n24596 ) | ( n16047 & n52458 ) | ( ~n24596 & n52458 ) ;
  assign n52460 = n46434 ^ n36203 ^ 1'b0 ;
  assign n52461 = n23553 | n52460 ;
  assign n52462 = n3683 & ~n52461 ;
  assign n52463 = n52462 ^ n25138 ^ 1'b0 ;
  assign n52464 = ( n533 & n25151 ) | ( n533 & ~n51964 ) | ( n25151 & ~n51964 ) ;
  assign n52465 = n20389 ^ n16896 ^ 1'b0 ;
  assign n52466 = n52464 & n52465 ;
  assign n52467 = n51532 ^ n38401 ^ n26416 ;
  assign n52468 = ( n10346 & n20632 ) | ( n10346 & n27266 ) | ( n20632 & n27266 ) ;
  assign n52469 = n24381 ^ n3121 ^ n575 ;
  assign n52470 = ( ~n21571 & n52468 ) | ( ~n21571 & n52469 ) | ( n52468 & n52469 ) ;
  assign n52471 = n52470 ^ n29520 ^ n15095 ;
  assign n52472 = ( n3750 & n6476 ) | ( n3750 & n16702 ) | ( n6476 & n16702 ) ;
  assign n52473 = n52472 ^ n37265 ^ n8829 ;
  assign n52474 = n52094 ^ n48367 ^ n10271 ;
  assign n52475 = n13134 & ~n31081 ;
  assign n52476 = n52475 ^ n52067 ^ n17640 ;
  assign n52477 = ( n37641 & n46089 ) | ( n37641 & ~n50629 ) | ( n46089 & ~n50629 ) ;
  assign n52478 = n35782 ^ n8608 ^ 1'b0 ;
  assign n52479 = n52478 ^ n22482 ^ x125 ;
  assign n52480 = n52479 ^ n3696 ^ 1'b0 ;
  assign n52481 = n25584 ^ n18456 ^ n7755 ;
  assign n52482 = ( n7770 & n23265 ) | ( n7770 & n52481 ) | ( n23265 & n52481 ) ;
  assign n52483 = n16117 ^ n7544 ^ 1'b0 ;
  assign n52484 = n52482 | n52483 ;
  assign n52485 = n18415 ^ n2367 ^ 1'b0 ;
  assign n52486 = n3170 ^ n1631 ^ 1'b0 ;
  assign n52487 = ~n26823 & n52486 ;
  assign n52488 = n52487 ^ n45379 ^ n5632 ;
  assign n52489 = n52488 ^ n23955 ^ n1451 ;
  assign n52490 = n16104 ^ n9404 ^ 1'b0 ;
  assign n52491 = ( n7276 & ~n12842 ) | ( n7276 & n30457 ) | ( ~n12842 & n30457 ) ;
  assign n52492 = n52293 ^ n3005 ^ n662 ;
  assign n52493 = n52492 ^ n18604 ^ n12859 ;
  assign n52494 = ( ~n2028 & n20538 ) | ( ~n2028 & n52493 ) | ( n20538 & n52493 ) ;
  assign n52495 = n27090 ^ n26724 ^ n21361 ;
  assign n52496 = ( n23549 & ~n37132 ) | ( n23549 & n52495 ) | ( ~n37132 & n52495 ) ;
  assign n52497 = ( n691 & n8118 ) | ( n691 & n13439 ) | ( n8118 & n13439 ) ;
  assign n52498 = n11302 | n52497 ;
  assign n52499 = n52498 ^ n52119 ^ 1'b0 ;
  assign n52500 = n52499 ^ n36154 ^ n28617 ;
  assign n52501 = n52500 ^ n33518 ^ n5395 ;
  assign n52502 = n50397 ^ n3314 ^ 1'b0 ;
  assign n52503 = n21082 ^ n5634 ^ n3950 ;
  assign n52504 = n27679 ^ n14107 ^ n6558 ;
  assign n52505 = n8692 & n16430 ;
  assign n52506 = ~n52504 & n52505 ;
  assign n52507 = ( n19731 & ~n52503 ) | ( n19731 & n52506 ) | ( ~n52503 & n52506 ) ;
  assign n52508 = n26165 & n42187 ;
  assign n52509 = n2292 & n52508 ;
  assign n52510 = n8983 & ~n9057 ;
  assign n52511 = n52509 & n52510 ;
  assign n52512 = ( ~n7400 & n18263 ) | ( ~n7400 & n30767 ) | ( n18263 & n30767 ) ;
  assign n52513 = n1977 & ~n29928 ;
  assign n52514 = n52512 & n52513 ;
  assign n52515 = ( n27646 & ~n32998 ) | ( n27646 & n51653 ) | ( ~n32998 & n51653 ) ;
  assign n52516 = ( n3453 & ~n12801 ) | ( n3453 & n27368 ) | ( ~n12801 & n27368 ) ;
  assign n52517 = ( n21074 & n46577 ) | ( n21074 & ~n52516 ) | ( n46577 & ~n52516 ) ;
  assign n52518 = n44952 ^ n19956 ^ n8561 ;
  assign n52519 = n52518 ^ n18713 ^ 1'b0 ;
  assign n52521 = n28892 ^ n26119 ^ n24574 ;
  assign n52520 = ( n20349 & ~n25942 ) | ( n20349 & n48857 ) | ( ~n25942 & n48857 ) ;
  assign n52522 = n52521 ^ n52520 ^ n9681 ;
  assign n52523 = ( ~n2141 & n26250 ) | ( ~n2141 & n33550 ) | ( n26250 & n33550 ) ;
  assign n52524 = ( n563 & ~n11339 ) | ( n563 & n14654 ) | ( ~n11339 & n14654 ) ;
  assign n52525 = ( ~n2597 & n52523 ) | ( ~n2597 & n52524 ) | ( n52523 & n52524 ) ;
  assign n52526 = n37486 ^ n4874 ^ x253 ;
  assign n52527 = n35769 ^ n10086 ^ n4606 ;
  assign n52528 = ( n34824 & ~n48392 ) | ( n34824 & n52527 ) | ( ~n48392 & n52527 ) ;
  assign n52529 = ( ~n19621 & n22533 ) | ( ~n19621 & n36709 ) | ( n22533 & n36709 ) ;
  assign n52530 = n21926 | n28281 ;
  assign n52531 = n52530 ^ n18709 ^ 1'b0 ;
  assign n52532 = n22765 & ~n24602 ;
  assign n52533 = ~n19742 & n52532 ;
  assign n52534 = ( ~n2880 & n15430 ) | ( ~n2880 & n27986 ) | ( n15430 & n27986 ) ;
  assign n52535 = ( n18614 & ~n52533 ) | ( n18614 & n52534 ) | ( ~n52533 & n52534 ) ;
  assign n52536 = ( n18572 & n21028 ) | ( n18572 & ~n44236 ) | ( n21028 & ~n44236 ) ;
  assign n52537 = ( n18670 & n19610 ) | ( n18670 & n52536 ) | ( n19610 & n52536 ) ;
  assign n52538 = n34323 ^ n27141 ^ n4646 ;
  assign n52539 = ( n292 & n38293 ) | ( n292 & ~n48669 ) | ( n38293 & ~n48669 ) ;
  assign n52540 = n52539 ^ n45894 ^ n891 ;
  assign n52541 = n35736 ^ n22521 ^ x227 ;
  assign n52542 = n19475 ^ n16975 ^ n9686 ;
  assign n52543 = ( ~x216 & n3888 ) | ( ~x216 & n31180 ) | ( n3888 & n31180 ) ;
  assign n52545 = ( ~n4197 & n5149 ) | ( ~n4197 & n28954 ) | ( n5149 & n28954 ) ;
  assign n52546 = ( n4867 & n18451 ) | ( n4867 & ~n19235 ) | ( n18451 & ~n19235 ) ;
  assign n52547 = n52546 ^ n15057 ^ n4321 ;
  assign n52548 = ( n30392 & ~n52545 ) | ( n30392 & n52547 ) | ( ~n52545 & n52547 ) ;
  assign n52544 = n39504 ^ n14813 ^ n13637 ;
  assign n52549 = n52548 ^ n52544 ^ n24221 ;
  assign n52550 = n4174 | n7042 ;
  assign n52551 = n35426 | n52550 ;
  assign n52552 = n991 & n18867 ;
  assign n52553 = n52552 ^ n30547 ^ 1'b0 ;
  assign n52554 = n52553 ^ n40566 ^ n36777 ;
  assign n52555 = ( n8234 & ~n25322 ) | ( n8234 & n29385 ) | ( ~n25322 & n29385 ) ;
  assign n52556 = ( n8157 & n46638 ) | ( n8157 & n52555 ) | ( n46638 & n52555 ) ;
  assign n52557 = n40707 ^ n34052 ^ n18741 ;
  assign n52558 = n52557 ^ n40906 ^ n36471 ;
  assign n52559 = ( n18123 & n20561 ) | ( n18123 & n41863 ) | ( n20561 & n41863 ) ;
  assign n52560 = ( n891 & ~n44936 ) | ( n891 & n52559 ) | ( ~n44936 & n52559 ) ;
  assign n52561 = ( ~n25937 & n52558 ) | ( ~n25937 & n52560 ) | ( n52558 & n52560 ) ;
  assign n52562 = n18229 ^ n5509 ^ 1'b0 ;
  assign n52563 = ~n7046 & n52562 ;
  assign n52564 = ( n16732 & n23385 ) | ( n16732 & n52563 ) | ( n23385 & n52563 ) ;
  assign n52565 = ( x199 & ~n5403 ) | ( x199 & n10316 ) | ( ~n5403 & n10316 ) ;
  assign n52566 = n22464 & n37502 ;
  assign n52567 = ~n2630 & n3937 ;
  assign n52568 = n52567 ^ n7640 ^ 1'b0 ;
  assign n52569 = ( n26405 & n46093 ) | ( n26405 & n52568 ) | ( n46093 & n52568 ) ;
  assign n52570 = ( n863 & n16239 ) | ( n863 & ~n17204 ) | ( n16239 & ~n17204 ) ;
  assign n52571 = ( n10244 & ~n22840 ) | ( n10244 & n52570 ) | ( ~n22840 & n52570 ) ;
  assign n52575 = ~n14993 & n28327 ;
  assign n52572 = n41473 ^ n33388 ^ 1'b0 ;
  assign n52573 = ( ~n17046 & n46459 ) | ( ~n17046 & n52572 ) | ( n46459 & n52572 ) ;
  assign n52574 = n52573 ^ n35726 ^ n27648 ;
  assign n52576 = n52575 ^ n52574 ^ n23963 ;
  assign n52577 = n31953 ^ n20928 ^ n603 ;
  assign n52578 = n18173 ^ n17139 ^ n11821 ;
  assign n52579 = ( n16709 & n52577 ) | ( n16709 & ~n52578 ) | ( n52577 & ~n52578 ) ;
  assign n52580 = n45436 ^ n11812 ^ n11301 ;
  assign n52581 = ( n21916 & ~n28891 ) | ( n21916 & n40159 ) | ( ~n28891 & n40159 ) ;
  assign n52582 = ( n9885 & n52580 ) | ( n9885 & n52581 ) | ( n52580 & n52581 ) ;
  assign n52583 = ( ~n19376 & n49381 ) | ( ~n19376 & n52582 ) | ( n49381 & n52582 ) ;
  assign n52584 = n39906 ^ n30664 ^ n11051 ;
  assign n52585 = ( n13761 & ~n20267 ) | ( n13761 & n52584 ) | ( ~n20267 & n52584 ) ;
  assign n52586 = n1799 | n16383 ;
  assign n52587 = n52586 ^ n36091 ^ n14599 ;
  assign n52588 = n50977 ^ n30615 ^ n22235 ;
  assign n52589 = n50788 ^ n30853 ^ n2831 ;
  assign n52590 = n52589 ^ n32493 ^ 1'b0 ;
  assign n52591 = n31768 & ~n52590 ;
  assign n52596 = n36751 ^ n3365 ^ n2003 ;
  assign n52593 = n31439 ^ n21820 ^ 1'b0 ;
  assign n52594 = n9509 & n52593 ;
  assign n52592 = n30393 & n41999 ;
  assign n52595 = n52594 ^ n52592 ^ 1'b0 ;
  assign n52597 = n52596 ^ n52595 ^ n6829 ;
  assign n52598 = n34162 ^ n31021 ^ n12198 ;
  assign n52599 = n52598 ^ n28455 ^ 1'b0 ;
  assign n52600 = ( n3214 & ~n50852 ) | ( n3214 & n52599 ) | ( ~n50852 & n52599 ) ;
  assign n52601 = n9387 | n52600 ;
  assign n52602 = n52597 & ~n52601 ;
  assign n52604 = ( ~n25111 & n31272 ) | ( ~n25111 & n45856 ) | ( n31272 & n45856 ) ;
  assign n52603 = n1046 & n18706 ;
  assign n52605 = n52604 ^ n52603 ^ n40219 ;
  assign n52606 = n27757 & n42974 ;
  assign n52607 = n52606 ^ n35073 ^ n7997 ;
  assign n52608 = ( ~n13449 & n19519 ) | ( ~n13449 & n38577 ) | ( n19519 & n38577 ) ;
  assign n52609 = ( n10167 & n17347 ) | ( n10167 & n24657 ) | ( n17347 & n24657 ) ;
  assign n52610 = ( n3246 & n48620 ) | ( n3246 & n52609 ) | ( n48620 & n52609 ) ;
  assign n52611 = n38589 ^ n21324 ^ n10509 ;
  assign n52612 = ( ~n10294 & n52610 ) | ( ~n10294 & n52611 ) | ( n52610 & n52611 ) ;
  assign n52613 = n18066 ^ n4053 ^ n2606 ;
  assign n52615 = ( n14768 & n23032 ) | ( n14768 & n28983 ) | ( n23032 & n28983 ) ;
  assign n52614 = ( n14537 & n38358 ) | ( n14537 & n49864 ) | ( n38358 & n49864 ) ;
  assign n52616 = n52615 ^ n52614 ^ n9817 ;
  assign n52617 = ( ~n38428 & n40419 ) | ( ~n38428 & n52616 ) | ( n40419 & n52616 ) ;
  assign n52618 = ( n4134 & ~n42502 ) | ( n4134 & n48704 ) | ( ~n42502 & n48704 ) ;
  assign n52619 = n36170 ^ n33358 ^ n10711 ;
  assign n52620 = n43660 ^ n14158 ^ n1503 ;
  assign n52621 = n9283 & n31497 ;
  assign n52622 = n52620 & n52621 ;
  assign n52623 = ( n15100 & n52619 ) | ( n15100 & ~n52622 ) | ( n52619 & ~n52622 ) ;
  assign n52624 = ( ~x55 & n2054 ) | ( ~x55 & n20901 ) | ( n2054 & n20901 ) ;
  assign n52625 = ( n5396 & n24507 ) | ( n5396 & n52624 ) | ( n24507 & n52624 ) ;
  assign n52626 = n51729 ^ n4598 ^ 1'b0 ;
  assign n52627 = ~n52625 & n52626 ;
  assign n52628 = n19513 ^ n14635 ^ n8678 ;
  assign n52629 = n52628 ^ n20050 ^ x195 ;
  assign n52630 = n16669 & ~n26249 ;
  assign n52631 = ( ~n3194 & n47637 ) | ( ~n3194 & n52630 ) | ( n47637 & n52630 ) ;
  assign n52632 = n43670 ^ n39533 ^ 1'b0 ;
  assign n52633 = n2982 & ~n15279 ;
  assign n52634 = ~n37613 & n52633 ;
  assign n52635 = n52634 ^ n10869 ^ x52 ;
  assign n52636 = n17240 & n33901 ;
  assign n52637 = ~n6703 & n52636 ;
  assign n52638 = ( n4728 & n17990 ) | ( n4728 & n52637 ) | ( n17990 & n52637 ) ;
  assign n52640 = n19264 ^ n12828 ^ n8499 ;
  assign n52641 = ( n37629 & n48885 ) | ( n37629 & n52640 ) | ( n48885 & n52640 ) ;
  assign n52639 = ( ~n18713 & n26003 ) | ( ~n18713 & n43140 ) | ( n26003 & n43140 ) ;
  assign n52642 = n52641 ^ n52639 ^ n5876 ;
  assign n52643 = ( n10606 & ~n12378 ) | ( n10606 & n28279 ) | ( ~n12378 & n28279 ) ;
  assign n52644 = ( ~n4085 & n27050 ) | ( ~n4085 & n47655 ) | ( n27050 & n47655 ) ;
  assign n52645 = n52644 ^ n42230 ^ n34081 ;
  assign n52646 = ( ~n3013 & n12170 ) | ( ~n3013 & n37583 ) | ( n12170 & n37583 ) ;
  assign n52647 = n52646 ^ n44576 ^ n17973 ;
  assign n52648 = ( ~n14787 & n33847 ) | ( ~n14787 & n52647 ) | ( n33847 & n52647 ) ;
  assign n52649 = ( n13884 & ~n14726 ) | ( n13884 & n21782 ) | ( ~n14726 & n21782 ) ;
  assign n52650 = n52649 ^ n41488 ^ n6832 ;
  assign n52651 = n40976 & n52650 ;
  assign n52652 = n52651 ^ n1414 ^ 1'b0 ;
  assign n52653 = n827 & n45574 ;
  assign n52654 = ( ~n4889 & n17932 ) | ( ~n4889 & n25410 ) | ( n17932 & n25410 ) ;
  assign n52655 = ( n7281 & n9617 ) | ( n7281 & ~n52654 ) | ( n9617 & ~n52654 ) ;
  assign n52656 = ( ~n21062 & n52653 ) | ( ~n21062 & n52655 ) | ( n52653 & n52655 ) ;
  assign n52657 = n41816 ^ n28302 ^ 1'b0 ;
  assign n52658 = n611 & n52657 ;
  assign n52659 = ( n449 & n10430 ) | ( n449 & n52658 ) | ( n10430 & n52658 ) ;
  assign n52660 = ( n15747 & n32583 ) | ( n15747 & ~n52659 ) | ( n32583 & ~n52659 ) ;
  assign n52661 = n1447 | n43180 ;
  assign n52662 = n27895 & ~n52661 ;
  assign n52663 = n52662 ^ n37994 ^ n13802 ;
  assign n52664 = n26448 ^ n14403 ^ n8254 ;
  assign n52665 = n52664 ^ n11624 ^ n729 ;
  assign n52666 = n52665 ^ n16249 ^ n2713 ;
  assign n52667 = n31060 ^ x215 ^ 1'b0 ;
  assign n52668 = ( n34728 & ~n34844 ) | ( n34728 & n52667 ) | ( ~n34844 & n52667 ) ;
  assign n52669 = ( n299 & n4614 ) | ( n299 & n7691 ) | ( n4614 & n7691 ) ;
  assign n52670 = ( ~n2007 & n37591 ) | ( ~n2007 & n52669 ) | ( n37591 & n52669 ) ;
  assign n52671 = ( n906 & ~n12235 ) | ( n906 & n24864 ) | ( ~n12235 & n24864 ) ;
  assign n52672 = ( ~n18908 & n30600 ) | ( ~n18908 & n52671 ) | ( n30600 & n52671 ) ;
  assign n52673 = n21140 ^ n14891 ^ n8835 ;
  assign n52674 = n52673 ^ n33160 ^ n21042 ;
  assign n52675 = n11852 & ~n18574 ;
  assign n52676 = ~n12792 & n52675 ;
  assign n52677 = ~n17205 & n45086 ;
  assign n52678 = ~n11090 & n52677 ;
  assign n52679 = n28202 ^ n18450 ^ n609 ;
  assign n52680 = n52679 ^ n43117 ^ n38209 ;
  assign n52681 = n29778 ^ n28415 ^ n18682 ;
  assign n52682 = n3514 & ~n20268 ;
  assign n52683 = ( n19060 & ~n30345 ) | ( n19060 & n40820 ) | ( ~n30345 & n40820 ) ;
  assign n52684 = n52683 ^ n50605 ^ n7574 ;
  assign n52685 = ~n24347 & n37104 ;
  assign n52689 = ( n1680 & ~n10277 ) | ( n1680 & n25317 ) | ( ~n10277 & n25317 ) ;
  assign n52686 = ( ~n3184 & n12192 ) | ( ~n3184 & n17402 ) | ( n12192 & n17402 ) ;
  assign n52687 = n52686 ^ n18498 ^ n9980 ;
  assign n52688 = ( n6509 & n19600 ) | ( n6509 & n52687 ) | ( n19600 & n52687 ) ;
  assign n52690 = n52689 ^ n52688 ^ x219 ;
  assign n52691 = ( n11937 & n20900 ) | ( n11937 & n44143 ) | ( n20900 & n44143 ) ;
  assign n52692 = n52691 ^ n22814 ^ n5813 ;
  assign n52693 = ( n17118 & n22018 ) | ( n17118 & ~n30918 ) | ( n22018 & ~n30918 ) ;
  assign n52694 = ( n19844 & n20180 ) | ( n19844 & n52693 ) | ( n20180 & n52693 ) ;
  assign n52695 = ( ~n6858 & n11899 ) | ( ~n6858 & n52694 ) | ( n11899 & n52694 ) ;
  assign n52696 = n7607 & n36395 ;
  assign n52697 = n52696 ^ n33604 ^ n26101 ;
  assign n52698 = ( n1877 & n28354 ) | ( n1877 & ~n31341 ) | ( n28354 & ~n31341 ) ;
  assign n52699 = ~n6000 & n52698 ;
  assign n52700 = n52699 ^ n18875 ^ 1'b0 ;
  assign n52701 = ( n11808 & n15806 ) | ( n11808 & ~n52700 ) | ( n15806 & ~n52700 ) ;
  assign n52702 = n52701 ^ n12175 ^ 1'b0 ;
  assign n52703 = n22550 & ~n52702 ;
  assign n52705 = n8325 ^ n4673 ^ n1002 ;
  assign n52704 = n27767 ^ n8849 ^ 1'b0 ;
  assign n52706 = n52705 ^ n52704 ^ n5733 ;
  assign n52707 = n25012 & ~n32233 ;
  assign n52708 = ~n52706 & n52707 ;
  assign n52709 = n31113 ^ n26794 ^ n21698 ;
  assign n52710 = n7894 & n12348 ;
  assign n52711 = ~n5725 & n52710 ;
  assign n52712 = n32916 | n52711 ;
  assign n52713 = n46849 | n52712 ;
  assign n52714 = ( n8598 & n51422 ) | ( n8598 & ~n52713 ) | ( n51422 & ~n52713 ) ;
  assign n52715 = ( ~n3569 & n51937 ) | ( ~n3569 & n52714 ) | ( n51937 & n52714 ) ;
  assign n52716 = ( n13157 & n22435 ) | ( n13157 & n48063 ) | ( n22435 & n48063 ) ;
  assign n52717 = ( x98 & n293 ) | ( x98 & n8552 ) | ( n293 & n8552 ) ;
  assign n52718 = ( n19848 & n35609 ) | ( n19848 & ~n38539 ) | ( n35609 & ~n38539 ) ;
  assign n52719 = ( n18224 & ~n24180 ) | ( n18224 & n33717 ) | ( ~n24180 & n33717 ) ;
  assign n52720 = ( ~n12830 & n34997 ) | ( ~n12830 & n52719 ) | ( n34997 & n52719 ) ;
  assign n52721 = n22896 ^ n20330 ^ n9081 ;
  assign n52722 = n14822 | n16243 ;
  assign n52723 = ( ~n8980 & n15627 ) | ( ~n8980 & n23497 ) | ( n15627 & n23497 ) ;
  assign n52724 = n2857 & n52723 ;
  assign n52725 = n33983 & n52724 ;
  assign n52726 = n23761 ^ n1617 ^ 1'b0 ;
  assign n52727 = n29488 ^ n27599 ^ n18444 ;
  assign n52728 = ( n32426 & ~n34810 ) | ( n32426 & n52727 ) | ( ~n34810 & n52727 ) ;
  assign n52729 = n35329 | n52728 ;
  assign n52730 = ( ~n3759 & n8219 ) | ( ~n3759 & n51316 ) | ( n8219 & n51316 ) ;
  assign n52731 = n37757 ^ n22649 ^ n15963 ;
  assign n52734 = n9638 & ~n36827 ;
  assign n52735 = n18243 | n45481 ;
  assign n52736 = n52735 ^ n24820 ^ 1'b0 ;
  assign n52737 = ( n11070 & n52734 ) | ( n11070 & ~n52736 ) | ( n52734 & ~n52736 ) ;
  assign n52732 = ( n14410 & n15007 ) | ( n14410 & ~n43023 ) | ( n15007 & ~n43023 ) ;
  assign n52733 = ( ~n32055 & n47668 ) | ( ~n32055 & n52732 ) | ( n47668 & n52732 ) ;
  assign n52738 = n52737 ^ n52733 ^ n897 ;
  assign n52739 = ( n21608 & n39549 ) | ( n21608 & n45854 ) | ( n39549 & n45854 ) ;
  assign n52740 = n13578 | n49741 ;
  assign n52741 = n43788 ^ n23108 ^ n11863 ;
  assign n52742 = n52577 ^ n20700 ^ n12462 ;
  assign n52747 = n5047 | n9138 ;
  assign n52744 = n13919 ^ n5214 ^ n2811 ;
  assign n52745 = ( ~n34029 & n37533 ) | ( ~n34029 & n52744 ) | ( n37533 & n52744 ) ;
  assign n52746 = ( n20069 & ~n28636 ) | ( n20069 & n52745 ) | ( ~n28636 & n52745 ) ;
  assign n52743 = ( n4570 & ~n36040 ) | ( n4570 & n45569 ) | ( ~n36040 & n45569 ) ;
  assign n52748 = n52747 ^ n52746 ^ n52743 ;
  assign n52749 = n20826 | n48899 ;
  assign n52750 = n39685 & ~n52749 ;
  assign n52751 = n31931 | n52750 ;
  assign n52752 = n52751 ^ n31834 ^ 1'b0 ;
  assign n52753 = n42337 ^ n30547 ^ n4043 ;
  assign n52754 = n32049 | n33236 ;
  assign n52755 = n13347 & ~n52754 ;
  assign n52756 = ( n21067 & ~n33743 ) | ( n21067 & n52755 ) | ( ~n33743 & n52755 ) ;
  assign n52757 = ( n773 & n37241 ) | ( n773 & ~n52756 ) | ( n37241 & ~n52756 ) ;
  assign n52758 = n45100 ^ n36894 ^ n12003 ;
  assign n52759 = n31293 ^ n26991 ^ n6072 ;
  assign n52760 = n31923 ^ n26984 ^ n6254 ;
  assign n52761 = n37753 ^ n30400 ^ 1'b0 ;
  assign n52762 = ( ~n6496 & n13259 ) | ( ~n6496 & n35272 ) | ( n13259 & n35272 ) ;
  assign n52763 = ( n35100 & n38298 ) | ( n35100 & ~n44911 ) | ( n38298 & ~n44911 ) ;
  assign n52765 = n10101 ^ n7869 ^ 1'b0 ;
  assign n52766 = n13134 | n52765 ;
  assign n52764 = n7296 | n36389 ;
  assign n52767 = n52766 ^ n52764 ^ n13370 ;
  assign n52768 = n8326 & ~n51335 ;
  assign n52769 = n52768 ^ n15056 ^ 1'b0 ;
  assign n52770 = ~n6576 & n52769 ;
  assign n52771 = ~n466 & n49231 ;
  assign n52772 = ~n52770 & n52771 ;
  assign n52773 = n7446 | n11795 ;
  assign n52774 = n29344 & ~n52773 ;
  assign n52775 = n12268 | n16545 ;
  assign n52776 = n52775 ^ n41791 ^ n11211 ;
  assign n52782 = n33255 ^ n15447 ^ n6473 ;
  assign n52777 = n22681 ^ n10094 ^ n987 ;
  assign n52778 = ( n15848 & n38916 ) | ( n15848 & n52777 ) | ( n38916 & n52777 ) ;
  assign n52779 = n27080 ^ n6457 ^ 1'b0 ;
  assign n52780 = ( n7253 & ~n39611 ) | ( n7253 & n52779 ) | ( ~n39611 & n52779 ) ;
  assign n52781 = n52778 | n52780 ;
  assign n52783 = n52782 ^ n52781 ^ n6827 ;
  assign n52784 = n17163 & n35735 ;
  assign n52785 = ( n11664 & ~n19541 ) | ( n11664 & n52098 ) | ( ~n19541 & n52098 ) ;
  assign n52786 = n24355 ^ n8311 ^ n6428 ;
  assign n52787 = n52786 ^ n23468 ^ n5290 ;
  assign n52788 = ( ~n4055 & n36498 ) | ( ~n4055 & n52787 ) | ( n36498 & n52787 ) ;
  assign n52789 = ( n602 & ~n8270 ) | ( n602 & n52788 ) | ( ~n8270 & n52788 ) ;
  assign n52790 = ( n8374 & n18659 ) | ( n8374 & n20215 ) | ( n18659 & n20215 ) ;
  assign n52791 = n33550 ^ n33064 ^ 1'b0 ;
  assign n52792 = n52791 ^ n45814 ^ n23982 ;
  assign n52793 = n35789 & ~n37528 ;
  assign n52794 = ~n3938 & n37924 ;
  assign n52795 = ( n2562 & n31534 ) | ( n2562 & ~n52794 ) | ( n31534 & ~n52794 ) ;
  assign n52796 = n1654 | n11651 ;
  assign n52797 = n1678 | n52796 ;
  assign n52798 = ( ~n2001 & n12188 ) | ( ~n2001 & n18588 ) | ( n12188 & n18588 ) ;
  assign n52799 = n52798 ^ n34472 ^ 1'b0 ;
  assign n52800 = n45150 & ~n52799 ;
  assign n52801 = ( n11009 & ~n12090 ) | ( n11009 & n15252 ) | ( ~n12090 & n15252 ) ;
  assign n52802 = n26935 | n52801 ;
  assign n52803 = n52802 ^ n50569 ^ n27595 ;
  assign n52804 = ( n912 & ~n13522 ) | ( n912 & n19672 ) | ( ~n13522 & n19672 ) ;
  assign n52805 = n1396 | n36937 ;
  assign n52806 = ( ~n6238 & n14268 ) | ( ~n6238 & n46503 ) | ( n14268 & n46503 ) ;
  assign n52807 = ( n2219 & ~n52805 ) | ( n2219 & n52806 ) | ( ~n52805 & n52806 ) ;
  assign n52808 = ( n18023 & ~n25637 ) | ( n18023 & n42159 ) | ( ~n25637 & n42159 ) ;
  assign n52809 = n8085 & n52808 ;
  assign n52810 = n17357 & n52809 ;
  assign n52811 = ( n20913 & n34659 ) | ( n20913 & ~n52810 ) | ( n34659 & ~n52810 ) ;
  assign n52812 = n52811 ^ n48232 ^ n31657 ;
  assign n52813 = ( n13354 & n25113 ) | ( n13354 & ~n45359 ) | ( n25113 & ~n45359 ) ;
  assign n52814 = ~n11074 & n21035 ;
  assign n52815 = ( n7430 & n8964 ) | ( n7430 & ~n41099 ) | ( n8964 & ~n41099 ) ;
  assign n52816 = n13222 ^ n2200 ^ 1'b0 ;
  assign n52817 = n52816 ^ n1205 ^ n720 ;
  assign n52818 = n52817 ^ n7126 ^ n5315 ;
  assign n52819 = n28764 & n31137 ;
  assign n52820 = n52819 ^ n48875 ^ 1'b0 ;
  assign n52821 = n11499 ^ n2653 ^ 1'b0 ;
  assign n52822 = n25017 | n52821 ;
  assign n52823 = ( n2498 & n20819 ) | ( n2498 & n39900 ) | ( n20819 & n39900 ) ;
  assign n52824 = ( n8585 & n25455 ) | ( n8585 & ~n52823 ) | ( n25455 & ~n52823 ) ;
  assign n52825 = ( n995 & ~n31658 ) | ( n995 & n47309 ) | ( ~n31658 & n47309 ) ;
  assign n52826 = ( ~x171 & n39491 ) | ( ~x171 & n52825 ) | ( n39491 & n52825 ) ;
  assign n52827 = ( ~n13682 & n52824 ) | ( ~n13682 & n52826 ) | ( n52824 & n52826 ) ;
  assign n52828 = ( n11926 & ~n18563 ) | ( n11926 & n45457 ) | ( ~n18563 & n45457 ) ;
  assign n52829 = n7736 ^ n7720 ^ n1495 ;
  assign n52830 = ( n37028 & n50508 ) | ( n37028 & ~n52829 ) | ( n50508 & ~n52829 ) ;
  assign n52832 = ( n1845 & n2603 ) | ( n1845 & n13627 ) | ( n2603 & n13627 ) ;
  assign n52831 = ( n13906 & n16302 ) | ( n13906 & ~n33592 ) | ( n16302 & ~n33592 ) ;
  assign n52833 = n52832 ^ n52831 ^ n36909 ;
  assign n52834 = n52833 ^ n43354 ^ n10429 ;
  assign n52835 = ( n15834 & n21910 ) | ( n15834 & ~n41364 ) | ( n21910 & ~n41364 ) ;
  assign n52836 = n7373 ^ n2783 ^ n1810 ;
  assign n52837 = n52836 ^ n15452 ^ n12384 ;
  assign n52838 = ( n25448 & n50956 ) | ( n25448 & n52837 ) | ( n50956 & n52837 ) ;
  assign n52842 = n14489 ^ n3090 ^ 1'b0 ;
  assign n52841 = ( n19864 & n32139 ) | ( n19864 & n44202 ) | ( n32139 & n44202 ) ;
  assign n52843 = n52842 ^ n52841 ^ n37850 ;
  assign n52839 = ( n3346 & ~n18983 ) | ( n3346 & n33940 ) | ( ~n18983 & n33940 ) ;
  assign n52840 = n52839 ^ n49439 ^ n42872 ;
  assign n52844 = n52843 ^ n52840 ^ n41292 ;
  assign n52845 = n20340 ^ n16085 ^ 1'b0 ;
  assign n52846 = ~n2378 & n52845 ;
  assign n52847 = n52846 ^ n34972 ^ n16702 ;
  assign n52848 = n28574 & n52847 ;
  assign n52849 = n16193 | n52848 ;
  assign n52850 = n52849 ^ n21463 ^ n18764 ;
  assign n52851 = n24275 ^ n14734 ^ n3954 ;
  assign n52852 = ( n17992 & n29988 ) | ( n17992 & ~n52851 ) | ( n29988 & ~n52851 ) ;
  assign n52853 = n1681 & ~n4950 ;
  assign n52854 = n566 & n52853 ;
  assign n52855 = n393 & ~n10359 ;
  assign n52856 = n52855 ^ n7879 ^ 1'b0 ;
  assign n52857 = n49749 ^ n45400 ^ n36313 ;
  assign n52858 = n52857 ^ n42768 ^ n11071 ;
  assign n52859 = n35792 ^ n1387 ^ 1'b0 ;
  assign n52860 = n52859 ^ n35701 ^ n11719 ;
  assign n52861 = n35230 ^ n3333 ^ n3223 ;
  assign n52862 = ( n20576 & n46726 ) | ( n20576 & n52861 ) | ( n46726 & n52861 ) ;
  assign n52863 = n47698 ^ n47464 ^ n30286 ;
  assign n52864 = ( n2677 & n17425 ) | ( n2677 & n33861 ) | ( n17425 & n33861 ) ;
  assign n52865 = n14331 ^ n6760 ^ 1'b0 ;
  assign n52866 = n24826 ^ n15847 ^ n8527 ;
  assign n52867 = n31791 & n39206 ;
  assign n52868 = ( n19130 & n52866 ) | ( n19130 & ~n52867 ) | ( n52866 & ~n52867 ) ;
  assign n52869 = n52416 ^ n39048 ^ n20618 ;
  assign n52870 = n52869 ^ n26050 ^ n20028 ;
  assign n52871 = ( x42 & ~n43000 ) | ( x42 & n43051 ) | ( ~n43000 & n43051 ) ;
  assign n52873 = n28646 ^ n3286 ^ 1'b0 ;
  assign n52874 = n21981 | n52873 ;
  assign n52872 = n825 & ~n14834 ;
  assign n52875 = n52874 ^ n52872 ^ 1'b0 ;
  assign n52878 = ( n1301 & ~n35335 ) | ( n1301 & n39460 ) | ( ~n35335 & n39460 ) ;
  assign n52876 = ~n10421 & n17369 ;
  assign n52877 = ~n30450 & n52876 ;
  assign n52879 = n52878 ^ n52877 ^ 1'b0 ;
  assign n52880 = n48809 ^ n768 ^ 1'b0 ;
  assign n52881 = n35954 & n52880 ;
  assign n52882 = n52881 ^ n33926 ^ n8163 ;
  assign n52883 = n48750 ^ n20665 ^ n16446 ;
  assign n52884 = n52883 ^ n39814 ^ n38120 ;
  assign n52885 = ~n16058 & n39829 ;
  assign n52886 = ( n1704 & n52628 ) | ( n1704 & ~n52885 ) | ( n52628 & ~n52885 ) ;
  assign n52887 = n8428 ^ n8199 ^ n6895 ;
  assign n52888 = n27484 ^ n7748 ^ 1'b0 ;
  assign n52889 = ( x103 & n5475 ) | ( x103 & n45444 ) | ( n5475 & n45444 ) ;
  assign n52890 = ( ~n4085 & n52888 ) | ( ~n4085 & n52889 ) | ( n52888 & n52889 ) ;
  assign n52891 = ( ~n22464 & n52887 ) | ( ~n22464 & n52890 ) | ( n52887 & n52890 ) ;
  assign n52892 = ( n5167 & n10865 ) | ( n5167 & ~n52891 ) | ( n10865 & ~n52891 ) ;
  assign n52893 = n52892 ^ n18434 ^ n9652 ;
  assign n52894 = ( n5853 & n10067 ) | ( n5853 & ~n30996 ) | ( n10067 & ~n30996 ) ;
  assign n52895 = ( n8969 & n34523 ) | ( n8969 & n52894 ) | ( n34523 & n52894 ) ;
  assign n52896 = n52895 ^ n29558 ^ n10300 ;
  assign n52897 = n46847 ^ n42802 ^ n42059 ;
  assign n52898 = n23651 ^ n15038 ^ n8666 ;
  assign n52899 = n52898 ^ n28882 ^ n19857 ;
  assign n52900 = ( n5774 & n19273 ) | ( n5774 & ~n24783 ) | ( n19273 & ~n24783 ) ;
  assign n52901 = n49732 ^ n31609 ^ n9533 ;
  assign n52902 = ( ~n22485 & n50724 ) | ( ~n22485 & n52901 ) | ( n50724 & n52901 ) ;
  assign n52903 = n22938 | n26925 ;
  assign n52904 = n4521 & ~n52903 ;
  assign n52905 = n31491 & n31927 ;
  assign n52906 = n52905 ^ n28999 ^ 1'b0 ;
  assign n52907 = n1601 & n52906 ;
  assign n52910 = n4210 ^ n1240 ^ 1'b0 ;
  assign n52911 = n286 & n52910 ;
  assign n52912 = ( ~n11239 & n24500 ) | ( ~n11239 & n52911 ) | ( n24500 & n52911 ) ;
  assign n52913 = ( n18589 & n18826 ) | ( n18589 & ~n52912 ) | ( n18826 & ~n52912 ) ;
  assign n52908 = n1085 & n38390 ;
  assign n52909 = ~n1573 & n52908 ;
  assign n52914 = n52913 ^ n52909 ^ 1'b0 ;
  assign n52915 = ( n17424 & ~n34755 ) | ( n17424 & n52914 ) | ( ~n34755 & n52914 ) ;
  assign n52916 = n17355 ^ n7465 ^ n747 ;
  assign n52917 = n52916 ^ n40607 ^ n32944 ;
  assign n52918 = n23002 ^ n16161 ^ n2853 ;
  assign n52919 = n52918 ^ n16857 ^ n6227 ;
  assign n52920 = ( n14627 & n19137 ) | ( n14627 & ~n44936 ) | ( n19137 & ~n44936 ) ;
  assign n52921 = n17350 ^ n10745 ^ n6857 ;
  assign n52922 = n52921 ^ n32575 ^ n6958 ;
  assign n52923 = ( n3180 & n44857 ) | ( n3180 & n52922 ) | ( n44857 & n52922 ) ;
  assign n52924 = n4435 | n32433 ;
  assign n52925 = n52924 ^ n32038 ^ 1'b0 ;
  assign n52926 = ( n6885 & ~n42130 ) | ( n6885 & n52925 ) | ( ~n42130 & n52925 ) ;
  assign n52927 = n28180 | n46910 ;
  assign n52928 = n11929 | n52927 ;
  assign n52929 = n52928 ^ n22766 ^ 1'b0 ;
  assign n52931 = ( n10024 & ~n38270 ) | ( n10024 & n39623 ) | ( ~n38270 & n39623 ) ;
  assign n52930 = ( n2370 & n33783 ) | ( n2370 & ~n44706 ) | ( n33783 & ~n44706 ) ;
  assign n52932 = n52931 ^ n52930 ^ n8582 ;
  assign n52933 = n29395 ^ n1352 ^ 1'b0 ;
  assign n52934 = ( ~n6831 & n18306 ) | ( ~n6831 & n31213 ) | ( n18306 & n31213 ) ;
  assign n52935 = n52934 ^ n37916 ^ n23998 ;
  assign n52936 = ~n26147 & n41436 ;
  assign n52937 = ~n15269 & n52936 ;
  assign n52938 = n52937 ^ n21943 ^ n12523 ;
  assign n52939 = ( ~n3465 & n11829 ) | ( ~n3465 & n24919 ) | ( n11829 & n24919 ) ;
  assign n52940 = ( n27239 & n51127 ) | ( n27239 & n52939 ) | ( n51127 & n52939 ) ;
  assign n52941 = ~n10152 & n52940 ;
  assign n52942 = ( ~n27785 & n29985 ) | ( ~n27785 & n30253 ) | ( n29985 & n30253 ) ;
  assign n52943 = ( n26679 & n27757 ) | ( n26679 & ~n52942 ) | ( n27757 & ~n52942 ) ;
  assign n52944 = n5705 & ~n5764 ;
  assign n52945 = n6132 | n17262 ;
  assign n52946 = ( n8102 & ~n10935 ) | ( n8102 & n52945 ) | ( ~n10935 & n52945 ) ;
  assign n52947 = n52946 ^ n49409 ^ n44322 ;
  assign n52948 = n52947 ^ n14960 ^ n6715 ;
  assign n52949 = ( n1254 & ~n10735 ) | ( n1254 & n33042 ) | ( ~n10735 & n33042 ) ;
  assign n52950 = n52949 ^ n15810 ^ n11113 ;
  assign n52951 = n30804 ^ n13852 ^ n13218 ;
  assign n52952 = n10189 ^ n6934 ^ n6823 ;
  assign n52953 = n22852 ^ n18765 ^ 1'b0 ;
  assign n52954 = n34011 & ~n52953 ;
  assign n52955 = ( ~n12662 & n31229 ) | ( ~n12662 & n43382 ) | ( n31229 & n43382 ) ;
  assign n52956 = ( ~n11081 & n19626 ) | ( ~n11081 & n49704 ) | ( n19626 & n49704 ) ;
  assign n52957 = n52956 ^ n29326 ^ 1'b0 ;
  assign n52958 = ( n30296 & n39500 ) | ( n30296 & n40695 ) | ( n39500 & n40695 ) ;
  assign n52959 = n52958 ^ n19093 ^ n16907 ;
  assign n52960 = ( n496 & n49755 ) | ( n496 & ~n52959 ) | ( n49755 & ~n52959 ) ;
  assign n52961 = ( ~n32971 & n40603 ) | ( ~n32971 & n47208 ) | ( n40603 & n47208 ) ;
  assign n52962 = ( n4020 & n12121 ) | ( n4020 & n27751 ) | ( n12121 & n27751 ) ;
  assign n52963 = ( n48128 & n50130 ) | ( n48128 & ~n52962 ) | ( n50130 & ~n52962 ) ;
  assign n52964 = ( n3770 & n24123 ) | ( n3770 & ~n38860 ) | ( n24123 & ~n38860 ) ;
  assign n52965 = ( n7397 & ~n13572 ) | ( n7397 & n34845 ) | ( ~n13572 & n34845 ) ;
  assign n52966 = ( n3130 & n32476 ) | ( n3130 & n52965 ) | ( n32476 & n52965 ) ;
  assign n52967 = ( n10367 & n23223 ) | ( n10367 & ~n30797 ) | ( n23223 & ~n30797 ) ;
  assign n52968 = n5923 & n9454 ;
  assign n52969 = ( n24450 & n49987 ) | ( n24450 & n52968 ) | ( n49987 & n52968 ) ;
  assign n52970 = ( n6668 & ~n39591 ) | ( n6668 & n52969 ) | ( ~n39591 & n52969 ) ;
  assign n52971 = n7872 | n52970 ;
  assign n52972 = n25348 ^ n20800 ^ 1'b0 ;
  assign n52973 = ~n24853 & n52972 ;
  assign n52974 = ( n6453 & n18299 ) | ( n6453 & ~n33821 ) | ( n18299 & ~n33821 ) ;
  assign n52975 = n52974 ^ n18837 ^ n3844 ;
  assign n52976 = n52975 ^ n31820 ^ n4823 ;
  assign n52977 = ( n10502 & n11263 ) | ( n10502 & ~n14158 ) | ( n11263 & ~n14158 ) ;
  assign n52978 = n11899 ^ n9517 ^ n2091 ;
  assign n52979 = ( n8584 & n34903 ) | ( n8584 & n52978 ) | ( n34903 & n52978 ) ;
  assign n52980 = ( ~n3287 & n15317 ) | ( ~n3287 & n47627 ) | ( n15317 & n47627 ) ;
  assign n52981 = n52980 ^ n34943 ^ n31289 ;
  assign n52982 = n30713 ^ n22005 ^ n1749 ;
  assign n52983 = n27701 ^ n26428 ^ n25496 ;
  assign n52984 = n31866 ^ n15050 ^ 1'b0 ;
  assign n52985 = ( n5886 & ~n20913 ) | ( n5886 & n52984 ) | ( ~n20913 & n52984 ) ;
  assign n52989 = n31280 ^ n24473 ^ n23367 ;
  assign n52990 = n52989 ^ n19247 ^ n14722 ;
  assign n52986 = ~n15345 & n32606 ;
  assign n52987 = ( n13469 & n14238 ) | ( n13469 & ~n52986 ) | ( n14238 & ~n52986 ) ;
  assign n52988 = n52987 ^ n49358 ^ n20152 ;
  assign n52991 = n52990 ^ n52988 ^ n24156 ;
  assign n52992 = ( ~n21195 & n35084 ) | ( ~n21195 & n52991 ) | ( n35084 & n52991 ) ;
  assign n52993 = n47483 ^ n39593 ^ n36004 ;
  assign n52994 = n3159 & ~n23603 ;
  assign n52995 = n3253 & n39638 ;
  assign n52996 = n9523 & n52995 ;
  assign n53000 = n29051 ^ n3357 ^ n2157 ;
  assign n52997 = n43137 ^ n32718 ^ 1'b0 ;
  assign n52998 = ~n37824 & n52997 ;
  assign n52999 = n52998 ^ n46402 ^ 1'b0 ;
  assign n53001 = n53000 ^ n52999 ^ n50171 ;
  assign n53002 = ( n22682 & n36340 ) | ( n22682 & n40707 ) | ( n36340 & n40707 ) ;
  assign n53003 = n53002 ^ n18782 ^ n12396 ;
  assign n53004 = n51894 ^ n40500 ^ n29169 ;
  assign n53005 = n47865 ^ n46953 ^ n26939 ;
  assign n53006 = ( n5476 & n35455 ) | ( n5476 & ~n53005 ) | ( n35455 & ~n53005 ) ;
  assign n53007 = n45430 ^ n31034 ^ n12344 ;
  assign n53008 = n43746 ^ n36376 ^ n25458 ;
  assign n53009 = n28569 ^ n10277 ^ 1'b0 ;
  assign n53010 = n52005 ^ n22320 ^ 1'b0 ;
  assign n53011 = n29928 & n49723 ;
  assign n53012 = n15209 | n34045 ;
  assign n53013 = n53012 ^ n33107 ^ 1'b0 ;
  assign n53014 = n33587 ^ n12975 ^ n5725 ;
  assign n53015 = n1868 | n24843 ;
  assign n53016 = n53014 & ~n53015 ;
  assign n53017 = n18660 ^ n16589 ^ n8500 ;
  assign n53018 = n35065 ^ n31198 ^ n8632 ;
  assign n53019 = ( n18498 & n21416 ) | ( n18498 & n53018 ) | ( n21416 & n53018 ) ;
  assign n53020 = n15533 & n39095 ;
  assign n53021 = n7484 & n53020 ;
  assign n53022 = n53021 ^ n11473 ^ n8168 ;
  assign n53023 = n53022 ^ n52598 ^ n29737 ;
  assign n53024 = n52067 ^ n38385 ^ n36170 ;
  assign n53025 = n53024 ^ n12086 ^ 1'b0 ;
  assign n53026 = n13622 ^ n8350 ^ 1'b0 ;
  assign n53027 = n53026 ^ n25318 ^ n6066 ;
  assign n53028 = ( n2799 & n6688 ) | ( n2799 & n53027 ) | ( n6688 & n53027 ) ;
  assign n53029 = n38099 ^ n24721 ^ n20728 ;
  assign n53030 = n53029 ^ n40186 ^ n10815 ;
  assign n53031 = n53030 ^ n42327 ^ n29374 ;
  assign n53032 = n37757 ^ n9496 ^ 1'b0 ;
  assign n53033 = ( n16808 & n21972 ) | ( n16808 & ~n53032 ) | ( n21972 & ~n53032 ) ;
  assign n53034 = ( ~n1250 & n8658 ) | ( ~n1250 & n35297 ) | ( n8658 & n35297 ) ;
  assign n53035 = ( n6053 & n30755 ) | ( n6053 & ~n53034 ) | ( n30755 & ~n53034 ) ;
  assign n53037 = n51290 ^ n3547 ^ n1904 ;
  assign n53036 = ( n44748 & n50686 ) | ( n44748 & ~n51417 ) | ( n50686 & ~n51417 ) ;
  assign n53038 = n53037 ^ n53036 ^ n12943 ;
  assign n53039 = ( x38 & n28595 ) | ( x38 & ~n49621 ) | ( n28595 & ~n49621 ) ;
  assign n53040 = n53039 ^ n41435 ^ n38447 ;
  assign n53041 = n19287 ^ n9069 ^ n4384 ;
  assign n53042 = n53041 ^ n29925 ^ n636 ;
  assign n53043 = ( n3381 & n12879 ) | ( n3381 & ~n53042 ) | ( n12879 & ~n53042 ) ;
  assign n53044 = n50405 ^ n49345 ^ n6386 ;
  assign n53049 = ( n2995 & n4344 ) | ( n2995 & n21168 ) | ( n4344 & n21168 ) ;
  assign n53045 = ( n2590 & n8564 ) | ( n2590 & ~n12047 ) | ( n8564 & ~n12047 ) ;
  assign n53046 = n6411 & ~n46428 ;
  assign n53047 = n53046 ^ x17 ^ 1'b0 ;
  assign n53048 = ( n3782 & ~n53045 ) | ( n3782 & n53047 ) | ( ~n53045 & n53047 ) ;
  assign n53050 = n53049 ^ n53048 ^ n10503 ;
  assign n53051 = ( n22262 & n53044 ) | ( n22262 & ~n53050 ) | ( n53044 & ~n53050 ) ;
  assign n53052 = n35097 ^ n20940 ^ n10094 ;
  assign n53053 = n20044 ^ n8325 ^ 1'b0 ;
  assign n53054 = n28882 | n49448 ;
  assign n53055 = n25105 & ~n53054 ;
  assign n53056 = ( n3858 & ~n29792 ) | ( n3858 & n34024 ) | ( ~n29792 & n34024 ) ;
  assign n53057 = ( n53053 & ~n53055 ) | ( n53053 & n53056 ) | ( ~n53055 & n53056 ) ;
  assign n53058 = ( n3903 & n39925 ) | ( n3903 & ~n42781 ) | ( n39925 & ~n42781 ) ;
  assign n53060 = n33750 ^ n32918 ^ n9484 ;
  assign n53059 = ( n18304 & n25217 ) | ( n18304 & n34149 ) | ( n25217 & n34149 ) ;
  assign n53061 = n53060 ^ n53059 ^ n52848 ;
  assign n53062 = n7634 & ~n26198 ;
  assign n53063 = n53062 ^ n49162 ^ 1'b0 ;
  assign n53064 = n23615 ^ n12440 ^ n9341 ;
  assign n53065 = n53064 ^ n1194 ^ 1'b0 ;
  assign n53066 = ( n18450 & n31430 ) | ( n18450 & n48520 ) | ( n31430 & n48520 ) ;
  assign n53067 = n35675 ^ n26940 ^ n18946 ;
  assign n53068 = n53067 ^ n22581 ^ n18158 ;
  assign n53069 = ( n37993 & n42899 ) | ( n37993 & ~n49278 ) | ( n42899 & ~n49278 ) ;
  assign n53070 = n53069 ^ n46902 ^ n14871 ;
  assign n53071 = ( n34875 & n39736 ) | ( n34875 & ~n45387 ) | ( n39736 & ~n45387 ) ;
  assign n53072 = ( ~n6512 & n40771 ) | ( ~n6512 & n53071 ) | ( n40771 & n53071 ) ;
  assign n53073 = n30383 ^ n2674 ^ 1'b0 ;
  assign n53074 = ( ~n11021 & n14478 ) | ( ~n11021 & n53073 ) | ( n14478 & n53073 ) ;
  assign n53075 = n2757 | n15729 ;
  assign n53076 = n3873 | n53075 ;
  assign n53077 = n5541 | n53076 ;
  assign n53078 = n53077 ^ n36384 ^ n34220 ;
  assign n53079 = n15656 ^ n4618 ^ 1'b0 ;
  assign n53080 = ~n24124 & n53079 ;
  assign n53081 = n53080 ^ n31075 ^ n2811 ;
  assign n53082 = ( n12857 & ~n14868 ) | ( n12857 & n16545 ) | ( ~n14868 & n16545 ) ;
  assign n53083 = n53082 ^ n19516 ^ n12553 ;
  assign n53084 = ( n1119 & n12031 ) | ( n1119 & ~n53083 ) | ( n12031 & ~n53083 ) ;
  assign n53085 = n53084 ^ n19053 ^ n14000 ;
  assign n53086 = n23755 ^ n15746 ^ 1'b0 ;
  assign n53087 = n53085 & n53086 ;
  assign n53088 = ( n10870 & ~n35372 ) | ( n10870 & n43071 ) | ( ~n35372 & n43071 ) ;
  assign n53089 = n38017 ^ n17588 ^ n12614 ;
  assign n53090 = n53089 ^ n49695 ^ n34095 ;
  assign n53091 = ( ~n10913 & n23417 ) | ( ~n10913 & n53090 ) | ( n23417 & n53090 ) ;
  assign n53092 = n38186 ^ n29121 ^ n26815 ;
  assign n53093 = ( ~n21740 & n35225 ) | ( ~n21740 & n44077 ) | ( n35225 & n44077 ) ;
  assign n53094 = ( n22881 & n26235 ) | ( n22881 & n53093 ) | ( n26235 & n53093 ) ;
  assign n53095 = n49315 ^ n28696 ^ n20467 ;
  assign n53096 = ( n18753 & n22051 ) | ( n18753 & n37097 ) | ( n22051 & n37097 ) ;
  assign n53097 = ( n750 & ~n53095 ) | ( n750 & n53096 ) | ( ~n53095 & n53096 ) ;
  assign n53098 = n51488 ^ n46199 ^ n32672 ;
  assign n53099 = n11786 & n48598 ;
  assign n53100 = n53099 ^ n42149 ^ 1'b0 ;
  assign n53101 = n4292 | n26935 ;
  assign n53102 = n45781 | n53101 ;
  assign n53103 = n2859 & n53102 ;
  assign n53104 = n53103 ^ n17722 ^ 1'b0 ;
  assign n53105 = n19262 | n43742 ;
  assign n53106 = n53105 ^ n44068 ^ 1'b0 ;
  assign n53107 = ( n9362 & n33718 ) | ( n9362 & n53106 ) | ( n33718 & n53106 ) ;
  assign n53108 = ( ~n3799 & n12037 ) | ( ~n3799 & n37770 ) | ( n12037 & n37770 ) ;
  assign n53109 = n53108 ^ n47904 ^ n37511 ;
  assign n53110 = n31691 ^ n9898 ^ 1'b0 ;
  assign n53111 = ~n5418 & n43677 ;
  assign n53112 = ~n41954 & n53111 ;
  assign n53113 = ( n3325 & n4352 ) | ( n3325 & ~n28084 ) | ( n4352 & ~n28084 ) ;
  assign n53114 = n53113 ^ n32985 ^ n4830 ;
  assign n53115 = n18143 & ~n38471 ;
  assign n53116 = ( ~n53112 & n53114 ) | ( ~n53112 & n53115 ) | ( n53114 & n53115 ) ;
  assign n53117 = n29654 ^ n26696 ^ n6332 ;
  assign n53118 = n28376 & ~n52596 ;
  assign n53119 = n33829 & n53118 ;
  assign n53120 = ( ~n51785 & n53117 ) | ( ~n51785 & n53119 ) | ( n53117 & n53119 ) ;
  assign n53121 = n46914 ^ n38234 ^ n5550 ;
  assign n53122 = n53121 ^ n17867 ^ n280 ;
  assign n53123 = n1143 & ~n16164 ;
  assign n53124 = ( n2100 & n23287 ) | ( n2100 & n53123 ) | ( n23287 & n53123 ) ;
  assign n53125 = n49315 ^ n22904 ^ n18980 ;
  assign n53126 = n53125 ^ n37462 ^ n6540 ;
  assign n53127 = ( n30509 & ~n53124 ) | ( n30509 & n53126 ) | ( ~n53124 & n53126 ) ;
  assign n53129 = ( n14884 & n15464 ) | ( n14884 & n26959 ) | ( n15464 & n26959 ) ;
  assign n53128 = ( n19140 & ~n23291 ) | ( n19140 & n44562 ) | ( ~n23291 & n44562 ) ;
  assign n53130 = n53129 ^ n53128 ^ 1'b0 ;
  assign n53131 = n53130 ^ n35700 ^ n9917 ;
  assign n53132 = ( ~n10227 & n11479 ) | ( ~n10227 & n48485 ) | ( n11479 & n48485 ) ;
  assign n53133 = n15262 ^ n13714 ^ n5570 ;
  assign n53134 = n53133 ^ n38684 ^ n22070 ;
  assign n53135 = ~n22523 & n52252 ;
  assign n53136 = n53134 & n53135 ;
  assign n53138 = ( n3340 & n12999 ) | ( n3340 & ~n29208 ) | ( n12999 & ~n29208 ) ;
  assign n53137 = n7574 & n49621 ;
  assign n53139 = n53138 ^ n53137 ^ 1'b0 ;
  assign n53140 = ( n5847 & n10735 ) | ( n5847 & ~n39685 ) | ( n10735 & ~n39685 ) ;
  assign n53141 = n53140 ^ n32789 ^ n27789 ;
  assign n53142 = n48329 ^ n29553 ^ 1'b0 ;
  assign n53143 = ( n7097 & ~n35756 ) | ( n7097 & n53142 ) | ( ~n35756 & n53142 ) ;
  assign n53144 = n16957 | n26788 ;
  assign n53145 = n17918 ^ n8569 ^ n6711 ;
  assign n53146 = n53145 ^ n14143 ^ n537 ;
  assign n53147 = ( ~n8658 & n14065 ) | ( ~n8658 & n28266 ) | ( n14065 & n28266 ) ;
  assign n53148 = ( n893 & n17087 ) | ( n893 & ~n53147 ) | ( n17087 & ~n53147 ) ;
  assign n53149 = n53113 ^ n18088 ^ n896 ;
  assign n53150 = ( n15063 & n53148 ) | ( n15063 & ~n53149 ) | ( n53148 & ~n53149 ) ;
  assign n53151 = ~n1602 & n21632 ;
  assign n53152 = ~n10849 & n53151 ;
  assign n53154 = n39458 ^ n25668 ^ n8083 ;
  assign n53153 = n45232 ^ n5996 ^ n4623 ;
  assign n53155 = n53154 ^ n53153 ^ n27991 ;
  assign n53156 = ( n11490 & ~n53152 ) | ( n11490 & n53155 ) | ( ~n53152 & n53155 ) ;
  assign n53157 = ( ~n3118 & n8756 ) | ( ~n3118 & n33570 ) | ( n8756 & n33570 ) ;
  assign n53158 = n53157 ^ n34569 ^ n26542 ;
  assign n53159 = ( n33037 & n45111 ) | ( n33037 & ~n45608 ) | ( n45111 & ~n45608 ) ;
  assign n53160 = n10264 ^ n6823 ^ 1'b0 ;
  assign n53161 = n45553 & ~n53160 ;
  assign n53162 = ~n33388 & n49456 ;
  assign n53163 = n21445 & n53162 ;
  assign n53164 = n18155 ^ n15647 ^ n6103 ;
  assign n53165 = ~n13307 & n53164 ;
  assign n53166 = ( x165 & ~n2893 ) | ( x165 & n37107 ) | ( ~n2893 & n37107 ) ;
  assign n53167 = ( ~n12787 & n27497 ) | ( ~n12787 & n53166 ) | ( n27497 & n53166 ) ;
  assign n53168 = n25343 ^ n11751 ^ 1'b0 ;
  assign n53169 = ~n504 & n53168 ;
  assign n53170 = n53169 ^ n27056 ^ n15431 ;
  assign n53171 = n53170 ^ n33185 ^ n28442 ;
  assign n53172 = ( ~n2085 & n35555 ) | ( ~n2085 & n36799 ) | ( n35555 & n36799 ) ;
  assign n53173 = n53172 ^ n46850 ^ n33260 ;
  assign n53175 = ( n9600 & n24733 ) | ( n9600 & n51892 ) | ( n24733 & n51892 ) ;
  assign n53176 = n53175 ^ n20472 ^ n6309 ;
  assign n53174 = n5884 & n24875 ;
  assign n53177 = n53176 ^ n53174 ^ 1'b0 ;
  assign n53178 = ( ~n7870 & n33143 ) | ( ~n7870 & n53177 ) | ( n33143 & n53177 ) ;
  assign n53180 = n33364 ^ n11479 ^ n451 ;
  assign n53179 = ( n16219 & ~n37740 ) | ( n16219 & n45740 ) | ( ~n37740 & n45740 ) ;
  assign n53181 = n53180 ^ n53179 ^ n48915 ;
  assign n53182 = n11610 | n13071 ;
  assign n53183 = ( n37032 & n53181 ) | ( n37032 & ~n53182 ) | ( n53181 & ~n53182 ) ;
  assign n53184 = ~n1463 & n6005 ;
  assign n53185 = n35494 & n53184 ;
  assign n53186 = n53185 ^ n48204 ^ n15866 ;
  assign n53189 = n50671 ^ n28660 ^ n17320 ;
  assign n53187 = ( n1259 & n16091 ) | ( n1259 & n27407 ) | ( n16091 & n27407 ) ;
  assign n53188 = ~n16915 & n53187 ;
  assign n53190 = n53189 ^ n53188 ^ 1'b0 ;
  assign n53191 = ( ~n12421 & n41955 ) | ( ~n12421 & n53190 ) | ( n41955 & n53190 ) ;
  assign n53192 = ( n7652 & n16470 ) | ( n7652 & ~n16753 ) | ( n16470 & ~n16753 ) ;
  assign n53193 = n53192 ^ n41460 ^ n27871 ;
  assign n53194 = ~n48176 & n49996 ;
  assign n53195 = n37252 ^ n7686 ^ 1'b0 ;
  assign n53196 = ~n53194 & n53195 ;
  assign n53202 = n3893 | n16074 ;
  assign n53203 = n2437 | n53202 ;
  assign n53197 = n19119 ^ n1858 ^ 1'b0 ;
  assign n53198 = n25944 & ~n53197 ;
  assign n53199 = ( n29616 & ~n44667 ) | ( n29616 & n53198 ) | ( ~n44667 & n53198 ) ;
  assign n53200 = ( n2225 & n42877 ) | ( n2225 & n53199 ) | ( n42877 & n53199 ) ;
  assign n53201 = n52923 & n53200 ;
  assign n53204 = n53203 ^ n53201 ^ 1'b0 ;
  assign n53205 = n18371 ^ n10074 ^ n5622 ;
  assign n53206 = n9444 & n53205 ;
  assign n53207 = n51488 ^ n38112 ^ n11995 ;
  assign n53208 = ( ~n9295 & n34124 ) | ( ~n9295 & n39846 ) | ( n34124 & n39846 ) ;
  assign n53209 = ( n9473 & n13565 ) | ( n9473 & n14711 ) | ( n13565 & n14711 ) ;
  assign n53210 = ( n7484 & n53208 ) | ( n7484 & ~n53209 ) | ( n53208 & ~n53209 ) ;
  assign n53211 = n4373 ^ n1942 ^ 1'b0 ;
  assign n53212 = n53211 ^ n14684 ^ 1'b0 ;
  assign n53213 = ( n23850 & ~n53180 ) | ( n23850 & n53212 ) | ( ~n53180 & n53212 ) ;
  assign n53214 = ( n3994 & n9234 ) | ( n3994 & n47918 ) | ( n9234 & n47918 ) ;
  assign n53215 = n53214 ^ n32704 ^ n7176 ;
  assign n53216 = n53215 ^ n26821 ^ n9222 ;
  assign n53217 = ~n10541 & n53216 ;
  assign n53218 = n33983 ^ n28804 ^ n26759 ;
  assign n53219 = ( ~n19436 & n35295 ) | ( ~n19436 & n52610 ) | ( n35295 & n52610 ) ;
  assign n53220 = n26963 ^ n6207 ^ n868 ;
  assign n53221 = n42929 ^ n30184 ^ n10081 ;
  assign n53225 = n36996 ^ n28002 ^ x175 ;
  assign n53222 = n8580 & ~n31222 ;
  assign n53223 = ~n10681 & n53222 ;
  assign n53224 = n53223 ^ n34875 ^ n34098 ;
  assign n53226 = n53225 ^ n53224 ^ n21860 ;
  assign n53227 = n34912 ^ n12230 ^ 1'b0 ;
  assign n53228 = n8804 ^ n2687 ^ n1636 ;
  assign n53229 = ( n22673 & n38363 ) | ( n22673 & n53228 ) | ( n38363 & n53228 ) ;
  assign n53230 = ( ~n762 & n33598 ) | ( ~n762 & n53229 ) | ( n33598 & n53229 ) ;
  assign n53231 = ( n25687 & ~n34773 ) | ( n25687 & n47454 ) | ( ~n34773 & n47454 ) ;
  assign n53232 = n53231 ^ n12064 ^ n1406 ;
  assign n53239 = n36621 ^ n21175 ^ n10224 ;
  assign n53240 = ( n11905 & ~n37325 ) | ( n11905 & n53239 ) | ( ~n37325 & n53239 ) ;
  assign n53236 = n15974 ^ n9384 ^ n8015 ;
  assign n53237 = ( ~n4264 & n12342 ) | ( ~n4264 & n53236 ) | ( n12342 & n53236 ) ;
  assign n53238 = ( n1567 & n15429 ) | ( n1567 & n53237 ) | ( n15429 & n53237 ) ;
  assign n53233 = n41964 ^ n28924 ^ n1304 ;
  assign n53234 = n9680 & n18683 ;
  assign n53235 = ~n53233 & n53234 ;
  assign n53241 = n53240 ^ n53238 ^ n53235 ;
  assign n53242 = ( ~n6389 & n6598 ) | ( ~n6389 & n49572 ) | ( n6598 & n49572 ) ;
  assign n53243 = n46205 ^ n25023 ^ n8301 ;
  assign n53244 = ( n2703 & n13648 ) | ( n2703 & ~n25753 ) | ( n13648 & ~n25753 ) ;
  assign n53245 = n53244 ^ n22517 ^ n18090 ;
  assign n53246 = n53245 ^ n22449 ^ n3814 ;
  assign n53247 = ( n25803 & n40081 ) | ( n25803 & n53246 ) | ( n40081 & n53246 ) ;
  assign n53252 = x201 | n52136 ;
  assign n53248 = ( ~n1094 & n7254 ) | ( ~n1094 & n16066 ) | ( n7254 & n16066 ) ;
  assign n53249 = n41495 ^ n3656 ^ 1'b0 ;
  assign n53250 = ~n53248 & n53249 ;
  assign n53251 = ( n10800 & n18415 ) | ( n10800 & n53250 ) | ( n18415 & n53250 ) ;
  assign n53253 = n53252 ^ n53251 ^ n33724 ;
  assign n53254 = n7136 & ~n13645 ;
  assign n53255 = ~n41179 & n53254 ;
  assign n53257 = n18112 ^ n12200 ^ n11715 ;
  assign n53256 = n28085 ^ n8722 ^ 1'b0 ;
  assign n53258 = n53257 ^ n53256 ^ n11810 ;
  assign n53259 = n8513 & n32610 ;
  assign n53260 = n6311 & n53259 ;
  assign n53261 = ( ~n1105 & n44159 ) | ( ~n1105 & n53260 ) | ( n44159 & n53260 ) ;
  assign n53262 = n3361 | n11341 ;
  assign n53263 = n53262 ^ n7004 ^ 1'b0 ;
  assign n53264 = ( ~n20299 & n52811 ) | ( ~n20299 & n53263 ) | ( n52811 & n53263 ) ;
  assign n53265 = n13365 & ~n23651 ;
  assign n53266 = n37548 ^ n23851 ^ n5862 ;
  assign n53267 = n11543 & n53266 ;
  assign n53268 = ( n19998 & ~n53265 ) | ( n19998 & n53267 ) | ( ~n53265 & n53267 ) ;
  assign n53269 = n20198 ^ n17561 ^ 1'b0 ;
  assign n53270 = n53269 ^ n33132 ^ n14817 ;
  assign n53271 = ( n3355 & ~n36203 ) | ( n3355 & n38681 ) | ( ~n36203 & n38681 ) ;
  assign n53273 = ( n13450 & ~n22644 ) | ( n13450 & n33371 ) | ( ~n22644 & n33371 ) ;
  assign n53272 = n36989 ^ n12325 ^ n7225 ;
  assign n53274 = n53273 ^ n53272 ^ n28633 ;
  assign n53275 = n53274 ^ n50094 ^ n4438 ;
  assign n53276 = ( n2815 & n14010 ) | ( n2815 & n53275 ) | ( n14010 & n53275 ) ;
  assign n53277 = n46215 ^ n7392 ^ n3058 ;
  assign n53278 = n13598 & ~n27891 ;
  assign n53279 = n11574 & n53278 ;
  assign n53280 = n28132 ^ n17353 ^ 1'b0 ;
  assign n53281 = n49581 & n53280 ;
  assign n53282 = n53281 ^ n32678 ^ n11596 ;
  assign n53283 = ( n16440 & n20270 ) | ( n16440 & ~n41157 ) | ( n20270 & ~n41157 ) ;
  assign n53285 = ( n4733 & n5028 ) | ( n4733 & ~n36881 ) | ( n5028 & ~n36881 ) ;
  assign n53284 = n35027 ^ n34402 ^ n2883 ;
  assign n53286 = n53285 ^ n53284 ^ n25411 ;
  assign n53289 = n14224 ^ n8374 ^ 1'b0 ;
  assign n53287 = n5729 ^ n1764 ^ 1'b0 ;
  assign n53288 = n9447 & n53287 ;
  assign n53290 = n53289 ^ n53288 ^ 1'b0 ;
  assign n53291 = ( n4216 & ~n34353 ) | ( n4216 & n44421 ) | ( ~n34353 & n44421 ) ;
  assign n53292 = ( n33508 & n48759 ) | ( n33508 & n53291 ) | ( n48759 & n53291 ) ;
  assign n53294 = n6347 ^ n1899 ^ 1'b0 ;
  assign n53293 = n34628 ^ n31697 ^ 1'b0 ;
  assign n53295 = n53294 ^ n53293 ^ n26016 ;
  assign n53296 = n53295 ^ n28596 ^ n28255 ;
  assign n53297 = n49708 ^ n11433 ^ n3834 ;
  assign n53298 = n49394 ^ n8709 ^ 1'b0 ;
  assign n53299 = ( n7387 & n34441 ) | ( n7387 & ~n53298 ) | ( n34441 & ~n53298 ) ;
  assign n53301 = ( ~n3180 & n7428 ) | ( ~n3180 & n22090 ) | ( n7428 & n22090 ) ;
  assign n53300 = n42161 ^ n40377 ^ n7225 ;
  assign n53302 = n53301 ^ n53300 ^ n28254 ;
  assign n53303 = ( n7113 & ~n12974 ) | ( n7113 & n53302 ) | ( ~n12974 & n53302 ) ;
  assign n53304 = n3596 & ~n12631 ;
  assign n53305 = n53304 ^ n43153 ^ 1'b0 ;
  assign n53306 = ( n5532 & n12446 ) | ( n5532 & n14362 ) | ( n12446 & n14362 ) ;
  assign n53307 = n5447 & ~n45212 ;
  assign n53308 = n53306 & n53307 ;
  assign n53309 = ( ~n13436 & n15830 ) | ( ~n13436 & n37443 ) | ( n15830 & n37443 ) ;
  assign n53313 = n20013 ^ n13551 ^ n3175 ;
  assign n53310 = ~n9860 & n17524 ;
  assign n53311 = n11824 & n53310 ;
  assign n53312 = n53311 ^ n13722 ^ n2093 ;
  assign n53314 = n53313 ^ n53312 ^ n30038 ;
  assign n53315 = n37327 ^ n8453 ^ n6713 ;
  assign n53316 = ( ~n2122 & n38201 ) | ( ~n2122 & n53315 ) | ( n38201 & n53315 ) ;
  assign n53317 = n53316 ^ n34792 ^ n31573 ;
  assign n53318 = ( ~n12809 & n15212 ) | ( ~n12809 & n19728 ) | ( n15212 & n19728 ) ;
  assign n53319 = ( ~n16966 & n31767 ) | ( ~n16966 & n53318 ) | ( n31767 & n53318 ) ;
  assign n53320 = ( n6772 & n34111 ) | ( n6772 & n53319 ) | ( n34111 & n53319 ) ;
  assign n53321 = n48534 ^ n12121 ^ n11869 ;
  assign n53322 = n16533 ^ n15229 ^ n753 ;
  assign n53323 = n17953 ^ n16310 ^ n9395 ;
  assign n53324 = n53323 ^ n6100 ^ n883 ;
  assign n53325 = n30397 ^ n28204 ^ n6008 ;
  assign n53326 = n34316 ^ n2298 ^ 1'b0 ;
  assign n53327 = ( ~n5105 & n53325 ) | ( ~n5105 & n53326 ) | ( n53325 & n53326 ) ;
  assign n53328 = ( n13128 & n20719 ) | ( n13128 & n47424 ) | ( n20719 & n47424 ) ;
  assign n53329 = n53328 ^ n9879 ^ 1'b0 ;
  assign n53330 = n11802 | n53329 ;
  assign n53331 = n9761 & ~n36830 ;
  assign n53332 = ~n2639 & n53331 ;
  assign n53333 = ( n1257 & n13894 ) | ( n1257 & n19830 ) | ( n13894 & n19830 ) ;
  assign n53334 = n53333 ^ n11349 ^ n7655 ;
  assign n53335 = ( n551 & n7921 ) | ( n551 & n16050 ) | ( n7921 & n16050 ) ;
  assign n53336 = n21728 & n27761 ;
  assign n53337 = n38969 ^ n29932 ^ n23758 ;
  assign n53338 = n53337 ^ n15477 ^ 1'b0 ;
  assign n53339 = n20926 & n53338 ;
  assign n53340 = ~n8566 & n53339 ;
  assign n53341 = n53340 ^ n8626 ^ 1'b0 ;
  assign n53342 = ~n4831 & n53341 ;
  assign n53343 = ~n8591 & n36080 ;
  assign n53344 = ~n50067 & n53343 ;
  assign n53345 = ( ~n19393 & n28158 ) | ( ~n19393 & n53344 ) | ( n28158 & n53344 ) ;
  assign n53346 = n53345 ^ n51458 ^ 1'b0 ;
  assign n53347 = ( n4974 & n53342 ) | ( n4974 & n53346 ) | ( n53342 & n53346 ) ;
  assign n53348 = ( n30131 & ~n45653 ) | ( n30131 & n46562 ) | ( ~n45653 & n46562 ) ;
  assign n53349 = n3147 | n21330 ;
  assign n53350 = n25022 ^ n16303 ^ 1'b0 ;
  assign n53351 = n53350 ^ n46265 ^ n18550 ;
  assign n53352 = n36648 ^ n27122 ^ n3604 ;
  assign n53353 = n13777 & ~n14056 ;
  assign n53354 = n53352 & n53353 ;
  assign n53355 = n31479 & ~n34580 ;
  assign n53356 = n6548 & ~n53355 ;
  assign n53357 = n49653 ^ n47222 ^ n7433 ;
  assign n53358 = ( n29290 & n31325 ) | ( n29290 & ~n31585 ) | ( n31325 & ~n31585 ) ;
  assign n53359 = ( ~n10318 & n28871 ) | ( ~n10318 & n42028 ) | ( n28871 & n42028 ) ;
  assign n53360 = n49318 ^ n33992 ^ n8916 ;
  assign n53361 = n53360 ^ n52339 ^ n45795 ;
  assign n53362 = n46982 ^ n16516 ^ n8464 ;
  assign n53363 = n21157 & ~n53362 ;
  assign n53364 = ~n37852 & n53363 ;
  assign n53365 = ( n7847 & n14784 ) | ( n7847 & n53364 ) | ( n14784 & n53364 ) ;
  assign n53366 = n1090 | n11748 ;
  assign n53367 = ( n17865 & ~n20657 ) | ( n17865 & n53366 ) | ( ~n20657 & n53366 ) ;
  assign n53368 = ~n28136 & n49700 ;
  assign n53369 = n24089 ^ n15901 ^ n5822 ;
  assign n53370 = n53369 ^ n45387 ^ n36303 ;
  assign n53371 = ( n3255 & ~n11833 ) | ( n3255 & n53370 ) | ( ~n11833 & n53370 ) ;
  assign n53373 = ( n2919 & n5327 ) | ( n2919 & n5399 ) | ( n5327 & n5399 ) ;
  assign n53374 = n53373 ^ n12689 ^ n8439 ;
  assign n53372 = n37010 | n53314 ;
  assign n53375 = n53374 ^ n53372 ^ 1'b0 ;
  assign n53376 = n44848 ^ n19494 ^ n8093 ;
  assign n53377 = n53376 ^ n37402 ^ n20690 ;
  assign n53378 = n46123 ^ n5594 ^ n4180 ;
  assign n53379 = ( n4234 & n12524 ) | ( n4234 & n32186 ) | ( n12524 & n32186 ) ;
  assign n53380 = ( n7438 & n12689 ) | ( n7438 & n29406 ) | ( n12689 & n29406 ) ;
  assign n53381 = ( n22581 & n34535 ) | ( n22581 & n38773 ) | ( n34535 & n38773 ) ;
  assign n53382 = ( ~n26170 & n31439 ) | ( ~n26170 & n46932 ) | ( n31439 & n46932 ) ;
  assign n53383 = n53382 ^ n38602 ^ 1'b0 ;
  assign n53384 = ~n47598 & n53383 ;
  assign n53385 = n53384 ^ n41999 ^ n7201 ;
  assign n53386 = ( ~n41390 & n44796 ) | ( ~n41390 & n48688 ) | ( n44796 & n48688 ) ;
  assign n53387 = ~n12069 & n50434 ;
  assign n53388 = n53387 ^ n52249 ^ 1'b0 ;
  assign n53389 = n43208 ^ n24987 ^ 1'b0 ;
  assign n53390 = n50104 ^ n48643 ^ n16612 ;
  assign n53391 = n23685 ^ n19552 ^ n19530 ;
  assign n53392 = ( n24116 & ~n24916 ) | ( n24116 & n26410 ) | ( ~n24916 & n26410 ) ;
  assign n53393 = n46397 ^ n16351 ^ 1'b0 ;
  assign n53394 = n16382 | n53393 ;
  assign n53395 = n53394 ^ n23291 ^ n17383 ;
  assign n53396 = ~n19553 & n36947 ;
  assign n53397 = ~n45223 & n53396 ;
  assign n53398 = ( n7925 & ~n28779 ) | ( n7925 & n53397 ) | ( ~n28779 & n53397 ) ;
  assign n53399 = n52750 ^ n24818 ^ n18938 ;
  assign n53400 = ( n28565 & ~n48158 ) | ( n28565 & n53399 ) | ( ~n48158 & n53399 ) ;
  assign n53401 = n52033 ^ n49359 ^ n11347 ;
  assign n53403 = ( ~n14052 & n35701 ) | ( ~n14052 & n48708 ) | ( n35701 & n48708 ) ;
  assign n53402 = n28595 ^ n26113 ^ n14382 ;
  assign n53404 = n53403 ^ n53402 ^ n35288 ;
  assign n53405 = n4123 ^ n2814 ^ 1'b0 ;
  assign n53406 = n6852 ^ n6725 ^ n5178 ;
  assign n53407 = ( n1245 & n32931 ) | ( n1245 & ~n48589 ) | ( n32931 & ~n48589 ) ;
  assign n53408 = n31561 & ~n53407 ;
  assign n53409 = n53406 & n53408 ;
  assign n53410 = n10232 | n19578 ;
  assign n53411 = n23128 | n53410 ;
  assign n53412 = n53411 ^ n24226 ^ n5740 ;
  assign n53413 = n53412 ^ n35157 ^ n2929 ;
  assign n53414 = n47307 ^ n33057 ^ n1783 ;
  assign n53415 = n34646 ^ n18723 ^ n8055 ;
  assign n53416 = ( n1542 & ~n4399 ) | ( n1542 & n53415 ) | ( ~n4399 & n53415 ) ;
  assign n53418 = ( n5756 & ~n13138 ) | ( n5756 & n30811 ) | ( ~n13138 & n30811 ) ;
  assign n53419 = n53418 ^ n35459 ^ n1760 ;
  assign n53417 = n27541 ^ n13054 ^ n7432 ;
  assign n53420 = n53419 ^ n53417 ^ n2980 ;
  assign n53421 = ( n13937 & n18848 ) | ( n13937 & ~n22374 ) | ( n18848 & ~n22374 ) ;
  assign n53422 = n53421 ^ n48845 ^ n40967 ;
  assign n53423 = ( n7725 & n19816 ) | ( n7725 & n28560 ) | ( n19816 & n28560 ) ;
  assign n53425 = ( n984 & n12286 ) | ( n984 & n22536 ) | ( n12286 & n22536 ) ;
  assign n53424 = ~n19406 & n25560 ;
  assign n53426 = n53425 ^ n53424 ^ 1'b0 ;
  assign n53427 = n53426 ^ n51504 ^ n4109 ;
  assign n53428 = ( ~n1861 & n10587 ) | ( ~n1861 & n53427 ) | ( n10587 & n53427 ) ;
  assign n53430 = ( n27177 & ~n50130 ) | ( n27177 & n51347 ) | ( ~n50130 & n51347 ) ;
  assign n53429 = ( n1801 & n5336 ) | ( n1801 & ~n15339 ) | ( n5336 & ~n15339 ) ;
  assign n53431 = n53430 ^ n53429 ^ n27565 ;
  assign n53432 = n53431 ^ n15557 ^ n276 ;
  assign n53433 = n24378 ^ n4228 ^ n2797 ;
  assign n53434 = n53433 ^ n9344 ^ n6908 ;
  assign n53435 = n53434 ^ n20051 ^ n5416 ;
  assign n53436 = ( n50721 & ~n53432 ) | ( n50721 & n53435 ) | ( ~n53432 & n53435 ) ;
  assign n53437 = n41308 ^ n16704 ^ 1'b0 ;
  assign n53439 = ( n7688 & n12157 ) | ( n7688 & n20987 ) | ( n12157 & n20987 ) ;
  assign n53438 = ~n3380 & n41436 ;
  assign n53440 = n53439 ^ n53438 ^ 1'b0 ;
  assign n53441 = ( n15847 & ~n31162 ) | ( n15847 & n33992 ) | ( ~n31162 & n33992 ) ;
  assign n53442 = ( n9785 & n38983 ) | ( n9785 & n51003 ) | ( n38983 & n51003 ) ;
  assign n53443 = ( n50882 & ~n52837 ) | ( n50882 & n53442 ) | ( ~n52837 & n53442 ) ;
  assign n53444 = n41519 ^ n21643 ^ n8045 ;
  assign n53445 = n17030 | n33405 ;
  assign n53446 = ( n14322 & n18695 ) | ( n14322 & ~n53445 ) | ( n18695 & ~n53445 ) ;
  assign n53447 = n30661 ^ n18937 ^ n18402 ;
  assign n53448 = n53447 ^ n38733 ^ n1079 ;
  assign n53449 = n21698 ^ n19506 ^ n15864 ;
  assign n53450 = n42654 ^ n35108 ^ n9074 ;
  assign n53451 = n53205 ^ n41978 ^ n33907 ;
  assign n53452 = n34638 ^ n16766 ^ n6464 ;
  assign n53453 = ( n11896 & n26175 ) | ( n11896 & n53452 ) | ( n26175 & n53452 ) ;
  assign n53454 = ( n6784 & n53451 ) | ( n6784 & ~n53453 ) | ( n53451 & ~n53453 ) ;
  assign n53455 = n14182 ^ n7841 ^ x118 ;
  assign n53456 = n34877 ^ n33523 ^ n7778 ;
  assign n53457 = n40330 ^ n21426 ^ 1'b0 ;
  assign n53458 = n53456 & n53457 ;
  assign n53459 = n6199 & n41500 ;
  assign n53463 = ( ~n881 & n9323 ) | ( ~n881 & n39272 ) | ( n9323 & n39272 ) ;
  assign n53461 = n13340 ^ n9316 ^ n4573 ;
  assign n53460 = n26307 ^ n19664 ^ n6746 ;
  assign n53462 = n53461 ^ n53460 ^ n26069 ;
  assign n53464 = n53463 ^ n53462 ^ n27534 ;
  assign n53465 = n18870 ^ n9807 ^ n8239 ;
  assign n53466 = n26770 ^ n23711 ^ n20114 ;
  assign n53467 = n22147 & ~n43772 ;
  assign n53468 = ( n18015 & n53466 ) | ( n18015 & n53467 ) | ( n53466 & n53467 ) ;
  assign n53469 = ( n4110 & n18900 ) | ( n4110 & ~n27901 ) | ( n18900 & ~n27901 ) ;
  assign n53470 = ( n17667 & n38225 ) | ( n17667 & n53469 ) | ( n38225 & n53469 ) ;
  assign n53471 = n19921 ^ n6995 ^ n1198 ;
  assign n53472 = n53471 ^ n14449 ^ 1'b0 ;
  assign n53473 = n36044 ^ n34838 ^ n34710 ;
  assign n53474 = n4319 | n33315 ;
  assign n53475 = n40772 ^ n38713 ^ 1'b0 ;
  assign n53476 = n5352 & ~n53475 ;
  assign n53478 = ( x105 & n11420 ) | ( x105 & ~n15234 ) | ( n11420 & ~n15234 ) ;
  assign n53479 = n53478 ^ n12021 ^ n6646 ;
  assign n53477 = n47543 ^ n9867 ^ n8718 ;
  assign n53480 = n53479 ^ n53477 ^ n1496 ;
  assign n53481 = n40674 ^ n16925 ^ 1'b0 ;
  assign n53482 = n29114 | n39696 ;
  assign n53485 = n18915 ^ n8142 ^ n6226 ;
  assign n53484 = n6579 ^ n3184 ^ 1'b0 ;
  assign n53483 = ( n24929 & ~n32363 ) | ( n24929 & n41495 ) | ( ~n32363 & n41495 ) ;
  assign n53486 = n53485 ^ n53484 ^ n53483 ;
  assign n53487 = ( x199 & n13904 ) | ( x199 & n24994 ) | ( n13904 & n24994 ) ;
  assign n53488 = ( n2659 & n3343 ) | ( n2659 & ~n53487 ) | ( n3343 & ~n53487 ) ;
  assign n53489 = n49477 ^ n43736 ^ n6805 ;
  assign n53490 = ( ~x46 & n11290 ) | ( ~x46 & n11767 ) | ( n11290 & n11767 ) ;
  assign n53491 = n19700 & n53490 ;
  assign n53492 = n53491 ^ n15892 ^ n8109 ;
  assign n53493 = ( ~n1077 & n16141 ) | ( ~n1077 & n28175 ) | ( n16141 & n28175 ) ;
  assign n53494 = n53493 ^ n30071 ^ n28841 ;
  assign n53495 = n35300 & ~n42172 ;
  assign n53496 = ( ~n8676 & n15840 ) | ( ~n8676 & n41507 ) | ( n15840 & n41507 ) ;
  assign n53497 = n53496 ^ n31105 ^ 1'b0 ;
  assign n53498 = n3712 & ~n53497 ;
  assign n53499 = ~n6050 & n17761 ;
  assign n53500 = n53499 ^ n47987 ^ 1'b0 ;
  assign n53501 = ~n23456 & n52181 ;
  assign n53502 = n9807 ^ n2866 ^ 1'b0 ;
  assign n53503 = ( n3667 & n22161 ) | ( n3667 & ~n34545 ) | ( n22161 & ~n34545 ) ;
  assign n53504 = n53503 ^ n17222 ^ n883 ;
  assign n53505 = ( ~n23223 & n52817 ) | ( ~n23223 & n53504 ) | ( n52817 & n53504 ) ;
  assign n53506 = n25960 | n42544 ;
  assign n53507 = ( n11586 & n28925 ) | ( n11586 & ~n51379 ) | ( n28925 & ~n51379 ) ;
  assign n53509 = ( n1982 & ~n2304 ) | ( n1982 & n8430 ) | ( ~n2304 & n8430 ) ;
  assign n53508 = ( n14803 & n23466 ) | ( n14803 & n27602 ) | ( n23466 & n27602 ) ;
  assign n53510 = n53509 ^ n53508 ^ n53209 ;
  assign n53515 = ( n8907 & ~n22514 ) | ( n8907 & n48805 ) | ( ~n22514 & n48805 ) ;
  assign n53512 = ( n7261 & n7658 ) | ( n7261 & n22121 ) | ( n7658 & n22121 ) ;
  assign n53513 = ( ~n17606 & n35420 ) | ( ~n17606 & n53512 ) | ( n35420 & n53512 ) ;
  assign n53511 = n33826 ^ n10372 ^ n5105 ;
  assign n53514 = n53513 ^ n53511 ^ n25753 ;
  assign n53516 = n53515 ^ n53514 ^ n31028 ;
  assign n53517 = n5138 & n19938 ;
  assign n53518 = n53274 & n53517 ;
  assign n53519 = n53518 ^ n19661 ^ n13192 ;
  assign n53520 = n43356 ^ n39087 ^ 1'b0 ;
  assign n53521 = n12491 | n53520 ;
  assign n53522 = n21728 & n22220 ;
  assign n53523 = ( n12359 & n28468 ) | ( n12359 & ~n53522 ) | ( n28468 & ~n53522 ) ;
  assign n53524 = ~n1701 & n53523 ;
  assign n53525 = ~n18422 & n53524 ;
  assign n53526 = n48280 ^ n28385 ^ n14967 ;
  assign n53527 = ( n15062 & ~n17890 ) | ( n15062 & n21759 ) | ( ~n17890 & n21759 ) ;
  assign n53528 = ( ~n5893 & n7643 ) | ( ~n5893 & n29058 ) | ( n7643 & n29058 ) ;
  assign n53529 = ( n10489 & ~n20493 ) | ( n10489 & n46492 ) | ( ~n20493 & n46492 ) ;
  assign n53530 = n53529 ^ n50256 ^ n38395 ;
  assign n53531 = ( n4517 & ~n39725 ) | ( n4517 & n43326 ) | ( ~n39725 & n43326 ) ;
  assign n53532 = n42100 ^ n35382 ^ n8072 ;
  assign n53533 = n46538 ^ n30616 ^ n6921 ;
  assign n53534 = ( n11199 & ~n17291 ) | ( n11199 & n35622 ) | ( ~n17291 & n35622 ) ;
  assign n53535 = n45518 ^ n38353 ^ 1'b0 ;
  assign n53536 = n19492 & ~n53535 ;
  assign n53537 = n35526 ^ n33823 ^ n28657 ;
  assign n53538 = n53537 ^ n45654 ^ 1'b0 ;
  assign n53539 = ~n31138 & n53538 ;
  assign n53540 = ~n9145 & n37051 ;
  assign n53541 = ~n30570 & n53540 ;
  assign n53542 = ( n10464 & n32700 ) | ( n10464 & n53541 ) | ( n32700 & n53541 ) ;
  assign n53543 = ( ~n22391 & n43055 ) | ( ~n22391 & n53542 ) | ( n43055 & n53542 ) ;
  assign n53544 = n46961 ^ n27148 ^ 1'b0 ;
  assign n53545 = n38748 ^ n23729 ^ n16659 ;
  assign n53546 = n53545 ^ n32509 ^ n345 ;
  assign n53547 = n6539 & n48623 ;
  assign n53548 = ( n5288 & ~n18039 ) | ( n5288 & n30384 ) | ( ~n18039 & n30384 ) ;
  assign n53549 = n47192 ^ n39399 ^ n29028 ;
  assign n53550 = n43040 ^ n27582 ^ n977 ;
  assign n53551 = n32641 ^ n22544 ^ n17584 ;
  assign n53552 = n4797 | n20106 ;
  assign n53553 = x215 | n53552 ;
  assign n53554 = n29493 ^ n14842 ^ 1'b0 ;
  assign n53555 = n10448 ^ n7892 ^ 1'b0 ;
  assign n53556 = ( n11120 & n53554 ) | ( n11120 & ~n53555 ) | ( n53554 & ~n53555 ) ;
  assign n53557 = n33622 ^ n27556 ^ n23722 ;
  assign n53558 = n33208 ^ n22721 ^ n20015 ;
  assign n53559 = ( n22453 & n53557 ) | ( n22453 & n53558 ) | ( n53557 & n53558 ) ;
  assign n53564 = ( n4058 & n35383 ) | ( n4058 & ~n49646 ) | ( n35383 & ~n49646 ) ;
  assign n53563 = n16819 ^ n16202 ^ n11579 ;
  assign n53565 = n53564 ^ n53563 ^ n33132 ;
  assign n53560 = ( n20908 & ~n23355 ) | ( n20908 & n30059 ) | ( ~n23355 & n30059 ) ;
  assign n53561 = n53560 ^ n45060 ^ n8867 ;
  assign n53562 = ( n11902 & n49993 ) | ( n11902 & ~n53561 ) | ( n49993 & ~n53561 ) ;
  assign n53566 = n53565 ^ n53562 ^ n41277 ;
  assign n53567 = n23811 ^ n12530 ^ 1'b0 ;
  assign n53568 = n2204 | n53567 ;
  assign n53570 = ~n19262 & n20728 ;
  assign n53571 = n53570 ^ n7423 ^ 1'b0 ;
  assign n53572 = ( n29058 & n36241 ) | ( n29058 & ~n53571 ) | ( n36241 & ~n53571 ) ;
  assign n53569 = n37173 ^ n26098 ^ n7654 ;
  assign n53573 = n53572 ^ n53569 ^ n2424 ;
  assign n53574 = ( ~n31270 & n53568 ) | ( ~n31270 & n53573 ) | ( n53568 & n53573 ) ;
  assign n53575 = ( n28804 & n36356 ) | ( n28804 & ~n53574 ) | ( n36356 & ~n53574 ) ;
  assign n53576 = ( n2884 & n24604 ) | ( n2884 & ~n29691 ) | ( n24604 & ~n29691 ) ;
  assign n53577 = n53576 ^ n6761 ^ x208 ;
  assign n53578 = ( n931 & n7833 ) | ( n931 & n10621 ) | ( n7833 & n10621 ) ;
  assign n53579 = n8850 ^ n4936 ^ 1'b0 ;
  assign n53580 = ( n1960 & n3336 ) | ( n1960 & ~n21910 ) | ( n3336 & ~n21910 ) ;
  assign n53581 = ( n21396 & ~n41709 ) | ( n21396 & n53580 ) | ( ~n41709 & n53580 ) ;
  assign n53582 = n21261 | n53581 ;
  assign n53583 = n12911 | n53582 ;
  assign n53584 = ( n16368 & ~n53579 ) | ( n16368 & n53583 ) | ( ~n53579 & n53583 ) ;
  assign n53585 = ( ~n28909 & n53578 ) | ( ~n28909 & n53584 ) | ( n53578 & n53584 ) ;
  assign n53586 = ( ~n2768 & n11198 ) | ( ~n2768 & n16867 ) | ( n11198 & n16867 ) ;
  assign n53587 = ( n4670 & n19974 ) | ( n4670 & n53586 ) | ( n19974 & n53586 ) ;
  assign n53588 = n34130 ^ n23540 ^ n10702 ;
  assign n53589 = n24273 ^ n6293 ^ n6118 ;
  assign n53590 = ( ~n36471 & n53588 ) | ( ~n36471 & n53589 ) | ( n53588 & n53589 ) ;
  assign n53600 = ( n624 & ~n3125 ) | ( n624 & n29850 ) | ( ~n3125 & n29850 ) ;
  assign n53598 = ( ~n23811 & n40997 ) | ( ~n23811 & n45619 ) | ( n40997 & n45619 ) ;
  assign n53592 = n39857 ^ n4751 ^ 1'b0 ;
  assign n53593 = n17905 ^ x195 ^ 1'b0 ;
  assign n53594 = n39268 & n53593 ;
  assign n53595 = ( ~n15704 & n53592 ) | ( ~n15704 & n53594 ) | ( n53592 & n53594 ) ;
  assign n53596 = ~n3784 & n53595 ;
  assign n53597 = n2570 & n53596 ;
  assign n53591 = n18592 ^ n2093 ^ 1'b0 ;
  assign n53599 = n53598 ^ n53597 ^ n53591 ;
  assign n53601 = n53600 ^ n53599 ^ n1170 ;
  assign n53602 = n34078 & ~n40995 ;
  assign n53603 = n1809 & n53602 ;
  assign n53604 = n44967 ^ n10828 ^ 1'b0 ;
  assign n53605 = n30914 & ~n40434 ;
  assign n53606 = n53605 ^ x190 ^ 1'b0 ;
  assign n53607 = ( n10773 & ~n11948 ) | ( n10773 & n53606 ) | ( ~n11948 & n53606 ) ;
  assign n53608 = ( n1581 & ~n23606 ) | ( n1581 & n49478 ) | ( ~n23606 & n49478 ) ;
  assign n53609 = ( n6985 & n25546 ) | ( n6985 & n37095 ) | ( n25546 & n37095 ) ;
  assign n53610 = ( ~n42657 & n46078 ) | ( ~n42657 & n53609 ) | ( n46078 & n53609 ) ;
  assign n53613 = ( n2497 & n16988 ) | ( n2497 & ~n31676 ) | ( n16988 & ~n31676 ) ;
  assign n53611 = ( ~n9572 & n14797 ) | ( ~n9572 & n43647 ) | ( n14797 & n43647 ) ;
  assign n53612 = n53611 ^ n28335 ^ n8048 ;
  assign n53614 = n53613 ^ n53612 ^ n52066 ;
  assign n53615 = n37126 ^ n11525 ^ n9024 ;
  assign n53616 = n53615 ^ n25230 ^ 1'b0 ;
  assign n53617 = n53616 ^ n41766 ^ n11645 ;
  assign n53618 = n53617 ^ n36351 ^ n12842 ;
  assign n53624 = ( n1986 & n8561 ) | ( n1986 & n24457 ) | ( n8561 & n24457 ) ;
  assign n53621 = x186 & ~n15940 ;
  assign n53622 = n53621 ^ n2411 ^ 1'b0 ;
  assign n53619 = ( x192 & x193 ) | ( x192 & n27141 ) | ( x193 & n27141 ) ;
  assign n53620 = n53619 ^ n20040 ^ n10613 ;
  assign n53623 = n53622 ^ n53620 ^ n20177 ;
  assign n53625 = n53624 ^ n53623 ^ n13090 ;
  assign n53626 = n41809 ^ n27339 ^ 1'b0 ;
  assign n53627 = n23468 & n53626 ;
  assign n53628 = n53627 ^ n9547 ^ n1270 ;
  assign n53629 = ( n8099 & n24041 ) | ( n8099 & n42694 ) | ( n24041 & n42694 ) ;
  assign n53630 = n9674 & n14672 ;
  assign n53631 = ~n13379 & n53630 ;
  assign n53632 = n3939 & n9538 ;
  assign n53633 = n21844 & n53632 ;
  assign n53634 = ( n9522 & n43642 ) | ( n9522 & ~n53633 ) | ( n43642 & ~n53633 ) ;
  assign n53635 = n12109 | n32070 ;
  assign n53636 = ( n7925 & n8682 ) | ( n7925 & n26108 ) | ( n8682 & n26108 ) ;
  assign n53637 = n53636 ^ n31190 ^ n8066 ;
  assign n53642 = ( n32522 & ~n43210 ) | ( n32522 & n49096 ) | ( ~n43210 & n49096 ) ;
  assign n53643 = ~n17589 & n31495 ;
  assign n53644 = n53642 & n53643 ;
  assign n53640 = n4414 ^ n4109 ^ 1'b0 ;
  assign n53641 = n51196 & ~n53640 ;
  assign n53645 = n53644 ^ n53641 ^ 1'b0 ;
  assign n53638 = n26414 ^ n15791 ^ n15658 ;
  assign n53639 = ( n21921 & ~n25194 ) | ( n21921 & n53638 ) | ( ~n25194 & n53638 ) ;
  assign n53646 = n53645 ^ n53639 ^ n16061 ;
  assign n53647 = n32962 ^ n27838 ^ n18235 ;
  assign n53648 = n16878 ^ n16195 ^ n11994 ;
  assign n53649 = n53648 ^ n21348 ^ n7334 ;
  assign n53652 = ( n5048 & ~n19073 ) | ( n5048 & n35156 ) | ( ~n19073 & n35156 ) ;
  assign n53650 = n43431 ^ n485 ^ 1'b0 ;
  assign n53651 = n21395 | n53650 ;
  assign n53653 = n53652 ^ n53651 ^ n9986 ;
  assign n53654 = n38326 ^ n8119 ^ n1539 ;
  assign n53655 = n39361 ^ n10017 ^ n2228 ;
  assign n53656 = n23234 ^ n12576 ^ 1'b0 ;
  assign n53657 = ~n21973 & n53656 ;
  assign n53658 = n43563 ^ n24759 ^ n10451 ;
  assign n53659 = n37293 ^ n27328 ^ n4980 ;
  assign n53660 = ~n48883 & n53659 ;
  assign n53661 = n19683 ^ n4744 ^ n3390 ;
  assign n53662 = ( n4221 & ~n30443 ) | ( n4221 & n53661 ) | ( ~n30443 & n53661 ) ;
  assign n53663 = ( n25744 & n25851 ) | ( n25744 & n53662 ) | ( n25851 & n53662 ) ;
  assign n53664 = ( n18153 & ~n21720 ) | ( n18153 & n23371 ) | ( ~n21720 & n23371 ) ;
  assign n53665 = n17868 ^ n13324 ^ n7135 ;
  assign n53666 = n53665 ^ n27060 ^ n11492 ;
  assign n53667 = n29012 ^ n5448 ^ n3343 ;
  assign n53668 = n53667 ^ n13762 ^ n5445 ;
  assign n53669 = n53668 ^ n47816 ^ n3849 ;
  assign n53670 = n28808 ^ n13186 ^ n4007 ;
  assign n53671 = n36504 ^ n12854 ^ n2143 ;
  assign n53672 = n24457 ^ n23714 ^ n16611 ;
  assign n53673 = ( n10167 & n21846 ) | ( n10167 & n22302 ) | ( n21846 & n22302 ) ;
  assign n53674 = n6382 & n52335 ;
  assign n53675 = ~n53673 & n53674 ;
  assign n53676 = ( n486 & ~n22085 ) | ( n486 & n23197 ) | ( ~n22085 & n23197 ) ;
  assign n53677 = ( n5082 & n7818 ) | ( n5082 & ~n53676 ) | ( n7818 & ~n53676 ) ;
  assign n53678 = n26682 | n53677 ;
  assign n53679 = ~n34099 & n53678 ;
  assign n53680 = n17162 & n53679 ;
  assign n53683 = n18552 ^ n12582 ^ 1'b0 ;
  assign n53681 = n10315 & n12170 ;
  assign n53682 = n24032 & n53681 ;
  assign n53684 = n53683 ^ n53682 ^ n13261 ;
  assign n53685 = n53684 ^ n39599 ^ n5146 ;
  assign n53691 = ( n3121 & n14200 ) | ( n3121 & ~n33251 ) | ( n14200 & ~n33251 ) ;
  assign n53690 = ( n10394 & ~n18427 ) | ( n10394 & n26122 ) | ( ~n18427 & n26122 ) ;
  assign n53688 = ( ~n1288 & n16507 ) | ( ~n1288 & n20521 ) | ( n16507 & n20521 ) ;
  assign n53686 = ~n23015 & n51988 ;
  assign n53687 = n19577 & n53686 ;
  assign n53689 = n53688 ^ n53687 ^ n37284 ;
  assign n53692 = n53691 ^ n53690 ^ n53689 ;
  assign n53693 = n48623 ^ n40030 ^ n8844 ;
  assign n53694 = ( n5834 & ~n9973 ) | ( n5834 & n29226 ) | ( ~n9973 & n29226 ) ;
  assign n53695 = n7415 & n19036 ;
  assign n53696 = n53695 ^ n5723 ^ 1'b0 ;
  assign n53697 = ( ~n19946 & n44807 ) | ( ~n19946 & n53696 ) | ( n44807 & n53696 ) ;
  assign n53698 = n53697 ^ n48770 ^ n12653 ;
  assign n53699 = n30628 ^ n7711 ^ n537 ;
  assign n53700 = ( n6362 & n7897 ) | ( n6362 & n9391 ) | ( n7897 & n9391 ) ;
  assign n53701 = ~n19142 & n41281 ;
  assign n53703 = n43881 ^ n39897 ^ n24779 ;
  assign n53702 = ( n4829 & ~n5737 ) | ( n4829 & n29043 ) | ( ~n5737 & n29043 ) ;
  assign n53704 = n53703 ^ n53702 ^ n11595 ;
  assign n53705 = ( n2895 & ~n41067 ) | ( n2895 & n53704 ) | ( ~n41067 & n53704 ) ;
  assign n53706 = n53705 ^ n51682 ^ n13105 ;
  assign n53707 = n50931 ^ n6940 ^ 1'b0 ;
  assign n53708 = n34140 & ~n53707 ;
  assign n53709 = n37812 ^ n23831 ^ n14847 ;
  assign n53710 = n8076 & ~n53709 ;
  assign n53711 = ( n10085 & ~n16335 ) | ( n10085 & n47020 ) | ( ~n16335 & n47020 ) ;
  assign n53712 = n23367 & ~n53711 ;
  assign n53713 = ~n53710 & n53712 ;
  assign n53714 = ( n6468 & n14544 ) | ( n6468 & n25661 ) | ( n14544 & n25661 ) ;
  assign n53715 = ( n39880 & n51596 ) | ( n39880 & n53714 ) | ( n51596 & n53714 ) ;
  assign n53716 = n21251 ^ n15102 ^ 1'b0 ;
  assign n53717 = ~n5458 & n53716 ;
  assign n53718 = ( n3501 & n27824 ) | ( n3501 & ~n53717 ) | ( n27824 & ~n53717 ) ;
  assign n53719 = ( n3475 & n9627 ) | ( n3475 & ~n53718 ) | ( n9627 & ~n53718 ) ;
  assign n53720 = n53403 ^ n23902 ^ n1275 ;
  assign n53721 = n38215 ^ n12064 ^ 1'b0 ;
  assign n53722 = n15413 & ~n53721 ;
  assign n53723 = n53722 ^ n1598 ^ 1'b0 ;
  assign n53724 = n38509 | n53723 ;
  assign n53725 = ~n53720 & n53724 ;
  assign n53726 = n16961 ^ n4439 ^ n2112 ;
  assign n53727 = ( ~n47005 & n47076 ) | ( ~n47005 & n53726 ) | ( n47076 & n53726 ) ;
  assign n53728 = ( n2962 & n9655 ) | ( n2962 & ~n14817 ) | ( n9655 & ~n14817 ) ;
  assign n53729 = n16031 ^ n13210 ^ n6988 ;
  assign n53730 = ( n2859 & n23756 ) | ( n2859 & n53729 ) | ( n23756 & n53729 ) ;
  assign n53731 = ( ~n7153 & n10562 ) | ( ~n7153 & n53730 ) | ( n10562 & n53730 ) ;
  assign n53732 = n53731 ^ n39411 ^ n3533 ;
  assign n53733 = n33582 ^ n16500 ^ n15909 ;
  assign n53734 = n53733 ^ n8363 ^ n6634 ;
  assign n53735 = n21283 & ~n53734 ;
  assign n53736 = ( ~n37163 & n37739 ) | ( ~n37163 & n43082 ) | ( n37739 & n43082 ) ;
  assign n53737 = n22346 ^ n20353 ^ n12891 ;
  assign n53738 = n13566 & ~n53737 ;
  assign n53739 = n53738 ^ n16441 ^ n14150 ;
  assign n53743 = ( ~n6643 & n9063 ) | ( ~n6643 & n22339 ) | ( n9063 & n22339 ) ;
  assign n53744 = n53743 ^ n18175 ^ n4104 ;
  assign n53740 = ~n11983 & n52939 ;
  assign n53741 = n53740 ^ n35631 ^ 1'b0 ;
  assign n53742 = n53741 ^ n26363 ^ n25204 ;
  assign n53745 = n53744 ^ n53742 ^ 1'b0 ;
  assign n53746 = n51759 ^ n46557 ^ n29995 ;
  assign n53747 = n4339 & n53746 ;
  assign n53748 = ~n53745 & n53747 ;
  assign n53749 = ~n750 & n28401 ;
  assign n53750 = ( n1619 & n30780 ) | ( n1619 & ~n43564 ) | ( n30780 & ~n43564 ) ;
  assign n53751 = ( n24581 & n25496 ) | ( n24581 & ~n42340 ) | ( n25496 & ~n42340 ) ;
  assign n53752 = ( n35477 & n36774 ) | ( n35477 & n53751 ) | ( n36774 & n53751 ) ;
  assign n53753 = n21872 & ~n22413 ;
  assign n53754 = n53753 ^ n29385 ^ 1'b0 ;
  assign n53755 = n46591 ^ n26280 ^ n25900 ;
  assign n53757 = ( n4151 & ~n23325 ) | ( n4151 & n39435 ) | ( ~n23325 & n39435 ) ;
  assign n53756 = n33089 ^ n12448 ^ n10592 ;
  assign n53758 = n53757 ^ n53756 ^ n47350 ;
  assign n53763 = n45822 ^ n4739 ^ n722 ;
  assign n53764 = ( n14997 & n17054 ) | ( n14997 & ~n53763 ) | ( n17054 & ~n53763 ) ;
  assign n53762 = n2448 & n8862 ;
  assign n53765 = n53764 ^ n53762 ^ 1'b0 ;
  assign n53759 = n12170 & n40516 ;
  assign n53760 = n53759 ^ n24527 ^ 1'b0 ;
  assign n53761 = ( n10907 & n20964 ) | ( n10907 & n53760 ) | ( n20964 & n53760 ) ;
  assign n53766 = n53765 ^ n53761 ^ n36536 ;
  assign n53767 = ( n17892 & n29404 ) | ( n17892 & ~n35432 ) | ( n29404 & ~n35432 ) ;
  assign n53768 = ( n45386 & n48302 ) | ( n45386 & n53767 ) | ( n48302 & n53767 ) ;
  assign n53769 = ( ~n25941 & n30518 ) | ( ~n25941 & n53768 ) | ( n30518 & n53768 ) ;
  assign n53770 = ( n47129 & ~n47171 ) | ( n47129 & n48633 ) | ( ~n47171 & n48633 ) ;
  assign n53771 = n3406 & ~n6959 ;
  assign n53772 = n53771 ^ n13201 ^ n11081 ;
  assign n53773 = ( n12958 & n31250 ) | ( n12958 & ~n39904 ) | ( n31250 & ~n39904 ) ;
  assign n53774 = ( n1120 & ~n11683 ) | ( n1120 & n15728 ) | ( ~n11683 & n15728 ) ;
  assign n53775 = n53774 ^ n51184 ^ n27703 ;
  assign n53776 = ( n11617 & n23909 ) | ( n11617 & n53775 ) | ( n23909 & n53775 ) ;
  assign n53777 = n40959 ^ n23487 ^ n3878 ;
  assign n53778 = n31293 ^ n13863 ^ n2713 ;
  assign n53779 = ( ~n2569 & n42066 ) | ( ~n2569 & n42502 ) | ( n42066 & n42502 ) ;
  assign n53780 = n44621 ^ n35492 ^ n1211 ;
  assign n53781 = ( n6178 & ~n30986 ) | ( n6178 & n53780 ) | ( ~n30986 & n53780 ) ;
  assign n53782 = ~n1581 & n33671 ;
  assign n53783 = n53782 ^ n38861 ^ n19840 ;
  assign n53784 = n53783 ^ n49695 ^ n12170 ;
  assign n53785 = n8905 ^ n5693 ^ 1'b0 ;
  assign n53786 = ~n11724 & n53785 ;
  assign n53789 = n2806 | n10158 ;
  assign n53790 = n5457 & ~n53789 ;
  assign n53787 = n28276 ^ n24752 ^ n18895 ;
  assign n53788 = n53787 ^ n19566 ^ n1746 ;
  assign n53791 = n53790 ^ n53788 ^ n19631 ;
  assign n53792 = ( n22661 & n31191 ) | ( n22661 & ~n35340 ) | ( n31191 & ~n35340 ) ;
  assign n53793 = ~n3184 & n18803 ;
  assign n53794 = ~n12858 & n53793 ;
  assign n53795 = n53794 ^ n32305 ^ n22965 ;
  assign n53796 = n31141 ^ n29904 ^ n17853 ;
  assign n53797 = ( n21691 & n37832 ) | ( n21691 & n53796 ) | ( n37832 & n53796 ) ;
  assign n53798 = ( n20160 & n42640 ) | ( n20160 & n51501 ) | ( n42640 & n51501 ) ;
  assign n53799 = ( n38671 & n51919 ) | ( n38671 & ~n53798 ) | ( n51919 & ~n53798 ) ;
  assign n53804 = n17831 ^ n5173 ^ 1'b0 ;
  assign n53805 = n5073 & n53804 ;
  assign n53801 = n36459 ^ n29085 ^ n12220 ;
  assign n53802 = n36982 ^ n15963 ^ 1'b0 ;
  assign n53803 = n53801 & n53802 ;
  assign n53800 = n5774 & ~n25928 ;
  assign n53806 = n53805 ^ n53803 ^ n53800 ;
  assign n53807 = n53806 ^ n16717 ^ n11021 ;
  assign n53808 = n468 | n47699 ;
  assign n53809 = n29814 & ~n53808 ;
  assign n53810 = n53809 ^ n39493 ^ 1'b0 ;
  assign n53811 = n33159 ^ n19991 ^ n4321 ;
  assign n53812 = ( n17611 & n22987 ) | ( n17611 & n33270 ) | ( n22987 & n33270 ) ;
  assign n53813 = n48085 ^ n10551 ^ 1'b0 ;
  assign n53814 = ~n11708 & n17187 ;
  assign n53815 = n299 & n53814 ;
  assign n53816 = ( n14505 & n20468 ) | ( n14505 & ~n31583 ) | ( n20468 & ~n31583 ) ;
  assign n53817 = n33644 ^ n25565 ^ n24116 ;
  assign n53818 = n53817 ^ n20316 ^ n3843 ;
  assign n53819 = ( ~n9355 & n53816 ) | ( ~n9355 & n53818 ) | ( n53816 & n53818 ) ;
  assign n53821 = ( n8758 & n48568 ) | ( n8758 & ~n53451 ) | ( n48568 & ~n53451 ) ;
  assign n53820 = ( ~n15452 & n21690 ) | ( ~n15452 & n51046 ) | ( n21690 & n51046 ) ;
  assign n53822 = n53821 ^ n53820 ^ n7494 ;
  assign n53823 = ( n5368 & ~n35431 ) | ( n5368 & n46818 ) | ( ~n35431 & n46818 ) ;
  assign n53824 = ( ~n18252 & n31021 ) | ( ~n18252 & n53823 ) | ( n31021 & n53823 ) ;
  assign n53825 = ( ~n25897 & n45117 ) | ( ~n25897 & n53824 ) | ( n45117 & n53824 ) ;
  assign n53826 = ( n2344 & n17718 ) | ( n2344 & ~n44628 ) | ( n17718 & ~n44628 ) ;
  assign n53827 = n53578 ^ n14195 ^ n1124 ;
  assign n53828 = n53827 ^ n45500 ^ n17478 ;
  assign n53829 = n40866 ^ n24487 ^ n8811 ;
  assign n53830 = ( ~n12638 & n23207 ) | ( ~n12638 & n53829 ) | ( n23207 & n53829 ) ;
  assign n53831 = n34914 ^ n14510 ^ n4551 ;
  assign n53832 = n26966 ^ n22081 ^ n20707 ;
  assign n53833 = ( ~n25389 & n33297 ) | ( ~n25389 & n53832 ) | ( n33297 & n53832 ) ;
  assign n53834 = ( ~n24958 & n47695 ) | ( ~n24958 & n53833 ) | ( n47695 & n53833 ) ;
  assign n53835 = n26639 ^ n23243 ^ n3577 ;
  assign n53836 = n5476 | n53835 ;
  assign n53837 = n17985 | n53836 ;
  assign n53838 = ( n19414 & n29841 ) | ( n19414 & ~n31231 ) | ( n29841 & ~n31231 ) ;
  assign n53839 = ( n493 & ~n14811 ) | ( n493 & n28804 ) | ( ~n14811 & n28804 ) ;
  assign n53840 = n53839 ^ n6588 ^ 1'b0 ;
  assign n53841 = ( n25481 & n46076 ) | ( n25481 & ~n53840 ) | ( n46076 & ~n53840 ) ;
  assign n53842 = n53841 ^ n10400 ^ 1'b0 ;
  assign n53849 = ( n9777 & n29656 ) | ( n9777 & n39178 ) | ( n29656 & n39178 ) ;
  assign n53843 = ( n4426 & ~n27456 ) | ( n4426 & n43337 ) | ( ~n27456 & n43337 ) ;
  assign n53844 = n53843 ^ n39703 ^ n30511 ;
  assign n53845 = n53844 ^ n24753 ^ n2453 ;
  assign n53846 = n53845 ^ n12638 ^ n1869 ;
  assign n53847 = ( n7080 & n8134 ) | ( n7080 & ~n53846 ) | ( n8134 & ~n53846 ) ;
  assign n53848 = n53847 ^ n33051 ^ n1225 ;
  assign n53850 = n53849 ^ n53848 ^ n23588 ;
  assign n53851 = n53850 ^ n19173 ^ n4743 ;
  assign n53852 = ~n14764 & n17201 ;
  assign n53853 = n53852 ^ n23999 ^ 1'b0 ;
  assign n53854 = ( n7297 & ~n51043 ) | ( n7297 & n53853 ) | ( ~n51043 & n53853 ) ;
  assign n53855 = n45761 ^ n10651 ^ 1'b0 ;
  assign n53856 = ~n14048 & n53855 ;
  assign n53857 = ( ~n16505 & n36646 ) | ( ~n16505 & n53856 ) | ( n36646 & n53856 ) ;
  assign n53858 = ( n16309 & n28616 ) | ( n16309 & ~n53857 ) | ( n28616 & ~n53857 ) ;
  assign n53859 = n19716 ^ n3175 ^ 1'b0 ;
  assign n53860 = ( n19181 & n33935 ) | ( n19181 & ~n50189 ) | ( n33935 & ~n50189 ) ;
  assign n53861 = ( n14984 & ~n22297 ) | ( n14984 & n40255 ) | ( ~n22297 & n40255 ) ;
  assign n53862 = n50581 ^ n36372 ^ n34928 ;
  assign n53863 = n17116 & ~n33438 ;
  assign n53864 = n39179 & n53863 ;
  assign n53865 = n8196 & ~n13556 ;
  assign n53866 = n30200 & n53865 ;
  assign n53867 = n4806 ^ n1318 ^ 1'b0 ;
  assign n53868 = n53866 | n53867 ;
  assign n53869 = n39962 & ~n43943 ;
  assign n53870 = n31251 & n53869 ;
  assign n53871 = n35702 ^ n19358 ^ n12403 ;
  assign n53872 = n53871 ^ n44958 ^ n16545 ;
  assign n53873 = ( n9781 & n19356 ) | ( n9781 & n21993 ) | ( n19356 & n21993 ) ;
  assign n53874 = n47608 ^ n22517 ^ n1566 ;
  assign n53875 = n53874 ^ n28290 ^ n26103 ;
  assign n53876 = ( n21508 & n53873 ) | ( n21508 & ~n53875 ) | ( n53873 & ~n53875 ) ;
  assign n53877 = ( n47138 & n53872 ) | ( n47138 & ~n53876 ) | ( n53872 & ~n53876 ) ;
  assign n53878 = ( n52669 & ~n53870 ) | ( n52669 & n53877 ) | ( ~n53870 & n53877 ) ;
  assign n53879 = n11854 & n20809 ;
  assign n53880 = n29731 ^ n12165 ^ n1732 ;
  assign n53881 = ( n7378 & ~n25101 ) | ( n7378 & n53880 ) | ( ~n25101 & n53880 ) ;
  assign n53882 = ( n10475 & ~n47436 ) | ( n10475 & n53881 ) | ( ~n47436 & n53881 ) ;
  assign n53883 = ( n4043 & ~n7685 ) | ( n4043 & n14491 ) | ( ~n7685 & n14491 ) ;
  assign n53884 = n20283 | n53883 ;
  assign n53885 = n10399 & ~n53884 ;
  assign n53886 = n53885 ^ n49862 ^ n4470 ;
  assign n53888 = n30428 ^ n27522 ^ n10682 ;
  assign n53887 = ( n2936 & n15088 ) | ( n2936 & ~n50175 ) | ( n15088 & ~n50175 ) ;
  assign n53889 = n53888 ^ n53887 ^ n6880 ;
  assign n53890 = ( n40326 & n53886 ) | ( n40326 & n53889 ) | ( n53886 & n53889 ) ;
  assign n53891 = n37425 ^ n19231 ^ n534 ;
  assign n53892 = n38925 ^ n38201 ^ n16712 ;
  assign n53893 = n53892 ^ n20503 ^ n14380 ;
  assign n53894 = n53893 ^ n43305 ^ n39453 ;
  assign n53895 = n13260 & n21522 ;
  assign n53896 = n53895 ^ n50355 ^ n12361 ;
  assign n53897 = n53148 ^ n21679 ^ 1'b0 ;
  assign n53898 = n53897 ^ n37534 ^ 1'b0 ;
  assign n53899 = ( n18802 & n24562 ) | ( n18802 & ~n26333 ) | ( n24562 & ~n26333 ) ;
  assign n53900 = n43432 ^ n20911 ^ n9521 ;
  assign n53901 = n8075 | n53900 ;
  assign n53902 = n53899 | n53901 ;
  assign n53903 = n38240 ^ n18742 ^ n4578 ;
  assign n53907 = n41133 ^ n29835 ^ n3358 ;
  assign n53908 = n53907 ^ n42378 ^ n1759 ;
  assign n53904 = n44156 ^ n30494 ^ n7045 ;
  assign n53905 = ( n1246 & n18173 ) | ( n1246 & ~n53904 ) | ( n18173 & ~n53904 ) ;
  assign n53906 = n53905 ^ n46920 ^ n43336 ;
  assign n53909 = n53908 ^ n53906 ^ 1'b0 ;
  assign n53910 = n23258 ^ n12223 ^ n11385 ;
  assign n53911 = n19886 & n53910 ;
  assign n53912 = ( ~n5072 & n25779 ) | ( ~n5072 & n34205 ) | ( n25779 & n34205 ) ;
  assign n53913 = n20380 ^ x11 ^ 1'b0 ;
  assign n53914 = n53913 ^ n49722 ^ n15940 ;
  assign n53915 = n21013 ^ n5376 ^ n3760 ;
  assign n53916 = n7655 & n53915 ;
  assign n53917 = ( ~n8620 & n17951 ) | ( ~n8620 & n28641 ) | ( n17951 & n28641 ) ;
  assign n53918 = ( ~n16293 & n36275 ) | ( ~n16293 & n53917 ) | ( n36275 & n53917 ) ;
  assign n53919 = ( n459 & n1518 ) | ( n459 & ~n53918 ) | ( n1518 & ~n53918 ) ;
  assign n53920 = n53328 ^ n47432 ^ n20495 ;
  assign n53921 = n6484 & n14940 ;
  assign n53922 = n53921 ^ n43770 ^ n37104 ;
  assign n53923 = n28417 & n49574 ;
  assign n53924 = n9174 & n53923 ;
  assign n53925 = n34841 | n35165 ;
  assign n53926 = n53925 ^ n31317 ^ n12948 ;
  assign n53927 = ( n1103 & n14784 ) | ( n1103 & ~n51581 ) | ( n14784 & ~n51581 ) ;
  assign n53928 = ( n7449 & ~n22515 ) | ( n7449 & n26278 ) | ( ~n22515 & n26278 ) ;
  assign n53929 = n53928 ^ n36260 ^ 1'b0 ;
  assign n53930 = ( n29520 & n53927 ) | ( n29520 & n53929 ) | ( n53927 & n53929 ) ;
  assign n53931 = n51107 ^ n47451 ^ n6528 ;
  assign n53932 = ( n12322 & n12676 ) | ( n12322 & ~n53931 ) | ( n12676 & ~n53931 ) ;
  assign n53933 = n39999 ^ n28254 ^ n24779 ;
  assign n53934 = ( n1969 & n33622 ) | ( n1969 & n53933 ) | ( n33622 & n53933 ) ;
  assign n53935 = n24289 & ~n36911 ;
  assign n53936 = ~n8543 & n53935 ;
  assign n53937 = ( n31728 & n47920 ) | ( n31728 & ~n53936 ) | ( n47920 & ~n53936 ) ;
  assign n53938 = ( n2611 & n10509 ) | ( n2611 & ~n26414 ) | ( n10509 & ~n26414 ) ;
  assign n53939 = n28897 ^ n12045 ^ n10774 ;
  assign n53940 = ( n22171 & ~n39986 ) | ( n22171 & n53939 ) | ( ~n39986 & n53939 ) ;
  assign n53941 = n53940 ^ n29817 ^ n28472 ;
  assign n53942 = n19478 | n40148 ;
  assign n53943 = n53942 ^ n36758 ^ n2533 ;
  assign n53944 = n53943 ^ n24634 ^ 1'b0 ;
  assign n53945 = n30519 & ~n53597 ;
  assign n53946 = n53945 ^ n5528 ^ 1'b0 ;
  assign n53947 = ( n7692 & n12698 ) | ( n7692 & ~n31457 ) | ( n12698 & ~n31457 ) ;
  assign n53948 = n32347 ^ n9289 ^ n414 ;
  assign n53949 = ( ~n27876 & n37738 ) | ( ~n27876 & n53948 ) | ( n37738 & n53948 ) ;
  assign n53950 = ( n5859 & n29449 ) | ( n5859 & n53949 ) | ( n29449 & n53949 ) ;
  assign n53951 = ( n39233 & ~n39668 ) | ( n39233 & n47701 ) | ( ~n39668 & n47701 ) ;
  assign n53952 = ( n15410 & ~n33302 ) | ( n15410 & n53951 ) | ( ~n33302 & n53951 ) ;
  assign n53953 = ( n23238 & ~n26044 ) | ( n23238 & n34223 ) | ( ~n26044 & n34223 ) ;
  assign n53954 = ( n3045 & ~n5194 ) | ( n3045 & n5435 ) | ( ~n5194 & n5435 ) ;
  assign n53955 = ( ~n5196 & n6296 ) | ( ~n5196 & n22602 ) | ( n6296 & n22602 ) ;
  assign n53956 = n53955 ^ n16846 ^ n5231 ;
  assign n53957 = ( n22211 & n53954 ) | ( n22211 & ~n53956 ) | ( n53954 & ~n53956 ) ;
  assign n53958 = n53957 ^ n37955 ^ n14745 ;
  assign n53959 = n7776 & n19213 ;
  assign n53960 = n32547 ^ n9000 ^ n7599 ;
  assign n53961 = n53960 ^ n36018 ^ n14909 ;
  assign n53962 = n42326 ^ n24422 ^ n1614 ;
  assign n53963 = n8203 | n20849 ;
  assign n53964 = n26729 | n53963 ;
  assign n53965 = ~n1477 & n52919 ;
  assign n53966 = n53965 ^ n20859 ^ 1'b0 ;
  assign n53967 = ( x61 & n21672 ) | ( x61 & ~n29323 ) | ( n21672 & ~n29323 ) ;
  assign n53968 = n53967 ^ n31256 ^ n22214 ;
  assign n53969 = n50264 ^ n40331 ^ n476 ;
  assign n53970 = ( ~n2349 & n35494 ) | ( ~n2349 & n53969 ) | ( n35494 & n53969 ) ;
  assign n53973 = ( n3150 & ~n4661 ) | ( n3150 & n8947 ) | ( ~n4661 & n8947 ) ;
  assign n53971 = n35986 ^ n35264 ^ n12722 ;
  assign n53972 = n53971 ^ n20505 ^ n7882 ;
  assign n53974 = n53973 ^ n53972 ^ n7598 ;
  assign n53975 = n18531 | n34284 ;
  assign n53976 = ~n52575 & n53975 ;
  assign n53977 = ( n14275 & n16528 ) | ( n14275 & ~n53976 ) | ( n16528 & ~n53976 ) ;
  assign n53978 = ( ~n2899 & n15513 ) | ( ~n2899 & n31173 ) | ( n15513 & n31173 ) ;
  assign n53979 = n23780 ^ n23250 ^ x244 ;
  assign n53980 = ( n19075 & n37456 ) | ( n19075 & n53979 ) | ( n37456 & n53979 ) ;
  assign n53981 = ( n7794 & n22844 ) | ( n7794 & ~n53767 ) | ( n22844 & ~n53767 ) ;
  assign n53982 = n14042 ^ n7260 ^ 1'b0 ;
  assign n53983 = n53982 ^ n27761 ^ n14949 ;
  assign n53984 = n34015 & n53983 ;
  assign n53985 = ( ~n24141 & n25119 ) | ( ~n24141 & n53907 ) | ( n25119 & n53907 ) ;
  assign n53986 = ( n26267 & n41019 ) | ( n26267 & n53985 ) | ( n41019 & n53985 ) ;
  assign n53988 = n22754 ^ n22417 ^ n1058 ;
  assign n53987 = ~n15926 & n17876 ;
  assign n53989 = n53988 ^ n53987 ^ 1'b0 ;
  assign n53990 = n1031 | n7683 ;
  assign n53991 = n53990 ^ n3866 ^ 1'b0 ;
  assign n53992 = n53991 ^ n8233 ^ 1'b0 ;
  assign n53993 = ( n1434 & n11873 ) | ( n1434 & n43787 ) | ( n11873 & n43787 ) ;
  assign n53994 = ( n13067 & n32524 ) | ( n13067 & ~n33858 ) | ( n32524 & ~n33858 ) ;
  assign n53995 = ( n1824 & ~n23505 ) | ( n1824 & n53994 ) | ( ~n23505 & n53994 ) ;
  assign n53996 = n53995 ^ n43926 ^ n7694 ;
  assign n53999 = ( n31886 & n35828 ) | ( n31886 & ~n35918 ) | ( n35828 & ~n35918 ) ;
  assign n53997 = ( ~x40 & n3393 ) | ( ~x40 & n24442 ) | ( n3393 & n24442 ) ;
  assign n53998 = n53997 ^ n48031 ^ 1'b0 ;
  assign n54000 = n53999 ^ n53998 ^ n19193 ;
  assign n54002 = n12836 ^ n10069 ^ n5647 ;
  assign n54001 = ( n9683 & n11231 ) | ( n9683 & ~n13538 ) | ( n11231 & ~n13538 ) ;
  assign n54003 = n54002 ^ n54001 ^ n12344 ;
  assign n54004 = n54003 ^ n42435 ^ n4474 ;
  assign n54005 = n46697 ^ n8710 ^ n8709 ;
  assign n54006 = ( ~n4025 & n23384 ) | ( ~n4025 & n26959 ) | ( n23384 & n26959 ) ;
  assign n54007 = n22772 ^ n11898 ^ n6880 ;
  assign n54008 = n54007 ^ n53847 ^ n42991 ;
  assign n54009 = n54008 ^ n16190 ^ n8457 ;
  assign n54010 = ( n4988 & n54006 ) | ( n4988 & ~n54009 ) | ( n54006 & ~n54009 ) ;
  assign n54011 = n54010 ^ n8179 ^ n4140 ;
  assign n54012 = ( n8714 & ~n16411 ) | ( n8714 & n26695 ) | ( ~n16411 & n26695 ) ;
  assign n54013 = ( n28523 & n53200 ) | ( n28523 & n54012 ) | ( n53200 & n54012 ) ;
  assign n54014 = n44135 ^ n38934 ^ n2867 ;
  assign n54015 = n23708 ^ n1797 ^ 1'b0 ;
  assign n54017 = ( ~n482 & n1783 ) | ( ~n482 & n11315 ) | ( n1783 & n11315 ) ;
  assign n54018 = ( n26330 & n42976 ) | ( n26330 & n54017 ) | ( n42976 & n54017 ) ;
  assign n54016 = n23936 & ~n44675 ;
  assign n54019 = n54018 ^ n54016 ^ 1'b0 ;
  assign n54020 = n560 & ~n40114 ;
  assign n54021 = ~n51771 & n54020 ;
  assign n54022 = ( n26963 & ~n27169 ) | ( n26963 & n28278 ) | ( ~n27169 & n28278 ) ;
  assign n54023 = ~n5489 & n54022 ;
  assign n54024 = ( n17327 & ~n17868 ) | ( n17327 & n38598 ) | ( ~n17868 & n38598 ) ;
  assign n54028 = n14275 | n31157 ;
  assign n54029 = n54028 ^ n33826 ^ 1'b0 ;
  assign n54026 = ( ~n3403 & n9516 ) | ( ~n3403 & n35485 ) | ( n9516 & n35485 ) ;
  assign n54025 = ( n8121 & n13432 ) | ( n8121 & ~n30628 ) | ( n13432 & ~n30628 ) ;
  assign n54027 = n54026 ^ n54025 ^ n15144 ;
  assign n54030 = n54029 ^ n54027 ^ n4088 ;
  assign n54031 = n938 & n1350 ;
  assign n54033 = ( n3656 & ~n16028 ) | ( n3656 & n29090 ) | ( ~n16028 & n29090 ) ;
  assign n54032 = ( n15856 & n28987 ) | ( n15856 & ~n49909 ) | ( n28987 & ~n49909 ) ;
  assign n54034 = n54033 ^ n54032 ^ n23851 ;
  assign n54035 = n54034 ^ n50795 ^ n19104 ;
  assign n54036 = n51160 ^ n44825 ^ n5064 ;
  assign n54037 = ( n21250 & n31317 ) | ( n21250 & ~n54036 ) | ( n31317 & ~n54036 ) ;
  assign n54038 = ( n922 & ~n6116 ) | ( n922 & n10910 ) | ( ~n6116 & n10910 ) ;
  assign n54039 = ( n35967 & n40270 ) | ( n35967 & n54038 ) | ( n40270 & n54038 ) ;
  assign n54040 = n54039 ^ n33774 ^ n13661 ;
  assign n54041 = n40105 ^ n4998 ^ n852 ;
  assign n54042 = n20887 ^ n10959 ^ n8735 ;
  assign n54043 = n774 | n37363 ;
  assign n54044 = n24833 & ~n54043 ;
  assign n54046 = ~n30508 & n43684 ;
  assign n54047 = n39907 & n54046 ;
  assign n54045 = ~n5177 & n25595 ;
  assign n54048 = n54047 ^ n54045 ^ 1'b0 ;
  assign n54049 = n36704 ^ n36136 ^ x221 ;
  assign n54050 = n54049 ^ n29619 ^ n29062 ;
  assign n54051 = ( n4739 & ~n51488 ) | ( n4739 & n54050 ) | ( ~n51488 & n54050 ) ;
  assign n54052 = n51018 ^ n20548 ^ n9024 ;
  assign n54053 = n52429 ^ n24093 ^ n15880 ;
  assign n54054 = ( n26435 & ~n40944 ) | ( n26435 & n44640 ) | ( ~n40944 & n44640 ) ;
  assign n54055 = n54054 ^ n47438 ^ n45081 ;
  assign n54056 = ( n1222 & ~n3568 ) | ( n1222 & n6902 ) | ( ~n3568 & n6902 ) ;
  assign n54057 = n14589 ^ n10399 ^ n937 ;
  assign n54058 = ( n3796 & n54056 ) | ( n3796 & n54057 ) | ( n54056 & n54057 ) ;
  assign n54059 = n31198 ^ n7567 ^ n3495 ;
  assign n54060 = n54059 ^ n23071 ^ n2495 ;
  assign n54061 = ~n3306 & n44844 ;
  assign n54062 = ~n6448 & n40449 ;
  assign n54063 = n6602 & n54062 ;
  assign n54064 = ( n4826 & n19876 ) | ( n4826 & ~n26473 ) | ( n19876 & ~n26473 ) ;
  assign n54065 = n54064 ^ n15918 ^ 1'b0 ;
  assign n54066 = n36171 & ~n54065 ;
  assign n54067 = ( ~n11506 & n17667 ) | ( ~n11506 & n25617 ) | ( n17667 & n25617 ) ;
  assign n54068 = n18329 & n47432 ;
  assign n54069 = ( n5224 & n45906 ) | ( n5224 & n54068 ) | ( n45906 & n54068 ) ;
  assign n54070 = ( ~n12621 & n21782 ) | ( ~n12621 & n30367 ) | ( n21782 & n30367 ) ;
  assign n54071 = n39682 ^ n14455 ^ n3155 ;
  assign n54072 = n54071 ^ n27090 ^ n5131 ;
  assign n54073 = n31398 ^ n7019 ^ n3276 ;
  assign n54074 = ( n16499 & n31011 ) | ( n16499 & n54073 ) | ( n31011 & n54073 ) ;
  assign n54077 = n38137 | n40243 ;
  assign n54075 = n550 & ~n38988 ;
  assign n54076 = n10005 & n54075 ;
  assign n54078 = n54077 ^ n54076 ^ n37243 ;
  assign n54079 = ~n3402 & n49212 ;
  assign n54080 = n54079 ^ n53667 ^ 1'b0 ;
  assign n54081 = n15128 & ~n17020 ;
  assign n54082 = ( n22319 & n23228 ) | ( n22319 & n53982 ) | ( n23228 & n53982 ) ;
  assign n54083 = n54082 ^ n26867 ^ n6655 ;
  assign n54084 = ( ~n32055 & n54081 ) | ( ~n32055 & n54083 ) | ( n54081 & n54083 ) ;
  assign n54085 = ( n26475 & n34887 ) | ( n26475 & ~n47521 ) | ( n34887 & ~n47521 ) ;
  assign n54086 = n52234 ^ n31088 ^ n17882 ;
  assign n54087 = n54086 ^ n31191 ^ 1'b0 ;
  assign n54088 = n23184 ^ n10420 ^ n3994 ;
  assign n54089 = n54088 ^ n26542 ^ n4191 ;
  assign n54090 = ( n3711 & n52970 ) | ( n3711 & ~n54089 ) | ( n52970 & ~n54089 ) ;
  assign n54091 = ( n27408 & n44474 ) | ( n27408 & ~n49401 ) | ( n44474 & ~n49401 ) ;
  assign n54092 = n53460 ^ n35787 ^ n21136 ;
  assign n54093 = n54092 ^ n38059 ^ n10249 ;
  assign n54094 = n34483 ^ n14049 ^ n4949 ;
  assign n54095 = ( n6157 & ~n20973 ) | ( n6157 & n32052 ) | ( ~n20973 & n32052 ) ;
  assign n54096 = ( n32575 & n53823 ) | ( n32575 & ~n54095 ) | ( n53823 & ~n54095 ) ;
  assign n54097 = n35527 ^ n19198 ^ 1'b0 ;
  assign n54098 = n28832 ^ n19004 ^ n460 ;
  assign n54099 = n54098 ^ n21958 ^ n5780 ;
  assign n54100 = n54099 ^ n9503 ^ 1'b0 ;
  assign n54101 = n40383 & n54100 ;
  assign n54102 = n31551 ^ n24740 ^ n4083 ;
  assign n54103 = n54102 ^ n742 ^ 1'b0 ;
  assign n54104 = ~n44816 & n54103 ;
  assign n54105 = ( n14477 & n34544 ) | ( n14477 & n40367 ) | ( n34544 & n40367 ) ;
  assign n54106 = ( n5944 & n32384 ) | ( n5944 & ~n53611 ) | ( n32384 & ~n53611 ) ;
  assign n54107 = ( n8810 & n13212 ) | ( n8810 & ~n16322 ) | ( n13212 & ~n16322 ) ;
  assign n54108 = n54107 ^ n53056 ^ n35777 ;
  assign n54111 = ( n7897 & n31204 ) | ( n7897 & n48109 ) | ( n31204 & n48109 ) ;
  assign n54109 = ~n11769 & n17353 ;
  assign n54110 = n54109 ^ n17644 ^ n11276 ;
  assign n54112 = n54111 ^ n54110 ^ n9580 ;
  assign n54113 = ( n12807 & n43410 ) | ( n12807 & n54112 ) | ( n43410 & n54112 ) ;
  assign n54114 = ( n14429 & n20414 ) | ( n14429 & n29242 ) | ( n20414 & n29242 ) ;
  assign n54115 = ( n2377 & n12468 ) | ( n2377 & ~n37845 ) | ( n12468 & ~n37845 ) ;
  assign n54116 = ( n3152 & n16528 ) | ( n3152 & n38430 ) | ( n16528 & n38430 ) ;
  assign n54117 = ( ~n13147 & n21919 ) | ( ~n13147 & n47897 ) | ( n21919 & n47897 ) ;
  assign n54118 = ( n1859 & n11664 ) | ( n1859 & ~n28024 ) | ( n11664 & ~n28024 ) ;
  assign n54119 = ( n21129 & ~n46308 ) | ( n21129 & n54118 ) | ( ~n46308 & n54118 ) ;
  assign n54120 = n32077 ^ n12530 ^ 1'b0 ;
  assign n54121 = n6595 | n54120 ;
  assign n54122 = n1691 | n54121 ;
  assign n54123 = n54122 ^ n53598 ^ 1'b0 ;
  assign n54124 = n30500 ^ n18673 ^ n1899 ;
  assign n54125 = n27738 ^ n3011 ^ x251 ;
  assign n54126 = ( n11124 & n25842 ) | ( n11124 & ~n54125 ) | ( n25842 & ~n54125 ) ;
  assign n54127 = ( ~n5848 & n54124 ) | ( ~n5848 & n54126 ) | ( n54124 & n54126 ) ;
  assign n54128 = ( n21523 & ~n30411 ) | ( n21523 & n39525 ) | ( ~n30411 & n39525 ) ;
  assign n54129 = ( ~n26934 & n27363 ) | ( ~n26934 & n49350 ) | ( n27363 & n49350 ) ;
  assign n54130 = n40738 ^ n21659 ^ n3405 ;
  assign n54131 = n52575 ^ n31987 ^ n30024 ;
  assign n54132 = ~n25258 & n54131 ;
  assign n54133 = n11413 ^ n3138 ^ x83 ;
  assign n54135 = n32234 ^ n16434 ^ n7590 ;
  assign n54134 = n2093 & ~n32232 ;
  assign n54136 = n54135 ^ n54134 ^ 1'b0 ;
  assign n54137 = ( n36425 & n45520 ) | ( n36425 & n54136 ) | ( n45520 & n54136 ) ;
  assign n54140 = ( n862 & n2204 ) | ( n862 & n8147 ) | ( n2204 & n8147 ) ;
  assign n54138 = n25975 | n46874 ;
  assign n54139 = n27366 | n54138 ;
  assign n54141 = n54140 ^ n54139 ^ n12644 ;
  assign n54142 = n54141 ^ n51612 ^ n46850 ;
  assign n54143 = ~n5523 & n20111 ;
  assign n54144 = n54143 ^ n6256 ^ 1'b0 ;
  assign n54145 = n8219 | n53301 ;
  assign n54146 = n49707 & ~n54145 ;
  assign n54147 = n34141 ^ n24557 ^ n16332 ;
  assign n54148 = ( n6790 & n12818 ) | ( n6790 & n41148 ) | ( n12818 & n41148 ) ;
  assign n54149 = n604 | n54148 ;
  assign n54150 = n43721 & ~n54149 ;
  assign n54151 = n54150 ^ n46840 ^ n43799 ;
  assign n54152 = n22082 ^ n18595 ^ n14356 ;
  assign n54153 = n54152 ^ n48998 ^ n9781 ;
  assign n54158 = n15503 ^ n3176 ^ n739 ;
  assign n54159 = ( n5002 & n45277 ) | ( n5002 & ~n54158 ) | ( n45277 & ~n54158 ) ;
  assign n54157 = ( ~n4495 & n23615 ) | ( ~n4495 & n32881 ) | ( n23615 & n32881 ) ;
  assign n54154 = ( ~n5687 & n5700 ) | ( ~n5687 & n9805 ) | ( n5700 & n9805 ) ;
  assign n54155 = n53337 ^ n37726 ^ n5774 ;
  assign n54156 = ( n41030 & ~n54154 ) | ( n41030 & n54155 ) | ( ~n54154 & n54155 ) ;
  assign n54160 = n54159 ^ n54157 ^ n54156 ;
  assign n54162 = n8023 & n23964 ;
  assign n54163 = n54162 ^ n10756 ^ 1'b0 ;
  assign n54164 = n54163 ^ n22852 ^ n18064 ;
  assign n54165 = ( n12489 & ~n47489 ) | ( n12489 & n54164 ) | ( ~n47489 & n54164 ) ;
  assign n54161 = ( n7288 & n17301 ) | ( n7288 & n31198 ) | ( n17301 & n31198 ) ;
  assign n54166 = n54165 ^ n54161 ^ n17727 ;
  assign n54167 = ( n3205 & n4689 ) | ( n3205 & n47991 ) | ( n4689 & n47991 ) ;
  assign n54168 = n38930 ^ n38816 ^ n28770 ;
  assign n54169 = ( n42746 & ~n47345 ) | ( n42746 & n49899 ) | ( ~n47345 & n49899 ) ;
  assign n54170 = ( ~n7339 & n13470 ) | ( ~n7339 & n19919 ) | ( n13470 & n19919 ) ;
  assign n54171 = ~n3439 & n32237 ;
  assign n54172 = n15506 & n54171 ;
  assign n54173 = n33440 ^ n4849 ^ 1'b0 ;
  assign n54174 = ~n41813 & n54173 ;
  assign n54175 = ( n1371 & ~n15003 ) | ( n1371 & n30033 ) | ( ~n15003 & n30033 ) ;
  assign n54176 = n39294 & n42921 ;
  assign n54177 = n54176 ^ n1598 ^ 1'b0 ;
  assign n54178 = ( n35929 & n54175 ) | ( n35929 & ~n54177 ) | ( n54175 & ~n54177 ) ;
  assign n54179 = ~n14443 & n42373 ;
  assign n54180 = n54179 ^ n28654 ^ 1'b0 ;
  assign n54181 = ( ~n11239 & n14633 ) | ( ~n11239 & n54180 ) | ( n14633 & n54180 ) ;
  assign n54182 = ( ~n4811 & n25824 ) | ( ~n4811 & n27206 ) | ( n25824 & n27206 ) ;
  assign n54183 = ( n21242 & ~n33089 ) | ( n21242 & n54182 ) | ( ~n33089 & n54182 ) ;
  assign n54184 = n54183 ^ n36239 ^ n2334 ;
  assign n54185 = n29596 ^ n18973 ^ 1'b0 ;
  assign n54186 = ( n5678 & ~n11688 ) | ( n5678 & n33628 ) | ( ~n11688 & n33628 ) ;
  assign n54187 = ( n7358 & ~n38344 ) | ( n7358 & n54186 ) | ( ~n38344 & n54186 ) ;
  assign n54188 = n19827 ^ n9233 ^ n7696 ;
  assign n54189 = ( n21055 & n25687 ) | ( n21055 & n48922 ) | ( n25687 & n48922 ) ;
  assign n54190 = n3457 | n28952 ;
  assign n54191 = n54190 ^ n8126 ^ n6398 ;
  assign n54192 = n52124 ^ n39408 ^ n33539 ;
  assign n54193 = n37305 ^ n17357 ^ 1'b0 ;
  assign n54194 = ~n30956 & n54193 ;
  assign n54195 = n18252 ^ n16815 ^ n4444 ;
  assign n54196 = n49961 ^ n28036 ^ n6595 ;
  assign n54197 = n54195 & n54196 ;
  assign n54198 = n54197 ^ n32961 ^ 1'b0 ;
  assign n54199 = ( n9617 & n14509 ) | ( n9617 & ~n25497 ) | ( n14509 & ~n25497 ) ;
  assign n54200 = n30733 & ~n35383 ;
  assign n54201 = ( n1622 & n11074 ) | ( n1622 & ~n31224 ) | ( n11074 & ~n31224 ) ;
  assign n54202 = n54201 ^ n27298 ^ n8302 ;
  assign n54203 = ( n13639 & n24733 ) | ( n13639 & n54202 ) | ( n24733 & n54202 ) ;
  assign n54205 = ( n1540 & n17135 ) | ( n1540 & n24517 ) | ( n17135 & n24517 ) ;
  assign n54204 = n37513 ^ n37328 ^ n25237 ;
  assign n54206 = n54205 ^ n54204 ^ n38872 ;
  assign n54207 = n19423 ^ n7945 ^ 1'b0 ;
  assign n54208 = n47134 | n54207 ;
  assign n54209 = n12060 ^ n7889 ^ n2351 ;
  assign n54210 = n47608 ^ n45789 ^ n41895 ;
  assign n54211 = ( n35967 & ~n42803 ) | ( n35967 & n54210 ) | ( ~n42803 & n54210 ) ;
  assign n54212 = n13669 & ~n54211 ;
  assign n54213 = n54212 ^ n11079 ^ n1594 ;
  assign n54214 = ( n54208 & n54209 ) | ( n54208 & n54213 ) | ( n54209 & n54213 ) ;
  assign n54215 = ( n990 & n4769 ) | ( n990 & ~n5056 ) | ( n4769 & ~n5056 ) ;
  assign n54216 = n54215 ^ n28322 ^ 1'b0 ;
  assign n54217 = n20341 & n54216 ;
  assign n54218 = ( n20808 & n46159 ) | ( n20808 & ~n54217 ) | ( n46159 & ~n54217 ) ;
  assign n54219 = n25323 & ~n33738 ;
  assign n54220 = n43446 ^ n43401 ^ 1'b0 ;
  assign n54221 = n3786 & n54220 ;
  assign n54222 = n54221 ^ n46427 ^ n40255 ;
  assign n54223 = ( n7499 & n13645 ) | ( n7499 & ~n38051 ) | ( n13645 & ~n38051 ) ;
  assign n54224 = n29593 & n37110 ;
  assign n54225 = ~n5515 & n54224 ;
  assign n54226 = n21038 | n54225 ;
  assign n54227 = n19747 & ~n54226 ;
  assign n54228 = n27230 ^ n19956 ^ n14635 ;
  assign n54229 = ( ~n1498 & n24734 ) | ( ~n1498 & n54228 ) | ( n24734 & n54228 ) ;
  assign n54237 = n9864 & ~n24332 ;
  assign n54230 = ( n3730 & n20788 ) | ( n3730 & n36917 ) | ( n20788 & n36917 ) ;
  assign n54234 = n35062 ^ n4052 ^ n1613 ;
  assign n54231 = n33559 ^ n13487 ^ 1'b0 ;
  assign n54232 = ( ~n11197 & n16473 ) | ( ~n11197 & n26343 ) | ( n16473 & n26343 ) ;
  assign n54233 = ( n27992 & n54231 ) | ( n27992 & ~n54232 ) | ( n54231 & ~n54232 ) ;
  assign n54235 = n54234 ^ n54233 ^ n35735 ;
  assign n54236 = ( n21316 & ~n54230 ) | ( n21316 & n54235 ) | ( ~n54230 & n54235 ) ;
  assign n54238 = n54237 ^ n54236 ^ n11037 ;
  assign n54239 = n19749 | n21717 ;
  assign n54240 = n39040 ^ n20652 ^ n17814 ;
  assign n54241 = ( n5576 & n37120 ) | ( n5576 & n47444 ) | ( n37120 & n47444 ) ;
  assign n54242 = n54240 | n54241 ;
  assign n54243 = n9455 ^ n372 ^ 1'b0 ;
  assign n54244 = n49345 | n54243 ;
  assign n54245 = ( n40750 & n54242 ) | ( n40750 & n54244 ) | ( n54242 & n54244 ) ;
  assign n54246 = n3396 & n9511 ;
  assign n54247 = n54246 ^ n44968 ^ n35929 ;
  assign n54248 = n31678 | n54247 ;
  assign n54249 = n29820 | n54248 ;
  assign n54250 = n54249 ^ n25956 ^ n15270 ;
  assign n54251 = n37468 ^ n14705 ^ 1'b0 ;
  assign n54252 = ( n47463 & n49529 ) | ( n47463 & ~n50103 ) | ( n49529 & ~n50103 ) ;
  assign n54253 = n10841 ^ n1868 ^ n273 ;
  assign n54254 = n41380 ^ n5163 ^ 1'b0 ;
  assign n54255 = n14400 & n45427 ;
  assign n54256 = n22330 ^ n19527 ^ 1'b0 ;
  assign n54257 = n3307 & n54256 ;
  assign n54258 = n54257 ^ n35520 ^ 1'b0 ;
  assign n54259 = ( ~n14313 & n17565 ) | ( ~n14313 & n50201 ) | ( n17565 & n50201 ) ;
  assign n54260 = n54259 ^ n36381 ^ n16967 ;
  assign n54261 = n11474 ^ n8580 ^ n4660 ;
  assign n54262 = n54261 ^ n23202 ^ n18485 ;
  assign n54263 = n17204 & ~n23748 ;
  assign n54264 = ~n38733 & n54263 ;
  assign n54265 = n54264 ^ n37320 ^ n16011 ;
  assign n54266 = n651 & n32704 ;
  assign n54267 = n54266 ^ n53832 ^ 1'b0 ;
  assign n54268 = n54267 ^ n41836 ^ n14748 ;
  assign n54269 = n30887 ^ n9192 ^ n6570 ;
  assign n54270 = n25253 ^ n9992 ^ 1'b0 ;
  assign n54271 = n54270 ^ n33841 ^ n2201 ;
  assign n54272 = n50625 ^ n18411 ^ n10837 ;
  assign n54273 = ( n1217 & n47989 ) | ( n1217 & n54272 ) | ( n47989 & n54272 ) ;
  assign n54274 = ~n11598 & n14668 ;
  assign n54275 = n6684 & n54274 ;
  assign n54276 = n17807 | n54275 ;
  assign n54277 = n30986 ^ n29123 ^ n15886 ;
  assign n54278 = ( ~n5938 & n31794 ) | ( ~n5938 & n54277 ) | ( n31794 & n54277 ) ;
  assign n54279 = ( n4831 & ~n5910 ) | ( n4831 & n52218 ) | ( ~n5910 & n52218 ) ;
  assign n54280 = n46733 ^ n5633 ^ n5605 ;
  assign n54281 = n40808 ^ n9219 ^ n3585 ;
  assign n54282 = n19111 ^ n11989 ^ n3126 ;
  assign n54283 = n2067 & n34279 ;
  assign n54284 = ( n11098 & ~n43198 ) | ( n11098 & n46371 ) | ( ~n43198 & n46371 ) ;
  assign n54285 = ( ~n32407 & n52885 ) | ( ~n32407 & n54284 ) | ( n52885 & n54284 ) ;
  assign n54286 = ( ~n11347 & n18296 ) | ( ~n11347 & n33460 ) | ( n18296 & n33460 ) ;
  assign n54287 = ( n296 & n49242 ) | ( n296 & ~n50399 ) | ( n49242 & ~n50399 ) ;
  assign n54288 = ( n14743 & ~n17974 ) | ( n14743 & n54287 ) | ( ~n17974 & n54287 ) ;
  assign n54289 = n31959 ^ n17225 ^ 1'b0 ;
  assign n54290 = ~n22603 & n54289 ;
  assign n54291 = n20014 | n43372 ;
  assign n54292 = n16468 ^ n8475 ^ n6709 ;
  assign n54293 = n36304 ^ n19950 ^ n3899 ;
  assign n54294 = n10602 | n54293 ;
  assign n54295 = ( n12198 & n54292 ) | ( n12198 & ~n54294 ) | ( n54292 & ~n54294 ) ;
  assign n54296 = ( ~n3331 & n9481 ) | ( ~n3331 & n54295 ) | ( n9481 & n54295 ) ;
  assign n54297 = ( n9508 & ~n43472 ) | ( n9508 & n49688 ) | ( ~n43472 & n49688 ) ;
  assign n54298 = ~n10127 & n32667 ;
  assign n54299 = ~n31639 & n54298 ;
  assign n54300 = ( n29240 & ~n36397 ) | ( n29240 & n54299 ) | ( ~n36397 & n54299 ) ;
  assign n54301 = ( n3983 & ~n16494 ) | ( n3983 & n49118 ) | ( ~n16494 & n49118 ) ;
  assign n54302 = n54301 ^ n48532 ^ 1'b0 ;
  assign n54303 = n46140 ^ n12154 ^ n4212 ;
  assign n54304 = ( n8434 & ~n13708 ) | ( n8434 & n54303 ) | ( ~n13708 & n54303 ) ;
  assign n54305 = ( n20537 & n43999 ) | ( n20537 & ~n54304 ) | ( n43999 & ~n54304 ) ;
  assign n54306 = ( n16718 & ~n29541 ) | ( n16718 & n39008 ) | ( ~n29541 & n39008 ) ;
  assign n54307 = n42883 ^ n22347 ^ n11617 ;
  assign n54308 = ( ~n8563 & n35111 ) | ( ~n8563 & n54307 ) | ( n35111 & n54307 ) ;
  assign n54309 = ( n11980 & ~n26298 ) | ( n11980 & n54308 ) | ( ~n26298 & n54308 ) ;
  assign n54310 = ( n32488 & n36352 ) | ( n32488 & n54309 ) | ( n36352 & n54309 ) ;
  assign n54311 = n52122 ^ n35256 ^ n31799 ;
  assign n54312 = n54311 ^ n43443 ^ n27338 ;
  assign n54313 = n54312 ^ n30364 ^ n29090 ;
  assign n54314 = ( n5843 & n15894 ) | ( n5843 & ~n27593 ) | ( n15894 & ~n27593 ) ;
  assign n54315 = n41735 ^ n6649 ^ 1'b0 ;
  assign n54316 = n40616 & ~n54315 ;
  assign n54317 = ( n2405 & n21393 ) | ( n2405 & ~n52931 ) | ( n21393 & ~n52931 ) ;
  assign n54318 = n22007 ^ n12238 ^ n1078 ;
  assign n54319 = ( n16935 & ~n21089 ) | ( n16935 & n28965 ) | ( ~n21089 & n28965 ) ;
  assign n54320 = n54319 ^ n37881 ^ n8246 ;
  assign n54321 = n54320 ^ n18926 ^ n5358 ;
  assign n54322 = n47616 ^ n39432 ^ n13861 ;
  assign n54323 = n36106 ^ n10140 ^ n1397 ;
  assign n54324 = n54092 ^ n48289 ^ n23047 ;
  assign n54325 = n33042 ^ n31822 ^ n17620 ;
  assign n54326 = ( n3153 & n4009 ) | ( n3153 & ~n14973 ) | ( n4009 & ~n14973 ) ;
  assign n54327 = n31382 ^ n17306 ^ 1'b0 ;
  assign n54328 = n4757 & ~n54327 ;
  assign n54329 = n27850 ^ n22954 ^ n16178 ;
  assign n54330 = ~n17483 & n54068 ;
  assign n54331 = ( n6241 & n54329 ) | ( n6241 & ~n54330 ) | ( n54329 & ~n54330 ) ;
  assign n54332 = n51418 ^ n37770 ^ 1'b0 ;
  assign n54333 = ( n25532 & ~n26758 ) | ( n25532 & n28180 ) | ( ~n26758 & n28180 ) ;
  assign n54334 = n31027 ^ n15270 ^ n1181 ;
  assign n54335 = n54334 ^ n26773 ^ n19545 ;
  assign n54336 = n25621 ^ n13661 ^ n12203 ;
  assign n54341 = ( ~n409 & n9778 ) | ( ~n409 & n12386 ) | ( n9778 & n12386 ) ;
  assign n54337 = n11901 & n33315 ;
  assign n54338 = ~n31625 & n54337 ;
  assign n54339 = ( n6701 & n38160 ) | ( n6701 & ~n54338 ) | ( n38160 & ~n54338 ) ;
  assign n54340 = ( n25580 & n26610 ) | ( n25580 & n54339 ) | ( n26610 & n54339 ) ;
  assign n54342 = n54341 ^ n54340 ^ n9588 ;
  assign n54343 = ( n10307 & ~n54336 ) | ( n10307 & n54342 ) | ( ~n54336 & n54342 ) ;
  assign n54344 = ( n2990 & ~n20978 ) | ( n2990 & n53633 ) | ( ~n20978 & n53633 ) ;
  assign n54345 = n54344 ^ n24791 ^ x127 ;
  assign n54346 = n6594 & ~n15940 ;
  assign n54347 = n54346 ^ n3509 ^ 1'b0 ;
  assign n54348 = n54347 ^ n36286 ^ n27397 ;
  assign n54349 = ( n27320 & ~n41661 ) | ( n27320 & n51349 ) | ( ~n41661 & n51349 ) ;
  assign n54350 = ( n5096 & n7910 ) | ( n5096 & ~n31144 ) | ( n7910 & ~n31144 ) ;
  assign n54351 = ( ~n12139 & n46007 ) | ( ~n12139 & n54350 ) | ( n46007 & n54350 ) ;
  assign n54352 = n2623 & ~n18815 ;
  assign n54353 = n54352 ^ n2927 ^ 1'b0 ;
  assign n54354 = n27687 ^ n27595 ^ n15805 ;
  assign n54355 = ~n51493 & n54354 ;
  assign n54356 = ~n1134 & n9564 ;
  assign n54357 = n17576 & n54356 ;
  assign n54358 = ( n6127 & n18473 ) | ( n6127 & n30503 ) | ( n18473 & n30503 ) ;
  assign n54359 = ( n16826 & n54357 ) | ( n16826 & ~n54358 ) | ( n54357 & ~n54358 ) ;
  assign n54360 = n54359 ^ n11749 ^ n7849 ;
  assign n54361 = n54360 ^ n48727 ^ n6802 ;
  assign n54362 = ( n13555 & n47804 ) | ( n13555 & n54361 ) | ( n47804 & n54361 ) ;
  assign n54363 = n13221 ^ n1309 ^ 1'b0 ;
  assign n54364 = n2615 & ~n54363 ;
  assign n54365 = ( n45866 & n54362 ) | ( n45866 & ~n54364 ) | ( n54362 & ~n54364 ) ;
  assign n54366 = ( ~n20206 & n25326 ) | ( ~n20206 & n37773 ) | ( n25326 & n37773 ) ;
  assign n54367 = n44924 ^ n10431 ^ n3930 ;
  assign n54368 = n50092 ^ n2633 ^ n578 ;
  assign n54369 = ( n1188 & n30204 ) | ( n1188 & n41723 ) | ( n30204 & n41723 ) ;
  assign n54370 = ( n2974 & ~n12985 ) | ( n2974 & n54369 ) | ( ~n12985 & n54369 ) ;
  assign n54371 = n54370 ^ n14152 ^ n4098 ;
  assign n54372 = ( ~n7723 & n13446 ) | ( ~n7723 & n30120 ) | ( n13446 & n30120 ) ;
  assign n54373 = n43670 ^ n41737 ^ n5242 ;
  assign n54374 = ( n13071 & n13564 ) | ( n13071 & ~n37921 ) | ( n13564 & ~n37921 ) ;
  assign n54375 = ( ~n54372 & n54373 ) | ( ~n54372 & n54374 ) | ( n54373 & n54374 ) ;
  assign n54376 = n22017 ^ n13822 ^ n2897 ;
  assign n54377 = n21486 ^ n18181 ^ n10268 ;
  assign n54378 = ( n11035 & ~n54376 ) | ( n11035 & n54377 ) | ( ~n54376 & n54377 ) ;
  assign n54379 = n46116 ^ n46115 ^ n17731 ;
  assign n54380 = ( ~n30590 & n37354 ) | ( ~n30590 & n54379 ) | ( n37354 & n54379 ) ;
  assign n54381 = n30117 ^ n22754 ^ n5826 ;
  assign n54382 = ( ~n11442 & n33446 ) | ( ~n11442 & n54381 ) | ( n33446 & n54381 ) ;
  assign n54384 = n39736 ^ n3614 ^ n1612 ;
  assign n54383 = ~n17526 & n22887 ;
  assign n54385 = n54384 ^ n54383 ^ 1'b0 ;
  assign n54386 = n54385 ^ n51961 ^ 1'b0 ;
  assign n54387 = n30729 | n54386 ;
  assign n54388 = n53848 ^ n40952 ^ n40772 ;
  assign n54389 = ( n355 & n9643 ) | ( n355 & n48833 ) | ( n9643 & n48833 ) ;
  assign n54390 = ( ~n13809 & n42167 ) | ( ~n13809 & n54389 ) | ( n42167 & n54389 ) ;
  assign n54391 = ( x65 & n24391 ) | ( x65 & n25164 ) | ( n24391 & n25164 ) ;
  assign n54392 = n54391 ^ n49135 ^ n4357 ;
  assign n54393 = ( n2870 & ~n5520 ) | ( n2870 & n32004 ) | ( ~n5520 & n32004 ) ;
  assign n54394 = n54393 ^ n14836 ^ n7088 ;
  assign n54395 = n8265 & ~n54394 ;
  assign n54396 = ( n17822 & n27510 ) | ( n17822 & n54395 ) | ( n27510 & n54395 ) ;
  assign n54397 = n54396 ^ n47690 ^ 1'b0 ;
  assign n54398 = ( n17838 & n21656 ) | ( n17838 & n25180 ) | ( n21656 & n25180 ) ;
  assign n54399 = n54398 ^ n13551 ^ 1'b0 ;
  assign n54400 = n54399 ^ n36306 ^ n25496 ;
  assign n54401 = n46129 ^ n45157 ^ 1'b0 ;
  assign n54402 = n14707 ^ n5719 ^ n2080 ;
  assign n54403 = ( n3591 & ~n16455 ) | ( n3591 & n36610 ) | ( ~n16455 & n36610 ) ;
  assign n54404 = n54403 ^ n50907 ^ n17381 ;
  assign n54405 = n50079 ^ n31190 ^ n30349 ;
  assign n54406 = n9651 | n16851 ;
  assign n54407 = n15963 & ~n54406 ;
  assign n54408 = ( n13345 & ~n41709 ) | ( n13345 & n42859 ) | ( ~n41709 & n42859 ) ;
  assign n54409 = n42888 ^ n28409 ^ n3442 ;
  assign n54410 = ( n17476 & n33524 ) | ( n17476 & ~n54341 ) | ( n33524 & ~n54341 ) ;
  assign n54411 = n8093 & n8910 ;
  assign n54412 = n54411 ^ n42490 ^ n9560 ;
  assign n54413 = n54412 ^ n26788 ^ n8054 ;
  assign n54414 = ( n5008 & n29176 ) | ( n5008 & n48701 ) | ( n29176 & n48701 ) ;
  assign n54415 = n47337 ^ n13763 ^ n10615 ;
  assign n54416 = ( n23542 & ~n54414 ) | ( n23542 & n54415 ) | ( ~n54414 & n54415 ) ;
  assign n54417 = n54416 ^ n50315 ^ n4802 ;
  assign n54418 = n48454 ^ n26674 ^ n25543 ;
  assign n54419 = ~n5036 & n24693 ;
  assign n54420 = ( n6654 & ~n17826 ) | ( n6654 & n18854 ) | ( ~n17826 & n18854 ) ;
  assign n54421 = ( ~n4058 & n16157 ) | ( ~n4058 & n31510 ) | ( n16157 & n31510 ) ;
  assign n54422 = n33037 ^ n18326 ^ n12913 ;
  assign n54423 = ( n15265 & n32717 ) | ( n15265 & n54422 ) | ( n32717 & n54422 ) ;
  assign n54424 = ( n28984 & n54421 ) | ( n28984 & ~n54423 ) | ( n54421 & ~n54423 ) ;
  assign n54425 = ( n27032 & ~n46391 ) | ( n27032 & n54424 ) | ( ~n46391 & n54424 ) ;
  assign n54427 = n8143 & n30459 ;
  assign n54426 = n7191 | n21996 ;
  assign n54428 = n54427 ^ n54426 ^ 1'b0 ;
  assign n54429 = n38578 ^ n30606 ^ n2453 ;
  assign n54430 = ( n8238 & ~n9022 ) | ( n8238 & n22708 ) | ( ~n9022 & n22708 ) ;
  assign n54431 = n16166 & n54430 ;
  assign n54432 = n54431 ^ n28726 ^ 1'b0 ;
  assign n54433 = n37750 ^ n26155 ^ n10829 ;
  assign n54434 = ( n13851 & n54432 ) | ( n13851 & n54433 ) | ( n54432 & n54433 ) ;
  assign n54435 = n54434 ^ n12990 ^ n10707 ;
  assign n54436 = ( ~n2039 & n6023 ) | ( ~n2039 & n9778 ) | ( n6023 & n9778 ) ;
  assign n54437 = n39463 | n40145 ;
  assign n54438 = n18982 ^ n11985 ^ n3969 ;
  assign n54439 = n54438 ^ n15553 ^ n421 ;
  assign n54440 = ( n7288 & ~n45597 ) | ( n7288 & n54439 ) | ( ~n45597 & n54439 ) ;
  assign n54441 = ( n923 & n42891 ) | ( n923 & ~n54440 ) | ( n42891 & ~n54440 ) ;
  assign n54442 = n15177 ^ n7916 ^ n2071 ;
  assign n54443 = n54442 ^ n8515 ^ 1'b0 ;
  assign n54444 = ( n17612 & ~n35967 ) | ( n17612 & n49078 ) | ( ~n35967 & n49078 ) ;
  assign n54445 = n5078 | n28721 ;
  assign n54446 = n54445 ^ n53513 ^ n4830 ;
  assign n54447 = ( n14705 & n20466 ) | ( n14705 & ~n44510 ) | ( n20466 & ~n44510 ) ;
  assign n54448 = n2475 & ~n10759 ;
  assign n54449 = ~n50775 & n54448 ;
  assign n54450 = n53783 ^ n53340 ^ n3183 ;
  assign n54451 = n34182 ^ n476 ^ 1'b0 ;
  assign n54452 = ( n1337 & ~n14046 ) | ( n1337 & n54451 ) | ( ~n14046 & n54451 ) ;
  assign n54453 = ( n10147 & ~n54450 ) | ( n10147 & n54452 ) | ( ~n54450 & n54452 ) ;
  assign n54454 = ( n20662 & ~n34454 ) | ( n20662 & n34798 ) | ( ~n34454 & n34798 ) ;
  assign n54455 = n54454 ^ n50374 ^ n16712 ;
  assign n54456 = n22037 ^ n16562 ^ n9997 ;
  assign n54457 = ( n1208 & n10824 ) | ( n1208 & n28684 ) | ( n10824 & n28684 ) ;
  assign n54458 = ( n8666 & n12830 ) | ( n8666 & n35534 ) | ( n12830 & n35534 ) ;
  assign n54459 = ( n4105 & ~n54457 ) | ( n4105 & n54458 ) | ( ~n54457 & n54458 ) ;
  assign n54460 = ( n8935 & n14819 ) | ( n8935 & ~n37443 ) | ( n14819 & ~n37443 ) ;
  assign n54461 = n53451 ^ n44048 ^ n28442 ;
  assign n54462 = ( n17817 & ~n48784 ) | ( n17817 & n54461 ) | ( ~n48784 & n54461 ) ;
  assign n54463 = ( ~n6405 & n10241 ) | ( ~n6405 & n54026 ) | ( n10241 & n54026 ) ;
  assign n54464 = n23708 ^ n17660 ^ n1687 ;
  assign n54465 = ( n19483 & ~n54463 ) | ( n19483 & n54464 ) | ( ~n54463 & n54464 ) ;
  assign n54466 = n48777 ^ n10181 ^ n607 ;
  assign n54467 = ( n7750 & n13448 ) | ( n7750 & n24606 ) | ( n13448 & n24606 ) ;
  assign n54468 = ( n6303 & ~n13600 ) | ( n6303 & n54467 ) | ( ~n13600 & n54467 ) ;
  assign n54469 = n36082 ^ n17302 ^ n10615 ;
  assign n54470 = ( n18856 & n33115 ) | ( n18856 & n54469 ) | ( n33115 & n54469 ) ;
  assign n54471 = n34380 ^ n32530 ^ n14738 ;
  assign n54472 = n26360 ^ n21478 ^ n2739 ;
  assign n54473 = n2147 | n17749 ;
  assign n54474 = n17542 & ~n24730 ;
  assign n54475 = n54474 ^ n8346 ^ 1'b0 ;
  assign n54476 = n54475 ^ n37224 ^ n4129 ;
  assign n54477 = x27 & n54476 ;
  assign n54478 = x212 & n28431 ;
  assign n54479 = n54478 ^ n20082 ^ n18412 ;
  assign n54481 = ( n9848 & n13400 ) | ( n9848 & ~n25390 ) | ( n13400 & ~n25390 ) ;
  assign n54480 = n36384 ^ n10558 ^ n8912 ;
  assign n54482 = n54481 ^ n54480 ^ 1'b0 ;
  assign n54483 = ( n4370 & n5769 ) | ( n4370 & n28286 ) | ( n5769 & n28286 ) ;
  assign n54484 = n33326 ^ n14061 ^ 1'b0 ;
  assign n54485 = n18000 | n45072 ;
  assign n54486 = n54485 ^ n28442 ^ 1'b0 ;
  assign n54488 = ( n565 & n2220 ) | ( n565 & n19964 ) | ( n2220 & n19964 ) ;
  assign n54489 = ~n11178 & n54488 ;
  assign n54490 = n40092 & n54489 ;
  assign n54491 = ( n20922 & ~n38026 ) | ( n20922 & n54490 ) | ( ~n38026 & n54490 ) ;
  assign n54492 = n54491 ^ n12152 ^ n5714 ;
  assign n54487 = ( n11906 & n12954 ) | ( n11906 & ~n13026 ) | ( n12954 & ~n13026 ) ;
  assign n54493 = n54492 ^ n54487 ^ n13583 ;
  assign n54494 = n43684 ^ n23268 ^ n20572 ;
  assign n54495 = n35286 ^ n23178 ^ n3210 ;
  assign n54496 = ( n13630 & ~n27191 ) | ( n13630 & n52885 ) | ( ~n27191 & n52885 ) ;
  assign n54497 = n52421 ^ n16019 ^ n5369 ;
  assign n54498 = ( n17432 & ~n35528 ) | ( n17432 & n45847 ) | ( ~n35528 & n45847 ) ;
  assign n54499 = ( n6088 & n44350 ) | ( n6088 & n54498 ) | ( n44350 & n54498 ) ;
  assign n54500 = n42557 ^ n32190 ^ n17408 ;
  assign n54501 = ~n40338 & n44021 ;
  assign n54502 = ( n49133 & n51349 ) | ( n49133 & ~n54501 ) | ( n51349 & ~n54501 ) ;
  assign n54503 = n11001 ^ n9451 ^ n8482 ;
  assign n54504 = n43954 ^ n32640 ^ n23888 ;
  assign n54505 = ~n47796 & n54504 ;
  assign n54506 = ( n14187 & ~n54503 ) | ( n14187 & n54505 ) | ( ~n54503 & n54505 ) ;
  assign n54507 = ( n13434 & ~n41626 ) | ( n13434 & n53345 ) | ( ~n41626 & n53345 ) ;
  assign n54508 = n43823 ^ n36450 ^ n20160 ;
  assign n54509 = n54508 ^ n20246 ^ 1'b0 ;
  assign n54510 = ~n54507 & n54509 ;
  assign n54511 = n46384 ^ n44749 ^ n11524 ;
  assign n54512 = ( n19793 & n26344 ) | ( n19793 & n29937 ) | ( n26344 & n29937 ) ;
  assign n54514 = n32606 ^ n8808 ^ n5422 ;
  assign n54513 = n40824 ^ n34366 ^ n15037 ;
  assign n54515 = n54514 ^ n54513 ^ n46790 ;
  assign n54518 = n14320 ^ n14162 ^ n5670 ;
  assign n54516 = ( n8554 & ~n13147 ) | ( n8554 & n23245 ) | ( ~n13147 & n23245 ) ;
  assign n54517 = n54516 ^ n49496 ^ n28799 ;
  assign n54519 = n54518 ^ n54517 ^ n8273 ;
  assign n54520 = n3675 & n46743 ;
  assign n54521 = n54520 ^ n11559 ^ n10788 ;
  assign n54522 = n22118 ^ n9965 ^ 1'b0 ;
  assign n54523 = ( n13857 & ~n41308 ) | ( n13857 & n54522 ) | ( ~n41308 & n54522 ) ;
  assign n54524 = ( n3585 & ~n23564 ) | ( n3585 & n26828 ) | ( ~n23564 & n26828 ) ;
  assign n54525 = ( n15391 & ~n38301 ) | ( n15391 & n54524 ) | ( ~n38301 & n54524 ) ;
  assign n54526 = n54241 ^ n27863 ^ n4789 ;
  assign n54527 = n50869 ^ n23720 ^ n7755 ;
  assign n54528 = ~n13046 & n34098 ;
  assign n54529 = n54528 ^ n48175 ^ 1'b0 ;
  assign n54530 = ( n1634 & n7265 ) | ( n1634 & n28283 ) | ( n7265 & n28283 ) ;
  assign n54531 = n10758 ^ n8815 ^ n4990 ;
  assign n54532 = ( n7719 & n54530 ) | ( n7719 & ~n54531 ) | ( n54530 & ~n54531 ) ;
  assign n54533 = n46266 ^ n45950 ^ n23419 ;
  assign n54534 = n54533 ^ n35397 ^ 1'b0 ;
  assign n54535 = n54532 & ~n54534 ;
  assign n54536 = n48910 ^ n18429 ^ n8153 ;
  assign n54537 = n54536 ^ n46221 ^ n6951 ;
  assign n54538 = ( ~n2937 & n6885 ) | ( ~n2937 & n29893 ) | ( n6885 & n29893 ) ;
  assign n54539 = ( n18060 & ~n30378 ) | ( n18060 & n54538 ) | ( ~n30378 & n54538 ) ;
  assign n54540 = ( n2616 & n4681 ) | ( n2616 & n37276 ) | ( n4681 & n37276 ) ;
  assign n54541 = ( n1811 & n54539 ) | ( n1811 & ~n54540 ) | ( n54539 & ~n54540 ) ;
  assign n54542 = n42597 ^ n20399 ^ n15502 ;
  assign n54543 = ( ~n17780 & n42616 ) | ( ~n17780 & n54542 ) | ( n42616 & n54542 ) ;
  assign n54544 = n54543 ^ n36779 ^ n9238 ;
  assign n54545 = ( n7287 & n14265 ) | ( n7287 & n16717 ) | ( n14265 & n16717 ) ;
  assign n54546 = ( n4105 & n8787 ) | ( n4105 & ~n26407 ) | ( n8787 & ~n26407 ) ;
  assign n54547 = n54546 ^ n26713 ^ n20635 ;
  assign n54548 = ( n54131 & n54545 ) | ( n54131 & n54547 ) | ( n54545 & n54547 ) ;
  assign n54549 = n54548 ^ n19631 ^ n19249 ;
  assign n54550 = ( ~n8521 & n31851 ) | ( ~n8521 & n35702 ) | ( n31851 & n35702 ) ;
  assign n54553 = n20316 ^ n10432 ^ n3475 ;
  assign n54552 = ( n9942 & n23426 ) | ( n9942 & ~n47641 ) | ( n23426 & ~n47641 ) ;
  assign n54551 = ( n9654 & n15410 ) | ( n9654 & ~n26815 ) | ( n15410 & ~n26815 ) ;
  assign n54554 = n54553 ^ n54552 ^ n54551 ;
  assign n54556 = n14712 ^ n5001 ^ n1667 ;
  assign n54555 = ( n3022 & n12995 ) | ( n3022 & ~n26102 ) | ( n12995 & ~n26102 ) ;
  assign n54557 = n54556 ^ n54555 ^ n33461 ;
  assign n54558 = n14253 ^ n12383 ^ 1'b0 ;
  assign n54559 = n23140 ^ n5763 ^ 1'b0 ;
  assign n54560 = n14560 ^ n14398 ^ 1'b0 ;
  assign n54561 = n54560 ^ n48171 ^ 1'b0 ;
  assign n54563 = n41820 ^ n30665 ^ n13393 ;
  assign n54562 = n31802 ^ n2681 ^ 1'b0 ;
  assign n54564 = n54563 ^ n54562 ^ n38463 ;
  assign n54565 = ( n15220 & n25179 ) | ( n15220 & ~n38709 ) | ( n25179 & ~n38709 ) ;
  assign n54566 = n5977 ^ n360 ^ 1'b0 ;
  assign n54567 = n54565 & ~n54566 ;
  assign n54568 = ( ~n8917 & n54564 ) | ( ~n8917 & n54567 ) | ( n54564 & n54567 ) ;
  assign n54569 = ( n26501 & ~n41013 ) | ( n26501 & n53998 ) | ( ~n41013 & n53998 ) ;
  assign n54570 = n43926 ^ n14332 ^ n5926 ;
  assign n54571 = ( n6540 & n20928 ) | ( n6540 & ~n54570 ) | ( n20928 & ~n54570 ) ;
  assign n54572 = n45961 ^ n716 ^ 1'b0 ;
  assign n54573 = n54572 ^ n8922 ^ n6821 ;
  assign n54574 = n49472 ^ n30827 ^ n289 ;
  assign n54575 = ( n20778 & n26684 ) | ( n20778 & n42580 ) | ( n26684 & n42580 ) ;
  assign n54576 = ( n1410 & n11554 ) | ( n1410 & ~n14566 ) | ( n11554 & ~n14566 ) ;
  assign n54577 = n19783 ^ n9479 ^ n1970 ;
  assign n54578 = n54577 ^ n44786 ^ n38068 ;
  assign n54579 = n8179 & n15798 ;
  assign n54580 = n54579 ^ n9771 ^ 1'b0 ;
  assign n54581 = n54580 ^ n17383 ^ n5122 ;
  assign n54583 = n22966 ^ n17808 ^ n12553 ;
  assign n54582 = ( n1997 & n11654 ) | ( n1997 & n44417 ) | ( n11654 & n44417 ) ;
  assign n54584 = n54583 ^ n54582 ^ n31434 ;
  assign n54585 = n46973 ^ n17707 ^ n5923 ;
  assign n54586 = ( ~n18014 & n18127 ) | ( ~n18014 & n47491 ) | ( n18127 & n47491 ) ;
  assign n54587 = n54586 ^ n33614 ^ 1'b0 ;
  assign n54588 = n37532 ^ n37020 ^ n21854 ;
  assign n54589 = n20585 ^ n2053 ^ n939 ;
  assign n54590 = n2493 & n20990 ;
  assign n54591 = n54589 & n54590 ;
  assign n54592 = ( ~n11488 & n32163 ) | ( ~n11488 & n54591 ) | ( n32163 & n54591 ) ;
  assign n54593 = n20697 ^ x66 ^ 1'b0 ;
  assign n54594 = ( ~n27053 & n37555 ) | ( ~n27053 & n53733 ) | ( n37555 & n53733 ) ;
  assign n54595 = ( n54592 & n54593 ) | ( n54592 & n54594 ) | ( n54593 & n54594 ) ;
  assign n54596 = n32463 ^ n5850 ^ n1833 ;
  assign n54597 = n54596 ^ n39537 ^ n2469 ;
  assign n54598 = ( n2702 & ~n7824 ) | ( n2702 & n24390 ) | ( ~n7824 & n24390 ) ;
  assign n54599 = ~n14643 & n23841 ;
  assign n54600 = n54599 ^ n33193 ^ 1'b0 ;
  assign n54601 = n20409 & n54600 ;
  assign n54602 = ( n6173 & n13059 ) | ( n6173 & ~n13304 ) | ( n13059 & ~n13304 ) ;
  assign n54603 = n41497 ^ n25937 ^ 1'b0 ;
  assign n54604 = n54602 & n54603 ;
  assign n54605 = n54307 ^ n40655 ^ n30797 ;
  assign n54606 = ( n17522 & n29730 ) | ( n17522 & n35153 ) | ( n29730 & n35153 ) ;
  assign n54607 = n32250 ^ n16228 ^ n15205 ;
  assign n54608 = ( ~n1078 & n18990 ) | ( ~n1078 & n54607 ) | ( n18990 & n54607 ) ;
  assign n54609 = ( ~n638 & n54606 ) | ( ~n638 & n54608 ) | ( n54606 & n54608 ) ;
  assign n54610 = n34659 ^ n10837 ^ n9369 ;
  assign n54611 = n54610 ^ n38534 ^ n3363 ;
  assign n54612 = n46448 & n54611 ;
  assign n54614 = ( n10491 & ~n21390 ) | ( n10491 & n27711 ) | ( ~n21390 & n27711 ) ;
  assign n54613 = ~n5601 & n23905 ;
  assign n54615 = n54614 ^ n54613 ^ 1'b0 ;
  assign n54616 = ~n2466 & n54615 ;
  assign n54617 = n54616 ^ n32328 ^ 1'b0 ;
  assign n54618 = n52123 ^ n17765 ^ n12676 ;
  assign n54619 = ( n2451 & n54617 ) | ( n2451 & ~n54618 ) | ( n54617 & ~n54618 ) ;
  assign n54622 = n5852 ^ n5483 ^ n3974 ;
  assign n54620 = ( ~n25541 & n26557 ) | ( ~n25541 & n28187 ) | ( n26557 & n28187 ) ;
  assign n54621 = n54620 ^ n44411 ^ n41034 ;
  assign n54623 = n54622 ^ n54621 ^ n2527 ;
  assign n54624 = n37305 ^ n36351 ^ n26164 ;
  assign n54625 = n31102 ^ n6778 ^ n1348 ;
  assign n54626 = n54625 ^ n53056 ^ n8654 ;
  assign n54627 = n26097 ^ n15953 ^ n9662 ;
  assign n54628 = n51420 ^ n45656 ^ n39066 ;
  assign n54629 = n11327 ^ n4288 ^ n4286 ;
  assign n54630 = ( n4308 & n15699 ) | ( n4308 & n39505 ) | ( n15699 & n39505 ) ;
  assign n54631 = ~n5516 & n54630 ;
  assign n54632 = ~n54629 & n54631 ;
  assign n54633 = ~n3409 & n23372 ;
  assign n54634 = n54633 ^ n7059 ^ 1'b0 ;
  assign n54635 = n48976 ^ n38943 ^ n5004 ;
  assign n54636 = n46319 ^ n16894 ^ n15041 ;
  assign n54637 = ( n23108 & ~n23287 ) | ( n23108 & n42505 ) | ( ~n23287 & n42505 ) ;
  assign n54638 = n25078 ^ n5290 ^ n420 ;
  assign n54639 = ( ~n10080 & n54637 ) | ( ~n10080 & n54638 ) | ( n54637 & n54638 ) ;
  assign n54640 = n54555 ^ n45435 ^ n32539 ;
  assign n54641 = n5002 & ~n49268 ;
  assign n54642 = n49732 ^ n23457 ^ n2188 ;
  assign n54647 = n12178 ^ n5991 ^ 1'b0 ;
  assign n54648 = n7084 | n54647 ;
  assign n54643 = ( ~n1509 & n4472 ) | ( ~n1509 & n32093 ) | ( n4472 & n32093 ) ;
  assign n54644 = ( n3282 & ~n28641 ) | ( n3282 & n54643 ) | ( ~n28641 & n54643 ) ;
  assign n54645 = n33332 ^ n8590 ^ n606 ;
  assign n54646 = ( n2233 & n54644 ) | ( n2233 & ~n54645 ) | ( n54644 & ~n54645 ) ;
  assign n54649 = n54648 ^ n54646 ^ n47323 ;
  assign n54650 = n2920 & ~n32611 ;
  assign n54651 = ( n7674 & n8040 ) | ( n7674 & n14677 ) | ( n8040 & n14677 ) ;
  assign n54652 = n13501 ^ n4212 ^ 1'b0 ;
  assign n54653 = ~n6879 & n32676 ;
  assign n54654 = n54653 ^ n47157 ^ 1'b0 ;
  assign n54655 = ( ~n12222 & n43752 ) | ( ~n12222 & n50178 ) | ( n43752 & n50178 ) ;
  assign n54656 = ( n7250 & n23088 ) | ( n7250 & ~n35373 ) | ( n23088 & ~n35373 ) ;
  assign n54657 = ( ~n8709 & n27646 ) | ( ~n8709 & n45249 ) | ( n27646 & n45249 ) ;
  assign n54658 = n54657 ^ n45833 ^ n7818 ;
  assign n54659 = n12355 & n47306 ;
  assign n54660 = ( n9193 & n13861 ) | ( n9193 & ~n54659 ) | ( n13861 & ~n54659 ) ;
  assign n54661 = ( ~n8452 & n33592 ) | ( ~n8452 & n38681 ) | ( n33592 & n38681 ) ;
  assign n54662 = ( n4447 & ~n19675 ) | ( n4447 & n36581 ) | ( ~n19675 & n36581 ) ;
  assign n54663 = n3197 & ~n44335 ;
  assign n54664 = n54663 ^ n6415 ^ 1'b0 ;
  assign n54665 = ( n709 & ~n12787 ) | ( n709 & n54664 ) | ( ~n12787 & n54664 ) ;
  assign n54666 = ( n19480 & n31198 ) | ( n19480 & ~n54665 ) | ( n31198 & ~n54665 ) ;
  assign n54669 = n9733 ^ n1596 ^ n534 ;
  assign n54668 = n1380 & ~n9278 ;
  assign n54670 = n54669 ^ n54668 ^ 1'b0 ;
  assign n54667 = n28740 ^ n10467 ^ n6993 ;
  assign n54671 = n54670 ^ n54667 ^ n52600 ;
  assign n54672 = n35391 ^ n10529 ^ n3065 ;
  assign n54673 = n39179 ^ n36065 ^ 1'b0 ;
  assign n54674 = ~n23691 & n54673 ;
  assign n54675 = n54674 ^ n18651 ^ n5056 ;
  assign n54676 = n15185 & ~n44495 ;
  assign n54677 = n54675 & n54676 ;
  assign n54678 = n25300 & ~n30514 ;
  assign n54679 = n54678 ^ n28172 ^ 1'b0 ;
  assign n54680 = n38742 ^ n31734 ^ n5590 ;
  assign n54681 = n54680 ^ n15900 ^ n14719 ;
  assign n54682 = ( n13065 & ~n26032 ) | ( n13065 & n37925 ) | ( ~n26032 & n37925 ) ;
  assign n54683 = n39962 ^ n11211 ^ n4566 ;
  assign n54684 = ( ~n12995 & n44210 ) | ( ~n12995 & n54683 ) | ( n44210 & n54683 ) ;
  assign n54685 = ( n25154 & n54682 ) | ( n25154 & ~n54684 ) | ( n54682 & ~n54684 ) ;
  assign n54686 = n24493 ^ n17153 ^ 1'b0 ;
  assign n54687 = n15095 & ~n54686 ;
  assign n54688 = n54687 ^ n15205 ^ n12689 ;
  assign n54689 = ( n6118 & n46554 ) | ( n6118 & n47451 ) | ( n46554 & n47451 ) ;
  assign n54690 = ( ~n48886 & n54688 ) | ( ~n48886 & n54689 ) | ( n54688 & n54689 ) ;
  assign n54691 = n729 & n28699 ;
  assign n54692 = n54691 ^ n23626 ^ n4581 ;
  assign n54693 = n24551 & ~n40441 ;
  assign n54694 = n54693 ^ n28461 ^ 1'b0 ;
  assign n54695 = ( n15317 & ~n29972 ) | ( n15317 & n35580 ) | ( ~n29972 & n35580 ) ;
  assign n54696 = ( n33424 & n54694 ) | ( n33424 & n54695 ) | ( n54694 & n54695 ) ;
  assign n54697 = ( n10203 & ~n22730 ) | ( n10203 & n54696 ) | ( ~n22730 & n54696 ) ;
  assign n54698 = n35563 ^ n21780 ^ n19545 ;
  assign n54699 = ( n5009 & n11035 ) | ( n5009 & ~n25442 ) | ( n11035 & ~n25442 ) ;
  assign n54700 = n28287 | n54699 ;
  assign n54701 = n21820 ^ n20751 ^ n9325 ;
  assign n54702 = ( n10007 & n22938 ) | ( n10007 & ~n54701 ) | ( n22938 & ~n54701 ) ;
  assign n54703 = n9954 & n54702 ;
  assign n54704 = n41988 & n54703 ;
  assign n54705 = ( n36355 & n43327 ) | ( n36355 & ~n54704 ) | ( n43327 & ~n54704 ) ;
  assign n54706 = ( n1927 & ~n5787 ) | ( n1927 & n16425 ) | ( ~n5787 & n16425 ) ;
  assign n54707 = n24313 ^ n18688 ^ 1'b0 ;
  assign n54708 = ( n25678 & n54706 ) | ( n25678 & n54707 ) | ( n54706 & n54707 ) ;
  assign n54709 = n1936 & ~n18899 ;
  assign n54710 = ( n8456 & n43660 ) | ( n8456 & n54709 ) | ( n43660 & n54709 ) ;
  assign n54711 = ~n2345 & n27759 ;
  assign n54712 = ~n41665 & n54711 ;
  assign n54713 = n54710 & n54712 ;
  assign n54714 = n32663 ^ n25559 ^ n6312 ;
  assign n54715 = n30955 ^ n13910 ^ 1'b0 ;
  assign n54716 = ~n54714 & n54715 ;
  assign n54717 = ~n2249 & n54716 ;
  assign n54718 = n54717 ^ n44195 ^ 1'b0 ;
  assign n54719 = ( n308 & n20090 ) | ( n308 & n48974 ) | ( n20090 & n48974 ) ;
  assign n54720 = n26848 ^ n16259 ^ 1'b0 ;
  assign n54721 = n15864 & n24194 ;
  assign n54722 = n54721 ^ n2557 ^ 1'b0 ;
  assign n54723 = n54722 ^ n39790 ^ n17695 ;
  assign n54724 = n54723 ^ n23240 ^ n4113 ;
  assign n54725 = n44532 ^ n33538 ^ n14967 ;
  assign n54726 = ( ~n23721 & n39625 ) | ( ~n23721 & n40699 ) | ( n39625 & n40699 ) ;
  assign n54727 = n54726 ^ n37615 ^ n18785 ;
  assign n54728 = n54727 ^ n3100 ^ 1'b0 ;
  assign n54729 = ~n3595 & n37914 ;
  assign n54734 = ( x66 & n2264 ) | ( x66 & ~n26944 ) | ( n2264 & ~n26944 ) ;
  assign n54731 = n43855 ^ n13159 ^ 1'b0 ;
  assign n54732 = ~n16056 & n54731 ;
  assign n54730 = ~n15385 & n31787 ;
  assign n54733 = n54732 ^ n54730 ^ n16631 ;
  assign n54735 = n54734 ^ n54733 ^ n44280 ;
  assign n54736 = n47125 ^ n28639 ^ 1'b0 ;
  assign n54737 = n3753 & n4034 ;
  assign n54738 = n54737 ^ n12863 ^ 1'b0 ;
  assign n54739 = n48669 ^ n44439 ^ 1'b0 ;
  assign n54740 = ( n48594 & ~n54738 ) | ( n48594 & n54739 ) | ( ~n54738 & n54739 ) ;
  assign n54741 = n22736 ^ n10357 ^ n5319 ;
  assign n54742 = n12163 | n54741 ;
  assign n54743 = ~n14702 & n54742 ;
  assign n54744 = n54743 ^ n8179 ^ 1'b0 ;
  assign n54745 = n8706 & ~n22097 ;
  assign n54746 = n20917 & n54745 ;
  assign n54747 = n54746 ^ n50019 ^ n4802 ;
  assign n54748 = ( n2204 & ~n12588 ) | ( n2204 & n27969 ) | ( ~n12588 & n27969 ) ;
  assign n54749 = n30290 ^ n15290 ^ n5008 ;
  assign n54750 = ( n33604 & n54748 ) | ( n33604 & n54749 ) | ( n54748 & n54749 ) ;
  assign n54751 = n54750 ^ n51281 ^ n41531 ;
  assign n54752 = ( n25312 & n38602 ) | ( n25312 & n40456 ) | ( n38602 & n40456 ) ;
  assign n54753 = n54752 ^ n37632 ^ n32866 ;
  assign n54754 = n19621 ^ n18475 ^ n4718 ;
  assign n54755 = ~n5433 & n54754 ;
  assign n54756 = n20842 & ~n54755 ;
  assign n54757 = ( n20397 & n28380 ) | ( n20397 & ~n54756 ) | ( n28380 & ~n54756 ) ;
  assign n54758 = n22596 ^ n10804 ^ n7997 ;
  assign n54759 = n54758 ^ n48755 ^ n5637 ;
  assign n54760 = n42366 ^ n28792 ^ n14540 ;
  assign n54761 = n50522 ^ n41301 ^ n5598 ;
  assign n54762 = ( ~n29490 & n54760 ) | ( ~n29490 & n54761 ) | ( n54760 & n54761 ) ;
  assign n54763 = n54762 ^ n40893 ^ n17278 ;
  assign n54764 = ( ~n21802 & n27012 ) | ( ~n21802 & n54763 ) | ( n27012 & n54763 ) ;
  assign n54767 = n25323 ^ n25132 ^ n18735 ;
  assign n54768 = ( n2995 & n35205 ) | ( n2995 & ~n54767 ) | ( n35205 & ~n54767 ) ;
  assign n54765 = n1041 ^ n1001 ^ 1'b0 ;
  assign n54766 = n3325 & n54765 ;
  assign n54769 = n54768 ^ n54766 ^ n2690 ;
  assign n54779 = ( n20144 & ~n20415 ) | ( n20144 & n24540 ) | ( ~n20415 & n24540 ) ;
  assign n54778 = n50527 ^ n20933 ^ n4174 ;
  assign n54770 = n30139 ^ n24262 ^ n6359 ;
  assign n54771 = n54770 ^ n8637 ^ 1'b0 ;
  assign n54775 = n19506 ^ n19126 ^ n5210 ;
  assign n54772 = n3576 | n13592 ;
  assign n54773 = n34171 ^ n23495 ^ n16520 ;
  assign n54774 = ( ~n37384 & n54772 ) | ( ~n37384 & n54773 ) | ( n54772 & n54773 ) ;
  assign n54776 = n54775 ^ n54774 ^ n41377 ;
  assign n54777 = ( n2911 & n54771 ) | ( n2911 & n54776 ) | ( n54771 & n54776 ) ;
  assign n54780 = n54779 ^ n54778 ^ n54777 ;
  assign n54781 = n9484 & ~n16281 ;
  assign n54782 = n54781 ^ n8734 ^ 1'b0 ;
  assign n54783 = n54782 ^ n35695 ^ n12644 ;
  assign n54784 = ~n22895 & n23638 ;
  assign n54785 = n54784 ^ n26466 ^ 1'b0 ;
  assign n54786 = n28569 ^ n28132 ^ n17659 ;
  assign n54787 = ( n32933 & n50964 ) | ( n32933 & n54786 ) | ( n50964 & n54786 ) ;
  assign n54788 = ( n8755 & n15944 ) | ( n8755 & ~n54787 ) | ( n15944 & ~n54787 ) ;
  assign n54789 = n21335 ^ n12902 ^ n9799 ;
  assign n54790 = ( n944 & n11293 ) | ( n944 & n28556 ) | ( n11293 & n28556 ) ;
  assign n54791 = n54790 ^ n48204 ^ n45751 ;
  assign n54792 = ( x145 & n23445 ) | ( x145 & ~n39272 ) | ( n23445 & ~n39272 ) ;
  assign n54795 = ( n21951 & n27214 ) | ( n21951 & ~n37081 ) | ( n27214 & ~n37081 ) ;
  assign n54796 = n54795 ^ n13157 ^ n5151 ;
  assign n54793 = ( n33409 & n33614 ) | ( n33409 & n40176 ) | ( n33614 & n40176 ) ;
  assign n54794 = n39015 | n54793 ;
  assign n54797 = n54796 ^ n54794 ^ n52271 ;
  assign n54798 = n28938 ^ n4358 ^ n732 ;
  assign n54799 = ( n3357 & n8862 ) | ( n3357 & ~n44167 ) | ( n8862 & ~n44167 ) ;
  assign n54800 = ( n13941 & ~n54798 ) | ( n13941 & n54799 ) | ( ~n54798 & n54799 ) ;
  assign n54803 = n36835 ^ n3903 ^ n1423 ;
  assign n54801 = n11655 ^ n10147 ^ n9712 ;
  assign n54802 = ( n11049 & n23869 ) | ( n11049 & n54801 ) | ( n23869 & n54801 ) ;
  assign n54804 = n54803 ^ n54802 ^ n31585 ;
  assign n54805 = n4751 | n33288 ;
  assign n54806 = ( n2140 & n16075 ) | ( n2140 & ~n34254 ) | ( n16075 & ~n34254 ) ;
  assign n54807 = n54806 ^ n31116 ^ n1205 ;
  assign n54809 = ~n4921 & n5334 ;
  assign n54810 = n54809 ^ n3851 ^ 1'b0 ;
  assign n54808 = n23430 & ~n47731 ;
  assign n54811 = n54810 ^ n54808 ^ n44863 ;
  assign n54812 = ( n9319 & n29166 ) | ( n9319 & ~n49099 ) | ( n29166 & ~n49099 ) ;
  assign n54813 = ( ~n19615 & n48962 ) | ( ~n19615 & n50534 ) | ( n48962 & n50534 ) ;
  assign n54814 = ( n3686 & n10314 ) | ( n3686 & n53152 ) | ( n10314 & n53152 ) ;
  assign n54815 = n54814 ^ n51940 ^ n12891 ;
  assign n54816 = n31857 ^ n23976 ^ 1'b0 ;
  assign n54817 = ~n3466 & n10180 ;
  assign n54818 = ~n7953 & n54817 ;
  assign n54819 = n54818 ^ n53145 ^ n39261 ;
  assign n54820 = n17377 & ~n20398 ;
  assign n54821 = n46355 ^ n26522 ^ 1'b0 ;
  assign n54822 = ~n22805 & n54821 ;
  assign n54823 = n54822 ^ n40657 ^ n8024 ;
  assign n54824 = ( n14588 & n17327 ) | ( n14588 & ~n34487 ) | ( n17327 & ~n34487 ) ;
  assign n54825 = n54824 ^ n16465 ^ 1'b0 ;
  assign n54826 = ~n31488 & n54825 ;
  assign n54827 = n45267 ^ n2443 ^ 1'b0 ;
  assign n54828 = n49465 & ~n54827 ;
  assign n54829 = n34374 ^ n33537 ^ n33531 ;
  assign n54830 = n17558 ^ n7231 ^ n5730 ;
  assign n54831 = n54830 ^ n30133 ^ n20373 ;
  assign n54832 = ( n16653 & ~n19602 ) | ( n16653 & n30904 ) | ( ~n19602 & n30904 ) ;
  assign n54835 = n35972 ^ n13036 ^ n3407 ;
  assign n54836 = n54835 ^ n34962 ^ n34294 ;
  assign n54833 = ( n6592 & n12946 ) | ( n6592 & n19653 ) | ( n12946 & n19653 ) ;
  assign n54834 = n54833 ^ n13507 ^ 1'b0 ;
  assign n54837 = n54836 ^ n54834 ^ n5424 ;
  assign n54838 = n40999 ^ n35325 ^ 1'b0 ;
  assign n54839 = n3952 | n23216 ;
  assign n54840 = ( n17304 & n35712 ) | ( n17304 & ~n52136 ) | ( n35712 & ~n52136 ) ;
  assign n54841 = n38795 ^ n15658 ^ n3112 ;
  assign n54842 = ( ~n11312 & n54840 ) | ( ~n11312 & n54841 ) | ( n54840 & n54841 ) ;
  assign n54843 = ( ~n30078 & n54839 ) | ( ~n30078 & n54842 ) | ( n54839 & n54842 ) ;
  assign n54844 = ( n814 & n6498 ) | ( n814 & n34441 ) | ( n6498 & n34441 ) ;
  assign n54845 = ( ~n22263 & n48229 ) | ( ~n22263 & n54844 ) | ( n48229 & n54844 ) ;
  assign n54846 = ( n11217 & n32168 ) | ( n11217 & n33317 ) | ( n32168 & n33317 ) ;
  assign n54847 = ( n5745 & n25030 ) | ( n5745 & ~n27203 ) | ( n25030 & ~n27203 ) ;
  assign n54848 = ( n12994 & n16087 ) | ( n12994 & n28504 ) | ( n16087 & n28504 ) ;
  assign n54849 = n45049 ^ n15160 ^ 1'b0 ;
  assign n54850 = n54848 & n54849 ;
  assign n54851 = ~n4647 & n26466 ;
  assign n54852 = n54851 ^ n5855 ^ 1'b0 ;
  assign n54853 = n44838 ^ n36316 ^ n11425 ;
  assign n54854 = n20079 ^ n19972 ^ n2000 ;
  assign n54855 = n54854 ^ n7658 ^ n6257 ;
  assign n54857 = n42130 ^ n37261 ^ 1'b0 ;
  assign n54856 = n46924 ^ n36872 ^ 1'b0 ;
  assign n54858 = n54857 ^ n54856 ^ n3550 ;
  assign n54859 = ( n10487 & ~n15553 ) | ( n10487 & n41821 ) | ( ~n15553 & n41821 ) ;
  assign n54860 = ( n2428 & n8031 ) | ( n2428 & n29135 ) | ( n8031 & n29135 ) ;
  assign n54861 = n16836 & n32270 ;
  assign n54862 = ~n36035 & n54861 ;
  assign n54863 = n54862 ^ n10395 ^ 1'b0 ;
  assign n54864 = n14270 ^ n1821 ^ n780 ;
  assign n54865 = ( n20292 & ~n22542 ) | ( n20292 & n54864 ) | ( ~n22542 & n54864 ) ;
  assign n54866 = ( ~n35917 & n45917 ) | ( ~n35917 & n49051 ) | ( n45917 & n49051 ) ;
  assign n54867 = ( ~n21933 & n41450 ) | ( ~n21933 & n43132 ) | ( n41450 & n43132 ) ;
  assign n54868 = n2428 & n24044 ;
  assign n54869 = n3721 & n54868 ;
  assign n54870 = n11107 ^ n5148 ^ 1'b0 ;
  assign n54871 = n23484 & n54870 ;
  assign n54879 = n10963 ^ n6194 ^ n3872 ;
  assign n54873 = n33520 ^ n6649 ^ n4202 ;
  assign n54874 = ( n13143 & ~n23341 ) | ( n13143 & n26933 ) | ( ~n23341 & n26933 ) ;
  assign n54875 = ( ~n32996 & n54873 ) | ( ~n32996 & n54874 ) | ( n54873 & n54874 ) ;
  assign n54876 = n54875 ^ n39019 ^ n8276 ;
  assign n54872 = ( ~n23634 & n41972 ) | ( ~n23634 & n43855 ) | ( n41972 & n43855 ) ;
  assign n54877 = n54876 ^ n54872 ^ n6272 ;
  assign n54878 = n54877 ^ n29966 ^ n3087 ;
  assign n54880 = n54879 ^ n54878 ^ n7424 ;
  assign n54882 = n33251 ^ n20776 ^ n15760 ;
  assign n54881 = ( n4863 & ~n7378 ) | ( n4863 & n8663 ) | ( ~n7378 & n8663 ) ;
  assign n54883 = n54882 ^ n54881 ^ n30259 ;
  assign n54884 = n20922 | n34210 ;
  assign n54885 = n54884 ^ n11511 ^ 1'b0 ;
  assign n54886 = n54885 ^ n36857 ^ n6121 ;
  assign n54887 = ( n11708 & n27390 ) | ( n11708 & ~n31508 ) | ( n27390 & ~n31508 ) ;
  assign n54888 = ( n10010 & n50581 ) | ( n10010 & n54887 ) | ( n50581 & n54887 ) ;
  assign n54889 = ( ~n24443 & n29972 ) | ( ~n24443 & n54888 ) | ( n29972 & n54888 ) ;
  assign n54890 = ( n21131 & n51722 ) | ( n21131 & n51938 ) | ( n51722 & n51938 ) ;
  assign n54891 = n9265 & n41508 ;
  assign n54892 = ( n16737 & ~n19468 ) | ( n16737 & n39092 ) | ( ~n19468 & n39092 ) ;
  assign n54893 = n5632 & ~n36232 ;
  assign n54894 = ~n54892 & n54893 ;
  assign n54895 = n54894 ^ n30693 ^ 1'b0 ;
  assign n54896 = n54895 ^ n52024 ^ n36286 ;
  assign n54899 = n36790 ^ n12045 ^ 1'b0 ;
  assign n54897 = n25389 & ~n45719 ;
  assign n54898 = n54897 ^ n29084 ^ 1'b0 ;
  assign n54900 = n54899 ^ n54898 ^ n8970 ;
  assign n54901 = n10475 & n26030 ;
  assign n54902 = n54901 ^ n3760 ^ 1'b0 ;
  assign n54903 = n37947 ^ n3333 ^ 1'b0 ;
  assign n54904 = n54903 ^ n21758 ^ n11674 ;
  assign n54908 = n22430 ^ n7393 ^ n7283 ;
  assign n54905 = ( ~n13559 & n16768 ) | ( ~n13559 & n23368 ) | ( n16768 & n23368 ) ;
  assign n54906 = n54905 ^ n25640 ^ n3437 ;
  assign n54907 = n54906 ^ n50493 ^ n1816 ;
  assign n54909 = n54908 ^ n54907 ^ n19709 ;
  assign n54910 = ~n27684 & n54909 ;
  assign n54911 = n6437 | n24612 ;
  assign n54912 = n24415 & ~n54911 ;
  assign n54913 = n54912 ^ n50329 ^ x216 ;
  assign n54915 = n50736 ^ n9604 ^ 1'b0 ;
  assign n54916 = n19249 | n54915 ;
  assign n54914 = n32505 ^ n26499 ^ n6819 ;
  assign n54917 = n54916 ^ n54914 ^ n1565 ;
  assign n54918 = n54917 ^ n25265 ^ n13377 ;
  assign n54919 = n54918 ^ n20339 ^ n20007 ;
  assign n54920 = ( ~n8301 & n18512 ) | ( ~n8301 & n43340 ) | ( n18512 & n43340 ) ;
  assign n54921 = ( ~n1596 & n3380 ) | ( ~n1596 & n40114 ) | ( n3380 & n40114 ) ;
  assign n54922 = n54921 ^ n15425 ^ n6096 ;
  assign n54923 = n20943 ^ n18506 ^ n4983 ;
  assign n54924 = ( n12603 & n17767 ) | ( n12603 & ~n54923 ) | ( n17767 & ~n54923 ) ;
  assign n54925 = ( ~n2646 & n8246 ) | ( ~n2646 & n50189 ) | ( n8246 & n50189 ) ;
  assign n54926 = ( n18633 & ~n20354 ) | ( n18633 & n22368 ) | ( ~n20354 & n22368 ) ;
  assign n54927 = n26447 ^ n3159 ^ n3131 ;
  assign n54928 = ( ~n48515 & n54926 ) | ( ~n48515 & n54927 ) | ( n54926 & n54927 ) ;
  assign n54929 = ( n12914 & n14921 ) | ( n12914 & n54928 ) | ( n14921 & n54928 ) ;
  assign n54930 = n20605 & ~n45821 ;
  assign n54931 = n54930 ^ n18561 ^ 1'b0 ;
  assign n54932 = ~n6536 & n23325 ;
  assign n54935 = ( ~n11178 & n18769 ) | ( ~n11178 & n19956 ) | ( n18769 & n19956 ) ;
  assign n54933 = n8860 ^ n5848 ^ n4160 ;
  assign n54934 = n54933 ^ n12651 ^ n5151 ;
  assign n54936 = n54935 ^ n54934 ^ n10667 ;
  assign n54937 = n43736 ^ n29167 ^ 1'b0 ;
  assign n54938 = ( n39314 & n45961 ) | ( n39314 & ~n54937 ) | ( n45961 & ~n54937 ) ;
  assign n54939 = n31771 ^ n29157 ^ n24567 ;
  assign n54940 = n45166 ^ n30207 ^ 1'b0 ;
  assign n54942 = n28161 ^ n14506 ^ n1873 ;
  assign n54941 = n32969 ^ x193 ^ x107 ;
  assign n54943 = n54942 ^ n54941 ^ n16990 ;
  assign n54944 = ( n6587 & ~n24596 ) | ( n6587 & n54943 ) | ( ~n24596 & n54943 ) ;
  assign n54945 = n28464 ^ n760 ^ 1'b0 ;
  assign n54946 = n21712 | n24196 ;
  assign n54947 = n50064 ^ n14861 ^ n8305 ;
  assign n54948 = n54947 ^ n39367 ^ n23079 ;
  assign n54949 = ( ~n8170 & n54946 ) | ( ~n8170 & n54948 ) | ( n54946 & n54948 ) ;
  assign n54950 = ( ~n21516 & n54945 ) | ( ~n21516 & n54949 ) | ( n54945 & n54949 ) ;
  assign n54951 = n40872 ^ n9692 ^ n8983 ;
  assign n54952 = ( n19401 & ~n29485 ) | ( n19401 & n45494 ) | ( ~n29485 & n45494 ) ;
  assign n54953 = ( n16926 & ~n54702 ) | ( n16926 & n54952 ) | ( ~n54702 & n54952 ) ;
  assign n54954 = n49722 ^ n10340 ^ 1'b0 ;
  assign n54955 = ~n8560 & n54954 ;
  assign n54956 = n38207 ^ n32295 ^ n28384 ;
  assign n54958 = n34535 ^ n15072 ^ 1'b0 ;
  assign n54957 = n23377 | n27762 ;
  assign n54959 = n54958 ^ n54957 ^ 1'b0 ;
  assign n54960 = n54959 ^ n41917 ^ 1'b0 ;
  assign n54961 = n54956 & n54960 ;
  assign n54962 = ( n4791 & ~n14228 ) | ( n4791 & n21711 ) | ( ~n14228 & n21711 ) ;
  assign n54963 = n32570 ^ n23161 ^ n5938 ;
  assign n54964 = ( n10612 & ~n14934 ) | ( n10612 & n54963 ) | ( ~n14934 & n54963 ) ;
  assign n54965 = n54964 ^ n51458 ^ n14025 ;
  assign n54966 = n36102 ^ n9635 ^ n2582 ;
  assign n54967 = ( n4737 & n7297 ) | ( n4737 & ~n35389 ) | ( n7297 & ~n35389 ) ;
  assign n54968 = n28043 ^ n26314 ^ n19606 ;
  assign n54969 = n50574 ^ n36636 ^ 1'b0 ;
  assign n54970 = ( n39181 & n54968 ) | ( n39181 & ~n54969 ) | ( n54968 & ~n54969 ) ;
  assign n54971 = ( n17266 & n25081 ) | ( n17266 & ~n54970 ) | ( n25081 & ~n54970 ) ;
  assign n54972 = n50702 ^ n44074 ^ n13258 ;
  assign n54973 = ( n17789 & ~n24018 ) | ( n17789 & n37354 ) | ( ~n24018 & n37354 ) ;
  assign n54974 = n1278 & ~n54973 ;
  assign n54975 = n6075 ^ n1341 ^ 1'b0 ;
  assign n54976 = n8228 | n54975 ;
  assign n54977 = n54976 ^ n20104 ^ 1'b0 ;
  assign n54978 = ( n8162 & n12164 ) | ( n8162 & ~n25633 ) | ( n12164 & ~n25633 ) ;
  assign n54979 = ( n38054 & n40808 ) | ( n38054 & n54978 ) | ( n40808 & n54978 ) ;
  assign n54980 = n25970 & ~n38933 ;
  assign n54981 = n53073 ^ n29937 ^ 1'b0 ;
  assign n54982 = n26342 & ~n54981 ;
  assign n54983 = n38137 ^ n36359 ^ n28766 ;
  assign n54984 = ( x216 & ~n52160 ) | ( x216 & n54983 ) | ( ~n52160 & n54983 ) ;
  assign n54985 = ~n2115 & n9328 ;
  assign n54986 = n54985 ^ n45665 ^ 1'b0 ;
  assign n54987 = ( n2954 & n3192 ) | ( n2954 & ~n37757 ) | ( n3192 & ~n37757 ) ;
  assign n54988 = n54987 ^ n24409 ^ n2517 ;
  assign n54989 = n37360 | n54988 ;
  assign n54990 = n20215 & ~n54989 ;
  assign n54991 = ( n15490 & n54986 ) | ( n15490 & ~n54990 ) | ( n54986 & ~n54990 ) ;
  assign n54992 = ( ~n14805 & n28801 ) | ( ~n14805 & n36425 ) | ( n28801 & n36425 ) ;
  assign n54993 = n54992 ^ n23010 ^ n2424 ;
  assign n54994 = n28411 ^ n446 ^ 1'b0 ;
  assign n54995 = ( n603 & ~n1880 ) | ( n603 & n48139 ) | ( ~n1880 & n48139 ) ;
  assign n54996 = n4902 & ~n22107 ;
  assign n54997 = n54996 ^ n4275 ^ 1'b0 ;
  assign n54998 = n54997 ^ n43352 ^ n30152 ;
  assign n55000 = ( n1245 & ~n2800 ) | ( n1245 & n16042 ) | ( ~n2800 & n16042 ) ;
  assign n54999 = n6598 & n8674 ;
  assign n55001 = n55000 ^ n54999 ^ n31202 ;
  assign n55002 = n27410 ^ n4598 ^ n361 ;
  assign n55003 = ( ~n1299 & n27646 ) | ( ~n1299 & n55002 ) | ( n27646 & n55002 ) ;
  assign n55004 = n15264 & n20737 ;
  assign n55005 = n55004 ^ n39478 ^ n14109 ;
  assign n55006 = n35369 ^ n21449 ^ n13474 ;
  assign n55009 = ( n6321 & ~n31876 ) | ( n6321 & n49078 ) | ( ~n31876 & n49078 ) ;
  assign n55007 = ~n7496 & n46197 ;
  assign n55008 = n55007 ^ n2573 ^ 1'b0 ;
  assign n55010 = n55009 ^ n55008 ^ n34985 ;
  assign n55011 = ( n16035 & ~n55006 ) | ( n16035 & n55010 ) | ( ~n55006 & n55010 ) ;
  assign n55012 = n12765 ^ n8818 ^ 1'b0 ;
  assign n55013 = n10055 & n55012 ;
  assign n55014 = n55013 ^ n48908 ^ n9958 ;
  assign n55015 = n14503 | n24002 ;
  assign n55017 = n14556 ^ n12854 ^ n11021 ;
  assign n55016 = n6551 ^ n5766 ^ n4759 ;
  assign n55018 = n55017 ^ n55016 ^ n30996 ;
  assign n55019 = n30756 & ~n38961 ;
  assign n55020 = n55019 ^ n30857 ^ 1'b0 ;
  assign n55021 = ( n25198 & ~n38447 ) | ( n25198 & n55020 ) | ( ~n38447 & n55020 ) ;
  assign n55022 = n55021 ^ n21114 ^ n20680 ;
  assign n55024 = n6795 & ~n15302 ;
  assign n55023 = n24525 ^ n22725 ^ n7155 ;
  assign n55025 = n55024 ^ n55023 ^ n21312 ;
  assign n55026 = ( n23355 & n28687 ) | ( n23355 & n55025 ) | ( n28687 & n55025 ) ;
  assign n55027 = ( ~n6902 & n22739 ) | ( ~n6902 & n31444 ) | ( n22739 & n31444 ) ;
  assign n55028 = ( n4488 & n43549 ) | ( n4488 & n55027 ) | ( n43549 & n55027 ) ;
  assign n55029 = n49965 & n55028 ;
  assign n55030 = n48063 ^ n8572 ^ n1930 ;
  assign n55031 = n39606 ^ n33792 ^ n15961 ;
  assign n55032 = n831 & n3265 ;
  assign n55033 = n55032 ^ n8349 ^ 1'b0 ;
  assign n55034 = ( ~n13144 & n24904 ) | ( ~n13144 & n55033 ) | ( n24904 & n55033 ) ;
  assign n55035 = ~n15221 & n55034 ;
  assign n55036 = n55035 ^ n41189 ^ 1'b0 ;
  assign n55037 = n48399 ^ n25063 ^ n13258 ;
  assign n55038 = ( n9864 & n11669 ) | ( n9864 & n55037 ) | ( n11669 & n55037 ) ;
  assign n55039 = n32895 ^ n11482 ^ 1'b0 ;
  assign n55040 = ( ~n17918 & n38509 ) | ( ~n17918 & n54530 ) | ( n38509 & n54530 ) ;
  assign n55041 = n20172 ^ n11385 ^ n6904 ;
  assign n55042 = n55041 ^ n27660 ^ n15030 ;
  assign n55043 = n55042 ^ n40591 ^ n24185 ;
  assign n55044 = n29837 ^ n26750 ^ 1'b0 ;
  assign n55045 = ( n18934 & n23332 ) | ( n18934 & ~n40505 ) | ( n23332 & ~n40505 ) ;
  assign n55046 = n55045 ^ n11533 ^ 1'b0 ;
  assign n55047 = n55046 ^ n16273 ^ n12570 ;
  assign n55050 = n44143 ^ n21245 ^ n15942 ;
  assign n55048 = n7493 & ~n20446 ;
  assign n55049 = n30216 & n55048 ;
  assign n55051 = n55050 ^ n55049 ^ n29013 ;
  assign n55052 = ( n40510 & n44469 ) | ( n40510 & n55051 ) | ( n44469 & n55051 ) ;
  assign n55053 = n50890 ^ n16412 ^ n3877 ;
  assign n55054 = n25253 & ~n55053 ;
  assign n55055 = n55054 ^ n49678 ^ n34005 ;
  assign n55056 = n55055 ^ n34751 ^ n6240 ;
  assign n55057 = n55056 ^ n21889 ^ n14907 ;
  assign n55058 = n48823 ^ n11216 ^ n706 ;
  assign n55059 = n17153 | n51418 ;
  assign n55060 = n45220 & ~n55059 ;
  assign n55062 = ( n16768 & n37906 ) | ( n16768 & n40536 ) | ( n37906 & n40536 ) ;
  assign n55061 = n1012 & ~n50739 ;
  assign n55063 = n55062 ^ n55061 ^ 1'b0 ;
  assign n55064 = ( n397 & n35347 ) | ( n397 & ~n35861 ) | ( n35347 & ~n35861 ) ;
  assign n55065 = ( ~n19013 & n37249 ) | ( ~n19013 & n50355 ) | ( n37249 & n50355 ) ;
  assign n55066 = ( n41950 & ~n55064 ) | ( n41950 & n55065 ) | ( ~n55064 & n55065 ) ;
  assign n55067 = ( n41438 & ~n51359 ) | ( n41438 & n55066 ) | ( ~n51359 & n55066 ) ;
  assign n55068 = ( n10605 & ~n31090 ) | ( n10605 & n33061 ) | ( ~n31090 & n33061 ) ;
  assign n55069 = ( ~n3535 & n16668 ) | ( ~n3535 & n24409 ) | ( n16668 & n24409 ) ;
  assign n55070 = ( ~n30530 & n36896 ) | ( ~n30530 & n45444 ) | ( n36896 & n45444 ) ;
  assign n55071 = ( n7239 & n51731 ) | ( n7239 & n55070 ) | ( n51731 & n55070 ) ;
  assign n55072 = n33098 ^ n25719 ^ n13361 ;
  assign n55073 = n765 | n32718 ;
  assign n55074 = n3999 & ~n55073 ;
  assign n55075 = ( ~n14267 & n48957 ) | ( ~n14267 & n55074 ) | ( n48957 & n55074 ) ;
  assign n55078 = n48755 ^ n15261 ^ 1'b0 ;
  assign n55079 = n36232 | n55078 ;
  assign n55076 = ( n22777 & n40547 ) | ( n22777 & ~n47624 ) | ( n40547 & ~n47624 ) ;
  assign n55077 = ( n28929 & n32398 ) | ( n28929 & ~n55076 ) | ( n32398 & ~n55076 ) ;
  assign n55080 = n55079 ^ n55077 ^ n38214 ;
  assign n55081 = n4211 & ~n25146 ;
  assign n55082 = n55081 ^ n21970 ^ n18586 ;
  assign n55083 = n2344 & n29054 ;
  assign n55084 = n55083 ^ n12668 ^ 1'b0 ;
  assign n55085 = n858 | n55084 ;
  assign n55086 = n16053 & ~n55085 ;
  assign n55087 = n38315 ^ n14687 ^ n2899 ;
  assign n55088 = n24688 ^ n18879 ^ 1'b0 ;
  assign n55089 = n9011 | n55088 ;
  assign n55090 = ( n55086 & ~n55087 ) | ( n55086 & n55089 ) | ( ~n55087 & n55089 ) ;
  assign n55091 = n19998 ^ n7536 ^ 1'b0 ;
  assign n55092 = n17282 & ~n55091 ;
  assign n55093 = n32754 ^ n1556 ^ 1'b0 ;
  assign n55094 = n35967 ^ n34540 ^ n32684 ;
  assign n55095 = n55094 ^ n3204 ^ 1'b0 ;
  assign n55096 = ( n12015 & ~n44931 ) | ( n12015 & n47283 ) | ( ~n44931 & n47283 ) ;
  assign n55097 = ( n38242 & n41752 ) | ( n38242 & n43742 ) | ( n41752 & n43742 ) ;
  assign n55098 = ( n8123 & ~n22320 ) | ( n8123 & n55097 ) | ( ~n22320 & n55097 ) ;
  assign n55099 = n52140 ^ n41975 ^ n11694 ;
  assign n55100 = ( n17562 & n25810 ) | ( n17562 & n45897 ) | ( n25810 & n45897 ) ;
  assign n55101 = n46657 ^ n41797 ^ n41387 ;
  assign n55102 = n46840 ^ n23627 ^ n9277 ;
  assign n55103 = n42098 & ~n54638 ;
  assign n55104 = ( n10845 & ~n21436 ) | ( n10845 & n55103 ) | ( ~n21436 & n55103 ) ;
  assign n55105 = n10252 ^ n342 ^ 1'b0 ;
  assign n55106 = n16146 & n55105 ;
  assign n55111 = n28801 ^ n18522 ^ n14549 ;
  assign n55112 = ( n5762 & n34691 ) | ( n5762 & n55111 ) | ( n34691 & n55111 ) ;
  assign n55107 = ( n8959 & n29357 ) | ( n8959 & n30841 ) | ( n29357 & n30841 ) ;
  assign n55108 = n55107 ^ n40807 ^ n27640 ;
  assign n55109 = ( n14165 & n35334 ) | ( n14165 & n55108 ) | ( n35334 & n55108 ) ;
  assign n55110 = n9418 | n55109 ;
  assign n55113 = n55112 ^ n55110 ^ 1'b0 ;
  assign n55114 = n16451 ^ n16045 ^ n282 ;
  assign n55115 = n45906 ^ n28439 ^ 1'b0 ;
  assign n55116 = ( n43643 & n55114 ) | ( n43643 & n55115 ) | ( n55114 & n55115 ) ;
  assign n55117 = ( n14949 & n41649 ) | ( n14949 & ~n51180 ) | ( n41649 & ~n51180 ) ;
  assign n55118 = n38127 ^ n31449 ^ 1'b0 ;
  assign n55119 = ( n6792 & n7672 ) | ( n6792 & n30860 ) | ( n7672 & n30860 ) ;
  assign n55120 = ( n16805 & n22087 ) | ( n16805 & n40103 ) | ( n22087 & n40103 ) ;
  assign n55121 = n49401 | n55120 ;
  assign n55122 = ( x91 & ~n10405 ) | ( x91 & n55121 ) | ( ~n10405 & n55121 ) ;
  assign n55123 = ( ~n11434 & n13198 ) | ( ~n11434 & n27306 ) | ( n13198 & n27306 ) ;
  assign n55124 = ( n35867 & n45057 ) | ( n35867 & ~n55123 ) | ( n45057 & ~n55123 ) ;
  assign n55125 = n35855 ^ n28378 ^ n5950 ;
  assign n55126 = n55125 ^ n52479 ^ n17487 ;
  assign n55127 = n38695 ^ n2288 ^ 1'b0 ;
  assign n55128 = n36356 ^ n21135 ^ n8701 ;
  assign n55129 = n36501 ^ n1507 ^ 1'b0 ;
  assign n55130 = n31896 | n55129 ;
  assign n55131 = ( ~n3300 & n17273 ) | ( ~n3300 & n17345 ) | ( n17273 & n17345 ) ;
  assign n55132 = ( ~n42153 & n44187 ) | ( ~n42153 & n55131 ) | ( n44187 & n55131 ) ;
  assign n55133 = n55132 ^ n15880 ^ n496 ;
  assign n55134 = n18891 ^ n9782 ^ n1817 ;
  assign n55135 = ~n6428 & n45978 ;
  assign n55136 = n9192 ^ n2795 ^ 1'b0 ;
  assign n55144 = n28384 ^ n19121 ^ n9923 ;
  assign n55145 = ( n1786 & n22596 ) | ( n1786 & ~n55144 ) | ( n22596 & ~n55144 ) ;
  assign n55140 = n7395 & n8783 ;
  assign n55141 = n55140 ^ n3957 ^ 1'b0 ;
  assign n55142 = ( n12337 & n32888 ) | ( n12337 & n55141 ) | ( n32888 & n55141 ) ;
  assign n55139 = ( n13813 & n15245 ) | ( n13813 & ~n34122 ) | ( n15245 & ~n34122 ) ;
  assign n55137 = n3622 & n41458 ;
  assign n55138 = n8452 & n55137 ;
  assign n55143 = n55142 ^ n55139 ^ n55138 ;
  assign n55146 = n55145 ^ n55143 ^ n6365 ;
  assign n55147 = n21966 ^ n6942 ^ 1'b0 ;
  assign n55148 = ( n33272 & ~n38370 ) | ( n33272 & n55147 ) | ( ~n38370 & n55147 ) ;
  assign n55149 = n20299 ^ n11427 ^ n3576 ;
  assign n55150 = n6803 & ~n11317 ;
  assign n55151 = n55150 ^ n9764 ^ 1'b0 ;
  assign n55152 = n55151 ^ n51614 ^ n12002 ;
  assign n55153 = ( n14047 & n16732 ) | ( n14047 & ~n25112 ) | ( n16732 & ~n25112 ) ;
  assign n55154 = n55153 ^ n30408 ^ n17401 ;
  assign n55155 = ( n9669 & ~n55152 ) | ( n9669 & n55154 ) | ( ~n55152 & n55154 ) ;
  assign n55156 = ( n5396 & n10257 ) | ( n5396 & ~n46655 ) | ( n10257 & ~n46655 ) ;
  assign n55157 = n55156 ^ n50483 ^ n17135 ;
  assign n55158 = ( n1705 & ~n12389 ) | ( n1705 & n38225 ) | ( ~n12389 & n38225 ) ;
  assign n55159 = n22729 | n44641 ;
  assign n55160 = ( n14794 & n17277 ) | ( n14794 & n51557 ) | ( n17277 & n51557 ) ;
  assign n55161 = n54488 ^ n28062 ^ n20397 ;
  assign n55162 = n55161 ^ n15293 ^ n646 ;
  assign n55163 = n29858 ^ n13300 ^ n4964 ;
  assign n55164 = n42602 & ~n49192 ;
  assign n55166 = n26048 ^ n12145 ^ n4811 ;
  assign n55165 = ( ~n27500 & n35518 ) | ( ~n27500 & n54782 ) | ( n35518 & n54782 ) ;
  assign n55167 = n55166 ^ n55165 ^ n34291 ;
  assign n55168 = n55167 ^ n47256 ^ n37049 ;
  assign n55169 = ( n6740 & ~n10893 ) | ( n6740 & n55168 ) | ( ~n10893 & n55168 ) ;
  assign n55170 = n31563 ^ n23703 ^ n12747 ;
  assign n55171 = n43775 ^ n35592 ^ n33339 ;
  assign n55172 = n2778 & n41417 ;
  assign n55173 = n55172 ^ n7815 ^ 1'b0 ;
  assign n55174 = n36713 ^ n35616 ^ n34943 ;
  assign n55175 = n30407 | n55174 ;
  assign n55176 = ~n14934 & n55175 ;
  assign n55177 = n52447 & n55176 ;
  assign n55178 = n52732 ^ n40929 ^ n2881 ;
  assign n55181 = n22045 ^ n5627 ^ n1506 ;
  assign n55179 = n46073 ^ n34325 ^ n28922 ;
  assign n55180 = ( ~x48 & n280 ) | ( ~x48 & n55179 ) | ( n280 & n55179 ) ;
  assign n55182 = n55181 ^ n55180 ^ n47090 ;
  assign n55183 = ( n34390 & n46601 ) | ( n34390 & n53880 ) | ( n46601 & n53880 ) ;
  assign n55184 = n23761 ^ x161 ^ 1'b0 ;
  assign n55185 = x207 | n55184 ;
  assign n55187 = ( n2056 & n29877 ) | ( n2056 & n49838 ) | ( n29877 & n49838 ) ;
  assign n55188 = n55187 ^ n44471 ^ n11816 ;
  assign n55186 = ~n5910 & n13949 ;
  assign n55189 = n55188 ^ n55186 ^ 1'b0 ;
  assign n55190 = ( ~n12344 & n44068 ) | ( ~n12344 & n55189 ) | ( n44068 & n55189 ) ;
  assign n55191 = n53149 ^ n34029 ^ n341 ;
  assign n55192 = ( n6931 & ~n13557 ) | ( n6931 & n30917 ) | ( ~n13557 & n30917 ) ;
  assign n55193 = n18408 ^ n5988 ^ n5918 ;
  assign n55194 = n38118 ^ n24418 ^ n4126 ;
  assign n55195 = n38086 ^ n25205 ^ n14353 ;
  assign n55196 = n55195 ^ n11854 ^ n8437 ;
  assign n55197 = ( n48665 & n55009 ) | ( n48665 & n55196 ) | ( n55009 & n55196 ) ;
  assign n55198 = ( ~n55193 & n55194 ) | ( ~n55193 & n55197 ) | ( n55194 & n55197 ) ;
  assign n55199 = n55198 ^ n8268 ^ n1887 ;
  assign n55200 = n52310 ^ n37842 ^ n10730 ;
  assign n55201 = n30715 & ~n51778 ;
  assign n55202 = ( ~n30642 & n37733 ) | ( ~n30642 & n42759 ) | ( n37733 & n42759 ) ;
  assign n55203 = n53704 ^ n30507 ^ n14663 ;
  assign n55204 = n29387 ^ n4784 ^ n3390 ;
  assign n55205 = ( n7522 & n11853 ) | ( n7522 & ~n44807 ) | ( n11853 & ~n44807 ) ;
  assign n55206 = n55205 ^ n26857 ^ 1'b0 ;
  assign n55207 = n11845 & n55206 ;
  assign n55208 = ( n9522 & n29523 ) | ( n9522 & n55207 ) | ( n29523 & n55207 ) ;
  assign n55209 = n52227 ^ n12060 ^ n2181 ;
  assign n55210 = n20034 ^ n11056 ^ 1'b0 ;
  assign n55213 = n19425 ^ n14708 ^ n14383 ;
  assign n55214 = n55213 ^ n33541 ^ n10957 ;
  assign n55211 = n13479 ^ n12871 ^ n3162 ;
  assign n55212 = ( ~n18701 & n33339 ) | ( ~n18701 & n55211 ) | ( n33339 & n55211 ) ;
  assign n55215 = n55214 ^ n55212 ^ n2046 ;
  assign n55216 = n29488 ^ n5083 ^ x229 ;
  assign n55217 = n52407 ^ n48712 ^ n3677 ;
  assign n55218 = n35407 ^ n1459 ^ 1'b0 ;
  assign n55219 = n9817 & n55218 ;
  assign n55220 = n49734 ^ n22864 ^ n499 ;
  assign n55221 = n52066 ^ n16139 ^ n15391 ;
  assign n55222 = n45589 ^ n43025 ^ 1'b0 ;
  assign n55223 = ( ~n39326 & n50695 ) | ( ~n39326 & n55222 ) | ( n50695 & n55222 ) ;
  assign n55224 = n38117 ^ n20271 ^ n4263 ;
  assign n55225 = n15586 | n55224 ;
  assign n55226 = n42602 ^ n27932 ^ n10290 ;
  assign n55227 = ( ~n39729 & n46081 ) | ( ~n39729 & n47440 ) | ( n46081 & n47440 ) ;
  assign n55228 = n7422 & ~n54196 ;
  assign n55229 = ( n3132 & ~n26306 ) | ( n3132 & n48151 ) | ( ~n26306 & n48151 ) ;
  assign n55230 = n51553 ^ n29372 ^ n28011 ;
  assign n55231 = n5015 | n7178 ;
  assign n55232 = ~n5220 & n52591 ;
  assign n55233 = n55232 ^ n50501 ^ 1'b0 ;
  assign n55234 = ( ~n1277 & n16495 ) | ( ~n1277 & n20022 ) | ( n16495 & n20022 ) ;
  assign n55235 = ( n605 & n10447 ) | ( n605 & ~n18786 ) | ( n10447 & ~n18786 ) ;
  assign n55236 = ( n12272 & n55234 ) | ( n12272 & ~n55235 ) | ( n55234 & ~n55235 ) ;
  assign n55237 = ( n8144 & n39062 ) | ( n8144 & ~n46896 ) | ( n39062 & ~n46896 ) ;
  assign n55238 = n55237 ^ n50558 ^ n17048 ;
  assign n55239 = n30962 ^ n22047 ^ n14805 ;
  assign n55240 = ( ~n6081 & n31534 ) | ( ~n6081 & n54607 ) | ( n31534 & n54607 ) ;
  assign n55241 = ( n20962 & n31748 ) | ( n20962 & n33393 ) | ( n31748 & n33393 ) ;
  assign n55242 = n46246 ^ n40110 ^ n10404 ;
  assign n55243 = ( n4844 & n55241 ) | ( n4844 & n55242 ) | ( n55241 & n55242 ) ;
  assign n55244 = n41391 ^ n36786 ^ n7044 ;
  assign n55245 = n8826 ^ n5218 ^ n4218 ;
  assign n55246 = n55245 ^ n49730 ^ n20928 ;
  assign n55247 = n55246 ^ n32393 ^ n584 ;
  assign n55250 = n19766 ^ n15632 ^ 1'b0 ;
  assign n55248 = n32165 ^ n11109 ^ n5170 ;
  assign n55249 = ( n5794 & n15055 ) | ( n5794 & n55248 ) | ( n15055 & n55248 ) ;
  assign n55251 = n55250 ^ n55249 ^ n1928 ;
  assign n55252 = ( n2093 & n6000 ) | ( n2093 & ~n9429 ) | ( n6000 & ~n9429 ) ;
  assign n55253 = n55252 ^ n11710 ^ n11494 ;
  assign n55254 = n55253 ^ n14563 ^ n9411 ;
  assign n55256 = ( ~n22941 & n34510 ) | ( ~n22941 & n35190 ) | ( n34510 & n35190 ) ;
  assign n55255 = ~n14828 & n16592 ;
  assign n55257 = n55256 ^ n55255 ^ 1'b0 ;
  assign n55258 = n46007 ^ n16991 ^ n6528 ;
  assign n55259 = ( ~n7354 & n13068 ) | ( ~n7354 & n55258 ) | ( n13068 & n55258 ) ;
  assign n55260 = ( n3841 & n26666 ) | ( n3841 & n44711 ) | ( n26666 & n44711 ) ;
  assign n55261 = ~n5949 & n29946 ;
  assign n55262 = ( n8065 & ~n18542 ) | ( n8065 & n40050 ) | ( ~n18542 & n40050 ) ;
  assign n55263 = n55262 ^ n47701 ^ n21974 ;
  assign n55264 = n7497 ^ n3334 ^ 1'b0 ;
  assign n55265 = ~n26859 & n55264 ;
  assign n55266 = n55265 ^ n19867 ^ n12262 ;
  assign n55267 = n41249 ^ n19806 ^ n11970 ;
  assign n55268 = ( n11037 & n27093 ) | ( n11037 & ~n51692 ) | ( n27093 & ~n51692 ) ;
  assign n55271 = n21730 ^ n19868 ^ n15559 ;
  assign n55272 = n55271 ^ n34005 ^ n11652 ;
  assign n55269 = n13953 ^ n3744 ^ n1833 ;
  assign n55270 = n55269 ^ n33956 ^ n4726 ;
  assign n55273 = n55272 ^ n55270 ^ n38989 ;
  assign n55274 = ~n10954 & n21804 ;
  assign n55275 = n17484 & n55274 ;
  assign n55276 = n55275 ^ n47420 ^ n17927 ;
  assign n55278 = n10809 & ~n25517 ;
  assign n55277 = n13770 & ~n46407 ;
  assign n55279 = n55278 ^ n55277 ^ 1'b0 ;
  assign n55280 = n25542 ^ n18461 ^ n4308 ;
  assign n55281 = ( ~n3728 & n16535 ) | ( ~n3728 & n28067 ) | ( n16535 & n28067 ) ;
  assign n55282 = n55281 ^ n54620 ^ n45319 ;
  assign n55283 = ~n29772 & n46871 ;
  assign n55284 = n48798 ^ n42237 ^ n28586 ;
  assign n55285 = ( n20470 & n37555 ) | ( n20470 & n52293 ) | ( n37555 & n52293 ) ;
  assign n55286 = n33862 ^ n2838 ^ 1'b0 ;
  assign n55287 = ( n6259 & n25371 ) | ( n6259 & ~n28096 ) | ( n25371 & ~n28096 ) ;
  assign n55288 = ( n12937 & n15241 ) | ( n12937 & n55287 ) | ( n15241 & n55287 ) ;
  assign n55289 = n28407 ^ n15062 ^ n7563 ;
  assign n55290 = n34131 ^ n25106 ^ n23825 ;
  assign n55291 = n55290 ^ n51460 ^ n18511 ;
  assign n55292 = ( n18494 & ~n19039 ) | ( n18494 & n55291 ) | ( ~n19039 & n55291 ) ;
  assign n55293 = n11040 & n24059 ;
  assign n55294 = n1741 & ~n6188 ;
  assign n55295 = ~n33619 & n55294 ;
  assign n55296 = n36450 ^ n25398 ^ n12481 ;
  assign n55297 = n37044 ^ n30961 ^ n16445 ;
  assign n55302 = n28596 ^ n18281 ^ n2657 ;
  assign n55298 = n6248 ^ n2344 ^ n290 ;
  assign n55299 = n50247 ^ n1148 ^ 1'b0 ;
  assign n55300 = ~n24334 & n55299 ;
  assign n55301 = ( ~n35874 & n55298 ) | ( ~n35874 & n55300 ) | ( n55298 & n55300 ) ;
  assign n55303 = n55302 ^ n55301 ^ n26894 ;
  assign n55304 = ( n3755 & n13349 ) | ( n3755 & n17708 ) | ( n13349 & n17708 ) ;
  assign n55305 = n33549 ^ n30374 ^ n10988 ;
  assign n55306 = ( n12138 & ~n52841 ) | ( n12138 & n55305 ) | ( ~n52841 & n55305 ) ;
  assign n55307 = ( n55303 & n55304 ) | ( n55303 & ~n55306 ) | ( n55304 & ~n55306 ) ;
  assign n55308 = n22294 ^ n11241 ^ n3322 ;
  assign n55309 = n55308 ^ n13529 ^ n5171 ;
  assign n55310 = n36884 ^ n19738 ^ 1'b0 ;
  assign n55311 = n14866 & n55310 ;
  assign n55312 = ( n26039 & ~n55309 ) | ( n26039 & n55311 ) | ( ~n55309 & n55311 ) ;
  assign n55314 = ( n1315 & n3240 ) | ( n1315 & ~n4378 ) | ( n3240 & ~n4378 ) ;
  assign n55315 = ( ~n41638 & n47599 ) | ( ~n41638 & n55314 ) | ( n47599 & n55314 ) ;
  assign n55313 = ( n18472 & ~n34302 ) | ( n18472 & n54688 ) | ( ~n34302 & n54688 ) ;
  assign n55316 = n55315 ^ n55313 ^ n17365 ;
  assign n55317 = ( n2018 & ~n38700 ) | ( n2018 & n47600 ) | ( ~n38700 & n47600 ) ;
  assign n55318 = n55317 ^ n10404 ^ 1'b0 ;
  assign n55319 = n41281 & n55318 ;
  assign n55320 = n55319 ^ n15844 ^ n12413 ;
  assign n55321 = n27924 ^ n16252 ^ n11982 ;
  assign n55322 = ( n15463 & n25377 ) | ( n15463 & ~n27568 ) | ( n25377 & ~n27568 ) ;
  assign n55323 = ( ~n23285 & n40844 ) | ( ~n23285 & n55322 ) | ( n40844 & n55322 ) ;
  assign n55324 = n55323 ^ n27686 ^ n21018 ;
  assign n55325 = ( n6824 & n16383 ) | ( n6824 & ~n44209 ) | ( n16383 & ~n44209 ) ;
  assign n55326 = n55325 ^ n13893 ^ n2652 ;
  assign n55327 = n16966 ^ n4914 ^ n3152 ;
  assign n55328 = ( ~n2148 & n28271 ) | ( ~n2148 & n42010 ) | ( n28271 & n42010 ) ;
  assign n55329 = n55328 ^ n15081 ^ 1'b0 ;
  assign n55330 = n55327 & ~n55329 ;
  assign n55331 = ( n22625 & n30615 ) | ( n22625 & n43205 ) | ( n30615 & n43205 ) ;
  assign n55332 = n26926 ^ n6037 ^ n2228 ;
  assign n55333 = n27322 ^ n4020 ^ n3809 ;
  assign n55334 = n38692 ^ n30872 ^ n2076 ;
  assign n55335 = n807 & n6937 ;
  assign n55336 = n55335 ^ n2867 ^ 1'b0 ;
  assign n55337 = ( n11364 & n28884 ) | ( n11364 & n52169 ) | ( n28884 & n52169 ) ;
  assign n55338 = ( n34860 & n55336 ) | ( n34860 & ~n55337 ) | ( n55336 & ~n55337 ) ;
  assign n55339 = n13437 ^ n9407 ^ 1'b0 ;
  assign n55340 = n24017 ^ n17327 ^ n1996 ;
  assign n55341 = ( n8515 & ~n46448 ) | ( n8515 & n55340 ) | ( ~n46448 & n55340 ) ;
  assign n55342 = ( ~n8803 & n55339 ) | ( ~n8803 & n55341 ) | ( n55339 & n55341 ) ;
  assign n55343 = n40991 ^ n36364 ^ n1153 ;
  assign n55344 = ( n6962 & ~n11267 ) | ( n6962 & n28236 ) | ( ~n11267 & n28236 ) ;
  assign n55345 = n55344 ^ n16589 ^ n7759 ;
  assign n55346 = n45096 ^ n22276 ^ 1'b0 ;
  assign n55347 = n2986 & ~n55346 ;
  assign n55348 = n55347 ^ n21888 ^ 1'b0 ;
  assign n55349 = n52321 ^ n39619 ^ n14230 ;
  assign n55350 = ( n16876 & ~n19746 ) | ( n16876 & n27176 ) | ( ~n19746 & n27176 ) ;
  assign n55351 = ( n28327 & n29495 ) | ( n28327 & ~n55350 ) | ( n29495 & ~n55350 ) ;
  assign n55355 = ( n2094 & ~n9197 ) | ( n2094 & n12933 ) | ( ~n9197 & n12933 ) ;
  assign n55356 = n55355 ^ n44157 ^ n33552 ;
  assign n55352 = ( n2944 & ~n3648 ) | ( n2944 & n28872 ) | ( ~n3648 & n28872 ) ;
  assign n55353 = n3241 | n55352 ;
  assign n55354 = n38846 & ~n55353 ;
  assign n55357 = n55356 ^ n55354 ^ n18105 ;
  assign n55358 = ( n5585 & n18904 ) | ( n5585 & n49839 ) | ( n18904 & n49839 ) ;
  assign n55360 = ( n10841 & n26288 ) | ( n10841 & ~n43078 ) | ( n26288 & ~n43078 ) ;
  assign n55359 = n2110 & n10434 ;
  assign n55361 = n55360 ^ n55359 ^ 1'b0 ;
  assign n55362 = n55361 ^ n9688 ^ n8485 ;
  assign n55363 = ( n21695 & n34761 ) | ( n21695 & ~n47400 ) | ( n34761 & ~n47400 ) ;
  assign n55364 = ( ~n2736 & n7797 ) | ( ~n2736 & n19440 ) | ( n7797 & n19440 ) ;
  assign n55365 = ( n39616 & n54927 ) | ( n39616 & n55364 ) | ( n54927 & n55364 ) ;
  assign n55366 = ~n358 & n28295 ;
  assign n55367 = n55366 ^ n46432 ^ 1'b0 ;
  assign n55368 = ( n15314 & n51132 ) | ( n15314 & n55367 ) | ( n51132 & n55367 ) ;
  assign y0 = x8 ;
  assign y1 = x9 ;
  assign y2 = x16 ;
  assign y3 = x34 ;
  assign y4 = x43 ;
  assign y5 = x70 ;
  assign y6 = x85 ;
  assign y7 = x87 ;
  assign y8 = x95 ;
  assign y9 = x105 ;
  assign y10 = x121 ;
  assign y11 = x129 ;
  assign y12 = x134 ;
  assign y13 = x153 ;
  assign y14 = x154 ;
  assign y15 = x177 ;
  assign y16 = x180 ;
  assign y17 = x182 ;
  assign y18 = x186 ;
  assign y19 = x188 ;
  assign y20 = x217 ;
  assign y21 = x218 ;
  assign y22 = x232 ;
  assign y23 = x234 ;
  assign y24 = x241 ;
  assign y25 = x244 ;
  assign y26 = n256 ;
  assign y27 = n260 ;
  assign y28 = n263 ;
  assign y29 = n265 ;
  assign y30 = ~n271 ;
  assign y31 = ~n275 ;
  assign y32 = ~n276 ;
  assign y33 = n278 ;
  assign y34 = n283 ;
  assign y35 = n284 ;
  assign y36 = ~n285 ;
  assign y37 = ~n291 ;
  assign y38 = ~n294 ;
  assign y39 = n297 ;
  assign y40 = ~n301 ;
  assign y41 = n305 ;
  assign y42 = n311 ;
  assign y43 = ~n314 ;
  assign y44 = ~n319 ;
  assign y45 = n325 ;
  assign y46 = n332 ;
  assign y47 = ~n336 ;
  assign y48 = n338 ;
  assign y49 = n342 ;
  assign y50 = n347 ;
  assign y51 = ~n349 ;
  assign y52 = n354 ;
  assign y53 = ~n358 ;
  assign y54 = ~1'b0 ;
  assign y55 = n365 ;
  assign y56 = n368 ;
  assign y57 = ~n372 ;
  assign y58 = n374 ;
  assign y59 = n375 ;
  assign y60 = ~n376 ;
  assign y61 = ~n382 ;
  assign y62 = ~n387 ;
  assign y63 = n400 ;
  assign y64 = n403 ;
  assign y65 = n415 ;
  assign y66 = ~n437 ;
  assign y67 = ~n448 ;
  assign y68 = ~n454 ;
  assign y69 = n463 ;
  assign y70 = ~n466 ;
  assign y71 = ~n468 ;
  assign y72 = n478 ;
  assign y73 = n480 ;
  assign y74 = ~n485 ;
  assign y75 = ~1'b0 ;
  assign y76 = ~n489 ;
  assign y77 = n497 ;
  assign y78 = ~n501 ;
  assign y79 = ~n515 ;
  assign y80 = ~n519 ;
  assign y81 = n521 ;
  assign y82 = ~n522 ;
  assign y83 = ~n548 ;
  assign y84 = n550 ;
  assign y85 = n554 ;
  assign y86 = ~n555 ;
  assign y87 = n560 ;
  assign y88 = n568 ;
  assign y89 = ~n582 ;
  assign y90 = ~1'b0 ;
  assign y91 = ~n585 ;
  assign y92 = n588 ;
  assign y93 = n599 ;
  assign y94 = ~n604 ;
  assign y95 = ~n623 ;
  assign y96 = n626 ;
  assign y97 = n632 ;
  assign y98 = ~n639 ;
  assign y99 = ~1'b0 ;
  assign y100 = ~n668 ;
  assign y101 = ~n679 ;
  assign y102 = ~n684 ;
  assign y103 = ~n691 ;
  assign y104 = ~n701 ;
  assign y105 = ~n703 ;
  assign y106 = n710 ;
  assign y107 = ~n716 ;
  assign y108 = n722 ;
  assign y109 = n728 ;
  assign y110 = n742 ;
  assign y111 = ~n743 ;
  assign y112 = ~n765 ;
  assign y113 = ~1'b0 ;
  assign y114 = ~n768 ;
  assign y115 = ~n774 ;
  assign y116 = n784 ;
  assign y117 = ~n794 ;
  assign y118 = ~n808 ;
  assign y119 = ~n812 ;
  assign y120 = n813 ;
  assign y121 = n815 ;
  assign y122 = n824 ;
  assign y123 = n825 ;
  assign y124 = n830 ;
  assign y125 = ~n831 ;
  assign y126 = n835 ;
  assign y127 = n836 ;
  assign y128 = ~n850 ;
  assign y129 = n851 ;
  assign y130 = ~n858 ;
  assign y131 = ~n860 ;
  assign y132 = n872 ;
  assign y133 = ~n878 ;
  assign y134 = n888 ;
  assign y135 = ~n902 ;
  assign y136 = n906 ;
  assign y137 = ~1'b0 ;
  assign y138 = ~n916 ;
  assign y139 = ~n926 ;
  assign y140 = ~n929 ;
  assign y141 = n935 ;
  assign y142 = n936 ;
  assign y143 = n975 ;
  assign y144 = n978 ;
  assign y145 = ~1'b0 ;
  assign y146 = ~n984 ;
  assign y147 = n1003 ;
  assign y148 = n1012 ;
  assign y149 = ~n1030 ;
  assign y150 = n1041 ;
  assign y151 = ~n1051 ;
  assign y152 = ~n1054 ;
  assign y153 = ~n1065 ;
  assign y154 = n1083 ;
  assign y155 = n1085 ;
  assign y156 = ~n1093 ;
  assign y157 = ~n1094 ;
  assign y158 = ~n1096 ;
  assign y159 = n1097 ;
  assign y160 = n1099 ;
  assign y161 = n1104 ;
  assign y162 = ~n1107 ;
  assign y163 = n1109 ;
  assign y164 = n1114 ;
  assign y165 = n1117 ;
  assign y166 = ~n1125 ;
  assign y167 = ~n1134 ;
  assign y168 = ~n1147 ;
  assign y169 = n1148 ;
  assign y170 = n1157 ;
  assign y171 = ~n1169 ;
  assign y172 = ~n1172 ;
  assign y173 = ~n1174 ;
  assign y174 = ~n1183 ;
  assign y175 = ~n1192 ;
  assign y176 = n1201 ;
  assign y177 = n1206 ;
  assign y178 = ~n1207 ;
  assign y179 = ~n1210 ;
  assign y180 = ~n1229 ;
  assign y181 = n1235 ;
  assign y182 = ~n1240 ;
  assign y183 = ~n1247 ;
  assign y184 = ~1'b0 ;
  assign y185 = n1258 ;
  assign y186 = ~n1260 ;
  assign y187 = ~n1271 ;
  assign y188 = ~1'b0 ;
  assign y189 = ~n1272 ;
  assign y190 = ~x66 ;
  assign y191 = ~n1281 ;
  assign y192 = n1287 ;
  assign y193 = ~n1290 ;
  assign y194 = n1303 ;
  assign y195 = ~n1312 ;
  assign y196 = ~n1327 ;
  assign y197 = n1335 ;
  assign y198 = ~1'b0 ;
  assign y199 = n1339 ;
  assign y200 = ~n1341 ;
  assign y201 = ~n1347 ;
  assign y202 = ~n1355 ;
  assign y203 = n1360 ;
  assign y204 = ~1'b0 ;
  assign y205 = n1364 ;
  assign y206 = n1375 ;
  assign y207 = n1389 ;
  assign y208 = n1398 ;
  assign y209 = ~n1399 ;
  assign y210 = n1404 ;
  assign y211 = ~n1407 ;
  assign y212 = ~n1425 ;
  assign y213 = ~n1447 ;
  assign y214 = n1449 ;
  assign y215 = ~n1456 ;
  assign y216 = ~n1463 ;
  assign y217 = ~n1470 ;
  assign y218 = ~n1476 ;
  assign y219 = ~n1492 ;
  assign y220 = ~n1495 ;
  assign y221 = ~n1507 ;
  assign y222 = ~n1510 ;
  assign y223 = ~n1529 ;
  assign y224 = n1541 ;
  assign y225 = ~1'b0 ;
  assign y226 = n1546 ;
  assign y227 = n1548 ;
  assign y228 = ~n1550 ;
  assign y229 = n1562 ;
  assign y230 = ~n1585 ;
  assign y231 = n1588 ;
  assign y232 = ~n1598 ;
  assign y233 = ~n1603 ;
  assign y234 = n1611 ;
  assign y235 = n1617 ;
  assign y236 = n1630 ;
  assign y237 = ~n1636 ;
  assign y238 = ~n1639 ;
  assign y239 = n1652 ;
  assign y240 = ~n1655 ;
  assign y241 = n1664 ;
  assign y242 = n1672 ;
  assign y243 = n1681 ;
  assign y244 = n1682 ;
  assign y245 = ~n1687 ;
  assign y246 = n1689 ;
  assign y247 = ~1'b0 ;
  assign y248 = ~n1691 ;
  assign y249 = ~n1701 ;
  assign y250 = n1727 ;
  assign y251 = ~n1734 ;
  assign y252 = ~1'b0 ;
  assign y253 = ~n1756 ;
  assign y254 = n1780 ;
  assign y255 = ~n1784 ;
  assign y256 = n1789 ;
  assign y257 = n1795 ;
  assign y258 = ~n1804 ;
  assign y259 = n1805 ;
  assign y260 = ~n1808 ;
  assign y261 = n1812 ;
  assign y262 = n1813 ;
  assign y263 = ~n1824 ;
  assign y264 = n1834 ;
  assign y265 = n1840 ;
  assign y266 = n1852 ;
  assign y267 = ~n1853 ;
  assign y268 = ~n1864 ;
  assign y269 = ~n1873 ;
  assign y270 = n1879 ;
  assign y271 = n1889 ;
  assign y272 = n1906 ;
  assign y273 = n1907 ;
  assign y274 = ~1'b0 ;
  assign y275 = ~n1933 ;
  assign y276 = ~n1934 ;
  assign y277 = ~n1938 ;
  assign y278 = n1944 ;
  assign y279 = ~n1945 ;
  assign y280 = n1949 ;
  assign y281 = ~n1965 ;
  assign y282 = n1972 ;
  assign y283 = n1976 ;
  assign y284 = n1982 ;
  assign y285 = n1986 ;
  assign y286 = n1987 ;
  assign y287 = ~n2000 ;
  assign y288 = n2010 ;
  assign y289 = n2026 ;
  assign y290 = n2029 ;
  assign y291 = ~n2035 ;
  assign y292 = ~n2055 ;
  assign y293 = n2061 ;
  assign y294 = n2064 ;
  assign y295 = ~n2074 ;
  assign y296 = n2077 ;
  assign y297 = ~n2087 ;
  assign y298 = ~n2104 ;
  assign y299 = n2124 ;
  assign y300 = n2129 ;
  assign y301 = ~n2130 ;
  assign y302 = ~n2134 ;
  assign y303 = n2139 ;
  assign y304 = n2166 ;
  assign y305 = ~n2167 ;
  assign y306 = ~1'b0 ;
  assign y307 = n2176 ;
  assign y308 = ~n2178 ;
  assign y309 = n2179 ;
  assign y310 = n2190 ;
  assign y311 = ~n2223 ;
  assign y312 = ~n2244 ;
  assign y313 = ~n2249 ;
  assign y314 = ~n2262 ;
  assign y315 = ~n2264 ;
  assign y316 = ~n2269 ;
  assign y317 = n2307 ;
  assign y318 = n2323 ;
  assign y319 = ~n2325 ;
  assign y320 = n2348 ;
  assign y321 = ~n2355 ;
  assign y322 = ~1'b0 ;
  assign y323 = n2388 ;
  assign y324 = ~n2392 ;
  assign y325 = ~n2408 ;
  assign y326 = n2412 ;
  assign y327 = ~n2415 ;
  assign y328 = n2426 ;
  assign y329 = ~n2434 ;
  assign y330 = ~n2440 ;
  assign y331 = ~n2443 ;
  assign y332 = n2448 ;
  assign y333 = n2454 ;
  assign y334 = n2461 ;
  assign y335 = ~n2466 ;
  assign y336 = ~n2467 ;
  assign y337 = n2475 ;
  assign y338 = n2498 ;
  assign y339 = n2500 ;
  assign y340 = n2502 ;
  assign y341 = n2507 ;
  assign y342 = ~n2513 ;
  assign y343 = ~n2516 ;
  assign y344 = n2518 ;
  assign y345 = n2524 ;
  assign y346 = ~1'b0 ;
  assign y347 = n2540 ;
  assign y348 = n2550 ;
  assign y349 = n2563 ;
  assign y350 = ~n2566 ;
  assign y351 = ~n2577 ;
  assign y352 = ~n2584 ;
  assign y353 = n2588 ;
  assign y354 = ~n2593 ;
  assign y355 = n2607 ;
  assign y356 = ~1'b0 ;
  assign y357 = ~n2609 ;
  assign y358 = ~n2616 ;
  assign y359 = n2631 ;
  assign y360 = ~n2636 ;
  assign y361 = n2641 ;
  assign y362 = ~n2645 ;
  assign y363 = n2653 ;
  assign y364 = ~n2664 ;
  assign y365 = n2671 ;
  assign y366 = n2684 ;
  assign y367 = n2685 ;
  assign y368 = ~n2688 ;
  assign y369 = ~n2697 ;
  assign y370 = ~n2708 ;
  assign y371 = ~n2712 ;
  assign y372 = n2729 ;
  assign y373 = ~n2753 ;
  assign y374 = ~n2756 ;
  assign y375 = ~n2764 ;
  assign y376 = n2778 ;
  assign y377 = n2787 ;
  assign y378 = ~n2788 ;
  assign y379 = n2791 ;
  assign y380 = ~n2806 ;
  assign y381 = n2808 ;
  assign y382 = ~n2814 ;
  assign y383 = ~n2820 ;
  assign y384 = n2841 ;
  assign y385 = ~n2846 ;
  assign y386 = ~n2852 ;
  assign y387 = n2857 ;
  assign y388 = n2859 ;
  assign y389 = ~n2868 ;
  assign y390 = n2887 ;
  assign y391 = n2897 ;
  assign y392 = n2901 ;
  assign y393 = n2909 ;
  assign y394 = n2918 ;
  assign y395 = n2923 ;
  assign y396 = n2933 ;
  assign y397 = n2947 ;
  assign y398 = ~n2948 ;
  assign y399 = n2954 ;
  assign y400 = ~n2964 ;
  assign y401 = n2965 ;
  assign y402 = n2970 ;
  assign y403 = n2976 ;
  assign y404 = n2986 ;
  assign y405 = n2999 ;
  assign y406 = n3020 ;
  assign y407 = ~n3030 ;
  assign y408 = n3032 ;
  assign y409 = n3039 ;
  assign y410 = ~1'b0 ;
  assign y411 = n3050 ;
  assign y412 = ~n3059 ;
  assign y413 = ~n3068 ;
  assign y414 = ~1'b0 ;
  assign y415 = n3075 ;
  assign y416 = n3078 ;
  assign y417 = ~n3087 ;
  assign y418 = n3093 ;
  assign y419 = n3104 ;
  assign y420 = ~n3107 ;
  assign y421 = n3114 ;
  assign y422 = ~n3118 ;
  assign y423 = n3121 ;
  assign y424 = ~n3129 ;
  assign y425 = ~n3137 ;
  assign y426 = ~n3150 ;
  assign y427 = n3155 ;
  assign y428 = n3158 ;
  assign y429 = n3160 ;
  assign y430 = n3170 ;
  assign y431 = ~n3182 ;
  assign y432 = ~n3189 ;
  assign y433 = n3197 ;
  assign y434 = n3209 ;
  assign y435 = ~n3215 ;
  assign y436 = n3227 ;
  assign y437 = n3229 ;
  assign y438 = ~n3239 ;
  assign y439 = ~n3241 ;
  assign y440 = n3253 ;
  assign y441 = n3254 ;
  assign y442 = n3257 ;
  assign y443 = ~n3267 ;
  assign y444 = n3271 ;
  assign y445 = n3274 ;
  assign y446 = ~n3278 ;
  assign y447 = ~n3281 ;
  assign y448 = n3291 ;
  assign y449 = n3298 ;
  assign y450 = n3313 ;
  assign y451 = ~n3327 ;
  assign y452 = ~n3334 ;
  assign y453 = ~n3344 ;
  assign y454 = n3349 ;
  assign y455 = ~n3354 ;
  assign y456 = ~1'b0 ;
  assign y457 = ~n3361 ;
  assign y458 = ~1'b0 ;
  assign y459 = n3370 ;
  assign y460 = ~n3371 ;
  assign y461 = ~n3380 ;
  assign y462 = ~n3386 ;
  assign y463 = ~1'b0 ;
  assign y464 = n3392 ;
  assign y465 = n3399 ;
  assign y466 = ~n3403 ;
  assign y467 = ~n3409 ;
  assign y468 = ~n3416 ;
  assign y469 = n3427 ;
  assign y470 = ~n3439 ;
  assign y471 = ~n3440 ;
  assign y472 = n3450 ;
  assign y473 = ~1'b0 ;
  assign y474 = n3456 ;
  assign y475 = n3473 ;
  assign y476 = n3476 ;
  assign y477 = n3493 ;
  assign y478 = n3495 ;
  assign y479 = ~n3499 ;
  assign y480 = ~n3505 ;
  assign y481 = ~n3506 ;
  assign y482 = n3507 ;
  assign y483 = n3510 ;
  assign y484 = n3521 ;
  assign y485 = n3528 ;
  assign y486 = n3545 ;
  assign y487 = n3549 ;
  assign y488 = ~n3555 ;
  assign y489 = n3557 ;
  assign y490 = ~n3562 ;
  assign y491 = n3568 ;
  assign y492 = ~n3582 ;
  assign y493 = ~n3587 ;
  assign y494 = ~n3591 ;
  assign y495 = ~n3597 ;
  assign y496 = ~n3607 ;
  assign y497 = n3608 ;
  assign y498 = ~n3610 ;
  assign y499 = n3622 ;
  assign y500 = n3624 ;
  assign y501 = n3637 ;
  assign y502 = n3642 ;
  assign y503 = ~n3665 ;
  assign y504 = ~n3681 ;
  assign y505 = n3683 ;
  assign y506 = n3690 ;
  assign y507 = ~n3738 ;
  assign y508 = ~n3741 ;
  assign y509 = ~n3784 ;
  assign y510 = ~n3787 ;
  assign y511 = n3800 ;
  assign y512 = n3808 ;
  assign y513 = ~1'b0 ;
  assign y514 = ~n3827 ;
  assign y515 = ~n3833 ;
  assign y516 = n3845 ;
  assign y517 = ~n3846 ;
  assign y518 = n3847 ;
  assign y519 = ~n3855 ;
  assign y520 = n3860 ;
  assign y521 = ~n3867 ;
  assign y522 = n3868 ;
  assign y523 = ~n3873 ;
  assign y524 = ~n3883 ;
  assign y525 = ~n3890 ;
  assign y526 = n3898 ;
  assign y527 = ~n3906 ;
  assign y528 = ~1'b0 ;
  assign y529 = n3916 ;
  assign y530 = n3926 ;
  assign y531 = n3929 ;
  assign y532 = n3937 ;
  assign y533 = ~1'b0 ;
  assign y534 = n3939 ;
  assign y535 = n3966 ;
  assign y536 = n3983 ;
  assign y537 = ~n3987 ;
  assign y538 = ~n3996 ;
  assign y539 = n4000 ;
  assign y540 = ~n4008 ;
  assign y541 = ~1'b0 ;
  assign y542 = ~n4021 ;
  assign y543 = n4028 ;
  assign y544 = ~n4033 ;
  assign y545 = n4047 ;
  assign y546 = n4078 ;
  assign y547 = n4103 ;
  assign y548 = n4122 ;
  assign y549 = ~n4125 ;
  assign y550 = ~n4135 ;
  assign y551 = n4137 ;
  assign y552 = ~n4142 ;
  assign y553 = n4153 ;
  assign y554 = ~n4155 ;
  assign y555 = ~n4157 ;
  assign y556 = ~n4166 ;
  assign y557 = ~n4185 ;
  assign y558 = n4203 ;
  assign y559 = n4207 ;
  assign y560 = n4211 ;
  assign y561 = ~n4221 ;
  assign y562 = ~n4229 ;
  assign y563 = ~n4243 ;
  assign y564 = n4256 ;
  assign y565 = n4264 ;
  assign y566 = ~n4269 ;
  assign y567 = n4274 ;
  assign y568 = n4279 ;
  assign y569 = n4290 ;
  assign y570 = n4305 ;
  assign y571 = n4312 ;
  assign y572 = ~n4315 ;
  assign y573 = n4318 ;
  assign y574 = ~n4327 ;
  assign y575 = ~n4335 ;
  assign y576 = n4339 ;
  assign y577 = ~n4343 ;
  assign y578 = ~n4346 ;
  assign y579 = ~n4356 ;
  assign y580 = n4363 ;
  assign y581 = n4369 ;
  assign y582 = n4374 ;
  assign y583 = ~n4379 ;
  assign y584 = n4384 ;
  assign y585 = n4386 ;
  assign y586 = n4407 ;
  assign y587 = n4414 ;
  assign y588 = ~n4425 ;
  assign y589 = ~n4435 ;
  assign y590 = n4437 ;
  assign y591 = n4442 ;
  assign y592 = n4478 ;
  assign y593 = n4499 ;
  assign y594 = ~n4506 ;
  assign y595 = ~n4513 ;
  assign y596 = ~n4515 ;
  assign y597 = n4516 ;
  assign y598 = ~n4519 ;
  assign y599 = ~n4531 ;
  assign y600 = n4532 ;
  assign y601 = ~n4534 ;
  assign y602 = n4535 ;
  assign y603 = ~n4548 ;
  assign y604 = n4558 ;
  assign y605 = ~n4569 ;
  assign y606 = n4587 ;
  assign y607 = ~n4592 ;
  assign y608 = ~n4603 ;
  assign y609 = n4607 ;
  assign y610 = n4618 ;
  assign y611 = ~n4642 ;
  assign y612 = ~n4653 ;
  assign y613 = n4662 ;
  assign y614 = n4674 ;
  assign y615 = ~n4683 ;
  assign y616 = ~n4684 ;
  assign y617 = n4695 ;
  assign y618 = ~n4697 ;
  assign y619 = n4699 ;
  assign y620 = ~n4703 ;
  assign y621 = ~n4711 ;
  assign y622 = n4713 ;
  assign y623 = n4721 ;
  assign y624 = ~n4723 ;
  assign y625 = ~1'b0 ;
  assign y626 = n4736 ;
  assign y627 = ~n4754 ;
  assign y628 = ~n4760 ;
  assign y629 = ~n4762 ;
  assign y630 = ~n4767 ;
  assign y631 = n4777 ;
  assign y632 = n4781 ;
  assign y633 = n4785 ;
  assign y634 = ~n4797 ;
  assign y635 = ~n4799 ;
  assign y636 = n4806 ;
  assign y637 = n4821 ;
  assign y638 = ~1'b0 ;
  assign y639 = ~n4827 ;
  assign y640 = n4844 ;
  assign y641 = ~n4845 ;
  assign y642 = n4849 ;
  assign y643 = n4854 ;
  assign y644 = ~n4873 ;
  assign y645 = n4883 ;
  assign y646 = n4888 ;
  assign y647 = n4894 ;
  assign y648 = ~n4901 ;
  assign y649 = ~n4912 ;
  assign y650 = ~n4921 ;
  assign y651 = ~n4927 ;
  assign y652 = n4938 ;
  assign y653 = n4942 ;
  assign y654 = ~n4957 ;
  assign y655 = n4963 ;
  assign y656 = ~n4968 ;
  assign y657 = ~n4975 ;
  assign y658 = ~n4996 ;
  assign y659 = n5001 ;
  assign y660 = ~n5012 ;
  assign y661 = ~n5015 ;
  assign y662 = n5037 ;
  assign y663 = ~n5042 ;
  assign y664 = n5068 ;
  assign y665 = ~n5077 ;
  assign y666 = n5079 ;
  assign y667 = n5081 ;
  assign y668 = ~n5088 ;
  assign y669 = ~n5099 ;
  assign y670 = ~n5111 ;
  assign y671 = n5120 ;
  assign y672 = n5125 ;
  assign y673 = ~n5129 ;
  assign y674 = n5133 ;
  assign y675 = n5138 ;
  assign y676 = ~n5154 ;
  assign y677 = n5157 ;
  assign y678 = n5166 ;
  assign y679 = ~1'b0 ;
  assign y680 = ~n5170 ;
  assign y681 = ~1'b0 ;
  assign y682 = ~n5173 ;
  assign y683 = n5174 ;
  assign y684 = ~1'b0 ;
  assign y685 = n5186 ;
  assign y686 = n5193 ;
  assign y687 = n5198 ;
  assign y688 = n5207 ;
  assign y689 = n5208 ;
  assign y690 = ~n5231 ;
  assign y691 = ~n5243 ;
  assign y692 = ~n5256 ;
  assign y693 = n5260 ;
  assign y694 = n5261 ;
  assign y695 = ~n5271 ;
  assign y696 = n5273 ;
  assign y697 = ~1'b0 ;
  assign y698 = ~n5281 ;
  assign y699 = n5282 ;
  assign y700 = n5295 ;
  assign y701 = ~n5318 ;
  assign y702 = ~n5325 ;
  assign y703 = n5328 ;
  assign y704 = n5348 ;
  assign y705 = n5353 ;
  assign y706 = ~n5354 ;
  assign y707 = ~n5360 ;
  assign y708 = ~n5363 ;
  assign y709 = n5364 ;
  assign y710 = n5365 ;
  assign y711 = n5373 ;
  assign y712 = ~n5385 ;
  assign y713 = n5400 ;
  assign y714 = ~n5402 ;
  assign y715 = ~n5404 ;
  assign y716 = ~n5406 ;
  assign y717 = ~n5409 ;
  assign y718 = ~n5412 ;
  assign y719 = ~n5418 ;
  assign y720 = ~n5423 ;
  assign y721 = n5425 ;
  assign y722 = ~n5441 ;
  assign y723 = n5451 ;
  assign y724 = ~n5458 ;
  assign y725 = n5465 ;
  assign y726 = n5472 ;
  assign y727 = n5473 ;
  assign y728 = ~n5476 ;
  assign y729 = ~n5487 ;
  assign y730 = ~n5509 ;
  assign y731 = ~n5513 ;
  assign y732 = ~n5516 ;
  assign y733 = ~n5523 ;
  assign y734 = n5524 ;
  assign y735 = ~n5538 ;
  assign y736 = n5541 ;
  assign y737 = ~n5549 ;
  assign y738 = n5557 ;
  assign y739 = n5575 ;
  assign y740 = n5590 ;
  assign y741 = ~n5596 ;
  assign y742 = ~n5606 ;
  assign y743 = ~n5623 ;
  assign y744 = ~1'b0 ;
  assign y745 = n5627 ;
  assign y746 = n5632 ;
  assign y747 = ~n5640 ;
  assign y748 = ~n5641 ;
  assign y749 = ~n5643 ;
  assign y750 = n5660 ;
  assign y751 = ~n5669 ;
  assign y752 = ~n5673 ;
  assign y753 = n5679 ;
  assign y754 = ~n5686 ;
  assign y755 = ~1'b0 ;
  assign y756 = ~n5698 ;
  assign y757 = n5717 ;
  assign y758 = ~n5729 ;
  assign y759 = n5732 ;
  assign y760 = ~n5765 ;
  assign y761 = n5781 ;
  assign y762 = n5785 ;
  assign y763 = ~n5788 ;
  assign y764 = ~n5793 ;
  assign y765 = n5806 ;
  assign y766 = n5815 ;
  assign y767 = n5820 ;
  assign y768 = n5827 ;
  assign y769 = ~n5844 ;
  assign y770 = n5854 ;
  assign y771 = ~1'b0 ;
  assign y772 = n5873 ;
  assign y773 = n5879 ;
  assign y774 = n5894 ;
  assign y775 = ~n5898 ;
  assign y776 = ~1'b0 ;
  assign y777 = n5903 ;
  assign y778 = ~1'b0 ;
  assign y779 = ~n5904 ;
  assign y780 = ~n5906 ;
  assign y781 = ~1'b0 ;
  assign y782 = ~n5909 ;
  assign y783 = n5924 ;
  assign y784 = ~n5928 ;
  assign y785 = n5936 ;
  assign y786 = n5943 ;
  assign y787 = n5950 ;
  assign y788 = ~n5975 ;
  assign y789 = n5977 ;
  assign y790 = n5986 ;
  assign y791 = ~n5988 ;
  assign y792 = n5991 ;
  assign y793 = ~n6000 ;
  assign y794 = n6005 ;
  assign y795 = ~n6015 ;
  assign y796 = n6031 ;
  assign y797 = ~n6045 ;
  assign y798 = n6047 ;
  assign y799 = n6058 ;
  assign y800 = ~n6060 ;
  assign y801 = ~n6065 ;
  assign y802 = n6069 ;
  assign y803 = ~n6073 ;
  assign y804 = n6098 ;
  assign y805 = n6102 ;
  assign y806 = n6109 ;
  assign y807 = ~n6130 ;
  assign y808 = ~n6140 ;
  assign y809 = ~n6151 ;
  assign y810 = ~n6157 ;
  assign y811 = n6181 ;
  assign y812 = ~n6182 ;
  assign y813 = ~n6188 ;
  assign y814 = n6195 ;
  assign y815 = ~n6209 ;
  assign y816 = ~n6211 ;
  assign y817 = n6220 ;
  assign y818 = ~1'b0 ;
  assign y819 = n6225 ;
  assign y820 = n6243 ;
  assign y821 = ~n6247 ;
  assign y822 = n6248 ;
  assign y823 = ~n6249 ;
  assign y824 = n6258 ;
  assign y825 = ~n6271 ;
  assign y826 = ~n6273 ;
  assign y827 = n6282 ;
  assign y828 = ~n6290 ;
  assign y829 = n6297 ;
  assign y830 = n6304 ;
  assign y831 = ~n6310 ;
  assign y832 = ~n6317 ;
  assign y833 = ~n6322 ;
  assign y834 = n6333 ;
  assign y835 = ~n6342 ;
  assign y836 = ~n6349 ;
  assign y837 = n6351 ;
  assign y838 = ~n6355 ;
  assign y839 = n6368 ;
  assign y840 = n6370 ;
  assign y841 = n6372 ;
  assign y842 = ~n6376 ;
  assign y843 = n6382 ;
  assign y844 = ~n6388 ;
  assign y845 = ~n6390 ;
  assign y846 = ~n6403 ;
  assign y847 = n6411 ;
  assign y848 = ~n6419 ;
  assign y849 = ~n6431 ;
  assign y850 = ~n6437 ;
  assign y851 = ~n6441 ;
  assign y852 = n6442 ;
  assign y853 = n6444 ;
  assign y854 = ~n6448 ;
  assign y855 = n6456 ;
  assign y856 = n6459 ;
  assign y857 = n6464 ;
  assign y858 = ~n6466 ;
  assign y859 = n6470 ;
  assign y860 = n6471 ;
  assign y861 = n6505 ;
  assign y862 = ~n6507 ;
  assign y863 = n6511 ;
  assign y864 = n6522 ;
  assign y865 = n6527 ;
  assign y866 = ~n6536 ;
  assign y867 = n6563 ;
  assign y868 = ~n6564 ;
  assign y869 = ~n6569 ;
  assign y870 = n6575 ;
  assign y871 = ~n6578 ;
  assign y872 = ~n6588 ;
  assign y873 = n6593 ;
  assign y874 = ~n6611 ;
  assign y875 = n6620 ;
  assign y876 = n6629 ;
  assign y877 = ~n6637 ;
  assign y878 = n6649 ;
  assign y879 = ~n6657 ;
  assign y880 = n6661 ;
  assign y881 = ~n6677 ;
  assign y882 = n6682 ;
  assign y883 = ~n6700 ;
  assign y884 = n6703 ;
  assign y885 = n6720 ;
  assign y886 = n6723 ;
  assign y887 = n6734 ;
  assign y888 = n6739 ;
  assign y889 = ~1'b0 ;
  assign y890 = n6749 ;
  assign y891 = ~n6755 ;
  assign y892 = ~n6756 ;
  assign y893 = n6757 ;
  assign y894 = ~n6785 ;
  assign y895 = ~n6795 ;
  assign y896 = ~n6796 ;
  assign y897 = ~n6800 ;
  assign y898 = ~n6809 ;
  assign y899 = n6810 ;
  assign y900 = n6812 ;
  assign y901 = ~n6823 ;
  assign y902 = n6844 ;
  assign y903 = n6850 ;
  assign y904 = n6855 ;
  assign y905 = ~n6860 ;
  assign y906 = ~n6872 ;
  assign y907 = ~n6879 ;
  assign y908 = n6882 ;
  assign y909 = n6887 ;
  assign y910 = n6888 ;
  assign y911 = n6893 ;
  assign y912 = n6896 ;
  assign y913 = n6904 ;
  assign y914 = ~n6927 ;
  assign y915 = n6937 ;
  assign y916 = n6943 ;
  assign y917 = n6948 ;
  assign y918 = ~n6949 ;
  assign y919 = n6954 ;
  assign y920 = n953 ;
  assign y921 = ~n6961 ;
  assign y922 = n6964 ;
  assign y923 = n6970 ;
  assign y924 = n6978 ;
  assign y925 = n6983 ;
  assign y926 = n6987 ;
  assign y927 = ~n6990 ;
  assign y928 = ~n6998 ;
  assign y929 = ~n7005 ;
  assign y930 = ~n7006 ;
  assign y931 = n7013 ;
  assign y932 = n7018 ;
  assign y933 = ~n7030 ;
  assign y934 = n7034 ;
  assign y935 = ~n7036 ;
  assign y936 = ~n7042 ;
  assign y937 = n7050 ;
  assign y938 = ~1'b0 ;
  assign y939 = ~n7053 ;
  assign y940 = ~n7058 ;
  assign y941 = n7068 ;
  assign y942 = n7075 ;
  assign y943 = n7081 ;
  assign y944 = ~n7084 ;
  assign y945 = ~n7099 ;
  assign y946 = ~n7106 ;
  assign y947 = ~n7109 ;
  assign y948 = n7136 ;
  assign y949 = ~n7144 ;
  assign y950 = ~1'b0 ;
  assign y951 = ~n7152 ;
  assign y952 = n7158 ;
  assign y953 = ~n7161 ;
  assign y954 = n7172 ;
  assign y955 = ~n7191 ;
  assign y956 = n7194 ;
  assign y957 = ~n7197 ;
  assign y958 = n7198 ;
  assign y959 = n7204 ;
  assign y960 = n7209 ;
  assign y961 = n7231 ;
  assign y962 = ~n7242 ;
  assign y963 = ~n7256 ;
  assign y964 = n7257 ;
  assign y965 = n7268 ;
  assign y966 = ~n7273 ;
  assign y967 = n7274 ;
  assign y968 = ~n7275 ;
  assign y969 = n7282 ;
  assign y970 = n7301 ;
  assign y971 = n7303 ;
  assign y972 = n7310 ;
  assign y973 = ~n7315 ;
  assign y974 = ~n7323 ;
  assign y975 = ~n7326 ;
  assign y976 = ~n7349 ;
  assign y977 = n7360 ;
  assign y978 = ~n7363 ;
  assign y979 = n7371 ;
  assign y980 = ~n7374 ;
  assign y981 = ~n7375 ;
  assign y982 = n7394 ;
  assign y983 = n7402 ;
  assign y984 = n7403 ;
  assign y985 = ~n7411 ;
  assign y986 = ~1'b0 ;
  assign y987 = n7415 ;
  assign y988 = n7420 ;
  assign y989 = ~n7427 ;
  assign y990 = n7431 ;
  assign y991 = ~1'b0 ;
  assign y992 = n7439 ;
  assign y993 = ~n7446 ;
  assign y994 = ~n7460 ;
  assign y995 = n7461 ;
  assign y996 = ~1'b0 ;
  assign y997 = ~n7479 ;
  assign y998 = n7493 ;
  assign y999 = n7503 ;
  assign y1000 = ~n7535 ;
  assign y1001 = n7544 ;
  assign y1002 = n7546 ;
  assign y1003 = ~n7547 ;
  assign y1004 = n7562 ;
  assign y1005 = n7564 ;
  assign y1006 = n7569 ;
  assign y1007 = n7571 ;
  assign y1008 = n7578 ;
  assign y1009 = ~n7601 ;
  assign y1010 = n7613 ;
  assign y1011 = ~n7614 ;
  assign y1012 = ~n7617 ;
  assign y1013 = ~n7628 ;
  assign y1014 = n7629 ;
  assign y1015 = n7636 ;
  assign y1016 = ~n7638 ;
  assign y1017 = ~1'b0 ;
  assign y1018 = n7651 ;
  assign y1019 = n7659 ;
  assign y1020 = n7662 ;
  assign y1021 = n7670 ;
  assign y1022 = n7677 ;
  assign y1023 = n7678 ;
  assign y1024 = ~n7681 ;
  assign y1025 = ~n7683 ;
  assign y1026 = ~n7697 ;
  assign y1027 = ~n7709 ;
  assign y1028 = n7718 ;
  assign y1029 = ~n7724 ;
  assign y1030 = n7730 ;
  assign y1031 = ~n7742 ;
  assign y1032 = ~n7744 ;
  assign y1033 = n7751 ;
  assign y1034 = ~n7761 ;
  assign y1035 = n7763 ;
  assign y1036 = n7768 ;
  assign y1037 = ~n7769 ;
  assign y1038 = n7775 ;
  assign y1039 = ~n7778 ;
  assign y1040 = ~1'b0 ;
  assign y1041 = ~n7788 ;
  assign y1042 = ~n7792 ;
  assign y1043 = n7793 ;
  assign y1044 = ~n7803 ;
  assign y1045 = ~n7805 ;
  assign y1046 = ~n7820 ;
  assign y1047 = n7821 ;
  assign y1048 = ~1'b0 ;
  assign y1049 = ~n7827 ;
  assign y1050 = ~n7831 ;
  assign y1051 = n7834 ;
  assign y1052 = n7840 ;
  assign y1053 = n7851 ;
  assign y1054 = n7856 ;
  assign y1055 = ~1'b0 ;
  assign y1056 = n7862 ;
  assign y1057 = ~n7868 ;
  assign y1058 = n7871 ;
  assign y1059 = ~n7874 ;
  assign y1060 = ~n7876 ;
  assign y1061 = n7881 ;
  assign y1062 = ~n7900 ;
  assign y1063 = n7902 ;
  assign y1064 = n7904 ;
  assign y1065 = n7915 ;
  assign y1066 = ~n7920 ;
  assign y1067 = n7928 ;
  assign y1068 = n7937 ;
  assign y1069 = n7942 ;
  assign y1070 = n7946 ;
  assign y1071 = ~n7949 ;
  assign y1072 = ~n7960 ;
  assign y1073 = ~n7961 ;
  assign y1074 = ~n7966 ;
  assign y1075 = n7975 ;
  assign y1076 = n7984 ;
  assign y1077 = ~n7986 ;
  assign y1078 = ~n7996 ;
  assign y1079 = n8001 ;
  assign y1080 = ~n8002 ;
  assign y1081 = ~n8015 ;
  assign y1082 = n8019 ;
  assign y1083 = n8020 ;
  assign y1084 = n8023 ;
  assign y1085 = ~n8027 ;
  assign y1086 = ~n8028 ;
  assign y1087 = ~n8029 ;
  assign y1088 = ~n8034 ;
  assign y1089 = ~n8039 ;
  assign y1090 = ~n8043 ;
  assign y1091 = ~n8049 ;
  assign y1092 = n8052 ;
  assign y1093 = ~n8062 ;
  assign y1094 = n8069 ;
  assign y1095 = ~n8075 ;
  assign y1096 = ~n8076 ;
  assign y1097 = n8082 ;
  assign y1098 = ~n8094 ;
  assign y1099 = ~n8114 ;
  assign y1100 = ~n8120 ;
  assign y1101 = n8124 ;
  assign y1102 = ~n8128 ;
  assign y1103 = n8132 ;
  assign y1104 = ~n8139 ;
  assign y1105 = ~n8145 ;
  assign y1106 = ~n8148 ;
  assign y1107 = ~n8151 ;
  assign y1108 = ~n8164 ;
  assign y1109 = n8169 ;
  assign y1110 = n8175 ;
  assign y1111 = ~n8176 ;
  assign y1112 = ~n8182 ;
  assign y1113 = ~n8197 ;
  assign y1114 = n8200 ;
  assign y1115 = ~n8211 ;
  assign y1116 = ~n8219 ;
  assign y1117 = n8235 ;
  assign y1118 = n8251 ;
  assign y1119 = n8262 ;
  assign y1120 = ~n8263 ;
  assign y1121 = ~n8276 ;
  assign y1122 = ~n8287 ;
  assign y1123 = ~n8288 ;
  assign y1124 = ~n8306 ;
  assign y1125 = ~n8310 ;
  assign y1126 = n8317 ;
  assign y1127 = ~n8318 ;
  assign y1128 = n8326 ;
  assign y1129 = n8334 ;
  assign y1130 = n8343 ;
  assign y1131 = n6927 ;
  assign y1132 = ~n8360 ;
  assign y1133 = n8367 ;
  assign y1134 = n8368 ;
  assign y1135 = ~1'b0 ;
  assign y1136 = ~n8371 ;
  assign y1137 = ~1'b0 ;
  assign y1138 = ~n8382 ;
  assign y1139 = ~n8384 ;
  assign y1140 = ~n8388 ;
  assign y1141 = ~n8403 ;
  assign y1142 = ~n8410 ;
  assign y1143 = ~n8411 ;
  assign y1144 = ~n8420 ;
  assign y1145 = ~n8423 ;
  assign y1146 = n8436 ;
  assign y1147 = n8439 ;
  assign y1148 = n8443 ;
  assign y1149 = ~n8461 ;
  assign y1150 = n8471 ;
  assign y1151 = ~n8477 ;
  assign y1152 = ~n8483 ;
  assign y1153 = ~n8486 ;
  assign y1154 = n8491 ;
  assign y1155 = n8493 ;
  assign y1156 = n8507 ;
  assign y1157 = n8511 ;
  assign y1158 = n8513 ;
  assign y1159 = n8516 ;
  assign y1160 = ~n8517 ;
  assign y1161 = n8520 ;
  assign y1162 = ~1'b0 ;
  assign y1163 = ~n8528 ;
  assign y1164 = n8540 ;
  assign y1165 = ~1'b0 ;
  assign y1166 = n8550 ;
  assign y1167 = ~n8570 ;
  assign y1168 = n8580 ;
  assign y1169 = ~n8583 ;
  assign y1170 = n8590 ;
  assign y1171 = ~n8591 ;
  assign y1172 = ~n8610 ;
  assign y1173 = ~n8612 ;
  assign y1174 = ~1'b0 ;
  assign y1175 = n8624 ;
  assign y1176 = ~n8626 ;
  assign y1177 = n8638 ;
  assign y1178 = ~n8644 ;
  assign y1179 = n8648 ;
  assign y1180 = n8649 ;
  assign y1181 = n8656 ;
  assign y1182 = n8659 ;
  assign y1183 = n8672 ;
  assign y1184 = n8692 ;
  assign y1185 = n8705 ;
  assign y1186 = n8708 ;
  assign y1187 = n8713 ;
  assign y1188 = n8717 ;
  assign y1189 = ~n8726 ;
  assign y1190 = ~n8729 ;
  assign y1191 = ~n8732 ;
  assign y1192 = ~n8745 ;
  assign y1193 = ~n8754 ;
  assign y1194 = ~n8764 ;
  assign y1195 = n8771 ;
  assign y1196 = ~n8774 ;
  assign y1197 = ~n8779 ;
  assign y1198 = ~n8780 ;
  assign y1199 = n8791 ;
  assign y1200 = n8797 ;
  assign y1201 = n8800 ;
  assign y1202 = ~n8812 ;
  assign y1203 = ~n8821 ;
  assign y1204 = ~1'b0 ;
  assign y1205 = n8828 ;
  assign y1206 = ~1'b0 ;
  assign y1207 = n8837 ;
  assign y1208 = ~n8840 ;
  assign y1209 = ~n8863 ;
  assign y1210 = ~n8875 ;
  assign y1211 = ~n8878 ;
  assign y1212 = n8889 ;
  assign y1213 = ~n8893 ;
  assign y1214 = n8898 ;
  assign y1215 = ~n8905 ;
  assign y1216 = n8909 ;
  assign y1217 = n8910 ;
  assign y1218 = n8915 ;
  assign y1219 = ~n8920 ;
  assign y1220 = n8934 ;
  assign y1221 = ~n8941 ;
  assign y1222 = ~n8942 ;
  assign y1223 = ~n8972 ;
  assign y1224 = ~1'b0 ;
  assign y1225 = n8989 ;
  assign y1226 = ~n8998 ;
  assign y1227 = n9005 ;
  assign y1228 = ~n9013 ;
  assign y1229 = ~n9018 ;
  assign y1230 = n9029 ;
  assign y1231 = ~n9039 ;
  assign y1232 = ~n9045 ;
  assign y1233 = ~n9047 ;
  assign y1234 = n9058 ;
  assign y1235 = ~n9062 ;
  assign y1236 = ~n9087 ;
  assign y1237 = n9093 ;
  assign y1238 = ~n9096 ;
  assign y1239 = ~n9108 ;
  assign y1240 = ~n9111 ;
  assign y1241 = ~n9113 ;
  assign y1242 = n9118 ;
  assign y1243 = ~n9120 ;
  assign y1244 = n9123 ;
  assign y1245 = ~n9127 ;
  assign y1246 = n9130 ;
  assign y1247 = n9149 ;
  assign y1248 = ~n9150 ;
  assign y1249 = ~n9157 ;
  assign y1250 = n9161 ;
  assign y1251 = ~n9168 ;
  assign y1252 = n9170 ;
  assign y1253 = n9187 ;
  assign y1254 = n9208 ;
  assign y1255 = n9214 ;
  assign y1256 = n9228 ;
  assign y1257 = ~n9231 ;
  assign y1258 = ~n9237 ;
  assign y1259 = ~n9240 ;
  assign y1260 = ~n9246 ;
  assign y1261 = ~n9271 ;
  assign y1262 = n9272 ;
  assign y1263 = n9273 ;
  assign y1264 = n9274 ;
  assign y1265 = ~n9276 ;
  assign y1266 = ~1'b0 ;
  assign y1267 = ~n9294 ;
  assign y1268 = n9297 ;
  assign y1269 = n9304 ;
  assign y1270 = ~n9307 ;
  assign y1271 = ~n9309 ;
  assign y1272 = n9312 ;
  assign y1273 = ~n9313 ;
  assign y1274 = ~n9314 ;
  assign y1275 = ~n9321 ;
  assign y1276 = n9323 ;
  assign y1277 = n9325 ;
  assign y1278 = ~n9326 ;
  assign y1279 = n9331 ;
  assign y1280 = n9339 ;
  assign y1281 = n9340 ;
  assign y1282 = n9342 ;
  assign y1283 = n9354 ;
  assign y1284 = ~n9360 ;
  assign y1285 = ~n9363 ;
  assign y1286 = ~n9371 ;
  assign y1287 = n9375 ;
  assign y1288 = n9385 ;
  assign y1289 = ~n9388 ;
  assign y1290 = n9393 ;
  assign y1291 = n9402 ;
  assign y1292 = ~n9418 ;
  assign y1293 = ~n1194 ;
  assign y1294 = ~n9431 ;
  assign y1295 = n9432 ;
  assign y1296 = ~n9437 ;
  assign y1297 = n9439 ;
  assign y1298 = ~n9443 ;
  assign y1299 = ~1'b0 ;
  assign y1300 = n9461 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = n9467 ;
  assign y1303 = n9468 ;
  assign y1304 = ~n9476 ;
  assign y1305 = ~n9479 ;
  assign y1306 = n9490 ;
  assign y1307 = ~n9495 ;
  assign y1308 = n9503 ;
  assign y1309 = n9505 ;
  assign y1310 = ~n9511 ;
  assign y1311 = ~n9512 ;
  assign y1312 = n9516 ;
  assign y1313 = n9527 ;
  assign y1314 = n9529 ;
  assign y1315 = ~n9531 ;
  assign y1316 = ~1'b0 ;
  assign y1317 = ~n9534 ;
  assign y1318 = ~n9545 ;
  assign y1319 = ~n9548 ;
  assign y1320 = ~n9551 ;
  assign y1321 = ~n9552 ;
  assign y1322 = n9567 ;
  assign y1323 = ~n9582 ;
  assign y1324 = ~n9595 ;
  assign y1325 = n9600 ;
  assign y1326 = n9604 ;
  assign y1327 = ~n9611 ;
  assign y1328 = ~n9616 ;
  assign y1329 = ~n9620 ;
  assign y1330 = n9631 ;
  assign y1331 = ~n9651 ;
  assign y1332 = n9661 ;
  assign y1333 = ~n9665 ;
  assign y1334 = n9671 ;
  assign y1335 = n9674 ;
  assign y1336 = n9676 ;
  assign y1337 = ~n9678 ;
  assign y1338 = ~n9691 ;
  assign y1339 = ~n9695 ;
  assign y1340 = ~n9722 ;
  assign y1341 = ~n9725 ;
  assign y1342 = n9732 ;
  assign y1343 = ~n9749 ;
  assign y1344 = n9751 ;
  assign y1345 = ~n9756 ;
  assign y1346 = n9761 ;
  assign y1347 = ~1'b0 ;
  assign y1348 = n9768 ;
  assign y1349 = ~n9779 ;
  assign y1350 = ~n9787 ;
  assign y1351 = n9788 ;
  assign y1352 = n9794 ;
  assign y1353 = ~n9804 ;
  assign y1354 = n9820 ;
  assign y1355 = ~n9822 ;
  assign y1356 = ~n9828 ;
  assign y1357 = ~n9837 ;
  assign y1358 = ~n9839 ;
  assign y1359 = ~n9853 ;
  assign y1360 = n9857 ;
  assign y1361 = ~n9859 ;
  assign y1362 = n9874 ;
  assign y1363 = n9878 ;
  assign y1364 = ~n9902 ;
  assign y1365 = n9904 ;
  assign y1366 = ~n9922 ;
  assign y1367 = ~n9923 ;
  assign y1368 = n9929 ;
  assign y1369 = ~n9944 ;
  assign y1370 = n9945 ;
  assign y1371 = ~n9947 ;
  assign y1372 = ~n9965 ;
  assign y1373 = ~n9971 ;
  assign y1374 = n9975 ;
  assign y1375 = ~n9977 ;
  assign y1376 = n9982 ;
  assign y1377 = n9989 ;
  assign y1378 = ~n9990 ;
  assign y1379 = ~n9994 ;
  assign y1380 = n10004 ;
  assign y1381 = n10018 ;
  assign y1382 = n10026 ;
  assign y1383 = n10032 ;
  assign y1384 = n10040 ;
  assign y1385 = n10048 ;
  assign y1386 = ~n10052 ;
  assign y1387 = ~1'b0 ;
  assign y1388 = n10053 ;
  assign y1389 = n10055 ;
  assign y1390 = ~n10057 ;
  assign y1391 = ~n10061 ;
  assign y1392 = ~n10068 ;
  assign y1393 = ~n10069 ;
  assign y1394 = n10074 ;
  assign y1395 = ~n10084 ;
  assign y1396 = n10086 ;
  assign y1397 = ~n10100 ;
  assign y1398 = n10117 ;
  assign y1399 = n10122 ;
  assign y1400 = n10141 ;
  assign y1401 = ~1'b0 ;
  assign y1402 = n10151 ;
  assign y1403 = n10153 ;
  assign y1404 = n10180 ;
  assign y1405 = ~1'b0 ;
  assign y1406 = ~n10196 ;
  assign y1407 = ~n10201 ;
  assign y1408 = ~n10206 ;
  assign y1409 = n10213 ;
  assign y1410 = ~n10232 ;
  assign y1411 = n10234 ;
  assign y1412 = n10238 ;
  assign y1413 = ~n10245 ;
  assign y1414 = n10259 ;
  assign y1415 = n10261 ;
  assign y1416 = ~n10279 ;
  assign y1417 = n10284 ;
  assign y1418 = ~n10288 ;
  assign y1419 = ~n10297 ;
  assign y1420 = ~n10299 ;
  assign y1421 = n10303 ;
  assign y1422 = n10321 ;
  assign y1423 = ~n10324 ;
  assign y1424 = ~n10332 ;
  assign y1425 = ~1'b0 ;
  assign y1426 = n10333 ;
  assign y1427 = ~n10340 ;
  assign y1428 = ~n10342 ;
  assign y1429 = ~n10353 ;
  assign y1430 = ~n10359 ;
  assign y1431 = ~n10369 ;
  assign y1432 = ~n10373 ;
  assign y1433 = n10376 ;
  assign y1434 = ~n10383 ;
  assign y1435 = ~n10385 ;
  assign y1436 = n10387 ;
  assign y1437 = ~n10393 ;
  assign y1438 = ~n10398 ;
  assign y1439 = ~n10406 ;
  assign y1440 = ~n10409 ;
  assign y1441 = n10413 ;
  assign y1442 = n10423 ;
  assign y1443 = n10425 ;
  assign y1444 = ~n10433 ;
  assign y1445 = n10434 ;
  assign y1446 = n10435 ;
  assign y1447 = ~n10456 ;
  assign y1448 = ~n10460 ;
  assign y1449 = n10471 ;
  assign y1450 = ~n10472 ;
  assign y1451 = ~n10486 ;
  assign y1452 = ~n10490 ;
  assign y1453 = ~1'b0 ;
  assign y1454 = ~n10500 ;
  assign y1455 = n10507 ;
  assign y1456 = n10514 ;
  assign y1457 = n10517 ;
  assign y1458 = n10526 ;
  assign y1459 = ~1'b0 ;
  assign y1460 = ~n10530 ;
  assign y1461 = n10543 ;
  assign y1462 = ~n10552 ;
  assign y1463 = n10553 ;
  assign y1464 = ~n10556 ;
  assign y1465 = n10561 ;
  assign y1466 = n10563 ;
  assign y1467 = ~n10569 ;
  assign y1468 = ~n10572 ;
  assign y1469 = n10576 ;
  assign y1470 = n10577 ;
  assign y1471 = n10588 ;
  assign y1472 = n10591 ;
  assign y1473 = n10608 ;
  assign y1474 = ~1'b0 ;
  assign y1475 = n10610 ;
  assign y1476 = n10616 ;
  assign y1477 = ~n10619 ;
  assign y1478 = ~n10622 ;
  assign y1479 = ~n10623 ;
  assign y1480 = ~n10638 ;
  assign y1481 = ~n10649 ;
  assign y1482 = ~n10655 ;
  assign y1483 = n10661 ;
  assign y1484 = ~n10670 ;
  assign y1485 = ~n10673 ;
  assign y1486 = ~n10685 ;
  assign y1487 = ~n10692 ;
  assign y1488 = ~n10693 ;
  assign y1489 = n10698 ;
  assign y1490 = ~n10715 ;
  assign y1491 = ~1'b0 ;
  assign y1492 = n10723 ;
  assign y1493 = n10733 ;
  assign y1494 = ~n10748 ;
  assign y1495 = ~n10749 ;
  assign y1496 = ~n10750 ;
  assign y1497 = ~n10754 ;
  assign y1498 = n10761 ;
  assign y1499 = n10768 ;
  assign y1500 = ~n10780 ;
  assign y1501 = ~n10789 ;
  assign y1502 = n10793 ;
  assign y1503 = n10796 ;
  assign y1504 = ~n10798 ;
  assign y1505 = n10802 ;
  assign y1506 = n10812 ;
  assign y1507 = ~n10813 ;
  assign y1508 = n10823 ;
  assign y1509 = n10830 ;
  assign y1510 = ~n10834 ;
  assign y1511 = n10847 ;
  assign y1512 = n10852 ;
  assign y1513 = ~n10854 ;
  assign y1514 = ~n10855 ;
  assign y1515 = ~n10858 ;
  assign y1516 = n10860 ;
  assign y1517 = ~n10868 ;
  assign y1518 = n10873 ;
  assign y1519 = ~n10876 ;
  assign y1520 = n10886 ;
  assign y1521 = ~n10887 ;
  assign y1522 = ~n10894 ;
  assign y1523 = n10911 ;
  assign y1524 = ~n10920 ;
  assign y1525 = ~n10929 ;
  assign y1526 = ~n10931 ;
  assign y1527 = n10933 ;
  assign y1528 = ~1'b0 ;
  assign y1529 = n10936 ;
  assign y1530 = ~n10944 ;
  assign y1531 = n10947 ;
  assign y1532 = ~n10954 ;
  assign y1533 = ~n10961 ;
  assign y1534 = n10966 ;
  assign y1535 = ~n10968 ;
  assign y1536 = ~n10970 ;
  assign y1537 = ~n10971 ;
  assign y1538 = ~n10982 ;
  assign y1539 = ~n10987 ;
  assign y1540 = n10992 ;
  assign y1541 = n10996 ;
  assign y1542 = ~n11004 ;
  assign y1543 = ~n11010 ;
  assign y1544 = n11011 ;
  assign y1545 = ~n11025 ;
  assign y1546 = ~1'b0 ;
  assign y1547 = ~n11033 ;
  assign y1548 = n11038 ;
  assign y1549 = n11042 ;
  assign y1550 = n11062 ;
  assign y1551 = ~n11072 ;
  assign y1552 = n11082 ;
  assign y1553 = n11086 ;
  assign y1554 = ~n11093 ;
  assign y1555 = ~n11096 ;
  assign y1556 = ~n11105 ;
  assign y1557 = ~n11107 ;
  assign y1558 = ~n11123 ;
  assign y1559 = n11132 ;
  assign y1560 = ~n11143 ;
  assign y1561 = n11146 ;
  assign y1562 = ~n11151 ;
  assign y1563 = ~n11166 ;
  assign y1564 = n11187 ;
  assign y1565 = ~n11192 ;
  assign y1566 = n11203 ;
  assign y1567 = ~n11218 ;
  assign y1568 = n11229 ;
  assign y1569 = n11236 ;
  assign y1570 = ~n11240 ;
  assign y1571 = ~n11259 ;
  assign y1572 = n11260 ;
  assign y1573 = n11271 ;
  assign y1574 = ~n11285 ;
  assign y1575 = n11290 ;
  assign y1576 = n11295 ;
  assign y1577 = ~n11302 ;
  assign y1578 = n11309 ;
  assign y1579 = n11320 ;
  assign y1580 = ~n11330 ;
  assign y1581 = n11331 ;
  assign y1582 = ~n11333 ;
  assign y1583 = n11355 ;
  assign y1584 = n11368 ;
  assign y1585 = n11372 ;
  assign y1586 = n11386 ;
  assign y1587 = ~n11399 ;
  assign y1588 = n11409 ;
  assign y1589 = ~n11412 ;
  assign y1590 = n11417 ;
  assign y1591 = n11421 ;
  assign y1592 = ~n11440 ;
  assign y1593 = n11445 ;
  assign y1594 = n11449 ;
  assign y1595 = n11456 ;
  assign y1596 = ~n11458 ;
  assign y1597 = n11461 ;
  assign y1598 = ~n11463 ;
  assign y1599 = ~1'b0 ;
  assign y1600 = ~n11466 ;
  assign y1601 = n11472 ;
  assign y1602 = ~n11496 ;
  assign y1603 = n11504 ;
  assign y1604 = n11512 ;
  assign y1605 = ~n11518 ;
  assign y1606 = ~n11519 ;
  assign y1607 = ~n11533 ;
  assign y1608 = ~n11536 ;
  assign y1609 = n11537 ;
  assign y1610 = n11540 ;
  assign y1611 = n11544 ;
  assign y1612 = n11547 ;
  assign y1613 = n11548 ;
  assign y1614 = ~1'b0 ;
  assign y1615 = n11560 ;
  assign y1616 = n11561 ;
  assign y1617 = ~n11565 ;
  assign y1618 = ~n11570 ;
  assign y1619 = n11572 ;
  assign y1620 = ~n11581 ;
  assign y1621 = ~n11584 ;
  assign y1622 = ~n11594 ;
  assign y1623 = ~n11598 ;
  assign y1624 = ~n11609 ;
  assign y1625 = ~n11616 ;
  assign y1626 = n11623 ;
  assign y1627 = ~n11626 ;
  assign y1628 = ~n11631 ;
  assign y1629 = n11638 ;
  assign y1630 = n11644 ;
  assign y1631 = ~n11651 ;
  assign y1632 = n11656 ;
  assign y1633 = n11670 ;
  assign y1634 = ~n11679 ;
  assign y1635 = ~n11684 ;
  assign y1636 = n11697 ;
  assign y1637 = ~n11702 ;
  assign y1638 = n11707 ;
  assign y1639 = ~n11708 ;
  assign y1640 = n11729 ;
  assign y1641 = ~n11730 ;
  assign y1642 = ~n11734 ;
  assign y1643 = n11738 ;
  assign y1644 = n11743 ;
  assign y1645 = ~n11747 ;
  assign y1646 = ~n11762 ;
  assign y1647 = ~n11768 ;
  assign y1648 = ~n11774 ;
  assign y1649 = ~n11778 ;
  assign y1650 = ~n11780 ;
  assign y1651 = ~n11788 ;
  assign y1652 = ~1'b0 ;
  assign y1653 = ~1'b0 ;
  assign y1654 = ~n11789 ;
  assign y1655 = ~n11790 ;
  assign y1656 = n11797 ;
  assign y1657 = ~n11799 ;
  assign y1658 = ~n11801 ;
  assign y1659 = n11809 ;
  assign y1660 = ~n11823 ;
  assign y1661 = ~n11834 ;
  assign y1662 = n11837 ;
  assign y1663 = ~n11838 ;
  assign y1664 = ~n11842 ;
  assign y1665 = n11852 ;
  assign y1666 = ~n11860 ;
  assign y1667 = n11861 ;
  assign y1668 = ~n11868 ;
  assign y1669 = n11879 ;
  assign y1670 = n11888 ;
  assign y1671 = ~n11890 ;
  assign y1672 = n11894 ;
  assign y1673 = n11903 ;
  assign y1674 = ~n11909 ;
  assign y1675 = ~n11920 ;
  assign y1676 = ~1'b0 ;
  assign y1677 = n11921 ;
  assign y1678 = n11931 ;
  assign y1679 = n11950 ;
  assign y1680 = ~n11952 ;
  assign y1681 = n11956 ;
  assign y1682 = n11960 ;
  assign y1683 = n11971 ;
  assign y1684 = ~n11977 ;
  assign y1685 = ~n11983 ;
  assign y1686 = ~n12001 ;
  assign y1687 = ~n12010 ;
  assign y1688 = n12018 ;
  assign y1689 = n12023 ;
  assign y1690 = ~n12025 ;
  assign y1691 = ~n12032 ;
  assign y1692 = n12043 ;
  assign y1693 = n12046 ;
  assign y1694 = ~n12051 ;
  assign y1695 = n12054 ;
  assign y1696 = n12055 ;
  assign y1697 = n12059 ;
  assign y1698 = ~n12063 ;
  assign y1699 = ~n12069 ;
  assign y1700 = ~n12071 ;
  assign y1701 = ~n12073 ;
  assign y1702 = ~n12075 ;
  assign y1703 = ~n12081 ;
  assign y1704 = n12093 ;
  assign y1705 = ~n12100 ;
  assign y1706 = ~n12105 ;
  assign y1707 = ~n12106 ;
  assign y1708 = ~n12107 ;
  assign y1709 = ~n12118 ;
  assign y1710 = n12134 ;
  assign y1711 = ~n12136 ;
  assign y1712 = n12137 ;
  assign y1713 = n12145 ;
  assign y1714 = ~n12148 ;
  assign y1715 = n12167 ;
  assign y1716 = ~n12173 ;
  assign y1717 = n12174 ;
  assign y1718 = ~n12175 ;
  assign y1719 = ~n12180 ;
  assign y1720 = n12196 ;
  assign y1721 = ~n12206 ;
  assign y1722 = n12208 ;
  assign y1723 = ~n12213 ;
  assign y1724 = n12217 ;
  assign y1725 = n12225 ;
  assign y1726 = n12229 ;
  assign y1727 = ~n12233 ;
  assign y1728 = ~n12253 ;
  assign y1729 = n12271 ;
  assign y1730 = n12276 ;
  assign y1731 = ~n12281 ;
  assign y1732 = ~n12291 ;
  assign y1733 = n12294 ;
  assign y1734 = ~n12307 ;
  assign y1735 = n12318 ;
  assign y1736 = n12334 ;
  assign y1737 = n12345 ;
  assign y1738 = n12351 ;
  assign y1739 = ~n12353 ;
  assign y1740 = n12354 ;
  assign y1741 = ~n12365 ;
  assign y1742 = ~n12368 ;
  assign y1743 = n12377 ;
  assign y1744 = n12382 ;
  assign y1745 = n12394 ;
  assign y1746 = ~n12402 ;
  assign y1747 = n12406 ;
  assign y1748 = n12412 ;
  assign y1749 = n12416 ;
  assign y1750 = n12419 ;
  assign y1751 = ~n12423 ;
  assign y1752 = n12430 ;
  assign y1753 = ~n12431 ;
  assign y1754 = n12450 ;
  assign y1755 = n12452 ;
  assign y1756 = ~n12469 ;
  assign y1757 = n12475 ;
  assign y1758 = ~n12480 ;
  assign y1759 = ~n12488 ;
  assign y1760 = n12499 ;
  assign y1761 = n12500 ;
  assign y1762 = ~n12501 ;
  assign y1763 = ~n12503 ;
  assign y1764 = n12511 ;
  assign y1765 = ~n12515 ;
  assign y1766 = ~n12518 ;
  assign y1767 = n12530 ;
  assign y1768 = n12534 ;
  assign y1769 = n12549 ;
  assign y1770 = ~n12554 ;
  assign y1771 = n12557 ;
  assign y1772 = n12562 ;
  assign y1773 = ~1'b0 ;
  assign y1774 = ~n12563 ;
  assign y1775 = ~n12568 ;
  assign y1776 = n12573 ;
  assign y1777 = n12574 ;
  assign y1778 = ~n12576 ;
  assign y1779 = ~n12581 ;
  assign y1780 = ~n12586 ;
  assign y1781 = n12592 ;
  assign y1782 = ~n12596 ;
  assign y1783 = n12599 ;
  assign y1784 = n12600 ;
  assign y1785 = n12604 ;
  assign y1786 = ~n12616 ;
  assign y1787 = ~n12617 ;
  assign y1788 = n12619 ;
  assign y1789 = ~n12620 ;
  assign y1790 = n12624 ;
  assign y1791 = n12629 ;
  assign y1792 = n12630 ;
  assign y1793 = ~1'b0 ;
  assign y1794 = ~n12631 ;
  assign y1795 = n12636 ;
  assign y1796 = n12637 ;
  assign y1797 = n12646 ;
  assign y1798 = n12650 ;
  assign y1799 = n12656 ;
  assign y1800 = n12661 ;
  assign y1801 = n12666 ;
  assign y1802 = ~n12669 ;
  assign y1803 = n12670 ;
  assign y1804 = ~n12678 ;
  assign y1805 = ~n12686 ;
  assign y1806 = ~n12690 ;
  assign y1807 = n12692 ;
  assign y1808 = ~n12696 ;
  assign y1809 = ~n12703 ;
  assign y1810 = n12709 ;
  assign y1811 = ~n12715 ;
  assign y1812 = ~n12722 ;
  assign y1813 = ~n12728 ;
  assign y1814 = n12730 ;
  assign y1815 = n12737 ;
  assign y1816 = n12741 ;
  assign y1817 = n12742 ;
  assign y1818 = ~n12746 ;
  assign y1819 = ~n12764 ;
  assign y1820 = n12774 ;
  assign y1821 = ~n12776 ;
  assign y1822 = n12778 ;
  assign y1823 = n12786 ;
  assign y1824 = n12790 ;
  assign y1825 = n12794 ;
  assign y1826 = ~n12800 ;
  assign y1827 = ~n12804 ;
  assign y1828 = ~n12805 ;
  assign y1829 = n12809 ;
  assign y1830 = n12826 ;
  assign y1831 = ~n12838 ;
  assign y1832 = ~n12845 ;
  assign y1833 = ~n12846 ;
  assign y1834 = n12853 ;
  assign y1835 = ~n12865 ;
  assign y1836 = ~1'b0 ;
  assign y1837 = ~n12870 ;
  assign y1838 = ~n12885 ;
  assign y1839 = n12886 ;
  assign y1840 = n12898 ;
  assign y1841 = ~n12910 ;
  assign y1842 = n12917 ;
  assign y1843 = n12920 ;
  assign y1844 = ~n12924 ;
  assign y1845 = ~n12939 ;
  assign y1846 = n12945 ;
  assign y1847 = ~n12959 ;
  assign y1848 = ~n12968 ;
  assign y1849 = n12970 ;
  assign y1850 = ~1'b0 ;
  assign y1851 = n12976 ;
  assign y1852 = n12981 ;
  assign y1853 = ~n12997 ;
  assign y1854 = ~n13000 ;
  assign y1855 = n13001 ;
  assign y1856 = ~n13008 ;
  assign y1857 = ~n13009 ;
  assign y1858 = n13011 ;
  assign y1859 = ~n13021 ;
  assign y1860 = ~n13028 ;
  assign y1861 = ~1'b0 ;
  assign y1862 = n13029 ;
  assign y1863 = n13032 ;
  assign y1864 = ~n13033 ;
  assign y1865 = ~n13041 ;
  assign y1866 = n13050 ;
  assign y1867 = n13055 ;
  assign y1868 = n13061 ;
  assign y1869 = ~n13062 ;
  assign y1870 = ~n13070 ;
  assign y1871 = n13080 ;
  assign y1872 = n13083 ;
  assign y1873 = ~n13091 ;
  assign y1874 = ~n13094 ;
  assign y1875 = n13102 ;
  assign y1876 = ~n13109 ;
  assign y1877 = ~n13125 ;
  assign y1878 = n13126 ;
  assign y1879 = ~1'b0 ;
  assign y1880 = ~n13131 ;
  assign y1881 = ~n13148 ;
  assign y1882 = ~n13150 ;
  assign y1883 = n13156 ;
  assign y1884 = n13161 ;
  assign y1885 = n13168 ;
  assign y1886 = ~n13172 ;
  assign y1887 = n13174 ;
  assign y1888 = n13183 ;
  assign y1889 = ~n13193 ;
  assign y1890 = n13197 ;
  assign y1891 = n13200 ;
  assign y1892 = n13205 ;
  assign y1893 = ~n13211 ;
  assign y1894 = ~n13221 ;
  assign y1895 = ~1'b0 ;
  assign y1896 = ~n13228 ;
  assign y1897 = n13237 ;
  assign y1898 = ~n13241 ;
  assign y1899 = n13250 ;
  assign y1900 = n13254 ;
  assign y1901 = n13263 ;
  assign y1902 = ~n13265 ;
  assign y1903 = n13267 ;
  assign y1904 = n13268 ;
  assign y1905 = n13270 ;
  assign y1906 = ~n13277 ;
  assign y1907 = ~n13278 ;
  assign y1908 = ~n13279 ;
  assign y1909 = ~1'b0 ;
  assign y1910 = ~n13280 ;
  assign y1911 = ~n13286 ;
  assign y1912 = ~n13289 ;
  assign y1913 = ~n13290 ;
  assign y1914 = n13295 ;
  assign y1915 = n13303 ;
  assign y1916 = n13305 ;
  assign y1917 = ~1'b0 ;
  assign y1918 = n13306 ;
  assign y1919 = ~n13326 ;
  assign y1920 = ~n13327 ;
  assign y1921 = ~n13332 ;
  assign y1922 = n13336 ;
  assign y1923 = ~n13339 ;
  assign y1924 = n13350 ;
  assign y1925 = n13362 ;
  assign y1926 = n13375 ;
  assign y1927 = n13380 ;
  assign y1928 = n13382 ;
  assign y1929 = ~n13404 ;
  assign y1930 = ~n13406 ;
  assign y1931 = n13414 ;
  assign y1932 = n13421 ;
  assign y1933 = ~n13426 ;
  assign y1934 = ~n13428 ;
  assign y1935 = n13433 ;
  assign y1936 = n13451 ;
  assign y1937 = n13452 ;
  assign y1938 = n13453 ;
  assign y1939 = ~n13456 ;
  assign y1940 = ~n13457 ;
  assign y1941 = n13461 ;
  assign y1942 = n13466 ;
  assign y1943 = ~n13471 ;
  assign y1944 = n13475 ;
  assign y1945 = n13480 ;
  assign y1946 = ~n13497 ;
  assign y1947 = ~n13514 ;
  assign y1948 = n13518 ;
  assign y1949 = n13524 ;
  assign y1950 = ~n13540 ;
  assign y1951 = ~n13543 ;
  assign y1952 = ~n13548 ;
  assign y1953 = n13552 ;
  assign y1954 = ~n13555 ;
  assign y1955 = ~n13556 ;
  assign y1956 = n13561 ;
  assign y1957 = ~n13571 ;
  assign y1958 = n13591 ;
  assign y1959 = ~n13594 ;
  assign y1960 = n13598 ;
  assign y1961 = ~n13604 ;
  assign y1962 = ~n13611 ;
  assign y1963 = ~n13613 ;
  assign y1964 = n13621 ;
  assign y1965 = ~n13624 ;
  assign y1966 = ~n13629 ;
  assign y1967 = ~n13642 ;
  assign y1968 = ~n13650 ;
  assign y1969 = n13652 ;
  assign y1970 = n13653 ;
  assign y1971 = n13656 ;
  assign y1972 = n13667 ;
  assign y1973 = n13674 ;
  assign y1974 = n13676 ;
  assign y1975 = ~n13688 ;
  assign y1976 = ~n13690 ;
  assign y1977 = n13699 ;
  assign y1978 = ~n13701 ;
  assign y1979 = ~1'b0 ;
  assign y1980 = n13702 ;
  assign y1981 = n13712 ;
  assign y1982 = ~n13721 ;
  assign y1983 = ~n13723 ;
  assign y1984 = n13732 ;
  assign y1985 = ~n13734 ;
  assign y1986 = ~n13739 ;
  assign y1987 = ~n13752 ;
  assign y1988 = n13756 ;
  assign y1989 = n13758 ;
  assign y1990 = ~n13759 ;
  assign y1991 = ~n13767 ;
  assign y1992 = ~n13774 ;
  assign y1993 = n13781 ;
  assign y1994 = n13786 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = n13787 ;
  assign y1997 = ~n13801 ;
  assign y1998 = n13828 ;
  assign y1999 = ~n13836 ;
  assign y2000 = n13858 ;
  assign y2001 = ~n13873 ;
  assign y2002 = ~n13879 ;
  assign y2003 = n13891 ;
  assign y2004 = ~n13910 ;
  assign y2005 = n13911 ;
  assign y2006 = ~n13915 ;
  assign y2007 = n13917 ;
  assign y2008 = n13922 ;
  assign y2009 = ~n13924 ;
  assign y2010 = n13928 ;
  assign y2011 = ~n13929 ;
  assign y2012 = ~n13931 ;
  assign y2013 = ~n13938 ;
  assign y2014 = n13945 ;
  assign y2015 = n13949 ;
  assign y2016 = n13963 ;
  assign y2017 = ~1'b0 ;
  assign y2018 = ~n13964 ;
  assign y2019 = ~n13968 ;
  assign y2020 = n13979 ;
  assign y2021 = ~n13989 ;
  assign y2022 = ~n13991 ;
  assign y2023 = n13993 ;
  assign y2024 = ~n13997 ;
  assign y2025 = n14005 ;
  assign y2026 = ~n14007 ;
  assign y2027 = ~n14023 ;
  assign y2028 = ~n14028 ;
  assign y2029 = n14035 ;
  assign y2030 = n14038 ;
  assign y2031 = n14045 ;
  assign y2032 = ~n14054 ;
  assign y2033 = ~n14056 ;
  assign y2034 = ~n14057 ;
  assign y2035 = ~n14070 ;
  assign y2036 = ~n14076 ;
  assign y2037 = ~1'b0 ;
  assign y2038 = ~n14078 ;
  assign y2039 = ~1'b0 ;
  assign y2040 = n14081 ;
  assign y2041 = n14082 ;
  assign y2042 = ~n14083 ;
  assign y2043 = n14093 ;
  assign y2044 = ~n14095 ;
  assign y2045 = n14111 ;
  assign y2046 = ~1'b0 ;
  assign y2047 = n14120 ;
  assign y2048 = ~n14121 ;
  assign y2049 = ~n14128 ;
  assign y2050 = ~n14133 ;
  assign y2051 = n14138 ;
  assign y2052 = n14146 ;
  assign y2053 = n14148 ;
  assign y2054 = n14151 ;
  assign y2055 = n14154 ;
  assign y2056 = ~n14157 ;
  assign y2057 = n14164 ;
  assign y2058 = ~n14176 ;
  assign y2059 = ~1'b0 ;
  assign y2060 = ~n14179 ;
  assign y2061 = ~n14188 ;
  assign y2062 = ~n14206 ;
  assign y2063 = ~n14208 ;
  assign y2064 = n14210 ;
  assign y2065 = ~n14217 ;
  assign y2066 = n14232 ;
  assign y2067 = n14236 ;
  assign y2068 = ~n14247 ;
  assign y2069 = n14260 ;
  assign y2070 = n14266 ;
  assign y2071 = ~n14272 ;
  assign y2072 = ~n14277 ;
  assign y2073 = n14282 ;
  assign y2074 = n14284 ;
  assign y2075 = ~n14290 ;
  assign y2076 = ~n14295 ;
  assign y2077 = ~n14300 ;
  assign y2078 = n14301 ;
  assign y2079 = n14308 ;
  assign y2080 = n14311 ;
  assign y2081 = ~n14314 ;
  assign y2082 = n14315 ;
  assign y2083 = n14318 ;
  assign y2084 = ~n14326 ;
  assign y2085 = n14329 ;
  assign y2086 = n14340 ;
  assign y2087 = ~n14342 ;
  assign y2088 = n14348 ;
  assign y2089 = n14351 ;
  assign y2090 = ~n14370 ;
  assign y2091 = ~n14373 ;
  assign y2092 = ~n14375 ;
  assign y2093 = n14389 ;
  assign y2094 = n14390 ;
  assign y2095 = n14393 ;
  assign y2096 = ~1'b0 ;
  assign y2097 = n14399 ;
  assign y2098 = ~n14404 ;
  assign y2099 = ~n14408 ;
  assign y2100 = ~n14415 ;
  assign y2101 = ~1'b0 ;
  assign y2102 = n14419 ;
  assign y2103 = ~1'b0 ;
  assign y2104 = ~n14425 ;
  assign y2105 = ~n14432 ;
  assign y2106 = n14434 ;
  assign y2107 = n14448 ;
  assign y2108 = ~n14453 ;
  assign y2109 = n14461 ;
  assign y2110 = n14465 ;
  assign y2111 = ~n14469 ;
  assign y2112 = n14472 ;
  assign y2113 = ~n14475 ;
  assign y2114 = n14481 ;
  assign y2115 = n14482 ;
  assign y2116 = n14493 ;
  assign y2117 = ~n14494 ;
  assign y2118 = ~n14496 ;
  assign y2119 = ~n14498 ;
  assign y2120 = ~n14500 ;
  assign y2121 = n14514 ;
  assign y2122 = n14515 ;
  assign y2123 = n14522 ;
  assign y2124 = ~n14529 ;
  assign y2125 = ~n14535 ;
  assign y2126 = ~n14546 ;
  assign y2127 = n14548 ;
  assign y2128 = ~n14552 ;
  assign y2129 = n14557 ;
  assign y2130 = n14562 ;
  assign y2131 = n14573 ;
  assign y2132 = n14574 ;
  assign y2133 = ~1'b0 ;
  assign y2134 = ~n14577 ;
  assign y2135 = ~n14580 ;
  assign y2136 = n14582 ;
  assign y2137 = ~n14583 ;
  assign y2138 = n14594 ;
  assign y2139 = n14597 ;
  assign y2140 = ~n14601 ;
  assign y2141 = ~n14605 ;
  assign y2142 = n14606 ;
  assign y2143 = ~1'b0 ;
  assign y2144 = ~n14607 ;
  assign y2145 = n14608 ;
  assign y2146 = ~n14610 ;
  assign y2147 = ~n14624 ;
  assign y2148 = ~n14626 ;
  assign y2149 = n14631 ;
  assign y2150 = ~n14634 ;
  assign y2151 = ~n14636 ;
  assign y2152 = n14637 ;
  assign y2153 = n14639 ;
  assign y2154 = ~n14641 ;
  assign y2155 = n14642 ;
  assign y2156 = n14644 ;
  assign y2157 = ~n14645 ;
  assign y2158 = n14648 ;
  assign y2159 = ~n14661 ;
  assign y2160 = ~n14678 ;
  assign y2161 = ~1'b0 ;
  assign y2162 = ~n14686 ;
  assign y2163 = ~n14693 ;
  assign y2164 = ~n14694 ;
  assign y2165 = n14696 ;
  assign y2166 = ~1'b0 ;
  assign y2167 = ~n14702 ;
  assign y2168 = n14703 ;
  assign y2169 = n14710 ;
  assign y2170 = n14713 ;
  assign y2171 = ~n14714 ;
  assign y2172 = ~n14718 ;
  assign y2173 = n14721 ;
  assign y2174 = ~n14737 ;
  assign y2175 = ~n14747 ;
  assign y2176 = n14750 ;
  assign y2177 = ~n14754 ;
  assign y2178 = ~n14755 ;
  assign y2179 = ~n14759 ;
  assign y2180 = n14760 ;
  assign y2181 = ~n14762 ;
  assign y2182 = ~n14772 ;
  assign y2183 = ~n14775 ;
  assign y2184 = n14781 ;
  assign y2185 = ~n14786 ;
  assign y2186 = ~n14792 ;
  assign y2187 = n14798 ;
  assign y2188 = n14801 ;
  assign y2189 = n14809 ;
  assign y2190 = ~n14810 ;
  assign y2191 = n14823 ;
  assign y2192 = ~n14828 ;
  assign y2193 = ~n14830 ;
  assign y2194 = ~n14831 ;
  assign y2195 = ~n14838 ;
  assign y2196 = n14841 ;
  assign y2197 = n14845 ;
  assign y2198 = n14855 ;
  assign y2199 = n14860 ;
  assign y2200 = ~1'b0 ;
  assign y2201 = n14863 ;
  assign y2202 = ~n14865 ;
  assign y2203 = n14872 ;
  assign y2204 = ~n14877 ;
  assign y2205 = n14880 ;
  assign y2206 = ~n14888 ;
  assign y2207 = ~n14893 ;
  assign y2208 = ~n14898 ;
  assign y2209 = ~1'b0 ;
  assign y2210 = n14910 ;
  assign y2211 = ~n14915 ;
  assign y2212 = ~n14918 ;
  assign y2213 = n14928 ;
  assign y2214 = n14931 ;
  assign y2215 = n14932 ;
  assign y2216 = ~n14934 ;
  assign y2217 = n14938 ;
  assign y2218 = n14956 ;
  assign y2219 = n14958 ;
  assign y2220 = ~n14962 ;
  assign y2221 = ~n14986 ;
  assign y2222 = n14988 ;
  assign y2223 = n14992 ;
  assign y2224 = n14996 ;
  assign y2225 = n14999 ;
  assign y2226 = ~n15005 ;
  assign y2227 = n15008 ;
  assign y2228 = n15009 ;
  assign y2229 = n15012 ;
  assign y2230 = ~n15019 ;
  assign y2231 = ~n15021 ;
  assign y2232 = ~n15023 ;
  assign y2233 = n15027 ;
  assign y2234 = ~n15043 ;
  assign y2235 = ~n15045 ;
  assign y2236 = n15052 ;
  assign y2237 = n15061 ;
  assign y2238 = ~n15071 ;
  assign y2239 = ~n15074 ;
  assign y2240 = ~n15077 ;
  assign y2241 = ~1'b0 ;
  assign y2242 = ~n15081 ;
  assign y2243 = ~n15086 ;
  assign y2244 = n15090 ;
  assign y2245 = n15094 ;
  assign y2246 = ~n15098 ;
  assign y2247 = ~n15099 ;
  assign y2248 = n15105 ;
  assign y2249 = n15107 ;
  assign y2250 = n15110 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = n15112 ;
  assign y2253 = n15123 ;
  assign y2254 = n15130 ;
  assign y2255 = ~n15131 ;
  assign y2256 = ~n15139 ;
  assign y2257 = ~n15143 ;
  assign y2258 = n15164 ;
  assign y2259 = ~n15166 ;
  assign y2260 = n15167 ;
  assign y2261 = n15168 ;
  assign y2262 = n15175 ;
  assign y2263 = n15185 ;
  assign y2264 = n15186 ;
  assign y2265 = n15198 ;
  assign y2266 = ~1'b0 ;
  assign y2267 = n15202 ;
  assign y2268 = ~n15209 ;
  assign y2269 = ~n15221 ;
  assign y2270 = ~n15227 ;
  assign y2271 = n15249 ;
  assign y2272 = ~n15253 ;
  assign y2273 = ~n15254 ;
  assign y2274 = ~n15261 ;
  assign y2275 = ~n15263 ;
  assign y2276 = n15277 ;
  assign y2277 = ~n15279 ;
  assign y2278 = ~n15283 ;
  assign y2279 = n15284 ;
  assign y2280 = ~n15291 ;
  assign y2281 = ~n15298 ;
  assign y2282 = n15300 ;
  assign y2283 = n15309 ;
  assign y2284 = n15311 ;
  assign y2285 = n15318 ;
  assign y2286 = n15320 ;
  assign y2287 = n15322 ;
  assign y2288 = ~n15331 ;
  assign y2289 = ~n15335 ;
  assign y2290 = ~n15338 ;
  assign y2291 = ~n15348 ;
  assign y2292 = n15352 ;
  assign y2293 = n15354 ;
  assign y2294 = n15358 ;
  assign y2295 = ~n15361 ;
  assign y2296 = n15362 ;
  assign y2297 = ~n15364 ;
  assign y2298 = ~n15372 ;
  assign y2299 = ~n15374 ;
  assign y2300 = ~n15375 ;
  assign y2301 = ~n15379 ;
  assign y2302 = ~n15382 ;
  assign y2303 = n15383 ;
  assign y2304 = n15384 ;
  assign y2305 = ~n15392 ;
  assign y2306 = ~n15396 ;
  assign y2307 = ~n15405 ;
  assign y2308 = n15409 ;
  assign y2309 = n15419 ;
  assign y2310 = n15424 ;
  assign y2311 = n15432 ;
  assign y2312 = n15434 ;
  assign y2313 = n15442 ;
  assign y2314 = ~n15445 ;
  assign y2315 = ~n15446 ;
  assign y2316 = ~n15448 ;
  assign y2317 = n15455 ;
  assign y2318 = n15458 ;
  assign y2319 = n15459 ;
  assign y2320 = ~n15461 ;
  assign y2321 = n15466 ;
  assign y2322 = ~n15473 ;
  assign y2323 = ~n15476 ;
  assign y2324 = ~n15480 ;
  assign y2325 = n15481 ;
  assign y2326 = n15491 ;
  assign y2327 = ~n15494 ;
  assign y2328 = ~1'b0 ;
  assign y2329 = ~n15495 ;
  assign y2330 = n15498 ;
  assign y2331 = ~n15503 ;
  assign y2332 = n15512 ;
  assign y2333 = ~1'b0 ;
  assign y2334 = ~n15514 ;
  assign y2335 = n15528 ;
  assign y2336 = ~n15531 ;
  assign y2337 = n15536 ;
  assign y2338 = ~n15538 ;
  assign y2339 = ~n15542 ;
  assign y2340 = ~n15545 ;
  assign y2341 = ~n15547 ;
  assign y2342 = ~n15551 ;
  assign y2343 = ~n15556 ;
  assign y2344 = n15571 ;
  assign y2345 = ~n15583 ;
  assign y2346 = n15588 ;
  assign y2347 = ~n15595 ;
  assign y2348 = ~1'b0 ;
  assign y2349 = ~n15604 ;
  assign y2350 = n15606 ;
  assign y2351 = ~1'b0 ;
  assign y2352 = n15607 ;
  assign y2353 = ~1'b0 ;
  assign y2354 = ~n15611 ;
  assign y2355 = ~n15616 ;
  assign y2356 = ~n15622 ;
  assign y2357 = n15627 ;
  assign y2358 = ~n15629 ;
  assign y2359 = ~n15636 ;
  assign y2360 = n15644 ;
  assign y2361 = ~n15645 ;
  assign y2362 = ~n15646 ;
  assign y2363 = ~n15650 ;
  assign y2364 = ~n15657 ;
  assign y2365 = ~n15662 ;
  assign y2366 = ~n15667 ;
  assign y2367 = ~n15680 ;
  assign y2368 = n15681 ;
  assign y2369 = n15688 ;
  assign y2370 = n15695 ;
  assign y2371 = ~n15701 ;
  assign y2372 = ~n15703 ;
  assign y2373 = ~n15716 ;
  assign y2374 = ~1'b0 ;
  assign y2375 = ~n15718 ;
  assign y2376 = ~n15721 ;
  assign y2377 = n15722 ;
  assign y2378 = ~n15726 ;
  assign y2379 = n15731 ;
  assign y2380 = ~n15733 ;
  assign y2381 = n15739 ;
  assign y2382 = ~n15742 ;
  assign y2383 = ~n15750 ;
  assign y2384 = n15754 ;
  assign y2385 = n15755 ;
  assign y2386 = ~n15756 ;
  assign y2387 = n15757 ;
  assign y2388 = ~n15759 ;
  assign y2389 = ~n15763 ;
  assign y2390 = ~n15766 ;
  assign y2391 = ~n15768 ;
  assign y2392 = ~n15771 ;
  assign y2393 = n15783 ;
  assign y2394 = ~n15785 ;
  assign y2395 = ~n15786 ;
  assign y2396 = n15795 ;
  assign y2397 = ~n15796 ;
  assign y2398 = n15798 ;
  assign y2399 = n15799 ;
  assign y2400 = n15802 ;
  assign y2401 = ~n15809 ;
  assign y2402 = ~n15814 ;
  assign y2403 = ~n15822 ;
  assign y2404 = ~n15825 ;
  assign y2405 = ~n15827 ;
  assign y2406 = ~n15831 ;
  assign y2407 = ~n15851 ;
  assign y2408 = ~n15858 ;
  assign y2409 = n15865 ;
  assign y2410 = ~n15869 ;
  assign y2411 = ~n15874 ;
  assign y2412 = ~n15883 ;
  assign y2413 = ~n15891 ;
  assign y2414 = ~n15893 ;
  assign y2415 = ~n15907 ;
  assign y2416 = ~n15910 ;
  assign y2417 = ~n15912 ;
  assign y2418 = ~n15914 ;
  assign y2419 = ~n15918 ;
  assign y2420 = ~1'b0 ;
  assign y2421 = n15928 ;
  assign y2422 = ~n15929 ;
  assign y2423 = ~n15930 ;
  assign y2424 = n15936 ;
  assign y2425 = n15950 ;
  assign y2426 = ~n15956 ;
  assign y2427 = n15962 ;
  assign y2428 = ~n15968 ;
  assign y2429 = ~n15971 ;
  assign y2430 = ~n15975 ;
  assign y2431 = ~n15987 ;
  assign y2432 = n15992 ;
  assign y2433 = ~n15993 ;
  assign y2434 = n15995 ;
  assign y2435 = ~n15999 ;
  assign y2436 = n16013 ;
  assign y2437 = n16033 ;
  assign y2438 = ~1'b0 ;
  assign y2439 = n16036 ;
  assign y2440 = n16041 ;
  assign y2441 = n16044 ;
  assign y2442 = ~n16064 ;
  assign y2443 = ~n16074 ;
  assign y2444 = ~n16078 ;
  assign y2445 = n16080 ;
  assign y2446 = ~n16083 ;
  assign y2447 = n16085 ;
  assign y2448 = ~n16088 ;
  assign y2449 = n16089 ;
  assign y2450 = n16107 ;
  assign y2451 = n16108 ;
  assign y2452 = ~n16113 ;
  assign y2453 = ~n16121 ;
  assign y2454 = ~n16127 ;
  assign y2455 = n16132 ;
  assign y2456 = ~n16147 ;
  assign y2457 = n16155 ;
  assign y2458 = ~n16163 ;
  assign y2459 = n16166 ;
  assign y2460 = n16174 ;
  assign y2461 = ~n16176 ;
  assign y2462 = n16182 ;
  assign y2463 = ~n16185 ;
  assign y2464 = n16200 ;
  assign y2465 = ~n16205 ;
  assign y2466 = n16206 ;
  assign y2467 = n16210 ;
  assign y2468 = ~n16214 ;
  assign y2469 = ~n16218 ;
  assign y2470 = n16229 ;
  assign y2471 = n16232 ;
  assign y2472 = n16238 ;
  assign y2473 = ~n16240 ;
  assign y2474 = n16241 ;
  assign y2475 = ~n16247 ;
  assign y2476 = n16255 ;
  assign y2477 = ~n16265 ;
  assign y2478 = n16266 ;
  assign y2479 = ~n16267 ;
  assign y2480 = n16276 ;
  assign y2481 = ~n16278 ;
  assign y2482 = n16279 ;
  assign y2483 = ~n16281 ;
  assign y2484 = ~n16294 ;
  assign y2485 = ~n16296 ;
  assign y2486 = n16317 ;
  assign y2487 = n16328 ;
  assign y2488 = n16331 ;
  assign y2489 = ~n16333 ;
  assign y2490 = ~n16349 ;
  assign y2491 = n16366 ;
  assign y2492 = n16373 ;
  assign y2493 = n16378 ;
  assign y2494 = n16384 ;
  assign y2495 = ~n16385 ;
  assign y2496 = ~n16387 ;
  assign y2497 = n16390 ;
  assign y2498 = n16394 ;
  assign y2499 = n16396 ;
  assign y2500 = ~n16399 ;
  assign y2501 = n16402 ;
  assign y2502 = ~n16405 ;
  assign y2503 = ~n16407 ;
  assign y2504 = n16417 ;
  assign y2505 = ~n16422 ;
  assign y2506 = n16426 ;
  assign y2507 = n16427 ;
  assign y2508 = n16431 ;
  assign y2509 = n16432 ;
  assign y2510 = ~n16437 ;
  assign y2511 = n16439 ;
  assign y2512 = ~n16444 ;
  assign y2513 = n16453 ;
  assign y2514 = ~1'b0 ;
  assign y2515 = ~n16456 ;
  assign y2516 = n16458 ;
  assign y2517 = n16465 ;
  assign y2518 = ~1'b0 ;
  assign y2519 = n16474 ;
  assign y2520 = ~n16486 ;
  assign y2521 = n16487 ;
  assign y2522 = ~1'b0 ;
  assign y2523 = ~n16502 ;
  assign y2524 = ~n16509 ;
  assign y2525 = ~n16521 ;
  assign y2526 = ~n16527 ;
  assign y2527 = ~n16532 ;
  assign y2528 = ~n16537 ;
  assign y2529 = ~n16539 ;
  assign y2530 = ~1'b0 ;
  assign y2531 = ~n16540 ;
  assign y2532 = ~n16551 ;
  assign y2533 = ~n16552 ;
  assign y2534 = n16553 ;
  assign y2535 = n16557 ;
  assign y2536 = ~n16559 ;
  assign y2537 = ~n16566 ;
  assign y2538 = ~n16573 ;
  assign y2539 = n16575 ;
  assign y2540 = ~n16588 ;
  assign y2541 = n16590 ;
  assign y2542 = ~n16594 ;
  assign y2543 = ~n16596 ;
  assign y2544 = n16597 ;
  assign y2545 = n16600 ;
  assign y2546 = ~1'b0 ;
  assign y2547 = ~n16613 ;
  assign y2548 = ~n16630 ;
  assign y2549 = n16633 ;
  assign y2550 = n16634 ;
  assign y2551 = ~n16637 ;
  assign y2552 = ~n16639 ;
  assign y2553 = ~n16642 ;
  assign y2554 = ~n16646 ;
  assign y2555 = n16649 ;
  assign y2556 = ~n16663 ;
  assign y2557 = n16664 ;
  assign y2558 = n16666 ;
  assign y2559 = ~n16667 ;
  assign y2560 = n16669 ;
  assign y2561 = n16671 ;
  assign y2562 = n16674 ;
  assign y2563 = n16677 ;
  assign y2564 = ~n16683 ;
  assign y2565 = n16688 ;
  assign y2566 = ~n16691 ;
  assign y2567 = n16695 ;
  assign y2568 = ~n16697 ;
  assign y2569 = n16704 ;
  assign y2570 = n16706 ;
  assign y2571 = n16715 ;
  assign y2572 = ~n16719 ;
  assign y2573 = n16728 ;
  assign y2574 = n16731 ;
  assign y2575 = n16735 ;
  assign y2576 = n16739 ;
  assign y2577 = n16742 ;
  assign y2578 = n16745 ;
  assign y2579 = n16752 ;
  assign y2580 = ~1'b0 ;
  assign y2581 = ~n16759 ;
  assign y2582 = n16776 ;
  assign y2583 = ~n16777 ;
  assign y2584 = ~n16778 ;
  assign y2585 = ~n16780 ;
  assign y2586 = ~n16781 ;
  assign y2587 = ~n16795 ;
  assign y2588 = n16798 ;
  assign y2589 = n16804 ;
  assign y2590 = n16807 ;
  assign y2591 = n16809 ;
  assign y2592 = ~n16813 ;
  assign y2593 = ~n16818 ;
  assign y2594 = n16831 ;
  assign y2595 = n16833 ;
  assign y2596 = n16837 ;
  assign y2597 = n16848 ;
  assign y2598 = ~n16852 ;
  assign y2599 = n16859 ;
  assign y2600 = n16862 ;
  assign y2601 = n16870 ;
  assign y2602 = ~n16871 ;
  assign y2603 = n16878 ;
  assign y2604 = ~n16889 ;
  assign y2605 = n16891 ;
  assign y2606 = ~n16897 ;
  assign y2607 = ~n16902 ;
  assign y2608 = n16903 ;
  assign y2609 = ~n16915 ;
  assign y2610 = n16921 ;
  assign y2611 = ~n16923 ;
  assign y2612 = n16928 ;
  assign y2613 = n16929 ;
  assign y2614 = n16931 ;
  assign y2615 = n16933 ;
  assign y2616 = ~n16937 ;
  assign y2617 = ~n16946 ;
  assign y2618 = ~n16949 ;
  assign y2619 = n16952 ;
  assign y2620 = ~n16953 ;
  assign y2621 = n16973 ;
  assign y2622 = ~n16981 ;
  assign y2623 = ~n16994 ;
  assign y2624 = ~n16996 ;
  assign y2625 = n17001 ;
  assign y2626 = ~n17003 ;
  assign y2627 = n17004 ;
  assign y2628 = ~n17008 ;
  assign y2629 = ~1'b0 ;
  assign y2630 = ~n17012 ;
  assign y2631 = n17013 ;
  assign y2632 = ~n17021 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = ~n17032 ;
  assign y2635 = ~n17035 ;
  assign y2636 = n17036 ;
  assign y2637 = n17038 ;
  assign y2638 = ~n17041 ;
  assign y2639 = ~n17044 ;
  assign y2640 = ~1'b0 ;
  assign y2641 = ~n17064 ;
  assign y2642 = n17070 ;
  assign y2643 = ~n17071 ;
  assign y2644 = n17081 ;
  assign y2645 = ~1'b0 ;
  assign y2646 = ~n17086 ;
  assign y2647 = ~n17089 ;
  assign y2648 = ~n17091 ;
  assign y2649 = n17093 ;
  assign y2650 = ~n17096 ;
  assign y2651 = n17102 ;
  assign y2652 = ~n17104 ;
  assign y2653 = n17106 ;
  assign y2654 = ~n17112 ;
  assign y2655 = ~n17113 ;
  assign y2656 = n17116 ;
  assign y2657 = ~n17126 ;
  assign y2658 = n17134 ;
  assign y2659 = n17144 ;
  assign y2660 = n17148 ;
  assign y2661 = n17152 ;
  assign y2662 = n17170 ;
  assign y2663 = n17176 ;
  assign y2664 = ~n17190 ;
  assign y2665 = n17191 ;
  assign y2666 = ~n17195 ;
  assign y2667 = ~1'b0 ;
  assign y2668 = n17196 ;
  assign y2669 = ~n17205 ;
  assign y2670 = n17206 ;
  assign y2671 = ~n17225 ;
  assign y2672 = n17229 ;
  assign y2673 = ~n17230 ;
  assign y2674 = ~1'b0 ;
  assign y2675 = n17235 ;
  assign y2676 = n17239 ;
  assign y2677 = n17240 ;
  assign y2678 = n17249 ;
  assign y2679 = ~n17250 ;
  assign y2680 = n17256 ;
  assign y2681 = n17257 ;
  assign y2682 = ~n17258 ;
  assign y2683 = ~n17260 ;
  assign y2684 = n17268 ;
  assign y2685 = n17272 ;
  assign y2686 = ~n17274 ;
  assign y2687 = n17296 ;
  assign y2688 = ~n17297 ;
  assign y2689 = n17300 ;
  assign y2690 = ~n17306 ;
  assign y2691 = ~n17316 ;
  assign y2692 = ~n17325 ;
  assign y2693 = n17329 ;
  assign y2694 = ~n17341 ;
  assign y2695 = ~n17342 ;
  assign y2696 = ~n17344 ;
  assign y2697 = n17352 ;
  assign y2698 = ~n17358 ;
  assign y2699 = ~n17361 ;
  assign y2700 = n17367 ;
  assign y2701 = ~n17368 ;
  assign y2702 = ~n17372 ;
  assign y2703 = n17384 ;
  assign y2704 = ~n17385 ;
  assign y2705 = ~n17391 ;
  assign y2706 = ~n17393 ;
  assign y2707 = ~n17396 ;
  assign y2708 = ~n17399 ;
  assign y2709 = n17400 ;
  assign y2710 = ~n17404 ;
  assign y2711 = n17428 ;
  assign y2712 = n17433 ;
  assign y2713 = n17437 ;
  assign y2714 = n17444 ;
  assign y2715 = ~n17448 ;
  assign y2716 = n17450 ;
  assign y2717 = n17455 ;
  assign y2718 = ~n17462 ;
  assign y2719 = ~1'b0 ;
  assign y2720 = n17466 ;
  assign y2721 = n17473 ;
  assign y2722 = ~n17483 ;
  assign y2723 = n17494 ;
  assign y2724 = ~n17500 ;
  assign y2725 = ~n17502 ;
  assign y2726 = ~n17506 ;
  assign y2727 = n17514 ;
  assign y2728 = ~n17523 ;
  assign y2729 = n17537 ;
  assign y2730 = ~n17538 ;
  assign y2731 = n17543 ;
  assign y2732 = n17550 ;
  assign y2733 = n17556 ;
  assign y2734 = ~n17557 ;
  assign y2735 = ~n17566 ;
  assign y2736 = n17573 ;
  assign y2737 = ~n17575 ;
  assign y2738 = ~n17589 ;
  assign y2739 = ~n17601 ;
  assign y2740 = ~n17607 ;
  assign y2741 = ~1'b0 ;
  assign y2742 = ~n17616 ;
  assign y2743 = ~n17619 ;
  assign y2744 = ~n17625 ;
  assign y2745 = n17630 ;
  assign y2746 = n17633 ;
  assign y2747 = ~n17638 ;
  assign y2748 = n17643 ;
  assign y2749 = ~n17664 ;
  assign y2750 = n17669 ;
  assign y2751 = ~n17675 ;
  assign y2752 = n17679 ;
  assign y2753 = ~n17686 ;
  assign y2754 = n17688 ;
  assign y2755 = ~n17689 ;
  assign y2756 = ~n17692 ;
  assign y2757 = n17694 ;
  assign y2758 = n17700 ;
  assign y2759 = ~n17703 ;
  assign y2760 = n17713 ;
  assign y2761 = n17725 ;
  assign y2762 = n17729 ;
  assign y2763 = n17730 ;
  assign y2764 = ~n17733 ;
  assign y2765 = n17736 ;
  assign y2766 = n17742 ;
  assign y2767 = ~n17744 ;
  assign y2768 = n17748 ;
  assign y2769 = n17750 ;
  assign y2770 = ~n17751 ;
  assign y2771 = ~n17752 ;
  assign y2772 = n17755 ;
  assign y2773 = ~n17757 ;
  assign y2774 = n17759 ;
  assign y2775 = n17761 ;
  assign y2776 = n17772 ;
  assign y2777 = n17773 ;
  assign y2778 = ~n17775 ;
  assign y2779 = ~n17778 ;
  assign y2780 = n17782 ;
  assign y2781 = ~n17783 ;
  assign y2782 = ~n17786 ;
  assign y2783 = n17796 ;
  assign y2784 = n17811 ;
  assign y2785 = ~n17812 ;
  assign y2786 = n17827 ;
  assign y2787 = ~n17842 ;
  assign y2788 = ~1'b0 ;
  assign y2789 = ~n17851 ;
  assign y2790 = n17852 ;
  assign y2791 = ~n17855 ;
  assign y2792 = ~n17856 ;
  assign y2793 = n17863 ;
  assign y2794 = n17870 ;
  assign y2795 = n17876 ;
  assign y2796 = n17878 ;
  assign y2797 = n17879 ;
  assign y2798 = n17883 ;
  assign y2799 = ~n17885 ;
  assign y2800 = n17892 ;
  assign y2801 = n17894 ;
  assign y2802 = ~n17898 ;
  assign y2803 = n17899 ;
  assign y2804 = ~n17904 ;
  assign y2805 = n17905 ;
  assign y2806 = ~n17906 ;
  assign y2807 = ~n17908 ;
  assign y2808 = ~n17910 ;
  assign y2809 = n17914 ;
  assign y2810 = ~n17915 ;
  assign y2811 = n17920 ;
  assign y2812 = ~n17921 ;
  assign y2813 = n17928 ;
  assign y2814 = ~n17929 ;
  assign y2815 = ~n17935 ;
  assign y2816 = ~n17941 ;
  assign y2817 = ~n17944 ;
  assign y2818 = n17945 ;
  assign y2819 = ~n17950 ;
  assign y2820 = n17956 ;
  assign y2821 = ~1'b0 ;
  assign y2822 = ~1'b0 ;
  assign y2823 = n17958 ;
  assign y2824 = n17962 ;
  assign y2825 = n17969 ;
  assign y2826 = ~n17970 ;
  assign y2827 = ~n17980 ;
  assign y2828 = ~n17993 ;
  assign y2829 = ~n17995 ;
  assign y2830 = ~n18000 ;
  assign y2831 = ~n18004 ;
  assign y2832 = n18010 ;
  assign y2833 = n18011 ;
  assign y2834 = ~n18013 ;
  assign y2835 = n18020 ;
  assign y2836 = ~n18024 ;
  assign y2837 = n18027 ;
  assign y2838 = n18028 ;
  assign y2839 = ~n18032 ;
  assign y2840 = n18035 ;
  assign y2841 = ~n18036 ;
  assign y2842 = n18037 ;
  assign y2843 = ~n18047 ;
  assign y2844 = n18049 ;
  assign y2845 = n18056 ;
  assign y2846 = n18062 ;
  assign y2847 = ~n18067 ;
  assign y2848 = ~n18070 ;
  assign y2849 = ~n18072 ;
  assign y2850 = n18076 ;
  assign y2851 = n18087 ;
  assign y2852 = ~n18095 ;
  assign y2853 = ~n18099 ;
  assign y2854 = ~n18108 ;
  assign y2855 = n18120 ;
  assign y2856 = ~n18122 ;
  assign y2857 = ~n18124 ;
  assign y2858 = ~n18130 ;
  assign y2859 = n18134 ;
  assign y2860 = n18135 ;
  assign y2861 = ~n18136 ;
  assign y2862 = ~n18138 ;
  assign y2863 = ~1'b0 ;
  assign y2864 = n18141 ;
  assign y2865 = n18143 ;
  assign y2866 = ~1'b0 ;
  assign y2867 = n18148 ;
  assign y2868 = ~1'b0 ;
  assign y2869 = n18164 ;
  assign y2870 = n18169 ;
  assign y2871 = ~n18174 ;
  assign y2872 = n18176 ;
  assign y2873 = n18179 ;
  assign y2874 = n18180 ;
  assign y2875 = ~n18185 ;
  assign y2876 = n18189 ;
  assign y2877 = ~n18190 ;
  assign y2878 = ~n18192 ;
  assign y2879 = ~n18194 ;
  assign y2880 = ~n18201 ;
  assign y2881 = n18204 ;
  assign y2882 = n18207 ;
  assign y2883 = ~n18208 ;
  assign y2884 = n18212 ;
  assign y2885 = ~n18220 ;
  assign y2886 = ~1'b0 ;
  assign y2887 = ~n18227 ;
  assign y2888 = n18233 ;
  assign y2889 = ~n18236 ;
  assign y2890 = ~n18243 ;
  assign y2891 = n18248 ;
  assign y2892 = n18250 ;
  assign y2893 = n18254 ;
  assign y2894 = ~n18258 ;
  assign y2895 = ~n18264 ;
  assign y2896 = n18265 ;
  assign y2897 = ~n18268 ;
  assign y2898 = ~n18278 ;
  assign y2899 = ~n18287 ;
  assign y2900 = n18289 ;
  assign y2901 = ~n18291 ;
  assign y2902 = n18297 ;
  assign y2903 = ~n18302 ;
  assign y2904 = ~n18308 ;
  assign y2905 = n18312 ;
  assign y2906 = n18316 ;
  assign y2907 = ~n18319 ;
  assign y2908 = ~n18320 ;
  assign y2909 = ~n18322 ;
  assign y2910 = ~n18323 ;
  assign y2911 = n18330 ;
  assign y2912 = ~n18335 ;
  assign y2913 = ~n18339 ;
  assign y2914 = ~n18340 ;
  assign y2915 = ~n18346 ;
  assign y2916 = ~n18350 ;
  assign y2917 = n18351 ;
  assign y2918 = ~n18354 ;
  assign y2919 = n18355 ;
  assign y2920 = n18357 ;
  assign y2921 = n18365 ;
  assign y2922 = ~1'b0 ;
  assign y2923 = ~n18366 ;
  assign y2924 = ~n18374 ;
  assign y2925 = n18379 ;
  assign y2926 = n18384 ;
  assign y2927 = ~1'b0 ;
  assign y2928 = n18387 ;
  assign y2929 = ~n18395 ;
  assign y2930 = ~n18398 ;
  assign y2931 = n18399 ;
  assign y2932 = n18400 ;
  assign y2933 = ~n18401 ;
  assign y2934 = n18407 ;
  assign y2935 = n18417 ;
  assign y2936 = n18421 ;
  assign y2937 = n18423 ;
  assign y2938 = ~n18424 ;
  assign y2939 = n18426 ;
  assign y2940 = n18428 ;
  assign y2941 = ~n18440 ;
  assign y2942 = n18446 ;
  assign y2943 = ~n18449 ;
  assign y2944 = ~n18452 ;
  assign y2945 = n18458 ;
  assign y2946 = n18465 ;
  assign y2947 = ~n18470 ;
  assign y2948 = n18476 ;
  assign y2949 = ~n18477 ;
  assign y2950 = ~n18481 ;
  assign y2951 = n18484 ;
  assign y2952 = ~1'b0 ;
  assign y2953 = ~n18497 ;
  assign y2954 = ~n18499 ;
  assign y2955 = ~n18508 ;
  assign y2956 = n18513 ;
  assign y2957 = ~n18515 ;
  assign y2958 = n18544 ;
  assign y2959 = n18551 ;
  assign y2960 = ~n18554 ;
  assign y2961 = n18555 ;
  assign y2962 = n18556 ;
  assign y2963 = n18559 ;
  assign y2964 = ~n18567 ;
  assign y2965 = ~n18568 ;
  assign y2966 = ~n18573 ;
  assign y2967 = ~n18579 ;
  assign y2968 = n18596 ;
  assign y2969 = ~n18599 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = n18600 ;
  assign y2972 = ~n18611 ;
  assign y2973 = ~n18613 ;
  assign y2974 = ~n18615 ;
  assign y2975 = n18617 ;
  assign y2976 = n18622 ;
  assign y2977 = ~n18623 ;
  assign y2978 = ~n18630 ;
  assign y2979 = n18631 ;
  assign y2980 = ~n18638 ;
  assign y2981 = n18639 ;
  assign y2982 = ~n18644 ;
  assign y2983 = n18649 ;
  assign y2984 = n18652 ;
  assign y2985 = ~n18655 ;
  assign y2986 = n18657 ;
  assign y2987 = n18661 ;
  assign y2988 = ~n18664 ;
  assign y2989 = ~n18669 ;
  assign y2990 = ~n18685 ;
  assign y2991 = n18694 ;
  assign y2992 = ~n18697 ;
  assign y2993 = ~n18698 ;
  assign y2994 = ~1'b0 ;
  assign y2995 = n18699 ;
  assign y2996 = n18704 ;
  assign y2997 = n18705 ;
  assign y2998 = n18708 ;
  assign y2999 = ~n18710 ;
  assign y3000 = ~n18712 ;
  assign y3001 = ~n18716 ;
  assign y3002 = n18731 ;
  assign y3003 = ~n18736 ;
  assign y3004 = ~n18748 ;
  assign y3005 = ~n18754 ;
  assign y3006 = ~n18757 ;
  assign y3007 = ~n18759 ;
  assign y3008 = n18761 ;
  assign y3009 = ~n18762 ;
  assign y3010 = ~n18763 ;
  assign y3011 = n18765 ;
  assign y3012 = n18770 ;
  assign y3013 = n18776 ;
  assign y3014 = ~n18783 ;
  assign y3015 = n18789 ;
  assign y3016 = ~n18793 ;
  assign y3017 = n18794 ;
  assign y3018 = ~n18798 ;
  assign y3019 = n18807 ;
  assign y3020 = ~n18810 ;
  assign y3021 = n18811 ;
  assign y3022 = n18814 ;
  assign y3023 = ~n18815 ;
  assign y3024 = ~n18826 ;
  assign y3025 = n18833 ;
  assign y3026 = ~n18840 ;
  assign y3027 = ~n18841 ;
  assign y3028 = n18844 ;
  assign y3029 = ~1'b0 ;
  assign y3030 = n18845 ;
  assign y3031 = ~n18847 ;
  assign y3032 = n18852 ;
  assign y3033 = ~n18858 ;
  assign y3034 = ~n18863 ;
  assign y3035 = n18865 ;
  assign y3036 = n18866 ;
  assign y3037 = n18867 ;
  assign y3038 = ~n18873 ;
  assign y3039 = ~n18879 ;
  assign y3040 = ~n18883 ;
  assign y3041 = ~n18885 ;
  assign y3042 = ~1'b0 ;
  assign y3043 = ~n18890 ;
  assign y3044 = n18899 ;
  assign y3045 = ~n18903 ;
  assign y3046 = n18909 ;
  assign y3047 = ~n18911 ;
  assign y3048 = n18914 ;
  assign y3049 = ~n18922 ;
  assign y3050 = n18955 ;
  assign y3051 = ~n18957 ;
  assign y3052 = ~n18977 ;
  assign y3053 = ~n18980 ;
  assign y3054 = ~n18985 ;
  assign y3055 = ~n18986 ;
  assign y3056 = n18991 ;
  assign y3057 = n18992 ;
  assign y3058 = n18997 ;
  assign y3059 = ~n19002 ;
  assign y3060 = n19006 ;
  assign y3061 = n19008 ;
  assign y3062 = n19011 ;
  assign y3063 = ~n19012 ;
  assign y3064 = ~n19016 ;
  assign y3065 = ~n19020 ;
  assign y3066 = n19024 ;
  assign y3067 = ~n19032 ;
  assign y3068 = n19033 ;
  assign y3069 = ~n19040 ;
  assign y3070 = ~1'b0 ;
  assign y3071 = n19045 ;
  assign y3072 = ~n19049 ;
  assign y3073 = n19058 ;
  assign y3074 = n19059 ;
  assign y3075 = n19072 ;
  assign y3076 = n19078 ;
  assign y3077 = n19083 ;
  assign y3078 = n19087 ;
  assign y3079 = ~n19109 ;
  assign y3080 = ~n19113 ;
  assign y3081 = ~n19114 ;
  assign y3082 = n19118 ;
  assign y3083 = ~n19125 ;
  assign y3084 = ~n19126 ;
  assign y3085 = n19128 ;
  assign y3086 = n19138 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = ~n19143 ;
  assign y3089 = ~n19154 ;
  assign y3090 = ~n19155 ;
  assign y3091 = ~n19157 ;
  assign y3092 = ~n19170 ;
  assign y3093 = n19171 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = n19174 ;
  assign y3096 = ~n19176 ;
  assign y3097 = n19177 ;
  assign y3098 = n19186 ;
  assign y3099 = n19187 ;
  assign y3100 = n19189 ;
  assign y3101 = ~n19191 ;
  assign y3102 = n19195 ;
  assign y3103 = n19200 ;
  assign y3104 = ~1'b0 ;
  assign y3105 = ~n19207 ;
  assign y3106 = ~n19208 ;
  assign y3107 = ~n19215 ;
  assign y3108 = ~n19216 ;
  assign y3109 = n19218 ;
  assign y3110 = ~n19221 ;
  assign y3111 = ~n19222 ;
  assign y3112 = ~n19223 ;
  assign y3113 = n19224 ;
  assign y3114 = ~n19226 ;
  assign y3115 = ~n19227 ;
  assign y3116 = n19234 ;
  assign y3117 = ~n19236 ;
  assign y3118 = ~n19241 ;
  assign y3119 = n19248 ;
  assign y3120 = n19254 ;
  assign y3121 = ~n19257 ;
  assign y3122 = n19259 ;
  assign y3123 = ~n19261 ;
  assign y3124 = n19269 ;
  assign y3125 = ~n19277 ;
  assign y3126 = ~n19283 ;
  assign y3127 = ~n19296 ;
  assign y3128 = ~n19298 ;
  assign y3129 = ~n19301 ;
  assign y3130 = ~n19304 ;
  assign y3131 = n19310 ;
  assign y3132 = n19311 ;
  assign y3133 = ~n19318 ;
  assign y3134 = n19327 ;
  assign y3135 = ~n19333 ;
  assign y3136 = ~n19337 ;
  assign y3137 = ~n19338 ;
  assign y3138 = ~n19348 ;
  assign y3139 = ~n19360 ;
  assign y3140 = ~n19362 ;
  assign y3141 = ~n19366 ;
  assign y3142 = ~n19368 ;
  assign y3143 = ~n19371 ;
  assign y3144 = n19374 ;
  assign y3145 = n19379 ;
  assign y3146 = ~n19382 ;
  assign y3147 = ~n19387 ;
  assign y3148 = n19391 ;
  assign y3149 = ~n19395 ;
  assign y3150 = ~n19396 ;
  assign y3151 = ~n19413 ;
  assign y3152 = ~1'b0 ;
  assign y3153 = ~1'b0 ;
  assign y3154 = n19417 ;
  assign y3155 = n19422 ;
  assign y3156 = ~n19423 ;
  assign y3157 = n19428 ;
  assign y3158 = ~n19431 ;
  assign y3159 = ~n19433 ;
  assign y3160 = n19439 ;
  assign y3161 = n19444 ;
  assign y3162 = ~1'b0 ;
  assign y3163 = ~n19446 ;
  assign y3164 = n19458 ;
  assign y3165 = ~n19461 ;
  assign y3166 = ~n19464 ;
  assign y3167 = n19465 ;
  assign y3168 = ~n19468 ;
  assign y3169 = ~n19473 ;
  assign y3170 = ~n19474 ;
  assign y3171 = ~1'b0 ;
  assign y3172 = ~n19476 ;
  assign y3173 = n19487 ;
  assign y3174 = n19489 ;
  assign y3175 = ~n19496 ;
  assign y3176 = n19503 ;
  assign y3177 = n19508 ;
  assign y3178 = n19515 ;
  assign y3179 = ~n19518 ;
  assign y3180 = ~n19524 ;
  assign y3181 = ~n19526 ;
  assign y3182 = ~n19531 ;
  assign y3183 = n19533 ;
  assign y3184 = n19536 ;
  assign y3185 = ~n19539 ;
  assign y3186 = n19550 ;
  assign y3187 = n19554 ;
  assign y3188 = ~n19560 ;
  assign y3189 = ~n19563 ;
  assign y3190 = ~n19569 ;
  assign y3191 = n19571 ;
  assign y3192 = ~n19574 ;
  assign y3193 = n19576 ;
  assign y3194 = n19580 ;
  assign y3195 = n19581 ;
  assign y3196 = ~n19584 ;
  assign y3197 = ~n19587 ;
  assign y3198 = ~n19599 ;
  assign y3199 = ~n19603 ;
  assign y3200 = ~n19605 ;
  assign y3201 = ~n19609 ;
  assign y3202 = n19611 ;
  assign y3203 = n19617 ;
  assign y3204 = n19622 ;
  assign y3205 = ~n19636 ;
  assign y3206 = ~n19638 ;
  assign y3207 = ~n19642 ;
  assign y3208 = n19644 ;
  assign y3209 = n19645 ;
  assign y3210 = n19647 ;
  assign y3211 = ~n19648 ;
  assign y3212 = ~1'b0 ;
  assign y3213 = ~1'b0 ;
  assign y3214 = ~n19651 ;
  assign y3215 = n19669 ;
  assign y3216 = n19671 ;
  assign y3217 = n19679 ;
  assign y3218 = n19687 ;
  assign y3219 = ~n19697 ;
  assign y3220 = ~n19699 ;
  assign y3221 = ~n19701 ;
  assign y3222 = n19705 ;
  assign y3223 = ~n19713 ;
  assign y3224 = n19715 ;
  assign y3225 = n19724 ;
  assign y3226 = n19725 ;
  assign y3227 = n19732 ;
  assign y3228 = n19738 ;
  assign y3229 = ~n19743 ;
  assign y3230 = n19750 ;
  assign y3231 = ~n19751 ;
  assign y3232 = n19755 ;
  assign y3233 = n19758 ;
  assign y3234 = n19764 ;
  assign y3235 = ~n19780 ;
  assign y3236 = ~n19784 ;
  assign y3237 = n19792 ;
  assign y3238 = n19795 ;
  assign y3239 = n19801 ;
  assign y3240 = ~n19807 ;
  assign y3241 = ~n19822 ;
  assign y3242 = n19837 ;
  assign y3243 = n19842 ;
  assign y3244 = ~n19852 ;
  assign y3245 = ~n19855 ;
  assign y3246 = n19856 ;
  assign y3247 = ~n19865 ;
  assign y3248 = ~n19873 ;
  assign y3249 = n19878 ;
  assign y3250 = n19879 ;
  assign y3251 = ~n19881 ;
  assign y3252 = ~n19882 ;
  assign y3253 = ~n19883 ;
  assign y3254 = n19884 ;
  assign y3255 = n19885 ;
  assign y3256 = ~n19890 ;
  assign y3257 = ~n19895 ;
  assign y3258 = n19896 ;
  assign y3259 = n19897 ;
  assign y3260 = n19899 ;
  assign y3261 = n19900 ;
  assign y3262 = n19902 ;
  assign y3263 = ~n19905 ;
  assign y3264 = ~n19908 ;
  assign y3265 = ~n19912 ;
  assign y3266 = ~n19915 ;
  assign y3267 = ~n19927 ;
  assign y3268 = ~n19928 ;
  assign y3269 = ~n19931 ;
  assign y3270 = ~1'b0 ;
  assign y3271 = n19933 ;
  assign y3272 = ~n19940 ;
  assign y3273 = n19943 ;
  assign y3274 = n19949 ;
  assign y3275 = n19958 ;
  assign y3276 = n19967 ;
  assign y3277 = ~n19973 ;
  assign y3278 = ~n19980 ;
  assign y3279 = n19992 ;
  assign y3280 = ~n19994 ;
  assign y3281 = n19998 ;
  assign y3282 = n19999 ;
  assign y3283 = n20012 ;
  assign y3284 = n20017 ;
  assign y3285 = n20023 ;
  assign y3286 = ~n20025 ;
  assign y3287 = ~n20036 ;
  assign y3288 = ~n20049 ;
  assign y3289 = n20056 ;
  assign y3290 = ~n20058 ;
  assign y3291 = n20064 ;
  assign y3292 = ~1'b0 ;
  assign y3293 = n20065 ;
  assign y3294 = n20067 ;
  assign y3295 = n20074 ;
  assign y3296 = n20077 ;
  assign y3297 = ~n20078 ;
  assign y3298 = ~n20080 ;
  assign y3299 = ~n20089 ;
  assign y3300 = ~n20093 ;
  assign y3301 = ~n20110 ;
  assign y3302 = n20115 ;
  assign y3303 = ~n20127 ;
  assign y3304 = n20129 ;
  assign y3305 = ~n20132 ;
  assign y3306 = ~n20134 ;
  assign y3307 = n20139 ;
  assign y3308 = n20142 ;
  assign y3309 = ~n20146 ;
  assign y3310 = ~n20147 ;
  assign y3311 = ~n20153 ;
  assign y3312 = ~n20155 ;
  assign y3313 = n20159 ;
  assign y3314 = ~n20161 ;
  assign y3315 = n20169 ;
  assign y3316 = ~n20173 ;
  assign y3317 = ~n20174 ;
  assign y3318 = n20178 ;
  assign y3319 = n20179 ;
  assign y3320 = n20185 ;
  assign y3321 = ~n20191 ;
  assign y3322 = n20197 ;
  assign y3323 = ~n20199 ;
  assign y3324 = ~n20205 ;
  assign y3325 = ~n20211 ;
  assign y3326 = n20215 ;
  assign y3327 = n20218 ;
  assign y3328 = n20221 ;
  assign y3329 = n20224 ;
  assign y3330 = n20230 ;
  assign y3331 = ~n20231 ;
  assign y3332 = n20237 ;
  assign y3333 = ~n20239 ;
  assign y3334 = n20245 ;
  assign y3335 = ~n20246 ;
  assign y3336 = ~n20250 ;
  assign y3337 = ~n20255 ;
  assign y3338 = n20260 ;
  assign y3339 = n20262 ;
  assign y3340 = ~n20265 ;
  assign y3341 = ~n20277 ;
  assign y3342 = ~n20279 ;
  assign y3343 = ~n20283 ;
  assign y3344 = n20285 ;
  assign y3345 = n20287 ;
  assign y3346 = ~n20301 ;
  assign y3347 = ~n20303 ;
  assign y3348 = n20306 ;
  assign y3349 = n20313 ;
  assign y3350 = ~1'b0 ;
  assign y3351 = n20317 ;
  assign y3352 = n20318 ;
  assign y3353 = n20321 ;
  assign y3354 = ~n20328 ;
  assign y3355 = n20331 ;
  assign y3356 = ~n20335 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = n20336 ;
  assign y3359 = ~n20337 ;
  assign y3360 = ~n20338 ;
  assign y3361 = ~n20348 ;
  assign y3362 = ~n12168 ;
  assign y3363 = n20355 ;
  assign y3364 = n20356 ;
  assign y3365 = ~n20358 ;
  assign y3366 = ~1'b0 ;
  assign y3367 = ~n20359 ;
  assign y3368 = ~n20362 ;
  assign y3369 = ~n20366 ;
  assign y3370 = ~n20371 ;
  assign y3371 = ~1'b0 ;
  assign y3372 = n20372 ;
  assign y3373 = ~n20382 ;
  assign y3374 = n20383 ;
  assign y3375 = n20385 ;
  assign y3376 = ~n20386 ;
  assign y3377 = n20389 ;
  assign y3378 = n20390 ;
  assign y3379 = ~n20392 ;
  assign y3380 = n20393 ;
  assign y3381 = n20396 ;
  assign y3382 = n20399 ;
  assign y3383 = ~n20404 ;
  assign y3384 = n20406 ;
  assign y3385 = ~1'b0 ;
  assign y3386 = n20408 ;
  assign y3387 = n20411 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = ~n20413 ;
  assign y3390 = ~n20422 ;
  assign y3391 = n20428 ;
  assign y3392 = n17505 ;
  assign y3393 = n20430 ;
  assign y3394 = n20435 ;
  assign y3395 = n20438 ;
  assign y3396 = n20443 ;
  assign y3397 = n20449 ;
  assign y3398 = ~n20452 ;
  assign y3399 = n20457 ;
  assign y3400 = n20462 ;
  assign y3401 = n20465 ;
  assign y3402 = ~n20471 ;
  assign y3403 = n20475 ;
  assign y3404 = n20477 ;
  assign y3405 = ~n20482 ;
  assign y3406 = ~n20489 ;
  assign y3407 = n20496 ;
  assign y3408 = ~n20499 ;
  assign y3409 = ~n20500 ;
  assign y3410 = ~n20502 ;
  assign y3411 = ~n20504 ;
  assign y3412 = ~n20516 ;
  assign y3413 = n20519 ;
  assign y3414 = ~n20520 ;
  assign y3415 = n20526 ;
  assign y3416 = ~1'b0 ;
  assign y3417 = ~n20527 ;
  assign y3418 = n20543 ;
  assign y3419 = ~n20552 ;
  assign y3420 = ~n20565 ;
  assign y3421 = n20566 ;
  assign y3422 = ~n20568 ;
  assign y3423 = n20569 ;
  assign y3424 = n20571 ;
  assign y3425 = ~n20579 ;
  assign y3426 = ~n20580 ;
  assign y3427 = ~n20581 ;
  assign y3428 = ~n20583 ;
  assign y3429 = ~n20595 ;
  assign y3430 = ~n20596 ;
  assign y3431 = n20603 ;
  assign y3432 = ~n20607 ;
  assign y3433 = ~n20612 ;
  assign y3434 = n20613 ;
  assign y3435 = ~n20616 ;
  assign y3436 = ~n20631 ;
  assign y3437 = ~n20637 ;
  assign y3438 = n20638 ;
  assign y3439 = ~n20642 ;
  assign y3440 = ~1'b0 ;
  assign y3441 = n20648 ;
  assign y3442 = ~n20655 ;
  assign y3443 = ~n20658 ;
  assign y3444 = ~n20664 ;
  assign y3445 = n20667 ;
  assign y3446 = ~n20669 ;
  assign y3447 = n20675 ;
  assign y3448 = n20677 ;
  assign y3449 = ~n20685 ;
  assign y3450 = n20687 ;
  assign y3451 = ~n20689 ;
  assign y3452 = n20693 ;
  assign y3453 = n20695 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = n20696 ;
  assign y3456 = ~n20698 ;
  assign y3457 = ~n20701 ;
  assign y3458 = ~n20704 ;
  assign y3459 = n20705 ;
  assign y3460 = ~n20706 ;
  assign y3461 = n20709 ;
  assign y3462 = n20711 ;
  assign y3463 = ~1'b0 ;
  assign y3464 = n20712 ;
  assign y3465 = ~n20713 ;
  assign y3466 = ~n20720 ;
  assign y3467 = n20727 ;
  assign y3468 = ~n20734 ;
  assign y3469 = n20739 ;
  assign y3470 = ~n20741 ;
  assign y3471 = ~n20742 ;
  assign y3472 = n20747 ;
  assign y3473 = n20755 ;
  assign y3474 = n20757 ;
  assign y3475 = ~n20758 ;
  assign y3476 = n20760 ;
  assign y3477 = ~n20767 ;
  assign y3478 = n20769 ;
  assign y3479 = n20779 ;
  assign y3480 = ~n20790 ;
  assign y3481 = ~n20793 ;
  assign y3482 = n20799 ;
  assign y3483 = ~n20805 ;
  assign y3484 = ~n20807 ;
  assign y3485 = ~n20820 ;
  assign y3486 = ~n20822 ;
  assign y3487 = ~n20831 ;
  assign y3488 = n20832 ;
  assign y3489 = ~n20849 ;
  assign y3490 = ~n20850 ;
  assign y3491 = n20852 ;
  assign y3492 = ~n20854 ;
  assign y3493 = ~n20855 ;
  assign y3494 = ~n20856 ;
  assign y3495 = n20861 ;
  assign y3496 = ~1'b0 ;
  assign y3497 = ~n20866 ;
  assign y3498 = n20871 ;
  assign y3499 = n20872 ;
  assign y3500 = n20873 ;
  assign y3501 = n20877 ;
  assign y3502 = ~n20878 ;
  assign y3503 = n20882 ;
  assign y3504 = n20889 ;
  assign y3505 = n20891 ;
  assign y3506 = ~n20899 ;
  assign y3507 = n20905 ;
  assign y3508 = ~n20909 ;
  assign y3509 = ~n20912 ;
  assign y3510 = n20919 ;
  assign y3511 = ~1'b0 ;
  assign y3512 = ~n20921 ;
  assign y3513 = n20926 ;
  assign y3514 = ~n20932 ;
  assign y3515 = ~n20948 ;
  assign y3516 = n20956 ;
  assign y3517 = ~1'b0 ;
  assign y3518 = n20958 ;
  assign y3519 = n20959 ;
  assign y3520 = ~n20966 ;
  assign y3521 = ~n20976 ;
  assign y3522 = ~n20979 ;
  assign y3523 = n20981 ;
  assign y3524 = ~n20983 ;
  assign y3525 = ~1'b0 ;
  assign y3526 = ~n20984 ;
  assign y3527 = n20993 ;
  assign y3528 = n21000 ;
  assign y3529 = n21001 ;
  assign y3530 = ~n21003 ;
  assign y3531 = n21014 ;
  assign y3532 = ~n21015 ;
  assign y3533 = n21033 ;
  assign y3534 = ~n21038 ;
  assign y3535 = n21041 ;
  assign y3536 = ~n21043 ;
  assign y3537 = ~n21046 ;
  assign y3538 = ~n21051 ;
  assign y3539 = n21054 ;
  assign y3540 = ~n21057 ;
  assign y3541 = n21058 ;
  assign y3542 = n21060 ;
  assign y3543 = n21064 ;
  assign y3544 = n21068 ;
  assign y3545 = n21075 ;
  assign y3546 = n21081 ;
  assign y3547 = n21084 ;
  assign y3548 = ~1'b0 ;
  assign y3549 = n21086 ;
  assign y3550 = n21090 ;
  assign y3551 = ~n21094 ;
  assign y3552 = ~n21102 ;
  assign y3553 = ~n21109 ;
  assign y3554 = n21121 ;
  assign y3555 = ~n21124 ;
  assign y3556 = n21137 ;
  assign y3557 = ~n21141 ;
  assign y3558 = n21147 ;
  assign y3559 = ~n21155 ;
  assign y3560 = n21157 ;
  assign y3561 = ~n21161 ;
  assign y3562 = ~n21165 ;
  assign y3563 = n21173 ;
  assign y3564 = ~n21174 ;
  assign y3565 = n21186 ;
  assign y3566 = ~n21188 ;
  assign y3567 = ~n21189 ;
  assign y3568 = ~n21197 ;
  assign y3569 = ~1'b0 ;
  assign y3570 = ~n21201 ;
  assign y3571 = ~n21203 ;
  assign y3572 = ~n21204 ;
  assign y3573 = ~1'b0 ;
  assign y3574 = ~n21205 ;
  assign y3575 = ~n21211 ;
  assign y3576 = n21216 ;
  assign y3577 = ~n21217 ;
  assign y3578 = n21229 ;
  assign y3579 = n21233 ;
  assign y3580 = ~n21235 ;
  assign y3581 = ~n21237 ;
  assign y3582 = n21259 ;
  assign y3583 = ~n21261 ;
  assign y3584 = ~n21263 ;
  assign y3585 = n21268 ;
  assign y3586 = ~n21290 ;
  assign y3587 = ~n21294 ;
  assign y3588 = ~n21295 ;
  assign y3589 = n21302 ;
  assign y3590 = ~n21304 ;
  assign y3591 = n21305 ;
  assign y3592 = ~n21306 ;
  assign y3593 = n21311 ;
  assign y3594 = ~n21318 ;
  assign y3595 = ~n21323 ;
  assign y3596 = ~n21331 ;
  assign y3597 = n21342 ;
  assign y3598 = n21344 ;
  assign y3599 = ~n21347 ;
  assign y3600 = n21350 ;
  assign y3601 = ~n21352 ;
  assign y3602 = ~n21358 ;
  assign y3603 = n21369 ;
  assign y3604 = n21372 ;
  assign y3605 = ~1'b0 ;
  assign y3606 = n21376 ;
  assign y3607 = n21378 ;
  assign y3608 = ~n21385 ;
  assign y3609 = n21387 ;
  assign y3610 = n21397 ;
  assign y3611 = ~n21400 ;
  assign y3612 = n21401 ;
  assign y3613 = n21406 ;
  assign y3614 = ~n21414 ;
  assign y3615 = n21417 ;
  assign y3616 = ~n21418 ;
  assign y3617 = ~n21420 ;
  assign y3618 = ~n21425 ;
  assign y3619 = ~n21426 ;
  assign y3620 = n21429 ;
  assign y3621 = n21435 ;
  assign y3622 = ~n21439 ;
  assign y3623 = n21443 ;
  assign y3624 = ~n21453 ;
  assign y3625 = ~n21455 ;
  assign y3626 = ~n21459 ;
  assign y3627 = ~n21461 ;
  assign y3628 = n21462 ;
  assign y3629 = n21464 ;
  assign y3630 = n21469 ;
  assign y3631 = ~n21473 ;
  assign y3632 = ~n21475 ;
  assign y3633 = ~n21476 ;
  assign y3634 = ~n21480 ;
  assign y3635 = n21481 ;
  assign y3636 = ~1'b0 ;
  assign y3637 = n21491 ;
  assign y3638 = ~n21492 ;
  assign y3639 = ~1'b0 ;
  assign y3640 = n21506 ;
  assign y3641 = n21509 ;
  assign y3642 = ~n21510 ;
  assign y3643 = ~n21512 ;
  assign y3644 = n21519 ;
  assign y3645 = n21520 ;
  assign y3646 = n21527 ;
  assign y3647 = ~n21528 ;
  assign y3648 = n21530 ;
  assign y3649 = ~n21532 ;
  assign y3650 = n21539 ;
  assign y3651 = n21544 ;
  assign y3652 = n21546 ;
  assign y3653 = ~n21549 ;
  assign y3654 = ~n21556 ;
  assign y3655 = ~n21561 ;
  assign y3656 = n21564 ;
  assign y3657 = ~n21569 ;
  assign y3658 = ~n21570 ;
  assign y3659 = ~n21581 ;
  assign y3660 = ~n21587 ;
  assign y3661 = ~n21596 ;
  assign y3662 = ~n21597 ;
  assign y3663 = ~n21601 ;
  assign y3664 = ~n21605 ;
  assign y3665 = ~n21609 ;
  assign y3666 = n21612 ;
  assign y3667 = ~n21615 ;
  assign y3668 = n21616 ;
  assign y3669 = n21627 ;
  assign y3670 = n21629 ;
  assign y3671 = n21644 ;
  assign y3672 = n21649 ;
  assign y3673 = ~n21654 ;
  assign y3674 = n21658 ;
  assign y3675 = n21671 ;
  assign y3676 = n21677 ;
  assign y3677 = n21683 ;
  assign y3678 = ~n21693 ;
  assign y3679 = ~n21694 ;
  assign y3680 = ~n21708 ;
  assign y3681 = n7038 ;
  assign y3682 = n21713 ;
  assign y3683 = n21716 ;
  assign y3684 = ~n21719 ;
  assign y3685 = n21723 ;
  assign y3686 = ~n21727 ;
  assign y3687 = n21737 ;
  assign y3688 = n21738 ;
  assign y3689 = n21739 ;
  assign y3690 = ~n21742 ;
  assign y3691 = ~n21745 ;
  assign y3692 = ~n21751 ;
  assign y3693 = n21756 ;
  assign y3694 = ~n21761 ;
  assign y3695 = n21763 ;
  assign y3696 = n21766 ;
  assign y3697 = ~n21767 ;
  assign y3698 = n21773 ;
  assign y3699 = ~n21779 ;
  assign y3700 = n21787 ;
  assign y3701 = n21798 ;
  assign y3702 = n21800 ;
  assign y3703 = n21807 ;
  assign y3704 = ~n21810 ;
  assign y3705 = n21813 ;
  assign y3706 = ~n21819 ;
  assign y3707 = ~1'b0 ;
  assign y3708 = n21825 ;
  assign y3709 = ~n21828 ;
  assign y3710 = n21830 ;
  assign y3711 = n21831 ;
  assign y3712 = n21832 ;
  assign y3713 = n21835 ;
  assign y3714 = ~n21836 ;
  assign y3715 = ~n21838 ;
  assign y3716 = ~n21840 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = n21841 ;
  assign y3719 = n21843 ;
  assign y3720 = ~n21848 ;
  assign y3721 = ~n21849 ;
  assign y3722 = n21855 ;
  assign y3723 = n21858 ;
  assign y3724 = n21865 ;
  assign y3725 = ~n21866 ;
  assign y3726 = ~n21868 ;
  assign y3727 = ~n21869 ;
  assign y3728 = ~n21876 ;
  assign y3729 = ~n21879 ;
  assign y3730 = ~n21882 ;
  assign y3731 = ~n21884 ;
  assign y3732 = ~n21889 ;
  assign y3733 = n21891 ;
  assign y3734 = n21895 ;
  assign y3735 = n21900 ;
  assign y3736 = n21903 ;
  assign y3737 = n21904 ;
  assign y3738 = ~n21911 ;
  assign y3739 = ~n21914 ;
  assign y3740 = ~n21915 ;
  assign y3741 = ~n21924 ;
  assign y3742 = ~n21926 ;
  assign y3743 = n21930 ;
  assign y3744 = ~n21935 ;
  assign y3745 = n21940 ;
  assign y3746 = ~n21945 ;
  assign y3747 = ~n21947 ;
  assign y3748 = n21948 ;
  assign y3749 = n21955 ;
  assign y3750 = ~1'b0 ;
  assign y3751 = ~1'b0 ;
  assign y3752 = ~n21956 ;
  assign y3753 = ~n21962 ;
  assign y3754 = ~n21969 ;
  assign y3755 = ~n21971 ;
  assign y3756 = ~n21975 ;
  assign y3757 = n21976 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = ~n21977 ;
  assign y3760 = n21982 ;
  assign y3761 = n21987 ;
  assign y3762 = n21988 ;
  assign y3763 = n21989 ;
  assign y3764 = ~n21991 ;
  assign y3765 = n21995 ;
  assign y3766 = ~n21998 ;
  assign y3767 = ~n21999 ;
  assign y3768 = n22003 ;
  assign y3769 = n22016 ;
  assign y3770 = ~n22021 ;
  assign y3771 = n22025 ;
  assign y3772 = ~n22032 ;
  assign y3773 = ~n22041 ;
  assign y3774 = n22044 ;
  assign y3775 = ~n22049 ;
  assign y3776 = n22050 ;
  assign y3777 = n22054 ;
  assign y3778 = ~n22058 ;
  assign y3779 = n22060 ;
  assign y3780 = n22062 ;
  assign y3781 = ~n22067 ;
  assign y3782 = n22079 ;
  assign y3783 = ~n22089 ;
  assign y3784 = ~n22093 ;
  assign y3785 = ~n22094 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = n22099 ;
  assign y3788 = ~n22100 ;
  assign y3789 = ~n22105 ;
  assign y3790 = n22108 ;
  assign y3791 = ~n22111 ;
  assign y3792 = n22113 ;
  assign y3793 = n22115 ;
  assign y3794 = ~n22123 ;
  assign y3795 = ~n22126 ;
  assign y3796 = n22134 ;
  assign y3797 = n22141 ;
  assign y3798 = ~n22144 ;
  assign y3799 = ~n22150 ;
  assign y3800 = n22159 ;
  assign y3801 = n22169 ;
  assign y3802 = ~n22177 ;
  assign y3803 = ~n22182 ;
  assign y3804 = n22187 ;
  assign y3805 = ~n22193 ;
  assign y3806 = n22199 ;
  assign y3807 = ~n22203 ;
  assign y3808 = n22206 ;
  assign y3809 = ~n22212 ;
  assign y3810 = ~1'b0 ;
  assign y3811 = n22213 ;
  assign y3812 = ~n22216 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = ~1'b0 ;
  assign y3815 = n22223 ;
  assign y3816 = ~n22227 ;
  assign y3817 = ~n22229 ;
  assign y3818 = n22231 ;
  assign y3819 = n22241 ;
  assign y3820 = n22258 ;
  assign y3821 = ~1'b0 ;
  assign y3822 = n22259 ;
  assign y3823 = ~n22266 ;
  assign y3824 = n22270 ;
  assign y3825 = ~n22272 ;
  assign y3826 = n22277 ;
  assign y3827 = ~n22280 ;
  assign y3828 = n22284 ;
  assign y3829 = ~n22287 ;
  assign y3830 = ~n22289 ;
  assign y3831 = ~n22291 ;
  assign y3832 = n22295 ;
  assign y3833 = ~1'b0 ;
  assign y3834 = n22298 ;
  assign y3835 = n22304 ;
  assign y3836 = n22309 ;
  assign y3837 = n22314 ;
  assign y3838 = ~n22315 ;
  assign y3839 = ~n22321 ;
  assign y3840 = ~n22325 ;
  assign y3841 = n22326 ;
  assign y3842 = ~n22327 ;
  assign y3843 = n22331 ;
  assign y3844 = ~n22333 ;
  assign y3845 = ~n22335 ;
  assign y3846 = ~n22341 ;
  assign y3847 = ~n22344 ;
  assign y3848 = n22351 ;
  assign y3849 = ~n22353 ;
  assign y3850 = ~n22354 ;
  assign y3851 = ~n22356 ;
  assign y3852 = ~n22364 ;
  assign y3853 = n22367 ;
  assign y3854 = ~n22370 ;
  assign y3855 = ~1'b0 ;
  assign y3856 = n22371 ;
  assign y3857 = ~n22376 ;
  assign y3858 = n22379 ;
  assign y3859 = n22381 ;
  assign y3860 = ~n22382 ;
  assign y3861 = ~n22385 ;
  assign y3862 = n22396 ;
  assign y3863 = ~n22403 ;
  assign y3864 = ~n22409 ;
  assign y3865 = ~n22420 ;
  assign y3866 = ~n22421 ;
  assign y3867 = n22428 ;
  assign y3868 = n22437 ;
  assign y3869 = n22438 ;
  assign y3870 = ~n22440 ;
  assign y3871 = n22441 ;
  assign y3872 = ~n22442 ;
  assign y3873 = ~n22444 ;
  assign y3874 = n22448 ;
  assign y3875 = ~1'b0 ;
  assign y3876 = ~n22450 ;
  assign y3877 = n22455 ;
  assign y3878 = ~1'b0 ;
  assign y3879 = ~n22470 ;
  assign y3880 = ~n22475 ;
  assign y3881 = n22478 ;
  assign y3882 = ~n22483 ;
  assign y3883 = ~n22487 ;
  assign y3884 = ~n22489 ;
  assign y3885 = ~n22499 ;
  assign y3886 = ~n22501 ;
  assign y3887 = ~n22507 ;
  assign y3888 = n22508 ;
  assign y3889 = n22513 ;
  assign y3890 = n22518 ;
  assign y3891 = ~n22520 ;
  assign y3892 = ~n22523 ;
  assign y3893 = ~n22526 ;
  assign y3894 = n22527 ;
  assign y3895 = ~1'b0 ;
  assign y3896 = n22540 ;
  assign y3897 = n22543 ;
  assign y3898 = ~n22545 ;
  assign y3899 = ~n22552 ;
  assign y3900 = ~n22553 ;
  assign y3901 = n22558 ;
  assign y3902 = n22570 ;
  assign y3903 = n22579 ;
  assign y3904 = n22589 ;
  assign y3905 = ~1'b0 ;
  assign y3906 = ~n22592 ;
  assign y3907 = n22594 ;
  assign y3908 = ~n22595 ;
  assign y3909 = n22607 ;
  assign y3910 = ~n22608 ;
  assign y3911 = ~n22610 ;
  assign y3912 = n22614 ;
  assign y3913 = n22623 ;
  assign y3914 = n22624 ;
  assign y3915 = ~n22635 ;
  assign y3916 = ~n22639 ;
  assign y3917 = ~n22642 ;
  assign y3918 = n22648 ;
  assign y3919 = n22650 ;
  assign y3920 = n22660 ;
  assign y3921 = n22663 ;
  assign y3922 = n22674 ;
  assign y3923 = ~n22675 ;
  assign y3924 = ~n22687 ;
  assign y3925 = n22704 ;
  assign y3926 = ~n22705 ;
  assign y3927 = n22707 ;
  assign y3928 = ~n22709 ;
  assign y3929 = n22711 ;
  assign y3930 = n22712 ;
  assign y3931 = n22716 ;
  assign y3932 = n22726 ;
  assign y3933 = n22733 ;
  assign y3934 = n22735 ;
  assign y3935 = n22737 ;
  assign y3936 = ~n22738 ;
  assign y3937 = ~n22744 ;
  assign y3938 = ~n22745 ;
  assign y3939 = n22747 ;
  assign y3940 = ~n22748 ;
  assign y3941 = ~n22751 ;
  assign y3942 = ~n22759 ;
  assign y3943 = ~n22760 ;
  assign y3944 = ~n22763 ;
  assign y3945 = n22765 ;
  assign y3946 = ~n22767 ;
  assign y3947 = ~n22771 ;
  assign y3948 = n22775 ;
  assign y3949 = n22776 ;
  assign y3950 = ~n22778 ;
  assign y3951 = n22782 ;
  assign y3952 = ~n22784 ;
  assign y3953 = n22787 ;
  assign y3954 = ~n22793 ;
  assign y3955 = n22795 ;
  assign y3956 = n22804 ;
  assign y3957 = n22807 ;
  assign y3958 = ~n22810 ;
  assign y3959 = ~n22811 ;
  assign y3960 = n22815 ;
  assign y3961 = n22820 ;
  assign y3962 = ~n22821 ;
  assign y3963 = n22823 ;
  assign y3964 = n22825 ;
  assign y3965 = n22829 ;
  assign y3966 = ~n22833 ;
  assign y3967 = ~n22836 ;
  assign y3968 = ~n22839 ;
  assign y3969 = n22843 ;
  assign y3970 = n22845 ;
  assign y3971 = ~n22848 ;
  assign y3972 = n22853 ;
  assign y3973 = n22854 ;
  assign y3974 = ~n22855 ;
  assign y3975 = ~n22857 ;
  assign y3976 = n22865 ;
  assign y3977 = n22872 ;
  assign y3978 = ~n22873 ;
  assign y3979 = ~n22878 ;
  assign y3980 = ~n22879 ;
  assign y3981 = ~n22882 ;
  assign y3982 = n22889 ;
  assign y3983 = n22890 ;
  assign y3984 = ~n22892 ;
  assign y3985 = ~n22893 ;
  assign y3986 = ~n22894 ;
  assign y3987 = ~n22897 ;
  assign y3988 = n22905 ;
  assign y3989 = n22906 ;
  assign y3990 = n22913 ;
  assign y3991 = ~n22916 ;
  assign y3992 = n22922 ;
  assign y3993 = n22923 ;
  assign y3994 = ~n22925 ;
  assign y3995 = n22926 ;
  assign y3996 = n22934 ;
  assign y3997 = ~n22938 ;
  assign y3998 = ~n22944 ;
  assign y3999 = n22946 ;
  assign y4000 = ~n22947 ;
  assign y4001 = n22948 ;
  assign y4002 = n22949 ;
  assign y4003 = n22958 ;
  assign y4004 = ~n22959 ;
  assign y4005 = ~n22962 ;
  assign y4006 = ~n22970 ;
  assign y4007 = n22976 ;
  assign y4008 = ~n22982 ;
  assign y4009 = ~n22984 ;
  assign y4010 = ~n22990 ;
  assign y4011 = ~n22995 ;
  assign y4012 = ~n23008 ;
  assign y4013 = ~n23011 ;
  assign y4014 = n23012 ;
  assign y4015 = n23013 ;
  assign y4016 = ~n23015 ;
  assign y4017 = n23025 ;
  assign y4018 = n23027 ;
  assign y4019 = n23029 ;
  assign y4020 = n23034 ;
  assign y4021 = n23036 ;
  assign y4022 = n23038 ;
  assign y4023 = n23041 ;
  assign y4024 = ~n23050 ;
  assign y4025 = ~n23063 ;
  assign y4026 = n23067 ;
  assign y4027 = ~n23072 ;
  assign y4028 = n23094 ;
  assign y4029 = n23095 ;
  assign y4030 = n23098 ;
  assign y4031 = ~n23104 ;
  assign y4032 = ~n23110 ;
  assign y4033 = n23111 ;
  assign y4034 = ~n23114 ;
  assign y4035 = ~n23116 ;
  assign y4036 = n23119 ;
  assign y4037 = ~n23120 ;
  assign y4038 = n23123 ;
  assign y4039 = n23131 ;
  assign y4040 = ~n23136 ;
  assign y4041 = ~n23141 ;
  assign y4042 = n23142 ;
  assign y4043 = ~n23146 ;
  assign y4044 = n23147 ;
  assign y4045 = n23148 ;
  assign y4046 = n23150 ;
  assign y4047 = n23151 ;
  assign y4048 = ~n23152 ;
  assign y4049 = ~n23155 ;
  assign y4050 = ~n23157 ;
  assign y4051 = ~n23158 ;
  assign y4052 = ~n23162 ;
  assign y4053 = n23165 ;
  assign y4054 = n23171 ;
  assign y4055 = n23193 ;
  assign y4056 = n23199 ;
  assign y4057 = ~n23205 ;
  assign y4058 = n23208 ;
  assign y4059 = ~n23210 ;
  assign y4060 = ~n23211 ;
  assign y4061 = n23217 ;
  assign y4062 = ~n23221 ;
  assign y4063 = ~1'b0 ;
  assign y4064 = n23229 ;
  assign y4065 = ~n23233 ;
  assign y4066 = ~n23235 ;
  assign y4067 = ~n23241 ;
  assign y4068 = n23246 ;
  assign y4069 = n23247 ;
  assign y4070 = n23252 ;
  assign y4071 = ~n23256 ;
  assign y4072 = ~n23260 ;
  assign y4073 = ~n23261 ;
  assign y4074 = n23262 ;
  assign y4075 = ~n23266 ;
  assign y4076 = ~n23272 ;
  assign y4077 = ~n23275 ;
  assign y4078 = ~n23278 ;
  assign y4079 = n23281 ;
  assign y4080 = n23289 ;
  assign y4081 = n23290 ;
  assign y4082 = ~n23298 ;
  assign y4083 = n23303 ;
  assign y4084 = ~n23306 ;
  assign y4085 = n23308 ;
  assign y4086 = n23311 ;
  assign y4087 = n23322 ;
  assign y4088 = ~n23331 ;
  assign y4089 = ~n23332 ;
  assign y4090 = ~n23335 ;
  assign y4091 = ~n23336 ;
  assign y4092 = n23338 ;
  assign y4093 = n23346 ;
  assign y4094 = ~1'b0 ;
  assign y4095 = ~n23352 ;
  assign y4096 = n23359 ;
  assign y4097 = n23363 ;
  assign y4098 = n23367 ;
  assign y4099 = ~n23373 ;
  assign y4100 = n23375 ;
  assign y4101 = n23382 ;
  assign y4102 = ~n23386 ;
  assign y4103 = n23392 ;
  assign y4104 = ~n23397 ;
  assign y4105 = ~1'b0 ;
  assign y4106 = n23398 ;
  assign y4107 = n23400 ;
  assign y4108 = ~n23402 ;
  assign y4109 = ~n23408 ;
  assign y4110 = ~n23415 ;
  assign y4111 = n23421 ;
  assign y4112 = n23422 ;
  assign y4113 = ~1'b0 ;
  assign y4114 = ~n23424 ;
  assign y4115 = n23432 ;
  assign y4116 = n23434 ;
  assign y4117 = ~n23435 ;
  assign y4118 = ~n23438 ;
  assign y4119 = ~n23440 ;
  assign y4120 = ~1'b0 ;
  assign y4121 = ~n23448 ;
  assign y4122 = ~n23450 ;
  assign y4123 = n23461 ;
  assign y4124 = n23471 ;
  assign y4125 = n23472 ;
  assign y4126 = ~n23493 ;
  assign y4127 = ~n23495 ;
  assign y4128 = n23496 ;
  assign y4129 = ~n23501 ;
  assign y4130 = ~n23510 ;
  assign y4131 = ~n23513 ;
  assign y4132 = ~1'b0 ;
  assign y4133 = n23515 ;
  assign y4134 = ~n23530 ;
  assign y4135 = n23531 ;
  assign y4136 = n23532 ;
  assign y4137 = ~n23535 ;
  assign y4138 = ~n23539 ;
  assign y4139 = ~n23541 ;
  assign y4140 = ~n23543 ;
  assign y4141 = n23545 ;
  assign y4142 = n23551 ;
  assign y4143 = ~1'b0 ;
  assign y4144 = n23561 ;
  assign y4145 = n23570 ;
  assign y4146 = ~n23573 ;
  assign y4147 = n23577 ;
  assign y4148 = n23582 ;
  assign y4149 = ~n23584 ;
  assign y4150 = ~n23591 ;
  assign y4151 = ~n23593 ;
  assign y4152 = n23595 ;
  assign y4153 = n23596 ;
  assign y4154 = ~n23599 ;
  assign y4155 = n23600 ;
  assign y4156 = ~n23602 ;
  assign y4157 = n23603 ;
  assign y4158 = ~n23607 ;
  assign y4159 = n23609 ;
  assign y4160 = ~n23613 ;
  assign y4161 = n23618 ;
  assign y4162 = ~n23621 ;
  assign y4163 = ~n23622 ;
  assign y4164 = ~n23625 ;
  assign y4165 = n23628 ;
  assign y4166 = ~n23629 ;
  assign y4167 = n23630 ;
  assign y4168 = n23632 ;
  assign y4169 = ~1'b0 ;
  assign y4170 = n23638 ;
  assign y4171 = n23640 ;
  assign y4172 = n23648 ;
  assign y4173 = ~n23664 ;
  assign y4174 = ~n23666 ;
  assign y4175 = ~n23667 ;
  assign y4176 = n23673 ;
  assign y4177 = n23675 ;
  assign y4178 = ~n23677 ;
  assign y4179 = ~n23679 ;
  assign y4180 = ~n23688 ;
  assign y4181 = n23693 ;
  assign y4182 = ~n23695 ;
  assign y4183 = ~n23698 ;
  assign y4184 = ~n23705 ;
  assign y4185 = ~n23710 ;
  assign y4186 = ~n23716 ;
  assign y4187 = n23726 ;
  assign y4188 = ~n23728 ;
  assign y4189 = n23732 ;
  assign y4190 = ~n23733 ;
  assign y4191 = n23736 ;
  assign y4192 = n23739 ;
  assign y4193 = n23743 ;
  assign y4194 = n23744 ;
  assign y4195 = ~n23745 ;
  assign y4196 = ~n23746 ;
  assign y4197 = ~n23751 ;
  assign y4198 = n23754 ;
  assign y4199 = n23755 ;
  assign y4200 = ~n23763 ;
  assign y4201 = ~n23768 ;
  assign y4202 = n23769 ;
  assign y4203 = n23787 ;
  assign y4204 = n23790 ;
  assign y4205 = ~n23792 ;
  assign y4206 = ~n23796 ;
  assign y4207 = n23798 ;
  assign y4208 = ~n23806 ;
  assign y4209 = n23808 ;
  assign y4210 = n23812 ;
  assign y4211 = n23819 ;
  assign y4212 = n23822 ;
  assign y4213 = ~n23827 ;
  assign y4214 = n23828 ;
  assign y4215 = n23830 ;
  assign y4216 = n23836 ;
  assign y4217 = ~n23838 ;
  assign y4218 = n23848 ;
  assign y4219 = ~1'b0 ;
  assign y4220 = ~1'b0 ;
  assign y4221 = ~n23849 ;
  assign y4222 = n23852 ;
  assign y4223 = ~n23858 ;
  assign y4224 = ~n23861 ;
  assign y4225 = ~n23868 ;
  assign y4226 = ~n23871 ;
  assign y4227 = ~n23889 ;
  assign y4228 = ~n23891 ;
  assign y4229 = n23892 ;
  assign y4230 = n23895 ;
  assign y4231 = ~n23904 ;
  assign y4232 = ~n23906 ;
  assign y4233 = ~n23907 ;
  assign y4234 = ~n23917 ;
  assign y4235 = ~n23920 ;
  assign y4236 = ~n23925 ;
  assign y4237 = ~n23928 ;
  assign y4238 = ~n23935 ;
  assign y4239 = n23937 ;
  assign y4240 = ~n23939 ;
  assign y4241 = ~n23941 ;
  assign y4242 = n23943 ;
  assign y4243 = ~n23945 ;
  assign y4244 = n23946 ;
  assign y4245 = n23947 ;
  assign y4246 = n23950 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = n23954 ;
  assign y4249 = ~n23956 ;
  assign y4250 = ~n23961 ;
  assign y4251 = n23973 ;
  assign y4252 = ~n23979 ;
  assign y4253 = n23980 ;
  assign y4254 = ~n23987 ;
  assign y4255 = n23988 ;
  assign y4256 = n23993 ;
  assign y4257 = ~n24001 ;
  assign y4258 = ~n24007 ;
  assign y4259 = ~n24010 ;
  assign y4260 = ~n24014 ;
  assign y4261 = ~n24023 ;
  assign y4262 = n24025 ;
  assign y4263 = ~n24027 ;
  assign y4264 = n24029 ;
  assign y4265 = n24037 ;
  assign y4266 = n24044 ;
  assign y4267 = n24049 ;
  assign y4268 = ~1'b0 ;
  assign y4269 = ~n24051 ;
  assign y4270 = n24053 ;
  assign y4271 = ~n24054 ;
  assign y4272 = ~n24055 ;
  assign y4273 = ~n24059 ;
  assign y4274 = ~n24064 ;
  assign y4275 = ~n24065 ;
  assign y4276 = n24069 ;
  assign y4277 = ~n24071 ;
  assign y4278 = n24073 ;
  assign y4279 = n24075 ;
  assign y4280 = n24076 ;
  assign y4281 = n24079 ;
  assign y4282 = n24084 ;
  assign y4283 = ~n24085 ;
  assign y4284 = ~1'b0 ;
  assign y4285 = ~n24088 ;
  assign y4286 = n24096 ;
  assign y4287 = n24097 ;
  assign y4288 = ~n24103 ;
  assign y4289 = ~n24106 ;
  assign y4290 = ~n24107 ;
  assign y4291 = ~n24112 ;
  assign y4292 = ~n24113 ;
  assign y4293 = ~n24121 ;
  assign y4294 = ~n24129 ;
  assign y4295 = n24136 ;
  assign y4296 = ~n24138 ;
  assign y4297 = ~n24157 ;
  assign y4298 = ~n24161 ;
  assign y4299 = ~n24164 ;
  assign y4300 = ~n24175 ;
  assign y4301 = n24186 ;
  assign y4302 = ~n24187 ;
  assign y4303 = n24188 ;
  assign y4304 = n24191 ;
  assign y4305 = ~n24198 ;
  assign y4306 = ~n24201 ;
  assign y4307 = n24204 ;
  assign y4308 = n24207 ;
  assign y4309 = n24208 ;
  assign y4310 = ~n24209 ;
  assign y4311 = ~n24210 ;
  assign y4312 = ~n24218 ;
  assign y4313 = n24230 ;
  assign y4314 = n24231 ;
  assign y4315 = ~n24233 ;
  assign y4316 = ~n24237 ;
  assign y4317 = n24238 ;
  assign y4318 = ~n24243 ;
  assign y4319 = n24245 ;
  assign y4320 = n24249 ;
  assign y4321 = n24255 ;
  assign y4322 = n24258 ;
  assign y4323 = ~n24259 ;
  assign y4324 = ~n24265 ;
  assign y4325 = ~n24267 ;
  assign y4326 = n24268 ;
  assign y4327 = n24274 ;
  assign y4328 = ~n24279 ;
  assign y4329 = ~n24281 ;
  assign y4330 = ~n24283 ;
  assign y4331 = ~1'b0 ;
  assign y4332 = ~n24287 ;
  assign y4333 = n24289 ;
  assign y4334 = n24290 ;
  assign y4335 = n24292 ;
  assign y4336 = ~1'b0 ;
  assign y4337 = n24294 ;
  assign y4338 = ~n24297 ;
  assign y4339 = n24302 ;
  assign y4340 = n24304 ;
  assign y4341 = ~n24305 ;
  assign y4342 = n24308 ;
  assign y4343 = n24310 ;
  assign y4344 = ~n24314 ;
  assign y4345 = ~n24322 ;
  assign y4346 = n24326 ;
  assign y4347 = n24333 ;
  assign y4348 = n24336 ;
  assign y4349 = ~1'b0 ;
  assign y4350 = ~n24339 ;
  assign y4351 = n24345 ;
  assign y4352 = ~n24351 ;
  assign y4353 = ~n24361 ;
  assign y4354 = n24362 ;
  assign y4355 = n24375 ;
  assign y4356 = n24376 ;
  assign y4357 = ~n24377 ;
  assign y4358 = n24381 ;
  assign y4359 = ~n24385 ;
  assign y4360 = n24387 ;
  assign y4361 = n24398 ;
  assign y4362 = ~n24399 ;
  assign y4363 = n24401 ;
  assign y4364 = n24402 ;
  assign y4365 = n24412 ;
  assign y4366 = n24413 ;
  assign y4367 = n24417 ;
  assign y4368 = n24421 ;
  assign y4369 = ~n24428 ;
  assign y4370 = ~n24433 ;
  assign y4371 = ~n24437 ;
  assign y4372 = ~n24440 ;
  assign y4373 = ~n24444 ;
  assign y4374 = n24449 ;
  assign y4375 = n24451 ;
  assign y4376 = ~n24453 ;
  assign y4377 = n24464 ;
  assign y4378 = ~n24471 ;
  assign y4379 = n24477 ;
  assign y4380 = n24479 ;
  assign y4381 = n24480 ;
  assign y4382 = ~n24481 ;
  assign y4383 = n24483 ;
  assign y4384 = ~n24486 ;
  assign y4385 = ~n24491 ;
  assign y4386 = ~n24505 ;
  assign y4387 = ~n24509 ;
  assign y4388 = ~n24510 ;
  assign y4389 = ~n24512 ;
  assign y4390 = ~n24518 ;
  assign y4391 = n24529 ;
  assign y4392 = ~n24530 ;
  assign y4393 = n24542 ;
  assign y4394 = ~n24545 ;
  assign y4395 = n24552 ;
  assign y4396 = n24564 ;
  assign y4397 = n24578 ;
  assign y4398 = n24583 ;
  assign y4399 = ~n24595 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = ~n24597 ;
  assign y4402 = ~n24598 ;
  assign y4403 = ~n24599 ;
  assign y4404 = ~n24607 ;
  assign y4405 = n24608 ;
  assign y4406 = n24614 ;
  assign y4407 = ~n24617 ;
  assign y4408 = ~n24618 ;
  assign y4409 = ~n24619 ;
  assign y4410 = n24621 ;
  assign y4411 = ~n24623 ;
  assign y4412 = n24630 ;
  assign y4413 = ~n24632 ;
  assign y4414 = n24638 ;
  assign y4415 = ~n24639 ;
  assign y4416 = ~n24644 ;
  assign y4417 = ~n24646 ;
  assign y4418 = ~n24648 ;
  assign y4419 = n24656 ;
  assign y4420 = n24662 ;
  assign y4421 = ~n24664 ;
  assign y4422 = ~n24669 ;
  assign y4423 = ~n24670 ;
  assign y4424 = ~n24683 ;
  assign y4425 = n24685 ;
  assign y4426 = ~n24686 ;
  assign y4427 = ~n24689 ;
  assign y4428 = ~n24690 ;
  assign y4429 = ~n24692 ;
  assign y4430 = ~n24695 ;
  assign y4431 = ~n24703 ;
  assign y4432 = ~1'b0 ;
  assign y4433 = ~n24716 ;
  assign y4434 = n24719 ;
  assign y4435 = n24724 ;
  assign y4436 = n24729 ;
  assign y4437 = ~n24737 ;
  assign y4438 = ~n24741 ;
  assign y4439 = n24747 ;
  assign y4440 = ~n24750 ;
  assign y4441 = n24755 ;
  assign y4442 = n24757 ;
  assign y4443 = n24761 ;
  assign y4444 = n24763 ;
  assign y4445 = ~1'b0 ;
  assign y4446 = ~n24770 ;
  assign y4447 = n24774 ;
  assign y4448 = ~n24780 ;
  assign y4449 = ~n24786 ;
  assign y4450 = ~n24787 ;
  assign y4451 = n24788 ;
  assign y4452 = n24795 ;
  assign y4453 = n24802 ;
  assign y4454 = ~n24805 ;
  assign y4455 = ~n24806 ;
  assign y4456 = n24808 ;
  assign y4457 = n24811 ;
  assign y4458 = ~n24813 ;
  assign y4459 = n24822 ;
  assign y4460 = n24824 ;
  assign y4461 = n24825 ;
  assign y4462 = n24831 ;
  assign y4463 = ~n24836 ;
  assign y4464 = n24838 ;
  assign y4465 = n24841 ;
  assign y4466 = ~n24842 ;
  assign y4467 = ~n24846 ;
  assign y4468 = n24855 ;
  assign y4469 = ~n24859 ;
  assign y4470 = n24863 ;
  assign y4471 = ~n24866 ;
  assign y4472 = n24870 ;
  assign y4473 = ~n24874 ;
  assign y4474 = n24875 ;
  assign y4475 = ~n24877 ;
  assign y4476 = n24879 ;
  assign y4477 = ~n24883 ;
  assign y4478 = n24886 ;
  assign y4479 = ~n24889 ;
  assign y4480 = ~n24890 ;
  assign y4481 = ~n24894 ;
  assign y4482 = ~n24896 ;
  assign y4483 = ~n24900 ;
  assign y4484 = ~n24901 ;
  assign y4485 = ~n24902 ;
  assign y4486 = ~n24903 ;
  assign y4487 = ~n24905 ;
  assign y4488 = n24906 ;
  assign y4489 = ~n24909 ;
  assign y4490 = ~n24914 ;
  assign y4491 = n24917 ;
  assign y4492 = ~n24918 ;
  assign y4493 = n24923 ;
  assign y4494 = n24925 ;
  assign y4495 = ~n24927 ;
  assign y4496 = ~n24930 ;
  assign y4497 = ~n24935 ;
  assign y4498 = n24938 ;
  assign y4499 = n24940 ;
  assign y4500 = n24941 ;
  assign y4501 = n24942 ;
  assign y4502 = ~1'b0 ;
  assign y4503 = ~n24946 ;
  assign y4504 = n24949 ;
  assign y4505 = ~n24962 ;
  assign y4506 = n24968 ;
  assign y4507 = ~n24970 ;
  assign y4508 = n24971 ;
  assign y4509 = ~n24974 ;
  assign y4510 = ~n24977 ;
  assign y4511 = ~n24980 ;
  assign y4512 = ~n24989 ;
  assign y4513 = n24992 ;
  assign y4514 = ~n24995 ;
  assign y4515 = ~n24997 ;
  assign y4516 = n25000 ;
  assign y4517 = ~n25009 ;
  assign y4518 = n25012 ;
  assign y4519 = ~n25013 ;
  assign y4520 = n25019 ;
  assign y4521 = n25027 ;
  assign y4522 = ~n25029 ;
  assign y4523 = n25033 ;
  assign y4524 = ~n25035 ;
  assign y4525 = ~n25036 ;
  assign y4526 = ~n25047 ;
  assign y4527 = n25051 ;
  assign y4528 = ~1'b0 ;
  assign y4529 = ~n25052 ;
  assign y4530 = ~n25060 ;
  assign y4531 = n25066 ;
  assign y4532 = ~n25068 ;
  assign y4533 = ~n25069 ;
  assign y4534 = ~n25070 ;
  assign y4535 = n25071 ;
  assign y4536 = n25073 ;
  assign y4537 = ~n25074 ;
  assign y4538 = n25075 ;
  assign y4539 = ~n25080 ;
  assign y4540 = n25084 ;
  assign y4541 = n25086 ;
  assign y4542 = ~1'b0 ;
  assign y4543 = n25093 ;
  assign y4544 = ~n25098 ;
  assign y4545 = ~n25100 ;
  assign y4546 = n25104 ;
  assign y4547 = ~n25107 ;
  assign y4548 = ~n25112 ;
  assign y4549 = n25115 ;
  assign y4550 = n25117 ;
  assign y4551 = n25118 ;
  assign y4552 = ~n25121 ;
  assign y4553 = n25122 ;
  assign y4554 = ~n25126 ;
  assign y4555 = n25133 ;
  assign y4556 = n25139 ;
  assign y4557 = n25144 ;
  assign y4558 = n25147 ;
  assign y4559 = n25159 ;
  assign y4560 = n25163 ;
  assign y4561 = ~n25168 ;
  assign y4562 = ~n25172 ;
  assign y4563 = n25178 ;
  assign y4564 = ~1'b0 ;
  assign y4565 = ~n25183 ;
  assign y4566 = ~n25185 ;
  assign y4567 = ~n25187 ;
  assign y4568 = ~n25190 ;
  assign y4569 = ~n25197 ;
  assign y4570 = ~n25211 ;
  assign y4571 = ~n25218 ;
  assign y4572 = ~n25221 ;
  assign y4573 = n25227 ;
  assign y4574 = n25240 ;
  assign y4575 = n25241 ;
  assign y4576 = ~1'b0 ;
  assign y4577 = n25242 ;
  assign y4578 = n25246 ;
  assign y4579 = n25247 ;
  assign y4580 = ~n25250 ;
  assign y4581 = ~n25262 ;
  assign y4582 = ~1'b0 ;
  assign y4583 = ~n25264 ;
  assign y4584 = n25272 ;
  assign y4585 = ~n25276 ;
  assign y4586 = ~n25284 ;
  assign y4587 = ~n25286 ;
  assign y4588 = n25288 ;
  assign y4589 = n25291 ;
  assign y4590 = n25295 ;
  assign y4591 = ~n25297 ;
  assign y4592 = n25306 ;
  assign y4593 = n25307 ;
  assign y4594 = n25313 ;
  assign y4595 = n25315 ;
  assign y4596 = ~n25324 ;
  assign y4597 = n25329 ;
  assign y4598 = n25330 ;
  assign y4599 = n25336 ;
  assign y4600 = ~n25339 ;
  assign y4601 = n25341 ;
  assign y4602 = n25342 ;
  assign y4603 = n25345 ;
  assign y4604 = n25346 ;
  assign y4605 = ~n25348 ;
  assign y4606 = n25349 ;
  assign y4607 = n25354 ;
  assign y4608 = ~n25356 ;
  assign y4609 = ~n25363 ;
  assign y4610 = n25364 ;
  assign y4611 = ~n25369 ;
  assign y4612 = n25370 ;
  assign y4613 = n25374 ;
  assign y4614 = ~n25384 ;
  assign y4615 = ~n25391 ;
  assign y4616 = ~n25394 ;
  assign y4617 = n25396 ;
  assign y4618 = n25403 ;
  assign y4619 = ~n25406 ;
  assign y4620 = n25415 ;
  assign y4621 = n25422 ;
  assign y4622 = ~n25430 ;
  assign y4623 = n25435 ;
  assign y4624 = n25438 ;
  assign y4625 = n25439 ;
  assign y4626 = ~n25440 ;
  assign y4627 = ~n25441 ;
  assign y4628 = n25444 ;
  assign y4629 = n25447 ;
  assign y4630 = n25450 ;
  assign y4631 = ~n25463 ;
  assign y4632 = ~n25464 ;
  assign y4633 = n25470 ;
  assign y4634 = ~n25476 ;
  assign y4635 = ~n25478 ;
  assign y4636 = n25483 ;
  assign y4637 = n25485 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = ~n25489 ;
  assign y4640 = ~n25491 ;
  assign y4641 = n12861 ;
  assign y4642 = ~n25492 ;
  assign y4643 = ~n25493 ;
  assign y4644 = n25499 ;
  assign y4645 = n25504 ;
  assign y4646 = n25506 ;
  assign y4647 = n25507 ;
  assign y4648 = n25509 ;
  assign y4649 = ~n25511 ;
  assign y4650 = ~n25512 ;
  assign y4651 = ~n25519 ;
  assign y4652 = n25522 ;
  assign y4653 = ~n25525 ;
  assign y4654 = n25531 ;
  assign y4655 = ~n25538 ;
  assign y4656 = ~n25544 ;
  assign y4657 = n25545 ;
  assign y4658 = n25550 ;
  assign y4659 = ~n25551 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = n25556 ;
  assign y4662 = n25560 ;
  assign y4663 = ~n25564 ;
  assign y4664 = n25567 ;
  assign y4665 = ~n25577 ;
  assign y4666 = ~1'b0 ;
  assign y4667 = n25578 ;
  assign y4668 = n25582 ;
  assign y4669 = ~n25585 ;
  assign y4670 = ~n25586 ;
  assign y4671 = ~n25588 ;
  assign y4672 = n25595 ;
  assign y4673 = n25601 ;
  assign y4674 = ~n25606 ;
  assign y4675 = ~n25609 ;
  assign y4676 = ~n25613 ;
  assign y4677 = ~n25625 ;
  assign y4678 = n25627 ;
  assign y4679 = ~n25635 ;
  assign y4680 = n25641 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = ~n25643 ;
  assign y4683 = n25646 ;
  assign y4684 = n25649 ;
  assign y4685 = ~n25654 ;
  assign y4686 = n25657 ;
  assign y4687 = ~n25659 ;
  assign y4688 = n25660 ;
  assign y4689 = n25662 ;
  assign y4690 = ~n25675 ;
  assign y4691 = ~n25693 ;
  assign y4692 = n25697 ;
  assign y4693 = n25700 ;
  assign y4694 = n25702 ;
  assign y4695 = n25707 ;
  assign y4696 = ~n25718 ;
  assign y4697 = ~n25727 ;
  assign y4698 = n25737 ;
  assign y4699 = n25746 ;
  assign y4700 = n25751 ;
  assign y4701 = n25756 ;
  assign y4702 = n25757 ;
  assign y4703 = ~n25764 ;
  assign y4704 = ~n25765 ;
  assign y4705 = ~n25768 ;
  assign y4706 = ~n25769 ;
  assign y4707 = ~n25771 ;
  assign y4708 = n25773 ;
  assign y4709 = n25774 ;
  assign y4710 = n25784 ;
  assign y4711 = ~n25787 ;
  assign y4712 = ~1'b0 ;
  assign y4713 = ~n25789 ;
  assign y4714 = ~n25794 ;
  assign y4715 = n25797 ;
  assign y4716 = n25800 ;
  assign y4717 = ~1'b0 ;
  assign y4718 = ~1'b0 ;
  assign y4719 = ~n25805 ;
  assign y4720 = n25807 ;
  assign y4721 = n25808 ;
  assign y4722 = n25814 ;
  assign y4723 = ~n25819 ;
  assign y4724 = n25826 ;
  assign y4725 = ~n25827 ;
  assign y4726 = ~n25833 ;
  assign y4727 = ~n25837 ;
  assign y4728 = ~n25838 ;
  assign y4729 = n25841 ;
  assign y4730 = n25845 ;
  assign y4731 = n25850 ;
  assign y4732 = ~n25854 ;
  assign y4733 = n25862 ;
  assign y4734 = ~n25866 ;
  assign y4735 = ~n25870 ;
  assign y4736 = ~n25872 ;
  assign y4737 = n25873 ;
  assign y4738 = n25875 ;
  assign y4739 = ~n25889 ;
  assign y4740 = n25898 ;
  assign y4741 = n25903 ;
  assign y4742 = ~n25909 ;
  assign y4743 = ~n25912 ;
  assign y4744 = ~n25913 ;
  assign y4745 = n25924 ;
  assign y4746 = n25925 ;
  assign y4747 = n25929 ;
  assign y4748 = n25932 ;
  assign y4749 = ~n25935 ;
  assign y4750 = n25945 ;
  assign y4751 = ~n25946 ;
  assign y4752 = ~n25948 ;
  assign y4753 = n25950 ;
  assign y4754 = n25951 ;
  assign y4755 = ~n25954 ;
  assign y4756 = n25955 ;
  assign y4757 = ~n25959 ;
  assign y4758 = ~n25961 ;
  assign y4759 = n25964 ;
  assign y4760 = n25972 ;
  assign y4761 = n25974 ;
  assign y4762 = ~n25976 ;
  assign y4763 = ~n25979 ;
  assign y4764 = ~n25980 ;
  assign y4765 = n25983 ;
  assign y4766 = ~n25985 ;
  assign y4767 = n25987 ;
  assign y4768 = ~1'b0 ;
  assign y4769 = n25989 ;
  assign y4770 = n25990 ;
  assign y4771 = n25991 ;
  assign y4772 = n25994 ;
  assign y4773 = n25998 ;
  assign y4774 = n25999 ;
  assign y4775 = ~n26004 ;
  assign y4776 = n26009 ;
  assign y4777 = n26014 ;
  assign y4778 = n26024 ;
  assign y4779 = n26030 ;
  assign y4780 = ~n26038 ;
  assign y4781 = ~n26043 ;
  assign y4782 = ~n26046 ;
  assign y4783 = ~n26047 ;
  assign y4784 = ~n26049 ;
  assign y4785 = ~n26060 ;
  assign y4786 = n26071 ;
  assign y4787 = n26078 ;
  assign y4788 = n26079 ;
  assign y4789 = n26086 ;
  assign y4790 = n26089 ;
  assign y4791 = ~n26090 ;
  assign y4792 = n26095 ;
  assign y4793 = n26096 ;
  assign y4794 = ~n26100 ;
  assign y4795 = n26112 ;
  assign y4796 = n26116 ;
  assign y4797 = n26121 ;
  assign y4798 = n26123 ;
  assign y4799 = n26125 ;
  assign y4800 = ~n26126 ;
  assign y4801 = ~n26128 ;
  assign y4802 = ~n26131 ;
  assign y4803 = ~n26132 ;
  assign y4804 = ~n26134 ;
  assign y4805 = n26135 ;
  assign y4806 = ~n26137 ;
  assign y4807 = ~1'b0 ;
  assign y4808 = n26138 ;
  assign y4809 = n26140 ;
  assign y4810 = ~n26151 ;
  assign y4811 = n26154 ;
  assign y4812 = ~n26157 ;
  assign y4813 = n26159 ;
  assign y4814 = ~n26162 ;
  assign y4815 = ~n26166 ;
  assign y4816 = ~n26169 ;
  assign y4817 = ~n26171 ;
  assign y4818 = ~n26173 ;
  assign y4819 = n26174 ;
  assign y4820 = ~n26177 ;
  assign y4821 = ~n26179 ;
  assign y4822 = ~n26191 ;
  assign y4823 = n26193 ;
  assign y4824 = ~n26197 ;
  assign y4825 = ~n26198 ;
  assign y4826 = ~n26203 ;
  assign y4827 = n26205 ;
  assign y4828 = n26212 ;
  assign y4829 = n26213 ;
  assign y4830 = n26215 ;
  assign y4831 = n26218 ;
  assign y4832 = n26221 ;
  assign y4833 = n26224 ;
  assign y4834 = n26233 ;
  assign y4835 = n26238 ;
  assign y4836 = ~n26242 ;
  assign y4837 = n26244 ;
  assign y4838 = ~1'b0 ;
  assign y4839 = n26256 ;
  assign y4840 = n26257 ;
  assign y4841 = ~n26260 ;
  assign y4842 = n26261 ;
  assign y4843 = ~n26266 ;
  assign y4844 = n26269 ;
  assign y4845 = ~n26272 ;
  assign y4846 = ~n26281 ;
  assign y4847 = ~n26283 ;
  assign y4848 = n26285 ;
  assign y4849 = n26290 ;
  assign y4850 = n26295 ;
  assign y4851 = ~n26299 ;
  assign y4852 = n26300 ;
  assign y4853 = n26301 ;
  assign y4854 = ~n26312 ;
  assign y4855 = ~n26313 ;
  assign y4856 = n26320 ;
  assign y4857 = ~n26321 ;
  assign y4858 = n26323 ;
  assign y4859 = n26324 ;
  assign y4860 = n26328 ;
  assign y4861 = n26332 ;
  assign y4862 = ~n26334 ;
  assign y4863 = ~n26347 ;
  assign y4864 = ~n26353 ;
  assign y4865 = ~n26355 ;
  assign y4866 = n26363 ;
  assign y4867 = ~n26364 ;
  assign y4868 = ~n26373 ;
  assign y4869 = n26377 ;
  assign y4870 = ~n26379 ;
  assign y4871 = ~n26380 ;
  assign y4872 = ~n26383 ;
  assign y4873 = n26387 ;
  assign y4874 = ~n26389 ;
  assign y4875 = n26392 ;
  assign y4876 = n26397 ;
  assign y4877 = ~n26403 ;
  assign y4878 = ~n26406 ;
  assign y4879 = ~n26408 ;
  assign y4880 = n26412 ;
  assign y4881 = ~1'b0 ;
  assign y4882 = n26417 ;
  assign y4883 = ~n26420 ;
  assign y4884 = ~n26427 ;
  assign y4885 = ~n26429 ;
  assign y4886 = ~n26433 ;
  assign y4887 = ~n26438 ;
  assign y4888 = n26441 ;
  assign y4889 = ~n26445 ;
  assign y4890 = n26449 ;
  assign y4891 = n26454 ;
  assign y4892 = ~n26458 ;
  assign y4893 = n26464 ;
  assign y4894 = n26466 ;
  assign y4895 = ~n26468 ;
  assign y4896 = n26469 ;
  assign y4897 = ~n26474 ;
  assign y4898 = ~n26478 ;
  assign y4899 = ~n26481 ;
  assign y4900 = ~n26487 ;
  assign y4901 = ~n26491 ;
  assign y4902 = ~n26495 ;
  assign y4903 = ~1'b0 ;
  assign y4904 = ~n26500 ;
  assign y4905 = n26502 ;
  assign y4906 = ~n26504 ;
  assign y4907 = ~n26506 ;
  assign y4908 = n26510 ;
  assign y4909 = n26511 ;
  assign y4910 = n26512 ;
  assign y4911 = ~n26513 ;
  assign y4912 = ~n26515 ;
  assign y4913 = ~n26516 ;
  assign y4914 = ~1'b0 ;
  assign y4915 = n26518 ;
  assign y4916 = ~n26521 ;
  assign y4917 = n26522 ;
  assign y4918 = n26531 ;
  assign y4919 = n26541 ;
  assign y4920 = n26545 ;
  assign y4921 = ~n26555 ;
  assign y4922 = n26556 ;
  assign y4923 = n26559 ;
  assign y4924 = n26565 ;
  assign y4925 = ~n26566 ;
  assign y4926 = n26567 ;
  assign y4927 = n26569 ;
  assign y4928 = ~n26570 ;
  assign y4929 = n26578 ;
  assign y4930 = ~n26581 ;
  assign y4931 = ~n26583 ;
  assign y4932 = ~n26584 ;
  assign y4933 = ~n26591 ;
  assign y4934 = ~n26596 ;
  assign y4935 = n26600 ;
  assign y4936 = n26606 ;
  assign y4937 = ~n26609 ;
  assign y4938 = n26617 ;
  assign y4939 = n26620 ;
  assign y4940 = n26624 ;
  assign y4941 = n26625 ;
  assign y4942 = ~n26627 ;
  assign y4943 = ~n26628 ;
  assign y4944 = n26629 ;
  assign y4945 = ~n26634 ;
  assign y4946 = ~n26645 ;
  assign y4947 = n26647 ;
  assign y4948 = ~n26652 ;
  assign y4949 = n26653 ;
  assign y4950 = n26656 ;
  assign y4951 = ~n26657 ;
  assign y4952 = ~n26660 ;
  assign y4953 = ~n26663 ;
  assign y4954 = n26667 ;
  assign y4955 = n26672 ;
  assign y4956 = n26683 ;
  assign y4957 = n26685 ;
  assign y4958 = ~1'b0 ;
  assign y4959 = ~n26686 ;
  assign y4960 = n26691 ;
  assign y4961 = n26707 ;
  assign y4962 = ~n26710 ;
  assign y4963 = ~1'b0 ;
  assign y4964 = ~n26715 ;
  assign y4965 = ~n26716 ;
  assign y4966 = n26718 ;
  assign y4967 = ~n26722 ;
  assign y4968 = ~n26723 ;
  assign y4969 = ~n26732 ;
  assign y4970 = n26735 ;
  assign y4971 = ~n26736 ;
  assign y4972 = n26746 ;
  assign y4973 = ~1'b0 ;
  assign y4974 = n26747 ;
  assign y4975 = ~n26748 ;
  assign y4976 = n26749 ;
  assign y4977 = ~n26761 ;
  assign y4978 = ~n26765 ;
  assign y4979 = ~n26766 ;
  assign y4980 = ~n26768 ;
  assign y4981 = ~1'b0 ;
  assign y4982 = ~n26776 ;
  assign y4983 = ~n26778 ;
  assign y4984 = ~n26782 ;
  assign y4985 = n26786 ;
  assign y4986 = ~n26787 ;
  assign y4987 = n26791 ;
  assign y4988 = n26802 ;
  assign y4989 = ~1'b0 ;
  assign y4990 = ~1'b0 ;
  assign y4991 = n26804 ;
  assign y4992 = ~n26805 ;
  assign y4993 = n26807 ;
  assign y4994 = ~n26809 ;
  assign y4995 = ~n26811 ;
  assign y4996 = ~n26816 ;
  assign y4997 = ~n26825 ;
  assign y4998 = ~n26833 ;
  assign y4999 = ~n26834 ;
  assign y5000 = ~n26837 ;
  assign y5001 = n26842 ;
  assign y5002 = n26852 ;
  assign y5003 = ~n26855 ;
  assign y5004 = n26871 ;
  assign y5005 = n26872 ;
  assign y5006 = ~n26875 ;
  assign y5007 = ~n26878 ;
  assign y5008 = ~1'b0 ;
  assign y5009 = ~n26879 ;
  assign y5010 = n26887 ;
  assign y5011 = ~n26892 ;
  assign y5012 = ~n26895 ;
  assign y5013 = ~n26900 ;
  assign y5014 = n26904 ;
  assign y5015 = n26910 ;
  assign y5016 = n26913 ;
  assign y5017 = n26928 ;
  assign y5018 = n26931 ;
  assign y5019 = ~n26946 ;
  assign y5020 = n26953 ;
  assign y5021 = ~n26955 ;
  assign y5022 = ~n26969 ;
  assign y5023 = n26973 ;
  assign y5024 = ~n26974 ;
  assign y5025 = ~n26976 ;
  assign y5026 = ~n26978 ;
  assign y5027 = ~n26982 ;
  assign y5028 = ~n26986 ;
  assign y5029 = n26990 ;
  assign y5030 = ~n26992 ;
  assign y5031 = ~n26995 ;
  assign y5032 = ~n26996 ;
  assign y5033 = n27004 ;
  assign y5034 = n27005 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = n27006 ;
  assign y5037 = ~n27009 ;
  assign y5038 = n27018 ;
  assign y5039 = n27021 ;
  assign y5040 = ~n27022 ;
  assign y5041 = n27028 ;
  assign y5042 = ~n27035 ;
  assign y5043 = n27037 ;
  assign y5044 = ~n27038 ;
  assign y5045 = ~n27039 ;
  assign y5046 = ~n27044 ;
  assign y5047 = ~n27047 ;
  assign y5048 = ~n27048 ;
  assign y5049 = ~n27049 ;
  assign y5050 = n27055 ;
  assign y5051 = ~n27057 ;
  assign y5052 = n27063 ;
  assign y5053 = ~n27067 ;
  assign y5054 = n27069 ;
  assign y5055 = ~n27072 ;
  assign y5056 = n27074 ;
  assign y5057 = n27077 ;
  assign y5058 = ~n27078 ;
  assign y5059 = n27082 ;
  assign y5060 = ~n27084 ;
  assign y5061 = ~n27089 ;
  assign y5062 = ~n27091 ;
  assign y5063 = ~n27092 ;
  assign y5064 = n27096 ;
  assign y5065 = n27098 ;
  assign y5066 = n27100 ;
  assign y5067 = n27105 ;
  assign y5068 = n27108 ;
  assign y5069 = n27112 ;
  assign y5070 = n27114 ;
  assign y5071 = ~n27120 ;
  assign y5072 = ~n10036 ;
  assign y5073 = n27123 ;
  assign y5074 = ~n27126 ;
  assign y5075 = ~n27128 ;
  assign y5076 = n27129 ;
  assign y5077 = ~n27136 ;
  assign y5078 = ~n27138 ;
  assign y5079 = ~n27139 ;
  assign y5080 = n27144 ;
  assign y5081 = ~n27146 ;
  assign y5082 = n27147 ;
  assign y5083 = ~n27149 ;
  assign y5084 = ~n27151 ;
  assign y5085 = n27152 ;
  assign y5086 = n27153 ;
  assign y5087 = ~n27156 ;
  assign y5088 = ~1'b0 ;
  assign y5089 = ~n27159 ;
  assign y5090 = ~n27160 ;
  assign y5091 = ~n27162 ;
  assign y5092 = n27163 ;
  assign y5093 = ~n27168 ;
  assign y5094 = ~n27171 ;
  assign y5095 = n27174 ;
  assign y5096 = n27179 ;
  assign y5097 = ~n27180 ;
  assign y5098 = n27182 ;
  assign y5099 = ~n27185 ;
  assign y5100 = n27190 ;
  assign y5101 = n27200 ;
  assign y5102 = n27205 ;
  assign y5103 = n27211 ;
  assign y5104 = ~n27212 ;
  assign y5105 = ~n27216 ;
  assign y5106 = ~n7048 ;
  assign y5107 = ~n27217 ;
  assign y5108 = ~n27226 ;
  assign y5109 = n27228 ;
  assign y5110 = n27229 ;
  assign y5111 = n27232 ;
  assign y5112 = n27235 ;
  assign y5113 = n27236 ;
  assign y5114 = ~n27244 ;
  assign y5115 = ~n27247 ;
  assign y5116 = ~n27250 ;
  assign y5117 = ~n27258 ;
  assign y5118 = n27259 ;
  assign y5119 = ~n27264 ;
  assign y5120 = n27273 ;
  assign y5121 = ~n27274 ;
  assign y5122 = ~n27277 ;
  assign y5123 = n27278 ;
  assign y5124 = n27280 ;
  assign y5125 = n27281 ;
  assign y5126 = ~n27289 ;
  assign y5127 = ~n27291 ;
  assign y5128 = ~n27296 ;
  assign y5129 = n27303 ;
  assign y5130 = n27304 ;
  assign y5131 = n27305 ;
  assign y5132 = n27310 ;
  assign y5133 = ~1'b0 ;
  assign y5134 = ~n27315 ;
  assign y5135 = ~1'b0 ;
  assign y5136 = n27318 ;
  assign y5137 = ~n27321 ;
  assign y5138 = ~n27324 ;
  assign y5139 = ~n27325 ;
  assign y5140 = n27333 ;
  assign y5141 = ~n27335 ;
  assign y5142 = ~n27336 ;
  assign y5143 = n27340 ;
  assign y5144 = n27341 ;
  assign y5145 = n27344 ;
  assign y5146 = ~1'b0 ;
  assign y5147 = n27345 ;
  assign y5148 = ~n27350 ;
  assign y5149 = ~n27355 ;
  assign y5150 = n27361 ;
  assign y5151 = ~n27378 ;
  assign y5152 = n27386 ;
  assign y5153 = ~n27394 ;
  assign y5154 = n27395 ;
  assign y5155 = n27402 ;
  assign y5156 = ~1'b0 ;
  assign y5157 = n27406 ;
  assign y5158 = ~n27409 ;
  assign y5159 = ~n27411 ;
  assign y5160 = n27417 ;
  assign y5161 = ~n27418 ;
  assign y5162 = ~n27421 ;
  assign y5163 = ~n27423 ;
  assign y5164 = ~n27429 ;
  assign y5165 = ~n27439 ;
  assign y5166 = n27444 ;
  assign y5167 = ~n27446 ;
  assign y5168 = n27455 ;
  assign y5169 = ~n27467 ;
  assign y5170 = ~n27471 ;
  assign y5171 = ~n27473 ;
  assign y5172 = ~n27474 ;
  assign y5173 = ~n27475 ;
  assign y5174 = n27482 ;
  assign y5175 = n27486 ;
  assign y5176 = n27487 ;
  assign y5177 = n27498 ;
  assign y5178 = ~n27503 ;
  assign y5179 = n27505 ;
  assign y5180 = ~n27508 ;
  assign y5181 = ~n27514 ;
  assign y5182 = ~n27516 ;
  assign y5183 = n27527 ;
  assign y5184 = ~n27530 ;
  assign y5185 = ~n27535 ;
  assign y5186 = n27537 ;
  assign y5187 = n27538 ;
  assign y5188 = ~1'b0 ;
  assign y5189 = ~n27539 ;
  assign y5190 = ~1'b0 ;
  assign y5191 = n27543 ;
  assign y5192 = ~n27548 ;
  assign y5193 = ~n27551 ;
  assign y5194 = ~1'b0 ;
  assign y5195 = ~n27553 ;
  assign y5196 = n27557 ;
  assign y5197 = ~n27559 ;
  assign y5198 = n27563 ;
  assign y5199 = ~n27571 ;
  assign y5200 = n27572 ;
  assign y5201 = n27573 ;
  assign y5202 = ~n27578 ;
  assign y5203 = ~n27584 ;
  assign y5204 = n27586 ;
  assign y5205 = n27587 ;
  assign y5206 = ~n27597 ;
  assign y5207 = n27600 ;
  assign y5208 = n27603 ;
  assign y5209 = ~n27604 ;
  assign y5210 = n27605 ;
  assign y5211 = n27608 ;
  assign y5212 = ~n27609 ;
  assign y5213 = n27610 ;
  assign y5214 = n27611 ;
  assign y5215 = n27614 ;
  assign y5216 = n27618 ;
  assign y5217 = ~n27621 ;
  assign y5218 = ~n27622 ;
  assign y5219 = ~n27628 ;
  assign y5220 = ~n27631 ;
  assign y5221 = ~n27633 ;
  assign y5222 = n27635 ;
  assign y5223 = ~n27641 ;
  assign y5224 = ~1'b0 ;
  assign y5225 = ~n27643 ;
  assign y5226 = n27645 ;
  assign y5227 = ~n27647 ;
  assign y5228 = ~n27649 ;
  assign y5229 = n27653 ;
  assign y5230 = ~n27656 ;
  assign y5231 = ~n27661 ;
  assign y5232 = n27665 ;
  assign y5233 = n27666 ;
  assign y5234 = n27670 ;
  assign y5235 = ~n27673 ;
  assign y5236 = n27676 ;
  assign y5237 = n27688 ;
  assign y5238 = n27689 ;
  assign y5239 = ~n27693 ;
  assign y5240 = n27698 ;
  assign y5241 = ~n27702 ;
  assign y5242 = ~n27705 ;
  assign y5243 = ~n27708 ;
  assign y5244 = n27712 ;
  assign y5245 = ~n27714 ;
  assign y5246 = n27717 ;
  assign y5247 = n27719 ;
  assign y5248 = ~n27722 ;
  assign y5249 = ~n27723 ;
  assign y5250 = n27725 ;
  assign y5251 = n27730 ;
  assign y5252 = n27734 ;
  assign y5253 = ~n27736 ;
  assign y5254 = n27739 ;
  assign y5255 = ~n27741 ;
  assign y5256 = n27743 ;
  assign y5257 = ~n27753 ;
  assign y5258 = ~n27755 ;
  assign y5259 = ~n27758 ;
  assign y5260 = ~n27762 ;
  assign y5261 = ~n27768 ;
  assign y5262 = ~n27776 ;
  assign y5263 = ~n27778 ;
  assign y5264 = ~n27779 ;
  assign y5265 = n27780 ;
  assign y5266 = ~n27781 ;
  assign y5267 = ~n27783 ;
  assign y5268 = ~n27787 ;
  assign y5269 = n27790 ;
  assign y5270 = n27791 ;
  assign y5271 = ~n27792 ;
  assign y5272 = n27793 ;
  assign y5273 = ~n27796 ;
  assign y5274 = ~n27804 ;
  assign y5275 = ~n27813 ;
  assign y5276 = n27820 ;
  assign y5277 = n27821 ;
  assign y5278 = n27826 ;
  assign y5279 = n27831 ;
  assign y5280 = ~n27832 ;
  assign y5281 = n27834 ;
  assign y5282 = ~n27835 ;
  assign y5283 = ~n27837 ;
  assign y5284 = n27839 ;
  assign y5285 = ~n27840 ;
  assign y5286 = n27844 ;
  assign y5287 = ~n27851 ;
  assign y5288 = n27855 ;
  assign y5289 = ~n27856 ;
  assign y5290 = n27864 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = ~n27866 ;
  assign y5293 = n27869 ;
  assign y5294 = n27874 ;
  assign y5295 = ~1'b0 ;
  assign y5296 = n27877 ;
  assign y5297 = n27879 ;
  assign y5298 = ~n27883 ;
  assign y5299 = ~n27884 ;
  assign y5300 = n27887 ;
  assign y5301 = n27889 ;
  assign y5302 = n27893 ;
  assign y5303 = ~n27899 ;
  assign y5304 = ~n27903 ;
  assign y5305 = ~n27906 ;
  assign y5306 = n27910 ;
  assign y5307 = ~n27919 ;
  assign y5308 = ~n27925 ;
  assign y5309 = n27926 ;
  assign y5310 = n27929 ;
  assign y5311 = ~n27936 ;
  assign y5312 = ~n27946 ;
  assign y5313 = n27953 ;
  assign y5314 = n27954 ;
  assign y5315 = n27964 ;
  assign y5316 = ~n27966 ;
  assign y5317 = n27967 ;
  assign y5318 = n27968 ;
  assign y5319 = n14936 ;
  assign y5320 = n27973 ;
  assign y5321 = ~n27978 ;
  assign y5322 = n27979 ;
  assign y5323 = ~n27986 ;
  assign y5324 = n27989 ;
  assign y5325 = ~n27993 ;
  assign y5326 = n27994 ;
  assign y5327 = ~n27998 ;
  assign y5328 = n28001 ;
  assign y5329 = ~n28005 ;
  assign y5330 = ~n28009 ;
  assign y5331 = n28015 ;
  assign y5332 = ~n28019 ;
  assign y5333 = n28028 ;
  assign y5334 = n28035 ;
  assign y5335 = n28045 ;
  assign y5336 = ~n28046 ;
  assign y5337 = n28047 ;
  assign y5338 = n28050 ;
  assign y5339 = ~n28054 ;
  assign y5340 = ~n28056 ;
  assign y5341 = n28058 ;
  assign y5342 = ~n28059 ;
  assign y5343 = n28060 ;
  assign y5344 = ~n28064 ;
  assign y5345 = ~n28070 ;
  assign y5346 = ~n28071 ;
  assign y5347 = ~n28075 ;
  assign y5348 = n28079 ;
  assign y5349 = ~n28089 ;
  assign y5350 = ~n28099 ;
  assign y5351 = ~n28100 ;
  assign y5352 = n28101 ;
  assign y5353 = ~n28105 ;
  assign y5354 = ~n28108 ;
  assign y5355 = n28109 ;
  assign y5356 = n28110 ;
  assign y5357 = ~n28113 ;
  assign y5358 = n28114 ;
  assign y5359 = n28122 ;
  assign y5360 = ~1'b0 ;
  assign y5361 = ~n28123 ;
  assign y5362 = ~n28128 ;
  assign y5363 = n28129 ;
  assign y5364 = n28130 ;
  assign y5365 = n28132 ;
  assign y5366 = n28135 ;
  assign y5367 = n28149 ;
  assign y5368 = n28150 ;
  assign y5369 = ~n28153 ;
  assign y5370 = n28154 ;
  assign y5371 = ~n28159 ;
  assign y5372 = n28163 ;
  assign y5373 = ~n28164 ;
  assign y5374 = n28166 ;
  assign y5375 = ~n28169 ;
  assign y5376 = ~n28171 ;
  assign y5377 = ~n28173 ;
  assign y5378 = n28174 ;
  assign y5379 = ~n28178 ;
  assign y5380 = ~n28182 ;
  assign y5381 = ~n28188 ;
  assign y5382 = ~n28190 ;
  assign y5383 = n28194 ;
  assign y5384 = n28199 ;
  assign y5385 = ~n28207 ;
  assign y5386 = n28217 ;
  assign y5387 = ~n28221 ;
  assign y5388 = n28227 ;
  assign y5389 = n28231 ;
  assign y5390 = ~n28234 ;
  assign y5391 = ~n28237 ;
  assign y5392 = ~1'b0 ;
  assign y5393 = ~n28244 ;
  assign y5394 = ~n28248 ;
  assign y5395 = n28249 ;
  assign y5396 = ~n28252 ;
  assign y5397 = n28253 ;
  assign y5398 = ~n28260 ;
  assign y5399 = n28265 ;
  assign y5400 = n28268 ;
  assign y5401 = n28271 ;
  assign y5402 = ~n28275 ;
  assign y5403 = n28282 ;
  assign y5404 = ~n28291 ;
  assign y5405 = ~n28292 ;
  assign y5406 = n28294 ;
  assign y5407 = ~1'b0 ;
  assign y5408 = ~1'b0 ;
  assign y5409 = ~n28296 ;
  assign y5410 = n28300 ;
  assign y5411 = n28303 ;
  assign y5412 = n28305 ;
  assign y5413 = ~n28307 ;
  assign y5414 = ~n28309 ;
  assign y5415 = ~n28310 ;
  assign y5416 = ~n28311 ;
  assign y5417 = ~n28316 ;
  assign y5418 = n28317 ;
  assign y5419 = ~n28319 ;
  assign y5420 = ~n28320 ;
  assign y5421 = n28321 ;
  assign y5422 = ~1'b0 ;
  assign y5423 = n28322 ;
  assign y5424 = ~n28325 ;
  assign y5425 = ~n28334 ;
  assign y5426 = n28336 ;
  assign y5427 = n28337 ;
  assign y5428 = ~n28342 ;
  assign y5429 = ~n28351 ;
  assign y5430 = ~n28352 ;
  assign y5431 = n28353 ;
  assign y5432 = n28357 ;
  assign y5433 = n28359 ;
  assign y5434 = n28362 ;
  assign y5435 = n28363 ;
  assign y5436 = n28372 ;
  assign y5437 = n28379 ;
  assign y5438 = n28383 ;
  assign y5439 = n28387 ;
  assign y5440 = n28388 ;
  assign y5441 = ~n28390 ;
  assign y5442 = ~n28393 ;
  assign y5443 = n28395 ;
  assign y5444 = n28399 ;
  assign y5445 = ~n28403 ;
  assign y5446 = ~n28406 ;
  assign y5447 = ~n28410 ;
  assign y5448 = ~n28414 ;
  assign y5449 = n28417 ;
  assign y5450 = n28422 ;
  assign y5451 = ~n28427 ;
  assign y5452 = n28428 ;
  assign y5453 = ~n28433 ;
  assign y5454 = ~n28434 ;
  assign y5455 = n28436 ;
  assign y5456 = n28440 ;
  assign y5457 = n28446 ;
  assign y5458 = ~n28452 ;
  assign y5459 = n28454 ;
  assign y5460 = n28457 ;
  assign y5461 = ~n28459 ;
  assign y5462 = n28463 ;
  assign y5463 = n28471 ;
  assign y5464 = ~n28478 ;
  assign y5465 = ~n28485 ;
  assign y5466 = ~n28488 ;
  assign y5467 = ~n1255 ;
  assign y5468 = ~n28493 ;
  assign y5469 = n28500 ;
  assign y5470 = ~n28509 ;
  assign y5471 = n28518 ;
  assign y5472 = ~n28519 ;
  assign y5473 = n28521 ;
  assign y5474 = ~1'b0 ;
  assign y5475 = ~n28526 ;
  assign y5476 = n28528 ;
  assign y5477 = ~n28529 ;
  assign y5478 = ~n28533 ;
  assign y5479 = ~n28536 ;
  assign y5480 = ~1'b0 ;
  assign y5481 = ~n28540 ;
  assign y5482 = n28541 ;
  assign y5483 = n28544 ;
  assign y5484 = n28545 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = ~n28547 ;
  assign y5487 = n28549 ;
  assign y5488 = n28559 ;
  assign y5489 = ~n28562 ;
  assign y5490 = n28564 ;
  assign y5491 = n28567 ;
  assign y5492 = n28568 ;
  assign y5493 = n28573 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = ~1'b0 ;
  assign y5496 = n28577 ;
  assign y5497 = n28587 ;
  assign y5498 = ~n28589 ;
  assign y5499 = n28590 ;
  assign y5500 = ~n28593 ;
  assign y5501 = ~n28599 ;
  assign y5502 = ~n28602 ;
  assign y5503 = ~n28603 ;
  assign y5504 = n28608 ;
  assign y5505 = n28610 ;
  assign y5506 = n28614 ;
  assign y5507 = ~n28618 ;
  assign y5508 = ~n28621 ;
  assign y5509 = n28622 ;
  assign y5510 = n28624 ;
  assign y5511 = ~n28626 ;
  assign y5512 = ~n28634 ;
  assign y5513 = n28635 ;
  assign y5514 = ~n28644 ;
  assign y5515 = n28645 ;
  assign y5516 = n28646 ;
  assign y5517 = ~n28648 ;
  assign y5518 = ~n28649 ;
  assign y5519 = n28652 ;
  assign y5520 = n28655 ;
  assign y5521 = ~n28661 ;
  assign y5522 = n28663 ;
  assign y5523 = n28665 ;
  assign y5524 = n28667 ;
  assign y5525 = n28668 ;
  assign y5526 = n28673 ;
  assign y5527 = n28674 ;
  assign y5528 = n28678 ;
  assign y5529 = ~n28682 ;
  assign y5530 = n28685 ;
  assign y5531 = ~n28693 ;
  assign y5532 = ~n28697 ;
  assign y5533 = n28701 ;
  assign y5534 = n28702 ;
  assign y5535 = n28703 ;
  assign y5536 = n28705 ;
  assign y5537 = ~n28708 ;
  assign y5538 = ~n28711 ;
  assign y5539 = n28717 ;
  assign y5540 = n28719 ;
  assign y5541 = ~n28723 ;
  assign y5542 = n28725 ;
  assign y5543 = ~1'b0 ;
  assign y5544 = ~n28727 ;
  assign y5545 = n28731 ;
  assign y5546 = n28734 ;
  assign y5547 = n28735 ;
  assign y5548 = ~n28736 ;
  assign y5549 = n28743 ;
  assign y5550 = ~n28746 ;
  assign y5551 = ~n28751 ;
  assign y5552 = ~n28754 ;
  assign y5553 = ~n28755 ;
  assign y5554 = ~n28758 ;
  assign y5555 = ~1'b0 ;
  assign y5556 = ~n28760 ;
  assign y5557 = n28765 ;
  assign y5558 = ~n28772 ;
  assign y5559 = ~n28776 ;
  assign y5560 = n28784 ;
  assign y5561 = ~n28786 ;
  assign y5562 = n28789 ;
  assign y5563 = n28796 ;
  assign y5564 = n28799 ;
  assign y5565 = n28800 ;
  assign y5566 = n28803 ;
  assign y5567 = n28807 ;
  assign y5568 = ~n28811 ;
  assign y5569 = n28812 ;
  assign y5570 = n28813 ;
  assign y5571 = n28817 ;
  assign y5572 = n28818 ;
  assign y5573 = ~n28823 ;
  assign y5574 = ~n28828 ;
  assign y5575 = n28829 ;
  assign y5576 = ~n28833 ;
  assign y5577 = n28835 ;
  assign y5578 = ~n28843 ;
  assign y5579 = n28854 ;
  assign y5580 = n28857 ;
  assign y5581 = n28861 ;
  assign y5582 = ~n28873 ;
  assign y5583 = n28874 ;
  assign y5584 = n28875 ;
  assign y5585 = n28881 ;
  assign y5586 = ~n28883 ;
  assign y5587 = ~1'b0 ;
  assign y5588 = n28895 ;
  assign y5589 = ~n28900 ;
  assign y5590 = n28907 ;
  assign y5591 = ~n28911 ;
  assign y5592 = n28914 ;
  assign y5593 = ~n28917 ;
  assign y5594 = n28935 ;
  assign y5595 = n28937 ;
  assign y5596 = n28941 ;
  assign y5597 = ~n28944 ;
  assign y5598 = ~n28946 ;
  assign y5599 = n28947 ;
  assign y5600 = n28949 ;
  assign y5601 = n28959 ;
  assign y5602 = ~n28969 ;
  assign y5603 = n28971 ;
  assign y5604 = ~n28977 ;
  assign y5605 = ~n28985 ;
  assign y5606 = n28989 ;
  assign y5607 = ~n28990 ;
  assign y5608 = ~n28992 ;
  assign y5609 = n28994 ;
  assign y5610 = n28999 ;
  assign y5611 = ~n29001 ;
  assign y5612 = n29005 ;
  assign y5613 = ~n29007 ;
  assign y5614 = n29010 ;
  assign y5615 = ~n29015 ;
  assign y5616 = ~n29018 ;
  assign y5617 = n29022 ;
  assign y5618 = n29023 ;
  assign y5619 = ~n29029 ;
  assign y5620 = n29032 ;
  assign y5621 = ~n29033 ;
  assign y5622 = ~n29037 ;
  assign y5623 = n29038 ;
  assign y5624 = n29046 ;
  assign y5625 = n29047 ;
  assign y5626 = n29048 ;
  assign y5627 = n29049 ;
  assign y5628 = ~n29052 ;
  assign y5629 = ~n29053 ;
  assign y5630 = n29054 ;
  assign y5631 = ~n29057 ;
  assign y5632 = n29060 ;
  assign y5633 = ~n29063 ;
  assign y5634 = ~n29065 ;
  assign y5635 = ~n29066 ;
  assign y5636 = ~n29067 ;
  assign y5637 = n29072 ;
  assign y5638 = ~n29075 ;
  assign y5639 = n29076 ;
  assign y5640 = n29078 ;
  assign y5641 = n29080 ;
  assign y5642 = n29081 ;
  assign y5643 = ~n29088 ;
  assign y5644 = n29091 ;
  assign y5645 = ~n29092 ;
  assign y5646 = ~n29094 ;
  assign y5647 = n29097 ;
  assign y5648 = ~n29106 ;
  assign y5649 = n29107 ;
  assign y5650 = n29108 ;
  assign y5651 = n29111 ;
  assign y5652 = ~n29113 ;
  assign y5653 = n29115 ;
  assign y5654 = ~n29116 ;
  assign y5655 = ~n29118 ;
  assign y5656 = n29129 ;
  assign y5657 = n29130 ;
  assign y5658 = n29140 ;
  assign y5659 = ~n29144 ;
  assign y5660 = n29145 ;
  assign y5661 = ~n29152 ;
  assign y5662 = ~n29155 ;
  assign y5663 = n29160 ;
  assign y5664 = ~n29163 ;
  assign y5665 = ~n29172 ;
  assign y5666 = n29173 ;
  assign y5667 = ~n29178 ;
  assign y5668 = n29182 ;
  assign y5669 = ~n29184 ;
  assign y5670 = n29185 ;
  assign y5671 = n29188 ;
  assign y5672 = ~n29192 ;
  assign y5673 = ~n29193 ;
  assign y5674 = ~n29194 ;
  assign y5675 = n29195 ;
  assign y5676 = ~n29197 ;
  assign y5677 = ~1'b0 ;
  assign y5678 = n29200 ;
  assign y5679 = ~n29201 ;
  assign y5680 = n29203 ;
  assign y5681 = n29206 ;
  assign y5682 = ~n29209 ;
  assign y5683 = n29216 ;
  assign y5684 = n29219 ;
  assign y5685 = ~1'b0 ;
  assign y5686 = ~n29223 ;
  assign y5687 = n29224 ;
  assign y5688 = ~n29225 ;
  assign y5689 = ~n29231 ;
  assign y5690 = n29238 ;
  assign y5691 = n29239 ;
  assign y5692 = n29241 ;
  assign y5693 = n29247 ;
  assign y5694 = ~1'b0 ;
  assign y5695 = ~n29254 ;
  assign y5696 = n29258 ;
  assign y5697 = n29260 ;
  assign y5698 = ~n29264 ;
  assign y5699 = ~1'b0 ;
  assign y5700 = n29265 ;
  assign y5701 = ~n29269 ;
  assign y5702 = ~n29275 ;
  assign y5703 = ~n29278 ;
  assign y5704 = ~n29279 ;
  assign y5705 = ~n29283 ;
  assign y5706 = n29286 ;
  assign y5707 = n29287 ;
  assign y5708 = ~n29303 ;
  assign y5709 = ~n29314 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = ~n29320 ;
  assign y5712 = n29321 ;
  assign y5713 = n29322 ;
  assign y5714 = n29325 ;
  assign y5715 = ~n29328 ;
  assign y5716 = n29346 ;
  assign y5717 = ~n29347 ;
  assign y5718 = n29351 ;
  assign y5719 = ~n29356 ;
  assign y5720 = ~n29359 ;
  assign y5721 = ~n29360 ;
  assign y5722 = n29363 ;
  assign y5723 = ~1'b0 ;
  assign y5724 = n29369 ;
  assign y5725 = n29373 ;
  assign y5726 = ~n29382 ;
  assign y5727 = n29386 ;
  assign y5728 = ~n29391 ;
  assign y5729 = ~n29396 ;
  assign y5730 = n29397 ;
  assign y5731 = ~n29400 ;
  assign y5732 = ~n29401 ;
  assign y5733 = n29402 ;
  assign y5734 = ~n29409 ;
  assign y5735 = ~n29410 ;
  assign y5736 = n29415 ;
  assign y5737 = n29422 ;
  assign y5738 = ~n29427 ;
  assign y5739 = ~n29431 ;
  assign y5740 = ~n29433 ;
  assign y5741 = n29440 ;
  assign y5742 = n29441 ;
  assign y5743 = n29446 ;
  assign y5744 = n29447 ;
  assign y5745 = ~n29455 ;
  assign y5746 = ~n29457 ;
  assign y5747 = ~n29460 ;
  assign y5748 = ~n29461 ;
  assign y5749 = n29464 ;
  assign y5750 = ~n29467 ;
  assign y5751 = ~n29468 ;
  assign y5752 = ~n29473 ;
  assign y5753 = n29476 ;
  assign y5754 = n29477 ;
  assign y5755 = n29479 ;
  assign y5756 = n29484 ;
  assign y5757 = ~n29486 ;
  assign y5758 = n29502 ;
  assign y5759 = ~n29504 ;
  assign y5760 = n29505 ;
  assign y5761 = n29507 ;
  assign y5762 = ~n29509 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = n29513 ;
  assign y5765 = ~n29524 ;
  assign y5766 = ~n29529 ;
  assign y5767 = n29532 ;
  assign y5768 = ~n29534 ;
  assign y5769 = n29535 ;
  assign y5770 = ~n29538 ;
  assign y5771 = ~n29546 ;
  assign y5772 = ~n29548 ;
  assign y5773 = ~n29549 ;
  assign y5774 = n29555 ;
  assign y5775 = ~n29562 ;
  assign y5776 = n29563 ;
  assign y5777 = n29564 ;
  assign y5778 = ~n29572 ;
  assign y5779 = ~1'b0 ;
  assign y5780 = ~n29574 ;
  assign y5781 = n29581 ;
  assign y5782 = n29584 ;
  assign y5783 = n29589 ;
  assign y5784 = n29590 ;
  assign y5785 = n29593 ;
  assign y5786 = ~n29594 ;
  assign y5787 = ~n29598 ;
  assign y5788 = ~n29599 ;
  assign y5789 = ~n29601 ;
  assign y5790 = n29605 ;
  assign y5791 = n29606 ;
  assign y5792 = ~n29609 ;
  assign y5793 = n29610 ;
  assign y5794 = ~n29613 ;
  assign y5795 = ~n29614 ;
  assign y5796 = n29615 ;
  assign y5797 = ~n29621 ;
  assign y5798 = ~1'b0 ;
  assign y5799 = ~n29626 ;
  assign y5800 = ~n29630 ;
  assign y5801 = n29633 ;
  assign y5802 = n29634 ;
  assign y5803 = ~n29635 ;
  assign y5804 = n29636 ;
  assign y5805 = ~1'b0 ;
  assign y5806 = n29638 ;
  assign y5807 = ~n29639 ;
  assign y5808 = ~n29642 ;
  assign y5809 = n29646 ;
  assign y5810 = ~n26476 ;
  assign y5811 = ~n29647 ;
  assign y5812 = ~n29648 ;
  assign y5813 = ~n29650 ;
  assign y5814 = n29655 ;
  assign y5815 = ~n29657 ;
  assign y5816 = ~n29663 ;
  assign y5817 = n29664 ;
  assign y5818 = ~n29667 ;
  assign y5819 = n29670 ;
  assign y5820 = n29676 ;
  assign y5821 = ~n29678 ;
  assign y5822 = n29679 ;
  assign y5823 = ~n29685 ;
  assign y5824 = ~n29687 ;
  assign y5825 = n29689 ;
  assign y5826 = n29690 ;
  assign y5827 = ~n29693 ;
  assign y5828 = n29702 ;
  assign y5829 = n29703 ;
  assign y5830 = ~n29706 ;
  assign y5831 = n29709 ;
  assign y5832 = ~n29711 ;
  assign y5833 = ~n29712 ;
  assign y5834 = ~n29722 ;
  assign y5835 = n29723 ;
  assign y5836 = ~n29725 ;
  assign y5837 = n29726 ;
  assign y5838 = ~n29728 ;
  assign y5839 = ~n29733 ;
  assign y5840 = ~n29739 ;
  assign y5841 = ~n29744 ;
  assign y5842 = ~n29751 ;
  assign y5843 = ~n29753 ;
  assign y5844 = ~n29756 ;
  assign y5845 = ~n29760 ;
  assign y5846 = ~n29767 ;
  assign y5847 = ~n29771 ;
  assign y5848 = n29777 ;
  assign y5849 = ~n29780 ;
  assign y5850 = ~n29784 ;
  assign y5851 = n29785 ;
  assign y5852 = n29793 ;
  assign y5853 = ~n29797 ;
  assign y5854 = ~1'b0 ;
  assign y5855 = n29802 ;
  assign y5856 = n29805 ;
  assign y5857 = n29807 ;
  assign y5858 = n29810 ;
  assign y5859 = ~n29815 ;
  assign y5860 = ~n29822 ;
  assign y5861 = ~n29823 ;
  assign y5862 = n29824 ;
  assign y5863 = n29830 ;
  assign y5864 = ~n29831 ;
  assign y5865 = n29833 ;
  assign y5866 = n29834 ;
  assign y5867 = ~n29844 ;
  assign y5868 = n29854 ;
  assign y5869 = ~n29855 ;
  assign y5870 = n29859 ;
  assign y5871 = ~n29862 ;
  assign y5872 = n29864 ;
  assign y5873 = ~n29865 ;
  assign y5874 = n29867 ;
  assign y5875 = ~n29869 ;
  assign y5876 = ~n29871 ;
  assign y5877 = n29873 ;
  assign y5878 = n29878 ;
  assign y5879 = ~n29880 ;
  assign y5880 = n29886 ;
  assign y5881 = n29887 ;
  assign y5882 = n29888 ;
  assign y5883 = n29890 ;
  assign y5884 = ~n29894 ;
  assign y5885 = ~n29895 ;
  assign y5886 = ~n29896 ;
  assign y5887 = n29898 ;
  assign y5888 = ~n29899 ;
  assign y5889 = ~n29901 ;
  assign y5890 = ~n29902 ;
  assign y5891 = ~n29903 ;
  assign y5892 = n29907 ;
  assign y5893 = ~n29913 ;
  assign y5894 = ~n29914 ;
  assign y5895 = ~n29916 ;
  assign y5896 = ~n29922 ;
  assign y5897 = ~n29924 ;
  assign y5898 = n29930 ;
  assign y5899 = n29931 ;
  assign y5900 = ~n29933 ;
  assign y5901 = ~n29937 ;
  assign y5902 = ~n29938 ;
  assign y5903 = ~n29943 ;
  assign y5904 = ~n29948 ;
  assign y5905 = n29951 ;
  assign y5906 = ~n29958 ;
  assign y5907 = n29959 ;
  assign y5908 = ~n29968 ;
  assign y5909 = n29969 ;
  assign y5910 = ~n29970 ;
  assign y5911 = ~n29971 ;
  assign y5912 = ~1'b0 ;
  assign y5913 = n29975 ;
  assign y5914 = n29981 ;
  assign y5915 = ~n29983 ;
  assign y5916 = n29985 ;
  assign y5917 = ~n29989 ;
  assign y5918 = ~n29990 ;
  assign y5919 = ~1'b0 ;
  assign y5920 = n29995 ;
  assign y5921 = ~n30000 ;
  assign y5922 = ~n30002 ;
  assign y5923 = n30003 ;
  assign y5924 = ~n30007 ;
  assign y5925 = n30010 ;
  assign y5926 = ~n30017 ;
  assign y5927 = n30026 ;
  assign y5928 = ~n30029 ;
  assign y5929 = n30031 ;
  assign y5930 = ~n30032 ;
  assign y5931 = n30034 ;
  assign y5932 = ~n30035 ;
  assign y5933 = ~n30037 ;
  assign y5934 = ~1'b0 ;
  assign y5935 = n30042 ;
  assign y5936 = n30043 ;
  assign y5937 = ~n30048 ;
  assign y5938 = ~n30057 ;
  assign y5939 = ~1'b0 ;
  assign y5940 = ~n30060 ;
  assign y5941 = n30061 ;
  assign y5942 = ~n30062 ;
  assign y5943 = n30067 ;
  assign y5944 = ~n30068 ;
  assign y5945 = ~n30073 ;
  assign y5946 = ~1'b0 ;
  assign y5947 = ~n30077 ;
  assign y5948 = ~n30085 ;
  assign y5949 = n30086 ;
  assign y5950 = ~n30087 ;
  assign y5951 = n30088 ;
  assign y5952 = n30098 ;
  assign y5953 = ~1'b0 ;
  assign y5954 = ~n30100 ;
  assign y5955 = ~1'b0 ;
  assign y5956 = ~1'b0 ;
  assign y5957 = ~n30108 ;
  assign y5958 = ~n30115 ;
  assign y5959 = ~n30121 ;
  assign y5960 = ~n30122 ;
  assign y5961 = ~n30124 ;
  assign y5962 = n30125 ;
  assign y5963 = ~n30126 ;
  assign y5964 = ~n30136 ;
  assign y5965 = ~n30142 ;
  assign y5966 = n30144 ;
  assign y5967 = n30146 ;
  assign y5968 = n30149 ;
  assign y5969 = n30153 ;
  assign y5970 = ~n30159 ;
  assign y5971 = ~n30164 ;
  assign y5972 = ~n30165 ;
  assign y5973 = ~n30174 ;
  assign y5974 = ~1'b0 ;
  assign y5975 = ~n30175 ;
  assign y5976 = n30176 ;
  assign y5977 = n30179 ;
  assign y5978 = ~n30181 ;
  assign y5979 = ~n30186 ;
  assign y5980 = n30188 ;
  assign y5981 = n30192 ;
  assign y5982 = ~n30201 ;
  assign y5983 = ~n30206 ;
  assign y5984 = ~n30211 ;
  assign y5985 = n30218 ;
  assign y5986 = n30219 ;
  assign y5987 = n30224 ;
  assign y5988 = ~1'b0 ;
  assign y5989 = n30228 ;
  assign y5990 = n30233 ;
  assign y5991 = ~n30235 ;
  assign y5992 = ~n30236 ;
  assign y5993 = ~n30237 ;
  assign y5994 = ~n30238 ;
  assign y5995 = n30239 ;
  assign y5996 = n30242 ;
  assign y5997 = n30246 ;
  assign y5998 = ~n30249 ;
  assign y5999 = ~n30250 ;
  assign y6000 = n30256 ;
  assign y6001 = n30257 ;
  assign y6002 = n30262 ;
  assign y6003 = ~n30270 ;
  assign y6004 = n30272 ;
  assign y6005 = n30273 ;
  assign y6006 = ~n30277 ;
  assign y6007 = ~1'b0 ;
  assign y6008 = n30278 ;
  assign y6009 = n30279 ;
  assign y6010 = ~n30288 ;
  assign y6011 = ~n30293 ;
  assign y6012 = ~n30295 ;
  assign y6013 = n30302 ;
  assign y6014 = n30303 ;
  assign y6015 = ~n30307 ;
  assign y6016 = n30310 ;
  assign y6017 = n30313 ;
  assign y6018 = ~n30314 ;
  assign y6019 = n30320 ;
  assign y6020 = n30322 ;
  assign y6021 = ~n30323 ;
  assign y6022 = n30325 ;
  assign y6023 = n30326 ;
  assign y6024 = n30330 ;
  assign y6025 = ~n30331 ;
  assign y6026 = n30332 ;
  assign y6027 = ~n30334 ;
  assign y6028 = ~n30336 ;
  assign y6029 = ~n30342 ;
  assign y6030 = ~n30344 ;
  assign y6031 = ~n30348 ;
  assign y6032 = n30355 ;
  assign y6033 = ~n30356 ;
  assign y6034 = ~n30360 ;
  assign y6035 = ~n30366 ;
  assign y6036 = ~n30369 ;
  assign y6037 = ~1'b0 ;
  assign y6038 = ~n30373 ;
  assign y6039 = ~n30377 ;
  assign y6040 = ~n30379 ;
  assign y6041 = n30380 ;
  assign y6042 = ~n30381 ;
  assign y6043 = n30386 ;
  assign y6044 = n30387 ;
  assign y6045 = ~n30388 ;
  assign y6046 = ~n30389 ;
  assign y6047 = n30391 ;
  assign y6048 = ~n30395 ;
  assign y6049 = n30402 ;
  assign y6050 = n30405 ;
  assign y6051 = ~n30412 ;
  assign y6052 = ~n30413 ;
  assign y6053 = ~n30415 ;
  assign y6054 = ~n30416 ;
  assign y6055 = ~n30417 ;
  assign y6056 = n30419 ;
  assign y6057 = ~n30420 ;
  assign y6058 = ~1'b0 ;
  assign y6059 = ~n30424 ;
  assign y6060 = n30427 ;
  assign y6061 = n30429 ;
  assign y6062 = n30431 ;
  assign y6063 = ~n30432 ;
  assign y6064 = ~n30433 ;
  assign y6065 = n30438 ;
  assign y6066 = ~n30444 ;
  assign y6067 = ~n30448 ;
  assign y6068 = ~n30450 ;
  assign y6069 = ~n30453 ;
  assign y6070 = n30454 ;
  assign y6071 = ~n30460 ;
  assign y6072 = n30461 ;
  assign y6073 = ~n30467 ;
  assign y6074 = n30468 ;
  assign y6075 = ~n30471 ;
  assign y6076 = n30474 ;
  assign y6077 = ~1'b0 ;
  assign y6078 = ~n30477 ;
  assign y6079 = n30481 ;
  assign y6080 = n30484 ;
  assign y6081 = ~n30485 ;
  assign y6082 = ~n30488 ;
  assign y6083 = ~n30491 ;
  assign y6084 = ~n30497 ;
  assign y6085 = ~n30501 ;
  assign y6086 = n30505 ;
  assign y6087 = ~1'b0 ;
  assign y6088 = ~n30510 ;
  assign y6089 = ~n30512 ;
  assign y6090 = ~n30514 ;
  assign y6091 = n30517 ;
  assign y6092 = n30519 ;
  assign y6093 = n30520 ;
  assign y6094 = ~n30524 ;
  assign y6095 = n30525 ;
  assign y6096 = ~n30526 ;
  assign y6097 = ~n30533 ;
  assign y6098 = n30546 ;
  assign y6099 = ~n30550 ;
  assign y6100 = n30553 ;
  assign y6101 = ~n30557 ;
  assign y6102 = ~n30560 ;
  assign y6103 = ~n30566 ;
  assign y6104 = n30568 ;
  assign y6105 = n30569 ;
  assign y6106 = ~n30572 ;
  assign y6107 = ~n30576 ;
  assign y6108 = n30578 ;
  assign y6109 = ~n30587 ;
  assign y6110 = ~n30589 ;
  assign y6111 = ~n30591 ;
  assign y6112 = ~n30598 ;
  assign y6113 = n30613 ;
  assign y6114 = n30614 ;
  assign y6115 = n30617 ;
  assign y6116 = n30619 ;
  assign y6117 = n30622 ;
  assign y6118 = n30623 ;
  assign y6119 = n30625 ;
  assign y6120 = n30626 ;
  assign y6121 = n30632 ;
  assign y6122 = ~n30637 ;
  assign y6123 = n30641 ;
  assign y6124 = n30645 ;
  assign y6125 = n30649 ;
  assign y6126 = ~n30652 ;
  assign y6127 = ~n30653 ;
  assign y6128 = n30657 ;
  assign y6129 = ~n30659 ;
  assign y6130 = ~n30662 ;
  assign y6131 = ~n30667 ;
  assign y6132 = n30674 ;
  assign y6133 = n30676 ;
  assign y6134 = n30677 ;
  assign y6135 = ~n30679 ;
  assign y6136 = ~n4751 ;
  assign y6137 = n30684 ;
  assign y6138 = n30685 ;
  assign y6139 = n30689 ;
  assign y6140 = n30696 ;
  assign y6141 = n30704 ;
  assign y6142 = n30705 ;
  assign y6143 = ~n30713 ;
  assign y6144 = ~n30718 ;
  assign y6145 = n30720 ;
  assign y6146 = n30721 ;
  assign y6147 = n30731 ;
  assign y6148 = n30734 ;
  assign y6149 = n30736 ;
  assign y6150 = n30738 ;
  assign y6151 = n30748 ;
  assign y6152 = ~n30751 ;
  assign y6153 = n30752 ;
  assign y6154 = ~n30757 ;
  assign y6155 = n30760 ;
  assign y6156 = n30762 ;
  assign y6157 = ~n30768 ;
  assign y6158 = n30770 ;
  assign y6159 = ~n30773 ;
  assign y6160 = n30775 ;
  assign y6161 = n30778 ;
  assign y6162 = n30781 ;
  assign y6163 = n30782 ;
  assign y6164 = ~n30785 ;
  assign y6165 = n30788 ;
  assign y6166 = n30789 ;
  assign y6167 = n30793 ;
  assign y6168 = n30794 ;
  assign y6169 = n30800 ;
  assign y6170 = ~n30802 ;
  assign y6171 = ~n30803 ;
  assign y6172 = n30809 ;
  assign y6173 = ~n30818 ;
  assign y6174 = n30821 ;
  assign y6175 = n30831 ;
  assign y6176 = n30835 ;
  assign y6177 = n30838 ;
  assign y6178 = n30842 ;
  assign y6179 = n30850 ;
  assign y6180 = ~n30856 ;
  assign y6181 = n30858 ;
  assign y6182 = ~n30862 ;
  assign y6183 = ~n30867 ;
  assign y6184 = n30871 ;
  assign y6185 = n30873 ;
  assign y6186 = ~n30874 ;
  assign y6187 = ~n30879 ;
  assign y6188 = ~n30880 ;
  assign y6189 = n30882 ;
  assign y6190 = n30889 ;
  assign y6191 = n30893 ;
  assign y6192 = n30894 ;
  assign y6193 = n30898 ;
  assign y6194 = n30900 ;
  assign y6195 = n30905 ;
  assign y6196 = ~n30908 ;
  assign y6197 = n30914 ;
  assign y6198 = ~n30919 ;
  assign y6199 = n30923 ;
  assign y6200 = ~n30924 ;
  assign y6201 = n30925 ;
  assign y6202 = ~n30926 ;
  assign y6203 = ~n30928 ;
  assign y6204 = ~n30932 ;
  assign y6205 = ~n30934 ;
  assign y6206 = n30943 ;
  assign y6207 = ~n30946 ;
  assign y6208 = n30947 ;
  assign y6209 = n30952 ;
  assign y6210 = n30958 ;
  assign y6211 = n30959 ;
  assign y6212 = n30968 ;
  assign y6213 = ~n30969 ;
  assign y6214 = ~n30970 ;
  assign y6215 = ~n30971 ;
  assign y6216 = n30972 ;
  assign y6217 = n30975 ;
  assign y6218 = n30980 ;
  assign y6219 = ~n30981 ;
  assign y6220 = n30984 ;
  assign y6221 = ~n30990 ;
  assign y6222 = ~n30992 ;
  assign y6223 = ~n30997 ;
  assign y6224 = n31008 ;
  assign y6225 = ~n31009 ;
  assign y6226 = n31013 ;
  assign y6227 = n31018 ;
  assign y6228 = ~n31019 ;
  assign y6229 = ~n31031 ;
  assign y6230 = ~n31032 ;
  assign y6231 = ~n31042 ;
  assign y6232 = n31044 ;
  assign y6233 = ~n31045 ;
  assign y6234 = ~n31054 ;
  assign y6235 = ~n31056 ;
  assign y6236 = ~n31061 ;
  assign y6237 = n31063 ;
  assign y6238 = ~n31064 ;
  assign y6239 = n31066 ;
  assign y6240 = n31071 ;
  assign y6241 = ~n31073 ;
  assign y6242 = ~n31074 ;
  assign y6243 = ~n31076 ;
  assign y6244 = n31077 ;
  assign y6245 = n31093 ;
  assign y6246 = ~n31094 ;
  assign y6247 = n31095 ;
  assign y6248 = n31098 ;
  assign y6249 = ~n31099 ;
  assign y6250 = ~n31104 ;
  assign y6251 = n31105 ;
  assign y6252 = ~n31106 ;
  assign y6253 = ~n31109 ;
  assign y6254 = n31111 ;
  assign y6255 = n31117 ;
  assign y6256 = n31119 ;
  assign y6257 = ~n31124 ;
  assign y6258 = n31129 ;
  assign y6259 = ~n31130 ;
  assign y6260 = ~n31131 ;
  assign y6261 = n31137 ;
  assign y6262 = n31139 ;
  assign y6263 = ~n31140 ;
  assign y6264 = n31148 ;
  assign y6265 = n31154 ;
  assign y6266 = ~n31155 ;
  assign y6267 = ~1'b0 ;
  assign y6268 = ~n31156 ;
  assign y6269 = ~n31164 ;
  assign y6270 = ~n31169 ;
  assign y6271 = ~n31172 ;
  assign y6272 = ~n31175 ;
  assign y6273 = n31179 ;
  assign y6274 = ~n31181 ;
  assign y6275 = ~n31182 ;
  assign y6276 = ~n31186 ;
  assign y6277 = ~n31189 ;
  assign y6278 = ~n31192 ;
  assign y6279 = n31193 ;
  assign y6280 = n31199 ;
  assign y6281 = n31201 ;
  assign y6282 = n31206 ;
  assign y6283 = ~n31215 ;
  assign y6284 = n31217 ;
  assign y6285 = ~n31226 ;
  assign y6286 = ~n31228 ;
  assign y6287 = ~n31230 ;
  assign y6288 = ~n31233 ;
  assign y6289 = ~1'b0 ;
  assign y6290 = ~n31237 ;
  assign y6291 = ~n31241 ;
  assign y6292 = n31244 ;
  assign y6293 = n31245 ;
  assign y6294 = n31247 ;
  assign y6295 = ~n31253 ;
  assign y6296 = ~n31255 ;
  assign y6297 = n31257 ;
  assign y6298 = n31262 ;
  assign y6299 = n31263 ;
  assign y6300 = n31267 ;
  assign y6301 = ~n31268 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = n31269 ;
  assign y6304 = n31276 ;
  assign y6305 = n31277 ;
  assign y6306 = ~n31279 ;
  assign y6307 = ~n31281 ;
  assign y6308 = ~n31287 ;
  assign y6309 = ~n31288 ;
  assign y6310 = n31290 ;
  assign y6311 = n31292 ;
  assign y6312 = ~n31295 ;
  assign y6313 = n31298 ;
  assign y6314 = n31302 ;
  assign y6315 = ~n31306 ;
  assign y6316 = ~n31308 ;
  assign y6317 = n31309 ;
  assign y6318 = ~n31310 ;
  assign y6319 = ~n31312 ;
  assign y6320 = ~n31313 ;
  assign y6321 = ~n31320 ;
  assign y6322 = ~n31321 ;
  assign y6323 = ~n31323 ;
  assign y6324 = n31330 ;
  assign y6325 = ~n31332 ;
  assign y6326 = n31337 ;
  assign y6327 = ~n31340 ;
  assign y6328 = ~n31342 ;
  assign y6329 = n31344 ;
  assign y6330 = n31346 ;
  assign y6331 = ~1'b0 ;
  assign y6332 = n31353 ;
  assign y6333 = ~n31355 ;
  assign y6334 = ~n31356 ;
  assign y6335 = n31358 ;
  assign y6336 = ~n31360 ;
  assign y6337 = n31370 ;
  assign y6338 = n31372 ;
  assign y6339 = ~n31375 ;
  assign y6340 = ~n31380 ;
  assign y6341 = n31384 ;
  assign y6342 = ~n31386 ;
  assign y6343 = ~n31391 ;
  assign y6344 = ~n31392 ;
  assign y6345 = n31394 ;
  assign y6346 = ~n31396 ;
  assign y6347 = ~n31399 ;
  assign y6348 = ~n31400 ;
  assign y6349 = n31402 ;
  assign y6350 = ~n31411 ;
  assign y6351 = n31413 ;
  assign y6352 = n31416 ;
  assign y6353 = ~n31421 ;
  assign y6354 = ~n31426 ;
  assign y6355 = ~1'b0 ;
  assign y6356 = ~n31433 ;
  assign y6357 = ~n31436 ;
  assign y6358 = n31442 ;
  assign y6359 = n31443 ;
  assign y6360 = n31447 ;
  assign y6361 = n31450 ;
  assign y6362 = ~n31452 ;
  assign y6363 = ~n31453 ;
  assign y6364 = ~n31455 ;
  assign y6365 = ~n31462 ;
  assign y6366 = n31463 ;
  assign y6367 = n31464 ;
  assign y6368 = n31468 ;
  assign y6369 = n31470 ;
  assign y6370 = n31479 ;
  assign y6371 = ~n31483 ;
  assign y6372 = ~n31485 ;
  assign y6373 = n31493 ;
  assign y6374 = n31494 ;
  assign y6375 = n31497 ;
  assign y6376 = ~n31501 ;
  assign y6377 = ~n31503 ;
  assign y6378 = ~n31505 ;
  assign y6379 = ~n31506 ;
  assign y6380 = n31521 ;
  assign y6381 = n31525 ;
  assign y6382 = ~n31531 ;
  assign y6383 = ~n1054 ;
  assign y6384 = n31535 ;
  assign y6385 = ~n31538 ;
  assign y6386 = n31540 ;
  assign y6387 = ~n31541 ;
  assign y6388 = ~n31542 ;
  assign y6389 = n31543 ;
  assign y6390 = ~n31548 ;
  assign y6391 = ~n31549 ;
  assign y6392 = ~n31553 ;
  assign y6393 = ~n31556 ;
  assign y6394 = ~1'b0 ;
  assign y6395 = n31561 ;
  assign y6396 = ~n31564 ;
  assign y6397 = ~n31565 ;
  assign y6398 = n31566 ;
  assign y6399 = n31571 ;
  assign y6400 = n31575 ;
  assign y6401 = ~n31579 ;
  assign y6402 = ~n31580 ;
  assign y6403 = n31584 ;
  assign y6404 = ~n31591 ;
  assign y6405 = n31593 ;
  assign y6406 = ~n31598 ;
  assign y6407 = ~n31605 ;
  assign y6408 = n31610 ;
  assign y6409 = n31611 ;
  assign y6410 = ~n31614 ;
  assign y6411 = ~n31620 ;
  assign y6412 = ~n31624 ;
  assign y6413 = n31628 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = n31632 ;
  assign y6416 = ~n31634 ;
  assign y6417 = n31636 ;
  assign y6418 = n31641 ;
  assign y6419 = ~n31643 ;
  assign y6420 = ~n31646 ;
  assign y6421 = n31651 ;
  assign y6422 = n31652 ;
  assign y6423 = n31656 ;
  assign y6424 = ~n31659 ;
  assign y6425 = ~n31663 ;
  assign y6426 = ~n31671 ;
  assign y6427 = ~n31674 ;
  assign y6428 = n31677 ;
  assign y6429 = ~n31678 ;
  assign y6430 = n31682 ;
  assign y6431 = n31686 ;
  assign y6432 = ~n31688 ;
  assign y6433 = ~n31695 ;
  assign y6434 = n31698 ;
  assign y6435 = n31700 ;
  assign y6436 = n31705 ;
  assign y6437 = n31710 ;
  assign y6438 = ~n31711 ;
  assign y6439 = ~n31714 ;
  assign y6440 = ~n31715 ;
  assign y6441 = ~n31723 ;
  assign y6442 = ~n31725 ;
  assign y6443 = ~n31731 ;
  assign y6444 = n31733 ;
  assign y6445 = ~1'b0 ;
  assign y6446 = ~n31740 ;
  assign y6447 = ~n31743 ;
  assign y6448 = n31749 ;
  assign y6449 = ~n31755 ;
  assign y6450 = n31756 ;
  assign y6451 = ~n31762 ;
  assign y6452 = ~n31763 ;
  assign y6453 = ~n31765 ;
  assign y6454 = n31766 ;
  assign y6455 = n31772 ;
  assign y6456 = ~n31777 ;
  assign y6457 = n31781 ;
  assign y6458 = n31785 ;
  assign y6459 = n31790 ;
  assign y6460 = n31795 ;
  assign y6461 = ~n31797 ;
  assign y6462 = ~n31801 ;
  assign y6463 = ~n31806 ;
  assign y6464 = ~n31809 ;
  assign y6465 = n31814 ;
  assign y6466 = ~n31817 ;
  assign y6467 = ~1'b0 ;
  assign y6468 = n31818 ;
  assign y6469 = ~n31826 ;
  assign y6470 = ~n31827 ;
  assign y6471 = n31828 ;
  assign y6472 = ~1'b0 ;
  assign y6473 = ~n31829 ;
  assign y6474 = ~n31831 ;
  assign y6475 = ~n31833 ;
  assign y6476 = ~n31835 ;
  assign y6477 = n31841 ;
  assign y6478 = ~n31842 ;
  assign y6479 = ~1'b0 ;
  assign y6480 = n31843 ;
  assign y6481 = n31845 ;
  assign y6482 = ~n31847 ;
  assign y6483 = n31850 ;
  assign y6484 = ~n31854 ;
  assign y6485 = ~n31859 ;
  assign y6486 = ~1'b0 ;
  assign y6487 = ~1'b0 ;
  assign y6488 = n31862 ;
  assign y6489 = ~n31867 ;
  assign y6490 = n31870 ;
  assign y6491 = ~n31873 ;
  assign y6492 = ~n31874 ;
  assign y6493 = n31877 ;
  assign y6494 = ~n31880 ;
  assign y6495 = n31885 ;
  assign y6496 = ~n31889 ;
  assign y6497 = n31891 ;
  assign y6498 = ~n31893 ;
  assign y6499 = ~n31894 ;
  assign y6500 = ~n31898 ;
  assign y6501 = n31900 ;
  assign y6502 = ~n31904 ;
  assign y6503 = n31906 ;
  assign y6504 = ~n31908 ;
  assign y6505 = n31910 ;
  assign y6506 = ~n31911 ;
  assign y6507 = n31913 ;
  assign y6508 = ~n31919 ;
  assign y6509 = n31926 ;
  assign y6510 = n31930 ;
  assign y6511 = ~n31931 ;
  assign y6512 = ~n31932 ;
  assign y6513 = n31939 ;
  assign y6514 = ~n31942 ;
  assign y6515 = n31943 ;
  assign y6516 = n31944 ;
  assign y6517 = ~n31945 ;
  assign y6518 = ~n31948 ;
  assign y6519 = ~n31952 ;
  assign y6520 = n31956 ;
  assign y6521 = n31967 ;
  assign y6522 = n31970 ;
  assign y6523 = n31974 ;
  assign y6524 = ~n31975 ;
  assign y6525 = ~n31981 ;
  assign y6526 = n31984 ;
  assign y6527 = n31990 ;
  assign y6528 = n31993 ;
  assign y6529 = ~n31995 ;
  assign y6530 = n32001 ;
  assign y6531 = ~n32007 ;
  assign y6532 = ~n32008 ;
  assign y6533 = ~1'b0 ;
  assign y6534 = ~n32010 ;
  assign y6535 = ~n32011 ;
  assign y6536 = n32013 ;
  assign y6537 = ~n32030 ;
  assign y6538 = ~n32032 ;
  assign y6539 = n32033 ;
  assign y6540 = n32034 ;
  assign y6541 = ~n32035 ;
  assign y6542 = ~n32037 ;
  assign y6543 = ~1'b0 ;
  assign y6544 = ~n32045 ;
  assign y6545 = ~n32048 ;
  assign y6546 = ~n32049 ;
  assign y6547 = n32058 ;
  assign y6548 = ~n32060 ;
  assign y6549 = n32061 ;
  assign y6550 = n32065 ;
  assign y6551 = ~1'b0 ;
  assign y6552 = n32067 ;
  assign y6553 = ~n32068 ;
  assign y6554 = n32071 ;
  assign y6555 = n32074 ;
  assign y6556 = ~1'b0 ;
  assign y6557 = ~n32078 ;
  assign y6558 = ~n32085 ;
  assign y6559 = ~n32088 ;
  assign y6560 = n32097 ;
  assign y6561 = ~n32103 ;
  assign y6562 = ~n32106 ;
  assign y6563 = ~1'b0 ;
  assign y6564 = n32109 ;
  assign y6565 = ~n32112 ;
  assign y6566 = ~n32117 ;
  assign y6567 = ~n32119 ;
  assign y6568 = ~1'b0 ;
  assign y6569 = n32121 ;
  assign y6570 = ~n32122 ;
  assign y6571 = ~n32126 ;
  assign y6572 = n32129 ;
  assign y6573 = n32132 ;
  assign y6574 = n32133 ;
  assign y6575 = n32135 ;
  assign y6576 = ~n32138 ;
  assign y6577 = n32141 ;
  assign y6578 = n32144 ;
  assign y6579 = n32146 ;
  assign y6580 = n32149 ;
  assign y6581 = n32155 ;
  assign y6582 = ~n32156 ;
  assign y6583 = n32157 ;
  assign y6584 = ~n32159 ;
  assign y6585 = ~n32164 ;
  assign y6586 = ~n32167 ;
  assign y6587 = ~n32171 ;
  assign y6588 = ~n32172 ;
  assign y6589 = ~n32173 ;
  assign y6590 = n32175 ;
  assign y6591 = n32176 ;
  assign y6592 = ~1'b0 ;
  assign y6593 = ~n32185 ;
  assign y6594 = n32187 ;
  assign y6595 = n32192 ;
  assign y6596 = n32193 ;
  assign y6597 = n32195 ;
  assign y6598 = ~1'b0 ;
  assign y6599 = ~n32199 ;
  assign y6600 = n32202 ;
  assign y6601 = n32205 ;
  assign y6602 = ~n32206 ;
  assign y6603 = ~n32208 ;
  assign y6604 = ~n32210 ;
  assign y6605 = ~n32214 ;
  assign y6606 = n32216 ;
  assign y6607 = n32218 ;
  assign y6608 = ~n32223 ;
  assign y6609 = n32229 ;
  assign y6610 = n32231 ;
  assign y6611 = ~n32247 ;
  assign y6612 = ~n32255 ;
  assign y6613 = ~n32261 ;
  assign y6614 = ~n32272 ;
  assign y6615 = ~n32274 ;
  assign y6616 = ~n32278 ;
  assign y6617 = ~n32279 ;
  assign y6618 = n32280 ;
  assign y6619 = n32284 ;
  assign y6620 = n32289 ;
  assign y6621 = n32291 ;
  assign y6622 = ~n32292 ;
  assign y6623 = ~n32297 ;
  assign y6624 = ~n32299 ;
  assign y6625 = n32302 ;
  assign y6626 = ~1'b0 ;
  assign y6627 = ~1'b0 ;
  assign y6628 = n32304 ;
  assign y6629 = ~n32308 ;
  assign y6630 = ~n32311 ;
  assign y6631 = ~n32313 ;
  assign y6632 = ~1'b0 ;
  assign y6633 = n32316 ;
  assign y6634 = n32317 ;
  assign y6635 = ~n32318 ;
  assign y6636 = n32319 ;
  assign y6637 = n32323 ;
  assign y6638 = ~n32325 ;
  assign y6639 = n32327 ;
  assign y6640 = n32332 ;
  assign y6641 = n32337 ;
  assign y6642 = ~n32338 ;
  assign y6643 = n32341 ;
  assign y6644 = n32344 ;
  assign y6645 = n32346 ;
  assign y6646 = ~n32353 ;
  assign y6647 = n32354 ;
  assign y6648 = n32355 ;
  assign y6649 = ~n32357 ;
  assign y6650 = ~n32365 ;
  assign y6651 = n32366 ;
  assign y6652 = ~n32371 ;
  assign y6653 = ~n32372 ;
  assign y6654 = n32374 ;
  assign y6655 = n32376 ;
  assign y6656 = ~n32383 ;
  assign y6657 = ~n32387 ;
  assign y6658 = n32389 ;
  assign y6659 = n32395 ;
  assign y6660 = ~n32399 ;
  assign y6661 = ~n32405 ;
  assign y6662 = n32406 ;
  assign y6663 = ~n32408 ;
  assign y6664 = ~n32410 ;
  assign y6665 = n32411 ;
  assign y6666 = n32413 ;
  assign y6667 = ~n32418 ;
  assign y6668 = n32423 ;
  assign y6669 = ~n32425 ;
  assign y6670 = n32427 ;
  assign y6671 = ~n32430 ;
  assign y6672 = ~n32431 ;
  assign y6673 = ~n32432 ;
  assign y6674 = n32437 ;
  assign y6675 = ~n32441 ;
  assign y6676 = n32446 ;
  assign y6677 = n32448 ;
  assign y6678 = n32450 ;
  assign y6679 = n32451 ;
  assign y6680 = n32454 ;
  assign y6681 = n32456 ;
  assign y6682 = ~n32457 ;
  assign y6683 = ~n32458 ;
  assign y6684 = n32459 ;
  assign y6685 = n32462 ;
  assign y6686 = ~n32464 ;
  assign y6687 = n32465 ;
  assign y6688 = ~n32467 ;
  assign y6689 = n32469 ;
  assign y6690 = n32470 ;
  assign y6691 = n32471 ;
  assign y6692 = n32474 ;
  assign y6693 = n32480 ;
  assign y6694 = ~n32484 ;
  assign y6695 = n32492 ;
  assign y6696 = n32493 ;
  assign y6697 = n32499 ;
  assign y6698 = n32501 ;
  assign y6699 = ~n32504 ;
  assign y6700 = n32512 ;
  assign y6701 = ~n32517 ;
  assign y6702 = n32519 ;
  assign y6703 = n32533 ;
  assign y6704 = ~n32534 ;
  assign y6705 = ~n32537 ;
  assign y6706 = ~n32540 ;
  assign y6707 = n32544 ;
  assign y6708 = ~n32558 ;
  assign y6709 = ~n32560 ;
  assign y6710 = n32561 ;
  assign y6711 = ~n32562 ;
  assign y6712 = ~n32563 ;
  assign y6713 = n32564 ;
  assign y6714 = n32569 ;
  assign y6715 = ~n32573 ;
  assign y6716 = n32578 ;
  assign y6717 = ~n32581 ;
  assign y6718 = ~n32582 ;
  assign y6719 = ~1'b0 ;
  assign y6720 = ~1'b0 ;
  assign y6721 = n32585 ;
  assign y6722 = n32586 ;
  assign y6723 = n32587 ;
  assign y6724 = ~1'b0 ;
  assign y6725 = ~n32590 ;
  assign y6726 = ~n32591 ;
  assign y6727 = ~n32592 ;
  assign y6728 = n32596 ;
  assign y6729 = n32599 ;
  assign y6730 = ~n32603 ;
  assign y6731 = ~n32604 ;
  assign y6732 = n32605 ;
  assign y6733 = n32612 ;
  assign y6734 = ~n32616 ;
  assign y6735 = n32623 ;
  assign y6736 = ~n32627 ;
  assign y6737 = n32633 ;
  assign y6738 = n32638 ;
  assign y6739 = ~1'b0 ;
  assign y6740 = ~n32642 ;
  assign y6741 = n32643 ;
  assign y6742 = n32646 ;
  assign y6743 = ~n32648 ;
  assign y6744 = ~n32651 ;
  assign y6745 = ~n32653 ;
  assign y6746 = ~n32660 ;
  assign y6747 = n32665 ;
  assign y6748 = ~n32670 ;
  assign y6749 = ~n32671 ;
  assign y6750 = ~n32675 ;
  assign y6751 = ~n32683 ;
  assign y6752 = n32685 ;
  assign y6753 = n32693 ;
  assign y6754 = n32695 ;
  assign y6755 = n32696 ;
  assign y6756 = ~n32699 ;
  assign y6757 = ~1'b0 ;
  assign y6758 = ~n32702 ;
  assign y6759 = n32706 ;
  assign y6760 = ~n32708 ;
  assign y6761 = n32709 ;
  assign y6762 = ~n32713 ;
  assign y6763 = n32715 ;
  assign y6764 = ~n32720 ;
  assign y6765 = n32724 ;
  assign y6766 = ~n32726 ;
  assign y6767 = n32727 ;
  assign y6768 = ~n32731 ;
  assign y6769 = n32732 ;
  assign y6770 = n32736 ;
  assign y6771 = n32739 ;
  assign y6772 = n32743 ;
  assign y6773 = n32751 ;
  assign y6774 = ~n32757 ;
  assign y6775 = n32759 ;
  assign y6776 = n32763 ;
  assign y6777 = n32765 ;
  assign y6778 = n32769 ;
  assign y6779 = n32770 ;
  assign y6780 = n32776 ;
  assign y6781 = ~n32777 ;
  assign y6782 = ~n32778 ;
  assign y6783 = n32782 ;
  assign y6784 = ~n32783 ;
  assign y6785 = ~n32784 ;
  assign y6786 = n32785 ;
  assign y6787 = n32787 ;
  assign y6788 = ~n32790 ;
  assign y6789 = ~n32791 ;
  assign y6790 = ~n32797 ;
  assign y6791 = n32804 ;
  assign y6792 = ~n32805 ;
  assign y6793 = ~n32810 ;
  assign y6794 = ~n32811 ;
  assign y6795 = n32813 ;
  assign y6796 = n32817 ;
  assign y6797 = n32823 ;
  assign y6798 = n32829 ;
  assign y6799 = n32832 ;
  assign y6800 = ~n32835 ;
  assign y6801 = n32836 ;
  assign y6802 = n32842 ;
  assign y6803 = n32843 ;
  assign y6804 = ~1'b0 ;
  assign y6805 = ~n32846 ;
  assign y6806 = ~n32850 ;
  assign y6807 = n32854 ;
  assign y6808 = n32855 ;
  assign y6809 = ~n32856 ;
  assign y6810 = n32861 ;
  assign y6811 = n32869 ;
  assign y6812 = ~n32871 ;
  assign y6813 = ~n32873 ;
  assign y6814 = ~n32878 ;
  assign y6815 = ~n32879 ;
  assign y6816 = ~n32880 ;
  assign y6817 = ~n32882 ;
  assign y6818 = n32885 ;
  assign y6819 = ~n32892 ;
  assign y6820 = ~n32894 ;
  assign y6821 = ~n32897 ;
  assign y6822 = ~n32899 ;
  assign y6823 = ~n32901 ;
  assign y6824 = ~n32902 ;
  assign y6825 = n32903 ;
  assign y6826 = ~n32905 ;
  assign y6827 = n32906 ;
  assign y6828 = ~n32908 ;
  assign y6829 = n32909 ;
  assign y6830 = ~n32912 ;
  assign y6831 = ~n32914 ;
  assign y6832 = ~n32921 ;
  assign y6833 = n32924 ;
  assign y6834 = ~n32929 ;
  assign y6835 = ~n32930 ;
  assign y6836 = n32934 ;
  assign y6837 = ~n32935 ;
  assign y6838 = ~1'b0 ;
  assign y6839 = ~n32937 ;
  assign y6840 = n32940 ;
  assign y6841 = n32943 ;
  assign y6842 = n32950 ;
  assign y6843 = n32954 ;
  assign y6844 = ~1'b0 ;
  assign y6845 = ~n32955 ;
  assign y6846 = n32957 ;
  assign y6847 = n32965 ;
  assign y6848 = ~n32966 ;
  assign y6849 = ~n32968 ;
  assign y6850 = n32975 ;
  assign y6851 = ~n32981 ;
  assign y6852 = ~n32982 ;
  assign y6853 = n32984 ;
  assign y6854 = ~n32987 ;
  assign y6855 = n32992 ;
  assign y6856 = n33003 ;
  assign y6857 = n33004 ;
  assign y6858 = n33005 ;
  assign y6859 = n33008 ;
  assign y6860 = n33012 ;
  assign y6861 = ~n33014 ;
  assign y6862 = ~n33017 ;
  assign y6863 = ~n33019 ;
  assign y6864 = n33027 ;
  assign y6865 = n33028 ;
  assign y6866 = n33030 ;
  assign y6867 = n33040 ;
  assign y6868 = ~n33043 ;
  assign y6869 = n33044 ;
  assign y6870 = ~n33050 ;
  assign y6871 = ~n33054 ;
  assign y6872 = ~n33059 ;
  assign y6873 = ~n33070 ;
  assign y6874 = n33073 ;
  assign y6875 = ~n33074 ;
  assign y6876 = ~n33078 ;
  assign y6877 = ~n33079 ;
  assign y6878 = n33080 ;
  assign y6879 = ~n33084 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = n33086 ;
  assign y6882 = ~n33097 ;
  assign y6883 = ~n33100 ;
  assign y6884 = n33106 ;
  assign y6885 = ~n33108 ;
  assign y6886 = ~n33109 ;
  assign y6887 = n33111 ;
  assign y6888 = n33117 ;
  assign y6889 = ~n33119 ;
  assign y6890 = ~n33125 ;
  assign y6891 = ~n33126 ;
  assign y6892 = ~1'b0 ;
  assign y6893 = n33131 ;
  assign y6894 = ~n33133 ;
  assign y6895 = ~n33138 ;
  assign y6896 = ~n33140 ;
  assign y6897 = n33142 ;
  assign y6898 = ~n33145 ;
  assign y6899 = n33148 ;
  assign y6900 = ~n33151 ;
  assign y6901 = n33153 ;
  assign y6902 = ~n33155 ;
  assign y6903 = n33158 ;
  assign y6904 = ~n33163 ;
  assign y6905 = n33164 ;
  assign y6906 = ~n33166 ;
  assign y6907 = ~n33168 ;
  assign y6908 = n33171 ;
  assign y6909 = ~n33174 ;
  assign y6910 = ~1'b0 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = n33176 ;
  assign y6913 = ~n33177 ;
  assign y6914 = ~n33189 ;
  assign y6915 = ~n33190 ;
  assign y6916 = n33192 ;
  assign y6917 = n33196 ;
  assign y6918 = n33198 ;
  assign y6919 = n33200 ;
  assign y6920 = n33202 ;
  assign y6921 = n33206 ;
  assign y6922 = n33209 ;
  assign y6923 = ~n33212 ;
  assign y6924 = n33215 ;
  assign y6925 = ~n33220 ;
  assign y6926 = ~n33223 ;
  assign y6927 = n33225 ;
  assign y6928 = ~n33227 ;
  assign y6929 = n33228 ;
  assign y6930 = n33229 ;
  assign y6931 = n33234 ;
  assign y6932 = ~n33237 ;
  assign y6933 = n33239 ;
  assign y6934 = ~1'b0 ;
  assign y6935 = n33243 ;
  assign y6936 = n33246 ;
  assign y6937 = ~n33252 ;
  assign y6938 = ~n33261 ;
  assign y6939 = n33262 ;
  assign y6940 = ~n33264 ;
  assign y6941 = ~n33266 ;
  assign y6942 = ~n33269 ;
  assign y6943 = ~n33274 ;
  assign y6944 = n33276 ;
  assign y6945 = ~n33279 ;
  assign y6946 = n33283 ;
  assign y6947 = n33286 ;
  assign y6948 = ~n33287 ;
  assign y6949 = n33293 ;
  assign y6950 = n33294 ;
  assign y6951 = n33296 ;
  assign y6952 = ~n33305 ;
  assign y6953 = n33307 ;
  assign y6954 = ~n33310 ;
  assign y6955 = ~n33312 ;
  assign y6956 = ~n33314 ;
  assign y6957 = ~n33318 ;
  assign y6958 = ~n33320 ;
  assign y6959 = ~1'b0 ;
  assign y6960 = n33325 ;
  assign y6961 = n33327 ;
  assign y6962 = n33338 ;
  assign y6963 = ~n33340 ;
  assign y6964 = n33343 ;
  assign y6965 = n33345 ;
  assign y6966 = n33351 ;
  assign y6967 = ~n33357 ;
  assign y6968 = ~n33369 ;
  assign y6969 = n33376 ;
  assign y6970 = n33377 ;
  assign y6971 = n33381 ;
  assign y6972 = ~n33383 ;
  assign y6973 = n33390 ;
  assign y6974 = n33394 ;
  assign y6975 = ~n33401 ;
  assign y6976 = ~1'b0 ;
  assign y6977 = ~n33406 ;
  assign y6978 = n33407 ;
  assign y6979 = ~n33412 ;
  assign y6980 = n33415 ;
  assign y6981 = ~n33417 ;
  assign y6982 = ~n33418 ;
  assign y6983 = ~n33419 ;
  assign y6984 = ~n33421 ;
  assign y6985 = ~n33425 ;
  assign y6986 = ~n33426 ;
  assign y6987 = ~n33427 ;
  assign y6988 = n33431 ;
  assign y6989 = n33435 ;
  assign y6990 = ~n33442 ;
  assign y6991 = ~n33445 ;
  assign y6992 = n33447 ;
  assign y6993 = n33450 ;
  assign y6994 = ~n33453 ;
  assign y6995 = n33454 ;
  assign y6996 = n33455 ;
  assign y6997 = ~1'b0 ;
  assign y6998 = n33456 ;
  assign y6999 = ~n33462 ;
  assign y7000 = n33464 ;
  assign y7001 = ~n33465 ;
  assign y7002 = ~n33467 ;
  assign y7003 = ~n33469 ;
  assign y7004 = n33471 ;
  assign y7005 = ~n33472 ;
  assign y7006 = n33475 ;
  assign y7007 = n33476 ;
  assign y7008 = n33482 ;
  assign y7009 = ~n33488 ;
  assign y7010 = ~n33489 ;
  assign y7011 = ~n33493 ;
  assign y7012 = ~n33496 ;
  assign y7013 = n33505 ;
  assign y7014 = ~n33509 ;
  assign y7015 = ~n33510 ;
  assign y7016 = n33513 ;
  assign y7017 = ~n33515 ;
  assign y7018 = n33525 ;
  assign y7019 = ~n33528 ;
  assign y7020 = ~n33529 ;
  assign y7021 = n33534 ;
  assign y7022 = ~n33551 ;
  assign y7023 = ~n33553 ;
  assign y7024 = ~n726 ;
  assign y7025 = n33556 ;
  assign y7026 = n33562 ;
  assign y7027 = n33565 ;
  assign y7028 = ~n33569 ;
  assign y7029 = n33572 ;
  assign y7030 = ~n33575 ;
  assign y7031 = ~n33576 ;
  assign y7032 = n33581 ;
  assign y7033 = ~n33585 ;
  assign y7034 = n33586 ;
  assign y7035 = n33589 ;
  assign y7036 = ~n33597 ;
  assign y7037 = n33599 ;
  assign y7038 = ~n33603 ;
  assign y7039 = ~n33606 ;
  assign y7040 = ~n33607 ;
  assign y7041 = ~n33611 ;
  assign y7042 = ~n33618 ;
  assign y7043 = ~n33620 ;
  assign y7044 = ~n33625 ;
  assign y7045 = ~n33627 ;
  assign y7046 = ~n33630 ;
  assign y7047 = n33636 ;
  assign y7048 = ~n33637 ;
  assign y7049 = n33638 ;
  assign y7050 = n33639 ;
  assign y7051 = n33642 ;
  assign y7052 = n33646 ;
  assign y7053 = n33650 ;
  assign y7054 = n33652 ;
  assign y7055 = ~n33656 ;
  assign y7056 = n33660 ;
  assign y7057 = ~n33662 ;
  assign y7058 = ~n33669 ;
  assign y7059 = ~n33670 ;
  assign y7060 = ~n33677 ;
  assign y7061 = ~n33680 ;
  assign y7062 = n33681 ;
  assign y7063 = n33683 ;
  assign y7064 = n33684 ;
  assign y7065 = ~n33687 ;
  assign y7066 = ~n33696 ;
  assign y7067 = n33701 ;
  assign y7068 = ~n33705 ;
  assign y7069 = n33714 ;
  assign y7070 = n33715 ;
  assign y7071 = n33722 ;
  assign y7072 = n33723 ;
  assign y7073 = n33729 ;
  assign y7074 = n33733 ;
  assign y7075 = ~n33735 ;
  assign y7076 = n33737 ;
  assign y7077 = n33740 ;
  assign y7078 = ~n33744 ;
  assign y7079 = ~n33746 ;
  assign y7080 = n33747 ;
  assign y7081 = ~n33748 ;
  assign y7082 = ~n33749 ;
  assign y7083 = ~n33751 ;
  assign y7084 = ~n33754 ;
  assign y7085 = n33756 ;
  assign y7086 = ~n33758 ;
  assign y7087 = n33762 ;
  assign y7088 = ~n33763 ;
  assign y7089 = n33767 ;
  assign y7090 = n33776 ;
  assign y7091 = ~n33778 ;
  assign y7092 = n33779 ;
  assign y7093 = ~n33784 ;
  assign y7094 = n33787 ;
  assign y7095 = n33788 ;
  assign y7096 = ~n33789 ;
  assign y7097 = n33791 ;
  assign y7098 = n33794 ;
  assign y7099 = n33797 ;
  assign y7100 = n33799 ;
  assign y7101 = n33801 ;
  assign y7102 = n33804 ;
  assign y7103 = ~n33807 ;
  assign y7104 = ~n33808 ;
  assign y7105 = n33813 ;
  assign y7106 = n33814 ;
  assign y7107 = n33816 ;
  assign y7108 = ~n33817 ;
  assign y7109 = n33824 ;
  assign y7110 = n33830 ;
  assign y7111 = n33831 ;
  assign y7112 = n33833 ;
  assign y7113 = ~n33835 ;
  assign y7114 = n33836 ;
  assign y7115 = ~n33837 ;
  assign y7116 = ~n33839 ;
  assign y7117 = ~n33842 ;
  assign y7118 = ~n33844 ;
  assign y7119 = n33845 ;
  assign y7120 = n33854 ;
  assign y7121 = n33868 ;
  assign y7122 = ~n33872 ;
  assign y7123 = ~n33874 ;
  assign y7124 = n33878 ;
  assign y7125 = ~n33884 ;
  assign y7126 = ~n33885 ;
  assign y7127 = n8837 ;
  assign y7128 = ~n33887 ;
  assign y7129 = ~n33888 ;
  assign y7130 = n33891 ;
  assign y7131 = ~n33893 ;
  assign y7132 = n33895 ;
  assign y7133 = n33897 ;
  assign y7134 = ~1'b0 ;
  assign y7135 = ~n33900 ;
  assign y7136 = ~n33904 ;
  assign y7137 = n33909 ;
  assign y7138 = n33910 ;
  assign y7139 = n33913 ;
  assign y7140 = ~n33915 ;
  assign y7141 = n33917 ;
  assign y7142 = ~n33925 ;
  assign y7143 = n33928 ;
  assign y7144 = n33931 ;
  assign y7145 = ~n33938 ;
  assign y7146 = ~n33939 ;
  assign y7147 = ~n33948 ;
  assign y7148 = ~n33952 ;
  assign y7149 = n33954 ;
  assign y7150 = ~n33957 ;
  assign y7151 = n33960 ;
  assign y7152 = ~n33962 ;
  assign y7153 = ~n33964 ;
  assign y7154 = ~1'b0 ;
  assign y7155 = ~n33965 ;
  assign y7156 = n33969 ;
  assign y7157 = n33975 ;
  assign y7158 = ~n33977 ;
  assign y7159 = n33980 ;
  assign y7160 = n33986 ;
  assign y7161 = ~n33989 ;
  assign y7162 = ~n33993 ;
  assign y7163 = ~n33996 ;
  assign y7164 = ~n33997 ;
  assign y7165 = n33998 ;
  assign y7166 = ~n33999 ;
  assign y7167 = ~n34006 ;
  assign y7168 = ~n34007 ;
  assign y7169 = ~n34012 ;
  assign y7170 = n34013 ;
  assign y7171 = n34016 ;
  assign y7172 = n34020 ;
  assign y7173 = ~n34021 ;
  assign y7174 = n34023 ;
  assign y7175 = ~n34026 ;
  assign y7176 = n34027 ;
  assign y7177 = ~n34033 ;
  assign y7178 = ~n34034 ;
  assign y7179 = n34036 ;
  assign y7180 = ~n34038 ;
  assign y7181 = n34048 ;
  assign y7182 = ~n34053 ;
  assign y7183 = ~n34056 ;
  assign y7184 = n34058 ;
  assign y7185 = n34059 ;
  assign y7186 = ~n34060 ;
  assign y7187 = ~n34062 ;
  assign y7188 = ~n34065 ;
  assign y7189 = ~n34067 ;
  assign y7190 = ~n34073 ;
  assign y7191 = ~n34075 ;
  assign y7192 = ~n34077 ;
  assign y7193 = n34079 ;
  assign y7194 = n34083 ;
  assign y7195 = n34086 ;
  assign y7196 = ~1'b0 ;
  assign y7197 = ~n34091 ;
  assign y7198 = ~n34093 ;
  assign y7199 = n34098 ;
  assign y7200 = ~n34099 ;
  assign y7201 = n34100 ;
  assign y7202 = ~1'b0 ;
  assign y7203 = n34102 ;
  assign y7204 = ~n34108 ;
  assign y7205 = n34112 ;
  assign y7206 = n34114 ;
  assign y7207 = n34116 ;
  assign y7208 = ~n34118 ;
  assign y7209 = ~n34121 ;
  assign y7210 = ~n34123 ;
  assign y7211 = n34125 ;
  assign y7212 = n34126 ;
  assign y7213 = ~n34128 ;
  assign y7214 = ~n34129 ;
  assign y7215 = ~n34133 ;
  assign y7216 = ~n34134 ;
  assign y7217 = ~n34136 ;
  assign y7218 = n34138 ;
  assign y7219 = ~n34142 ;
  assign y7220 = n34144 ;
  assign y7221 = n34150 ;
  assign y7222 = ~n34152 ;
  assign y7223 = ~n18187 ;
  assign y7224 = ~n34161 ;
  assign y7225 = n34165 ;
  assign y7226 = ~n34167 ;
  assign y7227 = n34169 ;
  assign y7228 = ~n34172 ;
  assign y7229 = ~n34176 ;
  assign y7230 = n34180 ;
  assign y7231 = n34184 ;
  assign y7232 = ~n34188 ;
  assign y7233 = n34189 ;
  assign y7234 = n34194 ;
  assign y7235 = ~n34195 ;
  assign y7236 = ~n34197 ;
  assign y7237 = ~n34203 ;
  assign y7238 = ~n34208 ;
  assign y7239 = ~n34209 ;
  assign y7240 = ~n34212 ;
  assign y7241 = n34216 ;
  assign y7242 = n34224 ;
  assign y7243 = ~n34225 ;
  assign y7244 = ~n34231 ;
  assign y7245 = ~n34232 ;
  assign y7246 = ~n34237 ;
  assign y7247 = ~n34239 ;
  assign y7248 = ~n34246 ;
  assign y7249 = ~n34248 ;
  assign y7250 = n34250 ;
  assign y7251 = ~n34251 ;
  assign y7252 = n34252 ;
  assign y7253 = ~n34255 ;
  assign y7254 = n34259 ;
  assign y7255 = ~n34262 ;
  assign y7256 = n34266 ;
  assign y7257 = n34270 ;
  assign y7258 = n34272 ;
  assign y7259 = n34273 ;
  assign y7260 = ~n34276 ;
  assign y7261 = ~n34282 ;
  assign y7262 = ~n34292 ;
  assign y7263 = n34297 ;
  assign y7264 = ~n34299 ;
  assign y7265 = n34303 ;
  assign y7266 = ~n34304 ;
  assign y7267 = ~n34306 ;
  assign y7268 = ~n34312 ;
  assign y7269 = ~n34313 ;
  assign y7270 = n34317 ;
  assign y7271 = n34319 ;
  assign y7272 = ~n34320 ;
  assign y7273 = n34321 ;
  assign y7274 = n34327 ;
  assign y7275 = ~n34328 ;
  assign y7276 = n34332 ;
  assign y7277 = ~n34333 ;
  assign y7278 = ~n34341 ;
  assign y7279 = n34346 ;
  assign y7280 = ~n34351 ;
  assign y7281 = n34362 ;
  assign y7282 = ~n34363 ;
  assign y7283 = n34364 ;
  assign y7284 = ~n34365 ;
  assign y7285 = ~n34367 ;
  assign y7286 = ~n34376 ;
  assign y7287 = ~1'b0 ;
  assign y7288 = n34378 ;
  assign y7289 = ~n34381 ;
  assign y7290 = ~n34382 ;
  assign y7291 = n34384 ;
  assign y7292 = ~n34385 ;
  assign y7293 = ~n34387 ;
  assign y7294 = ~n34394 ;
  assign y7295 = ~1'b0 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = ~n34396 ;
  assign y7298 = ~n34398 ;
  assign y7299 = n34406 ;
  assign y7300 = n34410 ;
  assign y7301 = ~n34413 ;
  assign y7302 = n34416 ;
  assign y7303 = ~n34420 ;
  assign y7304 = n34424 ;
  assign y7305 = ~n34425 ;
  assign y7306 = ~n34430 ;
  assign y7307 = ~n34433 ;
  assign y7308 = ~n34434 ;
  assign y7309 = n34439 ;
  assign y7310 = ~n34440 ;
  assign y7311 = n34443 ;
  assign y7312 = n34445 ;
  assign y7313 = ~n34448 ;
  assign y7314 = ~n34449 ;
  assign y7315 = n34450 ;
  assign y7316 = ~n34455 ;
  assign y7317 = n34461 ;
  assign y7318 = ~n34463 ;
  assign y7319 = ~n34465 ;
  assign y7320 = n34466 ;
  assign y7321 = ~n34472 ;
  assign y7322 = ~n34474 ;
  assign y7323 = n34477 ;
  assign y7324 = ~n34479 ;
  assign y7325 = ~n34486 ;
  assign y7326 = n34490 ;
  assign y7327 = ~n34492 ;
  assign y7328 = n34493 ;
  assign y7329 = ~n34495 ;
  assign y7330 = n34496 ;
  assign y7331 = ~n34498 ;
  assign y7332 = ~n34507 ;
  assign y7333 = n34512 ;
  assign y7334 = n34513 ;
  assign y7335 = ~n34516 ;
  assign y7336 = n34521 ;
  assign y7337 = ~n34522 ;
  assign y7338 = n34524 ;
  assign y7339 = ~n34526 ;
  assign y7340 = ~n34530 ;
  assign y7341 = ~n34533 ;
  assign y7342 = ~n34538 ;
  assign y7343 = ~n34539 ;
  assign y7344 = n34542 ;
  assign y7345 = n34546 ;
  assign y7346 = n34549 ;
  assign y7347 = n34550 ;
  assign y7348 = ~n34559 ;
  assign y7349 = n34563 ;
  assign y7350 = ~n34564 ;
  assign y7351 = ~n34565 ;
  assign y7352 = n34570 ;
  assign y7353 = ~n34571 ;
  assign y7354 = ~1'b0 ;
  assign y7355 = ~1'b0 ;
  assign y7356 = n34573 ;
  assign y7357 = n34576 ;
  assign y7358 = n34579 ;
  assign y7359 = ~n34583 ;
  assign y7360 = n34586 ;
  assign y7361 = ~n34587 ;
  assign y7362 = ~n34593 ;
  assign y7363 = ~n34597 ;
  assign y7364 = ~n34601 ;
  assign y7365 = ~n34605 ;
  assign y7366 = n34607 ;
  assign y7367 = ~n34611 ;
  assign y7368 = ~n34613 ;
  assign y7369 = ~1'b0 ;
  assign y7370 = ~1'b0 ;
  assign y7371 = ~n34616 ;
  assign y7372 = ~n34619 ;
  assign y7373 = n34620 ;
  assign y7374 = n34622 ;
  assign y7375 = n34623 ;
  assign y7376 = n34627 ;
  assign y7377 = ~1'b0 ;
  assign y7378 = ~n34635 ;
  assign y7379 = ~n34639 ;
  assign y7380 = ~n34640 ;
  assign y7381 = ~n34642 ;
  assign y7382 = n34649 ;
  assign y7383 = n34653 ;
  assign y7384 = ~1'b0 ;
  assign y7385 = ~n34655 ;
  assign y7386 = ~n34657 ;
  assign y7387 = n34663 ;
  assign y7388 = ~n34671 ;
  assign y7389 = ~n34674 ;
  assign y7390 = n34677 ;
  assign y7391 = ~n34679 ;
  assign y7392 = ~n34680 ;
  assign y7393 = n34683 ;
  assign y7394 = n34687 ;
  assign y7395 = ~n34690 ;
  assign y7396 = n34694 ;
  assign y7397 = ~n34697 ;
  assign y7398 = ~n34700 ;
  assign y7399 = ~n34701 ;
  assign y7400 = n34702 ;
  assign y7401 = n34704 ;
  assign y7402 = ~n34706 ;
  assign y7403 = n34707 ;
  assign y7404 = ~n34708 ;
  assign y7405 = ~n34711 ;
  assign y7406 = ~n34713 ;
  assign y7407 = ~n34714 ;
  assign y7408 = ~n34718 ;
  assign y7409 = n34723 ;
  assign y7410 = ~n34725 ;
  assign y7411 = n34727 ;
  assign y7412 = n34730 ;
  assign y7413 = ~n34731 ;
  assign y7414 = ~n34735 ;
  assign y7415 = n34737 ;
  assign y7416 = n34738 ;
  assign y7417 = n34747 ;
  assign y7418 = ~n34752 ;
  assign y7419 = ~n34756 ;
  assign y7420 = ~n34762 ;
  assign y7421 = ~n11803 ;
  assign y7422 = ~n34764 ;
  assign y7423 = ~n34767 ;
  assign y7424 = n34769 ;
  assign y7425 = n34772 ;
  assign y7426 = n34777 ;
  assign y7427 = n34780 ;
  assign y7428 = ~n34781 ;
  assign y7429 = n34782 ;
  assign y7430 = ~n34789 ;
  assign y7431 = ~n34793 ;
  assign y7432 = n34795 ;
  assign y7433 = ~n34799 ;
  assign y7434 = ~n34803 ;
  assign y7435 = n34808 ;
  assign y7436 = ~n34809 ;
  assign y7437 = ~n34811 ;
  assign y7438 = ~n34814 ;
  assign y7439 = n34818 ;
  assign y7440 = ~n34819 ;
  assign y7441 = n34820 ;
  assign y7442 = n34821 ;
  assign y7443 = n34822 ;
  assign y7444 = ~n34828 ;
  assign y7445 = n34831 ;
  assign y7446 = ~n34833 ;
  assign y7447 = ~n34835 ;
  assign y7448 = ~n34837 ;
  assign y7449 = n34840 ;
  assign y7450 = n34852 ;
  assign y7451 = ~1'b0 ;
  assign y7452 = n34856 ;
  assign y7453 = n34857 ;
  assign y7454 = n34859 ;
  assign y7455 = ~n34863 ;
  assign y7456 = ~n34864 ;
  assign y7457 = n34866 ;
  assign y7458 = ~n34868 ;
  assign y7459 = ~n34870 ;
  assign y7460 = ~n34871 ;
  assign y7461 = n34873 ;
  assign y7462 = ~n34876 ;
  assign y7463 = n34878 ;
  assign y7464 = n34880 ;
  assign y7465 = ~n34890 ;
  assign y7466 = n34891 ;
  assign y7467 = ~1'b0 ;
  assign y7468 = n34895 ;
  assign y7469 = ~n34897 ;
  assign y7470 = n34898 ;
  assign y7471 = ~n34899 ;
  assign y7472 = n34902 ;
  assign y7473 = ~n34904 ;
  assign y7474 = n34906 ;
  assign y7475 = n34908 ;
  assign y7476 = ~n34911 ;
  assign y7477 = n34919 ;
  assign y7478 = n34922 ;
  assign y7479 = ~n34925 ;
  assign y7480 = n34926 ;
  assign y7481 = ~n34931 ;
  assign y7482 = ~n34932 ;
  assign y7483 = ~n34934 ;
  assign y7484 = ~n34938 ;
  assign y7485 = ~n34940 ;
  assign y7486 = ~n34945 ;
  assign y7487 = ~n34950 ;
  assign y7488 = n34951 ;
  assign y7489 = n34953 ;
  assign y7490 = ~n34958 ;
  assign y7491 = n34959 ;
  assign y7492 = ~1'b0 ;
  assign y7493 = ~n34961 ;
  assign y7494 = ~n34964 ;
  assign y7495 = ~n34966 ;
  assign y7496 = ~n34967 ;
  assign y7497 = ~n34970 ;
  assign y7498 = ~n34974 ;
  assign y7499 = n34976 ;
  assign y7500 = n34978 ;
  assign y7501 = ~n34980 ;
  assign y7502 = n34982 ;
  assign y7503 = n34983 ;
  assign y7504 = ~n34992 ;
  assign y7505 = n34999 ;
  assign y7506 = n35005 ;
  assign y7507 = ~n35007 ;
  assign y7508 = n35008 ;
  assign y7509 = n35009 ;
  assign y7510 = n35011 ;
  assign y7511 = n35014 ;
  assign y7512 = ~n35017 ;
  assign y7513 = n35018 ;
  assign y7514 = n35022 ;
  assign y7515 = ~n35023 ;
  assign y7516 = ~n35024 ;
  assign y7517 = n35025 ;
  assign y7518 = n35032 ;
  assign y7519 = ~n35035 ;
  assign y7520 = ~1'b0 ;
  assign y7521 = n35037 ;
  assign y7522 = ~n35041 ;
  assign y7523 = ~n21550 ;
  assign y7524 = n35046 ;
  assign y7525 = n35049 ;
  assign y7526 = n35050 ;
  assign y7527 = ~n35051 ;
  assign y7528 = n35053 ;
  assign y7529 = ~n35055 ;
  assign y7530 = n35056 ;
  assign y7531 = n35058 ;
  assign y7532 = n35061 ;
  assign y7533 = n35064 ;
  assign y7534 = n35067 ;
  assign y7535 = n35068 ;
  assign y7536 = ~1'b0 ;
  assign y7537 = n35072 ;
  assign y7538 = n35074 ;
  assign y7539 = ~n35076 ;
  assign y7540 = n35078 ;
  assign y7541 = n35080 ;
  assign y7542 = n35081 ;
  assign y7543 = n35083 ;
  assign y7544 = ~n35088 ;
  assign y7545 = ~n35089 ;
  assign y7546 = ~n35091 ;
  assign y7547 = ~n35095 ;
  assign y7548 = ~n35098 ;
  assign y7549 = n35101 ;
  assign y7550 = n35103 ;
  assign y7551 = ~n35110 ;
  assign y7552 = ~n35113 ;
  assign y7553 = n35114 ;
  assign y7554 = ~n35117 ;
  assign y7555 = ~n35118 ;
  assign y7556 = ~n35120 ;
  assign y7557 = ~n35124 ;
  assign y7558 = ~n35125 ;
  assign y7559 = ~n35127 ;
  assign y7560 = n35129 ;
  assign y7561 = ~n35131 ;
  assign y7562 = n35133 ;
  assign y7563 = n35139 ;
  assign y7564 = ~1'b0 ;
  assign y7565 = n35141 ;
  assign y7566 = ~n35143 ;
  assign y7567 = n35147 ;
  assign y7568 = n35148 ;
  assign y7569 = ~n35149 ;
  assign y7570 = n35150 ;
  assign y7571 = n35152 ;
  assign y7572 = n35154 ;
  assign y7573 = ~n35158 ;
  assign y7574 = ~n35159 ;
  assign y7575 = ~n35162 ;
  assign y7576 = ~n7851 ;
  assign y7577 = n35171 ;
  assign y7578 = n35172 ;
  assign y7579 = ~n35173 ;
  assign y7580 = n35174 ;
  assign y7581 = ~n35176 ;
  assign y7582 = ~n35178 ;
  assign y7583 = n35181 ;
  assign y7584 = n35185 ;
  assign y7585 = n35189 ;
  assign y7586 = n35191 ;
  assign y7587 = n35194 ;
  assign y7588 = n35196 ;
  assign y7589 = n35197 ;
  assign y7590 = n35198 ;
  assign y7591 = n35200 ;
  assign y7592 = ~n35204 ;
  assign y7593 = ~n35206 ;
  assign y7594 = n35214 ;
  assign y7595 = ~n35215 ;
  assign y7596 = n35217 ;
  assign y7597 = n35220 ;
  assign y7598 = n35224 ;
  assign y7599 = n35226 ;
  assign y7600 = ~n35229 ;
  assign y7601 = n35233 ;
  assign y7602 = ~n35234 ;
  assign y7603 = ~n35238 ;
  assign y7604 = ~n35240 ;
  assign y7605 = n35242 ;
  assign y7606 = n35243 ;
  assign y7607 = ~n35246 ;
  assign y7608 = ~n35248 ;
  assign y7609 = ~n35252 ;
  assign y7610 = ~n35257 ;
  assign y7611 = n35258 ;
  assign y7612 = ~n35259 ;
  assign y7613 = ~n35262 ;
  assign y7614 = n35270 ;
  assign y7615 = ~n35274 ;
  assign y7616 = n35277 ;
  assign y7617 = ~n35278 ;
  assign y7618 = ~1'b0 ;
  assign y7619 = ~1'b0 ;
  assign y7620 = n35284 ;
  assign y7621 = ~n35285 ;
  assign y7622 = n35287 ;
  assign y7623 = n35294 ;
  assign y7624 = n35296 ;
  assign y7625 = ~n35301 ;
  assign y7626 = ~1'b0 ;
  assign y7627 = ~n35305 ;
  assign y7628 = n35308 ;
  assign y7629 = ~n35320 ;
  assign y7630 = ~n35322 ;
  assign y7631 = ~n35324 ;
  assign y7632 = ~n35328 ;
  assign y7633 = ~n35336 ;
  assign y7634 = n35338 ;
  assign y7635 = ~n35342 ;
  assign y7636 = n35345 ;
  assign y7637 = ~n35346 ;
  assign y7638 = ~n35348 ;
  assign y7639 = ~n35351 ;
  assign y7640 = ~1'b0 ;
  assign y7641 = n35352 ;
  assign y7642 = ~n35353 ;
  assign y7643 = n35354 ;
  assign y7644 = n35357 ;
  assign y7645 = n35360 ;
  assign y7646 = n35361 ;
  assign y7647 = ~n35363 ;
  assign y7648 = n35365 ;
  assign y7649 = ~n35366 ;
  assign y7650 = ~n35367 ;
  assign y7651 = n35374 ;
  assign y7652 = ~n35376 ;
  assign y7653 = ~n35385 ;
  assign y7654 = n35387 ;
  assign y7655 = n35388 ;
  assign y7656 = ~n35392 ;
  assign y7657 = ~n35395 ;
  assign y7658 = n35397 ;
  assign y7659 = n35402 ;
  assign y7660 = ~n35405 ;
  assign y7661 = n35407 ;
  assign y7662 = n35412 ;
  assign y7663 = ~n35414 ;
  assign y7664 = n35416 ;
  assign y7665 = ~n35418 ;
  assign y7666 = ~n35421 ;
  assign y7667 = ~n35427 ;
  assign y7668 = ~n35429 ;
  assign y7669 = ~n35436 ;
  assign y7670 = ~n35441 ;
  assign y7671 = n35446 ;
  assign y7672 = n35450 ;
  assign y7673 = ~n35453 ;
  assign y7674 = ~n35463 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~n35466 ;
  assign y7677 = ~n35470 ;
  assign y7678 = n35471 ;
  assign y7679 = ~n35473 ;
  assign y7680 = ~n35479 ;
  assign y7681 = n35483 ;
  assign y7682 = n35486 ;
  assign y7683 = ~n35487 ;
  assign y7684 = ~n35490 ;
  assign y7685 = n35493 ;
  assign y7686 = n35495 ;
  assign y7687 = ~n35497 ;
  assign y7688 = n35498 ;
  assign y7689 = ~n35507 ;
  assign y7690 = n35515 ;
  assign y7691 = n35516 ;
  assign y7692 = ~n35517 ;
  assign y7693 = n35521 ;
  assign y7694 = ~n35532 ;
  assign y7695 = ~n35535 ;
  assign y7696 = n35539 ;
  assign y7697 = ~n35545 ;
  assign y7698 = n35548 ;
  assign y7699 = ~n35550 ;
  assign y7700 = n35552 ;
  assign y7701 = ~n35557 ;
  assign y7702 = ~n35561 ;
  assign y7703 = n35564 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = ~n35567 ;
  assign y7706 = n35572 ;
  assign y7707 = ~n35574 ;
  assign y7708 = ~n35578 ;
  assign y7709 = ~n35581 ;
  assign y7710 = n35582 ;
  assign y7711 = n35597 ;
  assign y7712 = ~n35598 ;
  assign y7713 = ~n35599 ;
  assign y7714 = n35602 ;
  assign y7715 = n35611 ;
  assign y7716 = ~1'b0 ;
  assign y7717 = n35612 ;
  assign y7718 = n35615 ;
  assign y7719 = ~n35617 ;
  assign y7720 = ~n35618 ;
  assign y7721 = n35621 ;
  assign y7722 = ~n35624 ;
  assign y7723 = ~n35625 ;
  assign y7724 = n35626 ;
  assign y7725 = ~n35628 ;
  assign y7726 = ~n35629 ;
  assign y7727 = ~n35632 ;
  assign y7728 = n35636 ;
  assign y7729 = ~n35641 ;
  assign y7730 = ~n35644 ;
  assign y7731 = n35647 ;
  assign y7732 = ~n35654 ;
  assign y7733 = ~n35661 ;
  assign y7734 = ~n35667 ;
  assign y7735 = ~n35671 ;
  assign y7736 = n35673 ;
  assign y7737 = ~n35674 ;
  assign y7738 = n35676 ;
  assign y7739 = n35680 ;
  assign y7740 = ~n35683 ;
  assign y7741 = n35686 ;
  assign y7742 = n35687 ;
  assign y7743 = ~n35689 ;
  assign y7744 = ~n35692 ;
  assign y7745 = n35699 ;
  assign y7746 = n35704 ;
  assign y7747 = ~n35705 ;
  assign y7748 = ~n35710 ;
  assign y7749 = n35713 ;
  assign y7750 = n35718 ;
  assign y7751 = n35720 ;
  assign y7752 = n35723 ;
  assign y7753 = ~n35730 ;
  assign y7754 = n35734 ;
  assign y7755 = n35737 ;
  assign y7756 = ~1'b0 ;
  assign y7757 = ~n35743 ;
  assign y7758 = ~n35748 ;
  assign y7759 = n35749 ;
  assign y7760 = ~1'b0 ;
  assign y7761 = n35752 ;
  assign y7762 = n35754 ;
  assign y7763 = n35757 ;
  assign y7764 = n35759 ;
  assign y7765 = ~n35763 ;
  assign y7766 = ~n35765 ;
  assign y7767 = n35767 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = ~n35776 ;
  assign y7770 = ~n35783 ;
  assign y7771 = n35785 ;
  assign y7772 = n35788 ;
  assign y7773 = ~n35790 ;
  assign y7774 = n35794 ;
  assign y7775 = ~n35796 ;
  assign y7776 = ~n35799 ;
  assign y7777 = n35801 ;
  assign y7778 = ~n35805 ;
  assign y7779 = ~n35810 ;
  assign y7780 = n35813 ;
  assign y7781 = n35817 ;
  assign y7782 = ~n35820 ;
  assign y7783 = n35821 ;
  assign y7784 = ~n35822 ;
  assign y7785 = ~n35831 ;
  assign y7786 = n35833 ;
  assign y7787 = n35836 ;
  assign y7788 = n35837 ;
  assign y7789 = n35844 ;
  assign y7790 = n35845 ;
  assign y7791 = n35856 ;
  assign y7792 = n35858 ;
  assign y7793 = n35859 ;
  assign y7794 = ~1'b0 ;
  assign y7795 = ~n35862 ;
  assign y7796 = ~n35863 ;
  assign y7797 = ~n35864 ;
  assign y7798 = ~n35869 ;
  assign y7799 = n35878 ;
  assign y7800 = ~n35879 ;
  assign y7801 = ~n35882 ;
  assign y7802 = ~n35885 ;
  assign y7803 = ~n35886 ;
  assign y7804 = n35887 ;
  assign y7805 = ~1'b0 ;
  assign y7806 = n35893 ;
  assign y7807 = ~n35895 ;
  assign y7808 = n35897 ;
  assign y7809 = ~n35899 ;
  assign y7810 = n35900 ;
  assign y7811 = ~n35901 ;
  assign y7812 = n35904 ;
  assign y7813 = ~n35905 ;
  assign y7814 = ~n35909 ;
  assign y7815 = n35916 ;
  assign y7816 = ~n35919 ;
  assign y7817 = ~n35921 ;
  assign y7818 = n35923 ;
  assign y7819 = ~n35925 ;
  assign y7820 = n35927 ;
  assign y7821 = n35931 ;
  assign y7822 = ~n35934 ;
  assign y7823 = n35935 ;
  assign y7824 = n35948 ;
  assign y7825 = ~n35951 ;
  assign y7826 = ~n35952 ;
  assign y7827 = ~1'b0 ;
  assign y7828 = n35953 ;
  assign y7829 = n35957 ;
  assign y7830 = n35961 ;
  assign y7831 = n35965 ;
  assign y7832 = ~n35968 ;
  assign y7833 = ~n35975 ;
  assign y7834 = ~n35977 ;
  assign y7835 = n35981 ;
  assign y7836 = n35983 ;
  assign y7837 = n35984 ;
  assign y7838 = ~n35992 ;
  assign y7839 = n35999 ;
  assign y7840 = ~n36003 ;
  assign y7841 = ~n36007 ;
  assign y7842 = n36008 ;
  assign y7843 = n36010 ;
  assign y7844 = n36012 ;
  assign y7845 = ~n36020 ;
  assign y7846 = ~1'b0 ;
  assign y7847 = ~n36024 ;
  assign y7848 = n36025 ;
  assign y7849 = ~n36031 ;
  assign y7850 = n36037 ;
  assign y7851 = ~n36041 ;
  assign y7852 = n9002 ;
  assign y7853 = n36042 ;
  assign y7854 = n36043 ;
  assign y7855 = n36047 ;
  assign y7856 = n36049 ;
  assign y7857 = ~n36050 ;
  assign y7858 = ~n36052 ;
  assign y7859 = n36053 ;
  assign y7860 = ~n36055 ;
  assign y7861 = ~n36060 ;
  assign y7862 = ~n36064 ;
  assign y7863 = n36069 ;
  assign y7864 = ~n36070 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = n36071 ;
  assign y7867 = ~n36072 ;
  assign y7868 = ~n36073 ;
  assign y7869 = n36076 ;
  assign y7870 = n36077 ;
  assign y7871 = ~n36078 ;
  assign y7872 = ~1'b0 ;
  assign y7873 = n36081 ;
  assign y7874 = ~n36084 ;
  assign y7875 = ~n36089 ;
  assign y7876 = n36094 ;
  assign y7877 = n36098 ;
  assign y7878 = n36101 ;
  assign y7879 = n36103 ;
  assign y7880 = n36108 ;
  assign y7881 = n36111 ;
  assign y7882 = ~n36113 ;
  assign y7883 = ~n36114 ;
  assign y7884 = n36116 ;
  assign y7885 = n36117 ;
  assign y7886 = n36118 ;
  assign y7887 = ~n36119 ;
  assign y7888 = ~n36121 ;
  assign y7889 = n36128 ;
  assign y7890 = n36130 ;
  assign y7891 = n36141 ;
  assign y7892 = ~1'b0 ;
  assign y7893 = n36143 ;
  assign y7894 = ~n36146 ;
  assign y7895 = ~n36151 ;
  assign y7896 = n36156 ;
  assign y7897 = ~n36157 ;
  assign y7898 = ~n36160 ;
  assign y7899 = n36167 ;
  assign y7900 = n36169 ;
  assign y7901 = ~n36178 ;
  assign y7902 = ~n36183 ;
  assign y7903 = n36184 ;
  assign y7904 = n36185 ;
  assign y7905 = n36186 ;
  assign y7906 = n36187 ;
  assign y7907 = n36189 ;
  assign y7908 = ~n36190 ;
  assign y7909 = ~n36194 ;
  assign y7910 = ~n36199 ;
  assign y7911 = ~n36200 ;
  assign y7912 = ~1'b0 ;
  assign y7913 = ~n36204 ;
  assign y7914 = n36205 ;
  assign y7915 = ~n36210 ;
  assign y7916 = n36211 ;
  assign y7917 = n36213 ;
  assign y7918 = ~n36215 ;
  assign y7919 = ~n36216 ;
  assign y7920 = n36217 ;
  assign y7921 = ~n36220 ;
  assign y7922 = ~n36223 ;
  assign y7923 = ~n36226 ;
  assign y7924 = n36228 ;
  assign y7925 = n36230 ;
  assign y7926 = n36231 ;
  assign y7927 = n36236 ;
  assign y7928 = n36237 ;
  assign y7929 = n36242 ;
  assign y7930 = n36243 ;
  assign y7931 = ~n36244 ;
  assign y7932 = ~n36247 ;
  assign y7933 = ~1'b0 ;
  assign y7934 = n36248 ;
  assign y7935 = n36251 ;
  assign y7936 = n36254 ;
  assign y7937 = ~1'b0 ;
  assign y7938 = n36256 ;
  assign y7939 = ~n36258 ;
  assign y7940 = ~n36259 ;
  assign y7941 = n36260 ;
  assign y7942 = n36261 ;
  assign y7943 = ~n36266 ;
  assign y7944 = ~1'b0 ;
  assign y7945 = n36272 ;
  assign y7946 = ~n36273 ;
  assign y7947 = n36276 ;
  assign y7948 = n36281 ;
  assign y7949 = n36287 ;
  assign y7950 = ~n36289 ;
  assign y7951 = n36292 ;
  assign y7952 = n36293 ;
  assign y7953 = ~n36294 ;
  assign y7954 = ~n36297 ;
  assign y7955 = ~n36298 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = n36300 ;
  assign y7958 = ~n36301 ;
  assign y7959 = ~n36308 ;
  assign y7960 = ~n36314 ;
  assign y7961 = ~n36317 ;
  assign y7962 = n36322 ;
  assign y7963 = ~1'b0 ;
  assign y7964 = ~n36323 ;
  assign y7965 = n36325 ;
  assign y7966 = n36326 ;
  assign y7967 = ~n36328 ;
  assign y7968 = n36332 ;
  assign y7969 = n36341 ;
  assign y7970 = ~n36343 ;
  assign y7971 = ~n36346 ;
  assign y7972 = n36348 ;
  assign y7973 = ~n36349 ;
  assign y7974 = n36353 ;
  assign y7975 = ~n36361 ;
  assign y7976 = n36362 ;
  assign y7977 = ~n36370 ;
  assign y7978 = ~n36371 ;
  assign y7979 = ~n36379 ;
  assign y7980 = n36385 ;
  assign y7981 = ~n36387 ;
  assign y7982 = n36391 ;
  assign y7983 = n36394 ;
  assign y7984 = ~n36398 ;
  assign y7985 = ~n36401 ;
  assign y7986 = ~n36408 ;
  assign y7987 = ~n36409 ;
  assign y7988 = ~1'b0 ;
  assign y7989 = ~1'b0 ;
  assign y7990 = ~n36410 ;
  assign y7991 = ~n36412 ;
  assign y7992 = n36416 ;
  assign y7993 = ~n36417 ;
  assign y7994 = ~n36419 ;
  assign y7995 = ~n36421 ;
  assign y7996 = n36424 ;
  assign y7997 = n36427 ;
  assign y7998 = ~n36430 ;
  assign y7999 = ~n36435 ;
  assign y8000 = ~n36437 ;
  assign y8001 = n36443 ;
  assign y8002 = ~n36444 ;
  assign y8003 = n36448 ;
  assign y8004 = n36449 ;
  assign y8005 = ~n36452 ;
  assign y8006 = n36455 ;
  assign y8007 = n36457 ;
  assign y8008 = n36460 ;
  assign y8009 = ~n36464 ;
  assign y8010 = n36466 ;
  assign y8011 = n36469 ;
  assign y8012 = n36473 ;
  assign y8013 = ~n36476 ;
  assign y8014 = n36477 ;
  assign y8015 = n36482 ;
  assign y8016 = ~n36483 ;
  assign y8017 = ~n36485 ;
  assign y8018 = n36487 ;
  assign y8019 = ~n36493 ;
  assign y8020 = ~n36499 ;
  assign y8021 = ~n36500 ;
  assign y8022 = n36503 ;
  assign y8023 = n36506 ;
  assign y8024 = n36507 ;
  assign y8025 = n36515 ;
  assign y8026 = n36517 ;
  assign y8027 = ~n36518 ;
  assign y8028 = n36520 ;
  assign y8029 = ~n36521 ;
  assign y8030 = ~n36527 ;
  assign y8031 = n36529 ;
  assign y8032 = n36533 ;
  assign y8033 = n36535 ;
  assign y8034 = ~n36539 ;
  assign y8035 = ~n36540 ;
  assign y8036 = n36542 ;
  assign y8037 = ~n36545 ;
  assign y8038 = ~n36549 ;
  assign y8039 = n36554 ;
  assign y8040 = ~n36555 ;
  assign y8041 = ~n36558 ;
  assign y8042 = n36560 ;
  assign y8043 = n36563 ;
  assign y8044 = n36564 ;
  assign y8045 = ~n36565 ;
  assign y8046 = n36568 ;
  assign y8047 = n36571 ;
  assign y8048 = ~1'b0 ;
  assign y8049 = ~1'b0 ;
  assign y8050 = n36572 ;
  assign y8051 = ~n36576 ;
  assign y8052 = ~n36582 ;
  assign y8053 = ~n36584 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = ~1'b0 ;
  assign y8056 = ~n36585 ;
  assign y8057 = ~n36586 ;
  assign y8058 = n36593 ;
  assign y8059 = ~n36599 ;
  assign y8060 = n36601 ;
  assign y8061 = n36603 ;
  assign y8062 = ~n36607 ;
  assign y8063 = n36612 ;
  assign y8064 = n36613 ;
  assign y8065 = ~n36618 ;
  assign y8066 = n36619 ;
  assign y8067 = n36620 ;
  assign y8068 = ~n36624 ;
  assign y8069 = ~n36627 ;
  assign y8070 = n36628 ;
  assign y8071 = ~n36631 ;
  assign y8072 = ~n36633 ;
  assign y8073 = ~n36634 ;
  assign y8074 = ~n36638 ;
  assign y8075 = ~n36639 ;
  assign y8076 = n36642 ;
  assign y8077 = ~n36645 ;
  assign y8078 = n36649 ;
  assign y8079 = ~n36651 ;
  assign y8080 = ~1'b0 ;
  assign y8081 = ~n36652 ;
  assign y8082 = ~n36654 ;
  assign y8083 = n36655 ;
  assign y8084 = n36659 ;
  assign y8085 = ~n36661 ;
  assign y8086 = ~n36664 ;
  assign y8087 = ~n36667 ;
  assign y8088 = ~1'b0 ;
  assign y8089 = n36673 ;
  assign y8090 = ~n36677 ;
  assign y8091 = n36678 ;
  assign y8092 = ~n36682 ;
  assign y8093 = ~n36685 ;
  assign y8094 = ~n36688 ;
  assign y8095 = n36689 ;
  assign y8096 = ~n36692 ;
  assign y8097 = ~n36693 ;
  assign y8098 = ~1'b0 ;
  assign y8099 = ~n36694 ;
  assign y8100 = n36695 ;
  assign y8101 = n36698 ;
  assign y8102 = n36700 ;
  assign y8103 = n36702 ;
  assign y8104 = n36707 ;
  assign y8105 = ~n36708 ;
  assign y8106 = n36711 ;
  assign y8107 = ~n36718 ;
  assign y8108 = n36725 ;
  assign y8109 = n36726 ;
  assign y8110 = ~n36727 ;
  assign y8111 = n36729 ;
  assign y8112 = n36731 ;
  assign y8113 = n36733 ;
  assign y8114 = n36735 ;
  assign y8115 = n36736 ;
  assign y8116 = n36743 ;
  assign y8117 = ~n36744 ;
  assign y8118 = ~n36746 ;
  assign y8119 = n36747 ;
  assign y8120 = n36755 ;
  assign y8121 = n36762 ;
  assign y8122 = ~n36763 ;
  assign y8123 = ~n36767 ;
  assign y8124 = n36770 ;
  assign y8125 = n36775 ;
  assign y8126 = n36778 ;
  assign y8127 = n36785 ;
  assign y8128 = n36787 ;
  assign y8129 = ~n36788 ;
  assign y8130 = n36794 ;
  assign y8131 = n36796 ;
  assign y8132 = n36797 ;
  assign y8133 = ~n36798 ;
  assign y8134 = n36802 ;
  assign y8135 = n36805 ;
  assign y8136 = ~n36808 ;
  assign y8137 = ~n36810 ;
  assign y8138 = ~n36811 ;
  assign y8139 = ~n36812 ;
  assign y8140 = ~n36815 ;
  assign y8141 = n36818 ;
  assign y8142 = ~n36819 ;
  assign y8143 = ~n36825 ;
  assign y8144 = ~n36826 ;
  assign y8145 = ~n36834 ;
  assign y8146 = ~n36837 ;
  assign y8147 = ~n36839 ;
  assign y8148 = ~n36841 ;
  assign y8149 = ~n36842 ;
  assign y8150 = n36844 ;
  assign y8151 = ~n36849 ;
  assign y8152 = n36851 ;
  assign y8153 = ~n36854 ;
  assign y8154 = n36855 ;
  assign y8155 = n36858 ;
  assign y8156 = n36862 ;
  assign y8157 = n36869 ;
  assign y8158 = n36873 ;
  assign y8159 = ~n36877 ;
  assign y8160 = n36879 ;
  assign y8161 = ~n36880 ;
  assign y8162 = n36882 ;
  assign y8163 = ~n36887 ;
  assign y8164 = n36888 ;
  assign y8165 = ~n36889 ;
  assign y8166 = ~n36890 ;
  assign y8167 = ~n36893 ;
  assign y8168 = ~n36899 ;
  assign y8169 = ~n36900 ;
  assign y8170 = ~n36902 ;
  assign y8171 = n36903 ;
  assign y8172 = n36910 ;
  assign y8173 = n36912 ;
  assign y8174 = ~n36915 ;
  assign y8175 = ~1'b0 ;
  assign y8176 = ~n36923 ;
  assign y8177 = ~n36927 ;
  assign y8178 = n36933 ;
  assign y8179 = ~n36935 ;
  assign y8180 = ~n36939 ;
  assign y8181 = n36940 ;
  assign y8182 = n36946 ;
  assign y8183 = n36955 ;
  assign y8184 = n36960 ;
  assign y8185 = ~n36963 ;
  assign y8186 = n36966 ;
  assign y8187 = ~n36967 ;
  assign y8188 = ~n36969 ;
  assign y8189 = n36973 ;
  assign y8190 = ~n36975 ;
  assign y8191 = n36976 ;
  assign y8192 = n36977 ;
  assign y8193 = ~n36978 ;
  assign y8194 = n36980 ;
  assign y8195 = ~n36983 ;
  assign y8196 = ~1'b0 ;
  assign y8197 = n36984 ;
  assign y8198 = n36990 ;
  assign y8199 = n36998 ;
  assign y8200 = ~n37000 ;
  assign y8201 = ~n37006 ;
  assign y8202 = n37007 ;
  assign y8203 = ~n37012 ;
  assign y8204 = ~n37013 ;
  assign y8205 = ~n37016 ;
  assign y8206 = n37018 ;
  assign y8207 = ~n37024 ;
  assign y8208 = n37027 ;
  assign y8209 = n37030 ;
  assign y8210 = n37031 ;
  assign y8211 = ~n37034 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~n37036 ;
  assign y8214 = n37038 ;
  assign y8215 = n37039 ;
  assign y8216 = ~n37040 ;
  assign y8217 = n37045 ;
  assign y8218 = ~n37046 ;
  assign y8219 = ~n37047 ;
  assign y8220 = ~1'b0 ;
  assign y8221 = n37050 ;
  assign y8222 = ~n37052 ;
  assign y8223 = n37053 ;
  assign y8224 = ~n37054 ;
  assign y8225 = n37057 ;
  assign y8226 = ~n37060 ;
  assign y8227 = n37062 ;
  assign y8228 = ~1'b0 ;
  assign y8229 = n37064 ;
  assign y8230 = n37066 ;
  assign y8231 = n37069 ;
  assign y8232 = n37070 ;
  assign y8233 = n37076 ;
  assign y8234 = n37082 ;
  assign y8235 = n37089 ;
  assign y8236 = n37091 ;
  assign y8237 = ~n37092 ;
  assign y8238 = ~n37094 ;
  assign y8239 = ~n29547 ;
  assign y8240 = ~n37096 ;
  assign y8241 = n37103 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = n37105 ;
  assign y8244 = n37109 ;
  assign y8245 = n37112 ;
  assign y8246 = ~n37113 ;
  assign y8247 = ~n37116 ;
  assign y8248 = ~n37117 ;
  assign y8249 = n37118 ;
  assign y8250 = ~n37125 ;
  assign y8251 = n37127 ;
  assign y8252 = ~n37130 ;
  assign y8253 = n37131 ;
  assign y8254 = ~n37133 ;
  assign y8255 = ~n37139 ;
  assign y8256 = n37144 ;
  assign y8257 = n37145 ;
  assign y8258 = ~n37147 ;
  assign y8259 = ~n37148 ;
  assign y8260 = ~n37150 ;
  assign y8261 = ~1'b0 ;
  assign y8262 = n37152 ;
  assign y8263 = ~n37154 ;
  assign y8264 = n37155 ;
  assign y8265 = ~n37156 ;
  assign y8266 = n37157 ;
  assign y8267 = n37162 ;
  assign y8268 = n37164 ;
  assign y8269 = n37172 ;
  assign y8270 = ~n37177 ;
  assign y8271 = n37178 ;
  assign y8272 = n37181 ;
  assign y8273 = n37183 ;
  assign y8274 = ~n37184 ;
  assign y8275 = ~n37185 ;
  assign y8276 = ~n37188 ;
  assign y8277 = ~n37190 ;
  assign y8278 = ~n37192 ;
  assign y8279 = ~n37195 ;
  assign y8280 = ~n37197 ;
  assign y8281 = n37200 ;
  assign y8282 = n37201 ;
  assign y8283 = n37203 ;
  assign y8284 = ~n37205 ;
  assign y8285 = n37208 ;
  assign y8286 = ~n37210 ;
  assign y8287 = n37216 ;
  assign y8288 = n37220 ;
  assign y8289 = ~n37223 ;
  assign y8290 = ~n37226 ;
  assign y8291 = ~n37228 ;
  assign y8292 = n37230 ;
  assign y8293 = ~n37234 ;
  assign y8294 = n37235 ;
  assign y8295 = n37238 ;
  assign y8296 = ~n37239 ;
  assign y8297 = ~n37242 ;
  assign y8298 = ~n37244 ;
  assign y8299 = n37248 ;
  assign y8300 = n37251 ;
  assign y8301 = ~n37252 ;
  assign y8302 = n37254 ;
  assign y8303 = n37257 ;
  assign y8304 = ~n37258 ;
  assign y8305 = ~n37259 ;
  assign y8306 = n37266 ;
  assign y8307 = n37267 ;
  assign y8308 = ~n37270 ;
  assign y8309 = ~n37272 ;
  assign y8310 = n37273 ;
  assign y8311 = ~n37275 ;
  assign y8312 = ~n37278 ;
  assign y8313 = ~n37279 ;
  assign y8314 = ~n37283 ;
  assign y8315 = ~n37287 ;
  assign y8316 = n37289 ;
  assign y8317 = n37290 ;
  assign y8318 = n37295 ;
  assign y8319 = ~n37296 ;
  assign y8320 = n37297 ;
  assign y8321 = ~n37302 ;
  assign y8322 = n37304 ;
  assign y8323 = ~n37309 ;
  assign y8324 = n37316 ;
  assign y8325 = n37319 ;
  assign y8326 = ~n37321 ;
  assign y8327 = ~n37322 ;
  assign y8328 = ~n37324 ;
  assign y8329 = n37331 ;
  assign y8330 = ~n37335 ;
  assign y8331 = n37336 ;
  assign y8332 = ~n37337 ;
  assign y8333 = n37339 ;
  assign y8334 = n37343 ;
  assign y8335 = ~n37344 ;
  assign y8336 = ~n37345 ;
  assign y8337 = ~n37349 ;
  assign y8338 = ~1'b0 ;
  assign y8339 = n37350 ;
  assign y8340 = ~n37352 ;
  assign y8341 = n37356 ;
  assign y8342 = ~n37360 ;
  assign y8343 = n37362 ;
  assign y8344 = ~n37365 ;
  assign y8345 = ~n37367 ;
  assign y8346 = ~n37368 ;
  assign y8347 = n37376 ;
  assign y8348 = ~n37377 ;
  assign y8349 = ~n37379 ;
  assign y8350 = ~n37386 ;
  assign y8351 = ~n37388 ;
  assign y8352 = ~n37391 ;
  assign y8353 = ~n37393 ;
  assign y8354 = ~n37395 ;
  assign y8355 = ~n37396 ;
  assign y8356 = ~n37397 ;
  assign y8357 = n37398 ;
  assign y8358 = ~n37400 ;
  assign y8359 = n37403 ;
  assign y8360 = n37408 ;
  assign y8361 = ~n37409 ;
  assign y8362 = ~n37410 ;
  assign y8363 = ~n37411 ;
  assign y8364 = ~n37414 ;
  assign y8365 = ~n37417 ;
  assign y8366 = n37420 ;
  assign y8367 = ~1'b0 ;
  assign y8368 = ~n37424 ;
  assign y8369 = n37428 ;
  assign y8370 = n37430 ;
  assign y8371 = n37434 ;
  assign y8372 = n37437 ;
  assign y8373 = ~n37440 ;
  assign y8374 = n37441 ;
  assign y8375 = ~n37446 ;
  assign y8376 = ~n37448 ;
  assign y8377 = ~n37451 ;
  assign y8378 = ~n37453 ;
  assign y8379 = ~n37461 ;
  assign y8380 = n37464 ;
  assign y8381 = ~n37466 ;
  assign y8382 = ~n37467 ;
  assign y8383 = ~n37469 ;
  assign y8384 = n37472 ;
  assign y8385 = n37479 ;
  assign y8386 = n37480 ;
  assign y8387 = n37481 ;
  assign y8388 = ~1'b0 ;
  assign y8389 = n37483 ;
  assign y8390 = ~n37484 ;
  assign y8391 = ~n37491 ;
  assign y8392 = ~n37493 ;
  assign y8393 = n37498 ;
  assign y8394 = n37501 ;
  assign y8395 = ~n37504 ;
  assign y8396 = ~n37507 ;
  assign y8397 = n37509 ;
  assign y8398 = ~n37514 ;
  assign y8399 = n37516 ;
  assign y8400 = ~n37522 ;
  assign y8401 = ~n37527 ;
  assign y8402 = n37530 ;
  assign y8403 = n37535 ;
  assign y8404 = ~n37539 ;
  assign y8405 = n37541 ;
  assign y8406 = n37542 ;
  assign y8407 = ~n37543 ;
  assign y8408 = ~n37544 ;
  assign y8409 = ~n37545 ;
  assign y8410 = n37550 ;
  assign y8411 = n37554 ;
  assign y8412 = ~n37557 ;
  assign y8413 = n37558 ;
  assign y8414 = ~n37561 ;
  assign y8415 = ~n37565 ;
  assign y8416 = ~n37567 ;
  assign y8417 = n37568 ;
  assign y8418 = ~n37570 ;
  assign y8419 = n37572 ;
  assign y8420 = ~n37573 ;
  assign y8421 = n37577 ;
  assign y8422 = ~n37579 ;
  assign y8423 = ~n37580 ;
  assign y8424 = n37586 ;
  assign y8425 = n37589 ;
  assign y8426 = n37593 ;
  assign y8427 = ~n37594 ;
  assign y8428 = n37597 ;
  assign y8429 = ~n37598 ;
  assign y8430 = ~n37600 ;
  assign y8431 = n37602 ;
  assign y8432 = n37603 ;
  assign y8433 = n37612 ;
  assign y8434 = n37620 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~n37621 ;
  assign y8437 = n37626 ;
  assign y8438 = n37628 ;
  assign y8439 = ~n37633 ;
  assign y8440 = n37635 ;
  assign y8441 = ~n37638 ;
  assign y8442 = n37640 ;
  assign y8443 = n37644 ;
  assign y8444 = n37649 ;
  assign y8445 = ~n37651 ;
  assign y8446 = n37655 ;
  assign y8447 = n37661 ;
  assign y8448 = n37665 ;
  assign y8449 = ~n37668 ;
  assign y8450 = ~n37670 ;
  assign y8451 = ~n37674 ;
  assign y8452 = ~n37675 ;
  assign y8453 = n37681 ;
  assign y8454 = ~n37687 ;
  assign y8455 = ~n6822 ;
  assign y8456 = ~n37692 ;
  assign y8457 = ~1'b0 ;
  assign y8458 = ~n37693 ;
  assign y8459 = ~n37694 ;
  assign y8460 = ~n37695 ;
  assign y8461 = n37701 ;
  assign y8462 = n37702 ;
  assign y8463 = n37705 ;
  assign y8464 = ~n37706 ;
  assign y8465 = ~1'b0 ;
  assign y8466 = n37707 ;
  assign y8467 = ~n37708 ;
  assign y8468 = ~n37712 ;
  assign y8469 = ~n37713 ;
  assign y8470 = n37719 ;
  assign y8471 = ~n37723 ;
  assign y8472 = ~n37724 ;
  assign y8473 = ~n37725 ;
  assign y8474 = ~n37727 ;
  assign y8475 = n37728 ;
  assign y8476 = n37735 ;
  assign y8477 = ~n37743 ;
  assign y8478 = ~n37745 ;
  assign y8479 = n37747 ;
  assign y8480 = ~n37749 ;
  assign y8481 = ~1'b0 ;
  assign y8482 = n37755 ;
  assign y8483 = n37756 ;
  assign y8484 = ~n37759 ;
  assign y8485 = ~n37761 ;
  assign y8486 = ~n37762 ;
  assign y8487 = n37763 ;
  assign y8488 = ~n37765 ;
  assign y8489 = ~n37767 ;
  assign y8490 = n37771 ;
  assign y8491 = n37774 ;
  assign y8492 = n37775 ;
  assign y8493 = n37779 ;
  assign y8494 = n37783 ;
  assign y8495 = ~n37787 ;
  assign y8496 = ~n37788 ;
  assign y8497 = n37793 ;
  assign y8498 = ~n37794 ;
  assign y8499 = ~n37798 ;
  assign y8500 = n37799 ;
  assign y8501 = n37800 ;
  assign y8502 = ~n37801 ;
  assign y8503 = n37803 ;
  assign y8504 = ~n37810 ;
  assign y8505 = ~n37814 ;
  assign y8506 = n37820 ;
  assign y8507 = n37821 ;
  assign y8508 = ~n37823 ;
  assign y8509 = ~n37824 ;
  assign y8510 = n37827 ;
  assign y8511 = ~1'b0 ;
  assign y8512 = ~1'b0 ;
  assign y8513 = n37828 ;
  assign y8514 = n37829 ;
  assign y8515 = ~n37830 ;
  assign y8516 = n37831 ;
  assign y8517 = n37834 ;
  assign y8518 = ~n37843 ;
  assign y8519 = ~n37846 ;
  assign y8520 = ~1'b0 ;
  assign y8521 = ~n37849 ;
  assign y8522 = ~n37853 ;
  assign y8523 = n37854 ;
  assign y8524 = n37855 ;
  assign y8525 = ~n37859 ;
  assign y8526 = ~n37862 ;
  assign y8527 = n37864 ;
  assign y8528 = n37865 ;
  assign y8529 = n37873 ;
  assign y8530 = n37877 ;
  assign y8531 = ~n37878 ;
  assign y8532 = ~n37879 ;
  assign y8533 = ~n37880 ;
  assign y8534 = ~n37889 ;
  assign y8535 = n37890 ;
  assign y8536 = n37891 ;
  assign y8537 = ~n37893 ;
  assign y8538 = n37897 ;
  assign y8539 = ~n37900 ;
  assign y8540 = n37902 ;
  assign y8541 = ~n37904 ;
  assign y8542 = n37913 ;
  assign y8543 = n37917 ;
  assign y8544 = ~n37922 ;
  assign y8545 = ~n37923 ;
  assign y8546 = n37930 ;
  assign y8547 = ~n37932 ;
  assign y8548 = n37933 ;
  assign y8549 = n37935 ;
  assign y8550 = n37937 ;
  assign y8551 = ~n37938 ;
  assign y8552 = ~n37940 ;
  assign y8553 = n37944 ;
  assign y8554 = n37948 ;
  assign y8555 = n37953 ;
  assign y8556 = n37957 ;
  assign y8557 = n37960 ;
  assign y8558 = ~n37961 ;
  assign y8559 = ~n37965 ;
  assign y8560 = n37968 ;
  assign y8561 = ~n37972 ;
  assign y8562 = n37975 ;
  assign y8563 = n37977 ;
  assign y8564 = ~n37979 ;
  assign y8565 = ~n37980 ;
  assign y8566 = n37981 ;
  assign y8567 = n37982 ;
  assign y8568 = ~n37988 ;
  assign y8569 = n37995 ;
  assign y8570 = ~n37996 ;
  assign y8571 = ~1'b0 ;
  assign y8572 = n38003 ;
  assign y8573 = ~n38009 ;
  assign y8574 = ~n38010 ;
  assign y8575 = n38013 ;
  assign y8576 = ~n38014 ;
  assign y8577 = n38016 ;
  assign y8578 = ~n38023 ;
  assign y8579 = ~n38031 ;
  assign y8580 = n38034 ;
  assign y8581 = n38040 ;
  assign y8582 = ~n38046 ;
  assign y8583 = ~n38049 ;
  assign y8584 = ~n38055 ;
  assign y8585 = n38057 ;
  assign y8586 = ~n38061 ;
  assign y8587 = ~n38065 ;
  assign y8588 = n38066 ;
  assign y8589 = ~n38072 ;
  assign y8590 = n38073 ;
  assign y8591 = n38076 ;
  assign y8592 = ~1'b0 ;
  assign y8593 = ~n38079 ;
  assign y8594 = ~n38080 ;
  assign y8595 = ~n38081 ;
  assign y8596 = ~n38082 ;
  assign y8597 = n38084 ;
  assign y8598 = ~n38087 ;
  assign y8599 = ~n38092 ;
  assign y8600 = n38093 ;
  assign y8601 = ~n38104 ;
  assign y8602 = ~n38105 ;
  assign y8603 = ~n38108 ;
  assign y8604 = n38115 ;
  assign y8605 = ~n38121 ;
  assign y8606 = ~n38125 ;
  assign y8607 = n38129 ;
  assign y8608 = n38131 ;
  assign y8609 = n38132 ;
  assign y8610 = n38135 ;
  assign y8611 = n38138 ;
  assign y8612 = n38139 ;
  assign y8613 = n38142 ;
  assign y8614 = ~n38146 ;
  assign y8615 = n38149 ;
  assign y8616 = ~n38154 ;
  assign y8617 = n38157 ;
  assign y8618 = ~n38164 ;
  assign y8619 = n38165 ;
  assign y8620 = ~n38166 ;
  assign y8621 = n38167 ;
  assign y8622 = n38169 ;
  assign y8623 = ~n38170 ;
  assign y8624 = ~n38177 ;
  assign y8625 = ~n38179 ;
  assign y8626 = n38180 ;
  assign y8627 = ~n38183 ;
  assign y8628 = ~n38185 ;
  assign y8629 = n38187 ;
  assign y8630 = n38190 ;
  assign y8631 = ~n38191 ;
  assign y8632 = ~n38192 ;
  assign y8633 = ~n38194 ;
  assign y8634 = ~n38195 ;
  assign y8635 = n38202 ;
  assign y8636 = n38203 ;
  assign y8637 = n38219 ;
  assign y8638 = n38226 ;
  assign y8639 = n38230 ;
  assign y8640 = ~n38232 ;
  assign y8641 = ~n38236 ;
  assign y8642 = ~n38238 ;
  assign y8643 = n38239 ;
  assign y8644 = n38241 ;
  assign y8645 = ~n38245 ;
  assign y8646 = ~n38246 ;
  assign y8647 = n38247 ;
  assign y8648 = ~n38248 ;
  assign y8649 = n38251 ;
  assign y8650 = ~n38254 ;
  assign y8651 = ~n38264 ;
  assign y8652 = ~n38266 ;
  assign y8653 = ~n38269 ;
  assign y8654 = n38272 ;
  assign y8655 = n38274 ;
  assign y8656 = n38277 ;
  assign y8657 = ~n38280 ;
  assign y8658 = ~1'b0 ;
  assign y8659 = n38283 ;
  assign y8660 = n38285 ;
  assign y8661 = n38287 ;
  assign y8662 = ~n38288 ;
  assign y8663 = ~n38294 ;
  assign y8664 = n38296 ;
  assign y8665 = ~n38302 ;
  assign y8666 = ~n38303 ;
  assign y8667 = n38304 ;
  assign y8668 = ~n38311 ;
  assign y8669 = ~n38313 ;
  assign y8670 = ~n38316 ;
  assign y8671 = n38320 ;
  assign y8672 = ~n38322 ;
  assign y8673 = ~n38325 ;
  assign y8674 = n38327 ;
  assign y8675 = ~n38328 ;
  assign y8676 = n38331 ;
  assign y8677 = ~n38333 ;
  assign y8678 = ~n38335 ;
  assign y8679 = n38343 ;
  assign y8680 = n38345 ;
  assign y8681 = n38348 ;
  assign y8682 = ~n38349 ;
  assign y8683 = n38352 ;
  assign y8684 = ~n38353 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = ~n38355 ;
  assign y8687 = ~n38360 ;
  assign y8688 = n38365 ;
  assign y8689 = n38368 ;
  assign y8690 = n38369 ;
  assign y8691 = ~n38378 ;
  assign y8692 = ~n38380 ;
  assign y8693 = n38382 ;
  assign y8694 = ~n38383 ;
  assign y8695 = n38387 ;
  assign y8696 = n38391 ;
  assign y8697 = ~n38393 ;
  assign y8698 = ~n38394 ;
  assign y8699 = ~n38402 ;
  assign y8700 = n38405 ;
  assign y8701 = ~n38406 ;
  assign y8702 = ~n38416 ;
  assign y8703 = n38418 ;
  assign y8704 = ~n38420 ;
  assign y8705 = n38423 ;
  assign y8706 = ~n38429 ;
  assign y8707 = ~n38434 ;
  assign y8708 = ~n38435 ;
  assign y8709 = ~n38437 ;
  assign y8710 = n38442 ;
  assign y8711 = n38448 ;
  assign y8712 = ~n38452 ;
  assign y8713 = ~1'b0 ;
  assign y8714 = n38454 ;
  assign y8715 = ~n38458 ;
  assign y8716 = ~n38461 ;
  assign y8717 = ~n38462 ;
  assign y8718 = ~n38464 ;
  assign y8719 = n38468 ;
  assign y8720 = n38470 ;
  assign y8721 = n38472 ;
  assign y8722 = n38475 ;
  assign y8723 = ~n38478 ;
  assign y8724 = n38479 ;
  assign y8725 = n38481 ;
  assign y8726 = ~1'b0 ;
  assign y8727 = ~n38485 ;
  assign y8728 = ~n38489 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = n38492 ;
  assign y8731 = n38496 ;
  assign y8732 = n38498 ;
  assign y8733 = ~n38500 ;
  assign y8734 = ~n38505 ;
  assign y8735 = ~n38512 ;
  assign y8736 = n38514 ;
  assign y8737 = ~n38522 ;
  assign y8738 = ~n38523 ;
  assign y8739 = ~n38524 ;
  assign y8740 = ~n38525 ;
  assign y8741 = ~n38531 ;
  assign y8742 = n38532 ;
  assign y8743 = ~n38545 ;
  assign y8744 = ~n38547 ;
  assign y8745 = ~n6652 ;
  assign y8746 = ~n38550 ;
  assign y8747 = n38551 ;
  assign y8748 = ~n38560 ;
  assign y8749 = ~n38568 ;
  assign y8750 = n38570 ;
  assign y8751 = n38572 ;
  assign y8752 = ~n38573 ;
  assign y8753 = ~1'b0 ;
  assign y8754 = n38583 ;
  assign y8755 = n38587 ;
  assign y8756 = ~n38590 ;
  assign y8757 = ~n38592 ;
  assign y8758 = n38596 ;
  assign y8759 = n38601 ;
  assign y8760 = ~n38603 ;
  assign y8761 = n38605 ;
  assign y8762 = n38607 ;
  assign y8763 = n38609 ;
  assign y8764 = ~n38614 ;
  assign y8765 = n38615 ;
  assign y8766 = n38618 ;
  assign y8767 = ~n38621 ;
  assign y8768 = ~n38622 ;
  assign y8769 = ~n38623 ;
  assign y8770 = ~n38627 ;
  assign y8771 = ~n38635 ;
  assign y8772 = ~1'b0 ;
  assign y8773 = n38639 ;
  assign y8774 = n38640 ;
  assign y8775 = n38641 ;
  assign y8776 = n38644 ;
  assign y8777 = n38645 ;
  assign y8778 = ~n38649 ;
  assign y8779 = ~n38651 ;
  assign y8780 = ~n38654 ;
  assign y8781 = ~n38657 ;
  assign y8782 = n38663 ;
  assign y8783 = ~n38677 ;
  assign y8784 = ~n38679 ;
  assign y8785 = n38680 ;
  assign y8786 = n38691 ;
  assign y8787 = n38694 ;
  assign y8788 = n38696 ;
  assign y8789 = n38699 ;
  assign y8790 = ~n38703 ;
  assign y8791 = n38705 ;
  assign y8792 = n38706 ;
  assign y8793 = ~n38707 ;
  assign y8794 = n38711 ;
  assign y8795 = ~n38712 ;
  assign y8796 = n38716 ;
  assign y8797 = ~n38719 ;
  assign y8798 = n38721 ;
  assign y8799 = n38724 ;
  assign y8800 = n38726 ;
  assign y8801 = n38727 ;
  assign y8802 = n38730 ;
  assign y8803 = n38731 ;
  assign y8804 = ~n38734 ;
  assign y8805 = ~1'b0 ;
  assign y8806 = n38738 ;
  assign y8807 = n38744 ;
  assign y8808 = n38752 ;
  assign y8809 = n38755 ;
  assign y8810 = ~n38759 ;
  assign y8811 = n38761 ;
  assign y8812 = n38766 ;
  assign y8813 = ~n38772 ;
  assign y8814 = ~n38774 ;
  assign y8815 = ~n38781 ;
  assign y8816 = n38785 ;
  assign y8817 = n38790 ;
  assign y8818 = ~n38791 ;
  assign y8819 = ~n38792 ;
  assign y8820 = ~n38794 ;
  assign y8821 = n38797 ;
  assign y8822 = n38801 ;
  assign y8823 = ~n38802 ;
  assign y8824 = n38803 ;
  assign y8825 = ~n38812 ;
  assign y8826 = ~n38813 ;
  assign y8827 = ~n38815 ;
  assign y8828 = n38825 ;
  assign y8829 = n38828 ;
  assign y8830 = n38830 ;
  assign y8831 = n38840 ;
  assign y8832 = n38843 ;
  assign y8833 = n38845 ;
  assign y8834 = n38848 ;
  assign y8835 = n38849 ;
  assign y8836 = ~n38850 ;
  assign y8837 = ~n38851 ;
  assign y8838 = ~n38855 ;
  assign y8839 = ~n38857 ;
  assign y8840 = ~n38865 ;
  assign y8841 = ~n38866 ;
  assign y8842 = n38867 ;
  assign y8843 = n38875 ;
  assign y8844 = n38877 ;
  assign y8845 = ~n38878 ;
  assign y8846 = n38879 ;
  assign y8847 = ~n38883 ;
  assign y8848 = n38884 ;
  assign y8849 = n38886 ;
  assign y8850 = n38888 ;
  assign y8851 = n38890 ;
  assign y8852 = n38893 ;
  assign y8853 = n38895 ;
  assign y8854 = ~n38896 ;
  assign y8855 = ~n38899 ;
  assign y8856 = n38901 ;
  assign y8857 = n38905 ;
  assign y8858 = n38907 ;
  assign y8859 = ~n38913 ;
  assign y8860 = ~n38921 ;
  assign y8861 = n38924 ;
  assign y8862 = n38928 ;
  assign y8863 = ~n38931 ;
  assign y8864 = n38937 ;
  assign y8865 = n38938 ;
  assign y8866 = ~n38940 ;
  assign y8867 = n38951 ;
  assign y8868 = ~n38953 ;
  assign y8869 = n38954 ;
  assign y8870 = n38957 ;
  assign y8871 = ~n38959 ;
  assign y8872 = n38963 ;
  assign y8873 = ~n38964 ;
  assign y8874 = n38966 ;
  assign y8875 = ~n38971 ;
  assign y8876 = n38973 ;
  assign y8877 = n38979 ;
  assign y8878 = ~n38982 ;
  assign y8879 = n38985 ;
  assign y8880 = ~n38992 ;
  assign y8881 = ~n38995 ;
  assign y8882 = n38998 ;
  assign y8883 = ~n38999 ;
  assign y8884 = ~n39000 ;
  assign y8885 = n39014 ;
  assign y8886 = n39017 ;
  assign y8887 = ~n39018 ;
  assign y8888 = ~n39020 ;
  assign y8889 = n39023 ;
  assign y8890 = ~n39024 ;
  assign y8891 = ~1'b0 ;
  assign y8892 = ~n39025 ;
  assign y8893 = n39026 ;
  assign y8894 = ~n39027 ;
  assign y8895 = ~n39028 ;
  assign y8896 = ~n39032 ;
  assign y8897 = n39039 ;
  assign y8898 = ~n39042 ;
  assign y8899 = ~n39043 ;
  assign y8900 = n39045 ;
  assign y8901 = ~1'b0 ;
  assign y8902 = ~n39047 ;
  assign y8903 = n39050 ;
  assign y8904 = ~n39052 ;
  assign y8905 = n39053 ;
  assign y8906 = ~n39059 ;
  assign y8907 = ~n39060 ;
  assign y8908 = ~n39064 ;
  assign y8909 = n39068 ;
  assign y8910 = n39074 ;
  assign y8911 = n39078 ;
  assign y8912 = ~n39085 ;
  assign y8913 = n39087 ;
  assign y8914 = ~n39089 ;
  assign y8915 = ~1'b0 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = ~n39097 ;
  assign y8918 = ~n39099 ;
  assign y8919 = ~1'b0 ;
  assign y8920 = n39103 ;
  assign y8921 = n39107 ;
  assign y8922 = ~n39113 ;
  assign y8923 = ~n39118 ;
  assign y8924 = ~1'b0 ;
  assign y8925 = n39119 ;
  assign y8926 = n39120 ;
  assign y8927 = n39129 ;
  assign y8928 = ~n39132 ;
  assign y8929 = n39134 ;
  assign y8930 = n39135 ;
  assign y8931 = ~n39136 ;
  assign y8932 = n39139 ;
  assign y8933 = ~n39140 ;
  assign y8934 = ~n39144 ;
  assign y8935 = n39145 ;
  assign y8936 = ~n39147 ;
  assign y8937 = n39155 ;
  assign y8938 = n39160 ;
  assign y8939 = ~n39162 ;
  assign y8940 = ~1'b0 ;
  assign y8941 = n39167 ;
  assign y8942 = n39171 ;
  assign y8943 = n39172 ;
  assign y8944 = ~n39174 ;
  assign y8945 = n39176 ;
  assign y8946 = n39183 ;
  assign y8947 = ~n39187 ;
  assign y8948 = ~1'b0 ;
  assign y8949 = ~n39192 ;
  assign y8950 = ~n39198 ;
  assign y8951 = n39209 ;
  assign y8952 = n39211 ;
  assign y8953 = n39213 ;
  assign y8954 = n39219 ;
  assign y8955 = ~n39225 ;
  assign y8956 = ~n39227 ;
  assign y8957 = ~n21483 ;
  assign y8958 = n39228 ;
  assign y8959 = ~n39230 ;
  assign y8960 = n39244 ;
  assign y8961 = n39247 ;
  assign y8962 = n39249 ;
  assign y8963 = n39250 ;
  assign y8964 = n39252 ;
  assign y8965 = ~n39254 ;
  assign y8966 = ~n39255 ;
  assign y8967 = ~n39256 ;
  assign y8968 = ~n39260 ;
  assign y8969 = n39262 ;
  assign y8970 = n39265 ;
  assign y8971 = n39267 ;
  assign y8972 = ~n39276 ;
  assign y8973 = n39277 ;
  assign y8974 = ~n39278 ;
  assign y8975 = ~n39283 ;
  assign y8976 = ~n39287 ;
  assign y8977 = ~n39299 ;
  assign y8978 = n39301 ;
  assign y8979 = ~n39304 ;
  assign y8980 = n39308 ;
  assign y8981 = ~n39310 ;
  assign y8982 = n39311 ;
  assign y8983 = ~1'b0 ;
  assign y8984 = ~n39313 ;
  assign y8985 = n39315 ;
  assign y8986 = ~n39316 ;
  assign y8987 = n39318 ;
  assign y8988 = n39322 ;
  assign y8989 = n39323 ;
  assign y8990 = n39324 ;
  assign y8991 = ~n39329 ;
  assign y8992 = ~n39331 ;
  assign y8993 = n39334 ;
  assign y8994 = n39336 ;
  assign y8995 = n39339 ;
  assign y8996 = ~n39344 ;
  assign y8997 = ~n39347 ;
  assign y8998 = n39350 ;
  assign y8999 = ~n39352 ;
  assign y9000 = n39354 ;
  assign y9001 = n39355 ;
  assign y9002 = ~n39356 ;
  assign y9003 = ~n39359 ;
  assign y9004 = ~n39363 ;
  assign y9005 = ~n39365 ;
  assign y9006 = ~n39371 ;
  assign y9007 = n39372 ;
  assign y9008 = ~n39376 ;
  assign y9009 = n39378 ;
  assign y9010 = n39381 ;
  assign y9011 = n39382 ;
  assign y9012 = n39389 ;
  assign y9013 = n39390 ;
  assign y9014 = ~n39391 ;
  assign y9015 = ~n39396 ;
  assign y9016 = ~n39398 ;
  assign y9017 = n39401 ;
  assign y9018 = ~n39402 ;
  assign y9019 = ~n39405 ;
  assign y9020 = n39407 ;
  assign y9021 = ~n39410 ;
  assign y9022 = ~n39412 ;
  assign y9023 = ~n39413 ;
  assign y9024 = n39415 ;
  assign y9025 = ~n39417 ;
  assign y9026 = ~n39424 ;
  assign y9027 = ~n39433 ;
  assign y9028 = n39434 ;
  assign y9029 = n39436 ;
  assign y9030 = ~n39437 ;
  assign y9031 = ~n39442 ;
  assign y9032 = ~n39445 ;
  assign y9033 = n39452 ;
  assign y9034 = n39455 ;
  assign y9035 = n39456 ;
  assign y9036 = ~n39464 ;
  assign y9037 = ~n39465 ;
  assign y9038 = ~n39474 ;
  assign y9039 = n39475 ;
  assign y9040 = ~n39477 ;
  assign y9041 = ~1'b0 ;
  assign y9042 = n39485 ;
  assign y9043 = ~n39486 ;
  assign y9044 = n39488 ;
  assign y9045 = ~n39490 ;
  assign y9046 = n39492 ;
  assign y9047 = n39497 ;
  assign y9048 = n39499 ;
  assign y9049 = ~n39502 ;
  assign y9050 = ~n39506 ;
  assign y9051 = n39508 ;
  assign y9052 = n39512 ;
  assign y9053 = n39521 ;
  assign y9054 = ~n39522 ;
  assign y9055 = ~n39527 ;
  assign y9056 = ~n39529 ;
  assign y9057 = ~n39531 ;
  assign y9058 = ~n39535 ;
  assign y9059 = n39540 ;
  assign y9060 = ~n39546 ;
  assign y9061 = ~n39552 ;
  assign y9062 = n39553 ;
  assign y9063 = n39558 ;
  assign y9064 = ~n39566 ;
  assign y9065 = n39568 ;
  assign y9066 = ~n39569 ;
  assign y9067 = ~n39571 ;
  assign y9068 = n39572 ;
  assign y9069 = n39573 ;
  assign y9070 = ~n39577 ;
  assign y9071 = ~1'b0 ;
  assign y9072 = ~n39578 ;
  assign y9073 = n39580 ;
  assign y9074 = ~n39581 ;
  assign y9075 = n39583 ;
  assign y9076 = n39586 ;
  assign y9077 = ~n39589 ;
  assign y9078 = n39592 ;
  assign y9079 = ~n39594 ;
  assign y9080 = ~n39596 ;
  assign y9081 = ~n39597 ;
  assign y9082 = n39598 ;
  assign y9083 = ~n39604 ;
  assign y9084 = ~n39614 ;
  assign y9085 = ~n39618 ;
  assign y9086 = ~n39628 ;
  assign y9087 = ~n39634 ;
  assign y9088 = ~n39639 ;
  assign y9089 = n39643 ;
  assign y9090 = ~n39646 ;
  assign y9091 = n39649 ;
  assign y9092 = ~n39651 ;
  assign y9093 = ~n39654 ;
  assign y9094 = n39655 ;
  assign y9095 = ~n39657 ;
  assign y9096 = n39659 ;
  assign y9097 = ~n39662 ;
  assign y9098 = ~n39666 ;
  assign y9099 = n39669 ;
  assign y9100 = n39672 ;
  assign y9101 = ~1'b0 ;
  assign y9102 = n39673 ;
  assign y9103 = ~n39674 ;
  assign y9104 = ~n39675 ;
  assign y9105 = ~n39678 ;
  assign y9106 = ~n39681 ;
  assign y9107 = n39686 ;
  assign y9108 = n39689 ;
  assign y9109 = ~1'b0 ;
  assign y9110 = ~1'b0 ;
  assign y9111 = ~n39691 ;
  assign y9112 = ~n39694 ;
  assign y9113 = n39695 ;
  assign y9114 = n39700 ;
  assign y9115 = ~n39705 ;
  assign y9116 = n39710 ;
  assign y9117 = ~n39713 ;
  assign y9118 = n39718 ;
  assign y9119 = ~n39719 ;
  assign y9120 = n39720 ;
  assign y9121 = ~n39722 ;
  assign y9122 = ~n39723 ;
  assign y9123 = n39727 ;
  assign y9124 = n39731 ;
  assign y9125 = n39734 ;
  assign y9126 = ~n39735 ;
  assign y9127 = n39738 ;
  assign y9128 = n39739 ;
  assign y9129 = ~n39742 ;
  assign y9130 = ~n39746 ;
  assign y9131 = n39749 ;
  assign y9132 = ~n39754 ;
  assign y9133 = ~n39760 ;
  assign y9134 = ~n39762 ;
  assign y9135 = ~n39764 ;
  assign y9136 = ~n39768 ;
  assign y9137 = n39770 ;
  assign y9138 = ~1'b0 ;
  assign y9139 = n39772 ;
  assign y9140 = ~n39773 ;
  assign y9141 = ~n39776 ;
  assign y9142 = ~n39777 ;
  assign y9143 = n39778 ;
  assign y9144 = ~n39781 ;
  assign y9145 = n39783 ;
  assign y9146 = ~n39784 ;
  assign y9147 = ~n39794 ;
  assign y9148 = ~n39799 ;
  assign y9149 = n39801 ;
  assign y9150 = n39802 ;
  assign y9151 = ~n39804 ;
  assign y9152 = ~n39806 ;
  assign y9153 = n39807 ;
  assign y9154 = n39809 ;
  assign y9155 = n39812 ;
  assign y9156 = ~n39813 ;
  assign y9157 = n39818 ;
  assign y9158 = ~n39821 ;
  assign y9159 = n39823 ;
  assign y9160 = ~n39825 ;
  assign y9161 = n39827 ;
  assign y9162 = n39832 ;
  assign y9163 = ~n39833 ;
  assign y9164 = ~n39835 ;
  assign y9165 = ~n39840 ;
  assign y9166 = n39843 ;
  assign y9167 = ~n39845 ;
  assign y9168 = ~n39851 ;
  assign y9169 = ~n39852 ;
  assign y9170 = ~n39854 ;
  assign y9171 = ~n39862 ;
  assign y9172 = ~n39866 ;
  assign y9173 = ~n39867 ;
  assign y9174 = ~1'b0 ;
  assign y9175 = ~n39870 ;
  assign y9176 = n39872 ;
  assign y9177 = n39881 ;
  assign y9178 = ~n39882 ;
  assign y9179 = ~n39886 ;
  assign y9180 = n39895 ;
  assign y9181 = ~n39896 ;
  assign y9182 = ~n39899 ;
  assign y9183 = ~n39903 ;
  assign y9184 = n39905 ;
  assign y9185 = n39910 ;
  assign y9186 = ~n39912 ;
  assign y9187 = n39914 ;
  assign y9188 = ~n39916 ;
  assign y9189 = ~1'b0 ;
  assign y9190 = n39918 ;
  assign y9191 = ~n39921 ;
  assign y9192 = ~n39926 ;
  assign y9193 = n39927 ;
  assign y9194 = ~n39928 ;
  assign y9195 = n39930 ;
  assign y9196 = ~1'b0 ;
  assign y9197 = ~n39931 ;
  assign y9198 = ~n39935 ;
  assign y9199 = ~n39939 ;
  assign y9200 = ~n39940 ;
  assign y9201 = ~n39941 ;
  assign y9202 = ~n39944 ;
  assign y9203 = ~n39946 ;
  assign y9204 = ~n39950 ;
  assign y9205 = ~n39951 ;
  assign y9206 = n39953 ;
  assign y9207 = ~1'b0 ;
  assign y9208 = n39956 ;
  assign y9209 = n39959 ;
  assign y9210 = ~n39961 ;
  assign y9211 = ~n39963 ;
  assign y9212 = n39968 ;
  assign y9213 = ~n39971 ;
  assign y9214 = ~1'b0 ;
  assign y9215 = ~n39973 ;
  assign y9216 = ~n39975 ;
  assign y9217 = ~n39980 ;
  assign y9218 = ~n39981 ;
  assign y9219 = ~n39982 ;
  assign y9220 = ~n39985 ;
  assign y9221 = ~n39988 ;
  assign y9222 = ~n39990 ;
  assign y9223 = n39992 ;
  assign y9224 = n39993 ;
  assign y9225 = n39998 ;
  assign y9226 = n40006 ;
  assign y9227 = ~n40010 ;
  assign y9228 = n40015 ;
  assign y9229 = n40016 ;
  assign y9230 = ~n40021 ;
  assign y9231 = n40025 ;
  assign y9232 = n40029 ;
  assign y9233 = n40031 ;
  assign y9234 = ~1'b0 ;
  assign y9235 = n40033 ;
  assign y9236 = ~n40034 ;
  assign y9237 = n40036 ;
  assign y9238 = n40039 ;
  assign y9239 = n40046 ;
  assign y9240 = n40048 ;
  assign y9241 = n40051 ;
  assign y9242 = n40053 ;
  assign y9243 = n40054 ;
  assign y9244 = n40057 ;
  assign y9245 = n40062 ;
  assign y9246 = ~n40063 ;
  assign y9247 = ~n40070 ;
  assign y9248 = n40073 ;
  assign y9249 = ~n40075 ;
  assign y9250 = ~n40078 ;
  assign y9251 = ~n40079 ;
  assign y9252 = n40082 ;
  assign y9253 = n40087 ;
  assign y9254 = n40089 ;
  assign y9255 = ~n40090 ;
  assign y9256 = n40091 ;
  assign y9257 = ~n40095 ;
  assign y9258 = n40107 ;
  assign y9259 = ~n40111 ;
  assign y9260 = ~n40112 ;
  assign y9261 = ~n40118 ;
  assign y9262 = ~n40123 ;
  assign y9263 = ~n40124 ;
  assign y9264 = ~n40126 ;
  assign y9265 = n40130 ;
  assign y9266 = n40139 ;
  assign y9267 = ~n40146 ;
  assign y9268 = n40150 ;
  assign y9269 = ~n40152 ;
  assign y9270 = n40156 ;
  assign y9271 = ~1'b0 ;
  assign y9272 = n40157 ;
  assign y9273 = n40165 ;
  assign y9274 = ~n40166 ;
  assign y9275 = ~n40167 ;
  assign y9276 = ~n40171 ;
  assign y9277 = n40173 ;
  assign y9278 = ~n40180 ;
  assign y9279 = ~n40188 ;
  assign y9280 = n40192 ;
  assign y9281 = n40193 ;
  assign y9282 = n40197 ;
  assign y9283 = ~n40200 ;
  assign y9284 = ~n40201 ;
  assign y9285 = ~1'b0 ;
  assign y9286 = ~n40204 ;
  assign y9287 = ~n40205 ;
  assign y9288 = ~n40206 ;
  assign y9289 = ~n40208 ;
  assign y9290 = n40210 ;
  assign y9291 = ~n40211 ;
  assign y9292 = ~n40213 ;
  assign y9293 = n40216 ;
  assign y9294 = ~n40220 ;
  assign y9295 = n40222 ;
  assign y9296 = ~n40223 ;
  assign y9297 = ~n40229 ;
  assign y9298 = n40233 ;
  assign y9299 = n40237 ;
  assign y9300 = ~n40240 ;
  assign y9301 = ~n40241 ;
  assign y9302 = n40244 ;
  assign y9303 = n40254 ;
  assign y9304 = ~n40257 ;
  assign y9305 = n40258 ;
  assign y9306 = n40260 ;
  assign y9307 = n40262 ;
  assign y9308 = n40267 ;
  assign y9309 = ~n40268 ;
  assign y9310 = ~n40272 ;
  assign y9311 = n40275 ;
  assign y9312 = ~1'b0 ;
  assign y9313 = ~1'b0 ;
  assign y9314 = ~n40279 ;
  assign y9315 = ~n40280 ;
  assign y9316 = n40281 ;
  assign y9317 = ~n40283 ;
  assign y9318 = n40284 ;
  assign y9319 = ~n40288 ;
  assign y9320 = ~n40289 ;
  assign y9321 = n40294 ;
  assign y9322 = ~n40297 ;
  assign y9323 = n40298 ;
  assign y9324 = n40299 ;
  assign y9325 = n40301 ;
  assign y9326 = ~n40303 ;
  assign y9327 = n40315 ;
  assign y9328 = ~n40320 ;
  assign y9329 = ~n40322 ;
  assign y9330 = n40323 ;
  assign y9331 = ~n40324 ;
  assign y9332 = n40336 ;
  assign y9333 = n40339 ;
  assign y9334 = n40342 ;
  assign y9335 = ~n40344 ;
  assign y9336 = ~n40345 ;
  assign y9337 = n40346 ;
  assign y9338 = ~n40350 ;
  assign y9339 = n40352 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = ~n40355 ;
  assign y9342 = ~n40357 ;
  assign y9343 = n40359 ;
  assign y9344 = ~n40360 ;
  assign y9345 = n40361 ;
  assign y9346 = n40362 ;
  assign y9347 = n40364 ;
  assign y9348 = ~n40366 ;
  assign y9349 = n40369 ;
  assign y9350 = n40371 ;
  assign y9351 = ~n40372 ;
  assign y9352 = n40385 ;
  assign y9353 = ~n40386 ;
  assign y9354 = n40390 ;
  assign y9355 = n40396 ;
  assign y9356 = ~n40397 ;
  assign y9357 = n40399 ;
  assign y9358 = ~n40401 ;
  assign y9359 = ~n40402 ;
  assign y9360 = n40406 ;
  assign y9361 = ~n40407 ;
  assign y9362 = n40408 ;
  assign y9363 = ~n40410 ;
  assign y9364 = ~n40411 ;
  assign y9365 = n40413 ;
  assign y9366 = n40414 ;
  assign y9367 = n29465 ;
  assign y9368 = n40416 ;
  assign y9369 = ~n40418 ;
  assign y9370 = n40421 ;
  assign y9371 = n40424 ;
  assign y9372 = n40425 ;
  assign y9373 = n40429 ;
  assign y9374 = n40431 ;
  assign y9375 = ~n40432 ;
  assign y9376 = n40433 ;
  assign y9377 = n40437 ;
  assign y9378 = ~n40438 ;
  assign y9379 = n40440 ;
  assign y9380 = ~n40442 ;
  assign y9381 = ~n40445 ;
  assign y9382 = n40448 ;
  assign y9383 = ~n40451 ;
  assign y9384 = ~n40454 ;
  assign y9385 = ~n40460 ;
  assign y9386 = ~n40463 ;
  assign y9387 = n40471 ;
  assign y9388 = n40475 ;
  assign y9389 = ~n40477 ;
  assign y9390 = ~n40481 ;
  assign y9391 = n40482 ;
  assign y9392 = ~n40484 ;
  assign y9393 = ~n40486 ;
  assign y9394 = n40494 ;
  assign y9395 = ~n40495 ;
  assign y9396 = ~n40499 ;
  assign y9397 = ~n40501 ;
  assign y9398 = n40503 ;
  assign y9399 = n40507 ;
  assign y9400 = ~n40511 ;
  assign y9401 = n40516 ;
  assign y9402 = ~n40519 ;
  assign y9403 = ~n40521 ;
  assign y9404 = ~n40523 ;
  assign y9405 = ~n40526 ;
  assign y9406 = ~n40527 ;
  assign y9407 = n40530 ;
  assign y9408 = n40532 ;
  assign y9409 = n40538 ;
  assign y9410 = n40543 ;
  assign y9411 = ~n40546 ;
  assign y9412 = n40552 ;
  assign y9413 = ~1'b0 ;
  assign y9414 = n40553 ;
  assign y9415 = n40557 ;
  assign y9416 = n40562 ;
  assign y9417 = n40563 ;
  assign y9418 = n40565 ;
  assign y9419 = ~n40568 ;
  assign y9420 = ~1'b0 ;
  assign y9421 = ~n40572 ;
  assign y9422 = ~n40573 ;
  assign y9423 = ~n40574 ;
  assign y9424 = n40575 ;
  assign y9425 = ~n40580 ;
  assign y9426 = n40581 ;
  assign y9427 = n40585 ;
  assign y9428 = ~n40588 ;
  assign y9429 = n40590 ;
  assign y9430 = n40594 ;
  assign y9431 = n40595 ;
  assign y9432 = n40597 ;
  assign y9433 = ~n40598 ;
  assign y9434 = ~1'b0 ;
  assign y9435 = ~n40599 ;
  assign y9436 = n40610 ;
  assign y9437 = ~n40617 ;
  assign y9438 = n40620 ;
  assign y9439 = ~n40622 ;
  assign y9440 = n852 ;
  assign y9441 = ~n40630 ;
  assign y9442 = ~1'b0 ;
  assign y9443 = ~n40631 ;
  assign y9444 = n40633 ;
  assign y9445 = n40636 ;
  assign y9446 = ~n40637 ;
  assign y9447 = n40642 ;
  assign y9448 = ~n40645 ;
  assign y9449 = n40649 ;
  assign y9450 = n40661 ;
  assign y9451 = ~n40663 ;
  assign y9452 = ~n40664 ;
  assign y9453 = ~n40667 ;
  assign y9454 = n40673 ;
  assign y9455 = n40676 ;
  assign y9456 = n40678 ;
  assign y9457 = ~n40679 ;
  assign y9458 = n40680 ;
  assign y9459 = ~n40690 ;
  assign y9460 = ~n40691 ;
  assign y9461 = ~n40694 ;
  assign y9462 = ~n40698 ;
  assign y9463 = n40702 ;
  assign y9464 = ~n40704 ;
  assign y9465 = n40708 ;
  assign y9466 = ~n40710 ;
  assign y9467 = ~n40712 ;
  assign y9468 = n40714 ;
  assign y9469 = ~1'b0 ;
  assign y9470 = ~n40721 ;
  assign y9471 = ~n40723 ;
  assign y9472 = n40726 ;
  assign y9473 = n40733 ;
  assign y9474 = n40735 ;
  assign y9475 = n40736 ;
  assign y9476 = ~n40740 ;
  assign y9477 = ~1'b0 ;
  assign y9478 = n40744 ;
  assign y9479 = ~n40748 ;
  assign y9480 = n40753 ;
  assign y9481 = n40754 ;
  assign y9482 = ~n40756 ;
  assign y9483 = n40757 ;
  assign y9484 = n40764 ;
  assign y9485 = n40767 ;
  assign y9486 = n40769 ;
  assign y9487 = n40773 ;
  assign y9488 = ~n40775 ;
  assign y9489 = n40777 ;
  assign y9490 = ~n40779 ;
  assign y9491 = n40782 ;
  assign y9492 = ~n40788 ;
  assign y9493 = ~n40789 ;
  assign y9494 = ~n40799 ;
  assign y9495 = ~n40800 ;
  assign y9496 = ~n40802 ;
  assign y9497 = ~n40811 ;
  assign y9498 = ~n40813 ;
  assign y9499 = n40816 ;
  assign y9500 = n40825 ;
  assign y9501 = ~n40826 ;
  assign y9502 = n40829 ;
  assign y9503 = n40830 ;
  assign y9504 = ~n40833 ;
  assign y9505 = ~n40841 ;
  assign y9506 = ~n40845 ;
  assign y9507 = ~n40847 ;
  assign y9508 = ~n40851 ;
  assign y9509 = n40854 ;
  assign y9510 = ~n40856 ;
  assign y9511 = ~n40862 ;
  assign y9512 = n40863 ;
  assign y9513 = n40864 ;
  assign y9514 = ~n40868 ;
  assign y9515 = n40870 ;
  assign y9516 = ~1'b0 ;
  assign y9517 = n40871 ;
  assign y9518 = n40876 ;
  assign y9519 = ~n40878 ;
  assign y9520 = n40879 ;
  assign y9521 = n40880 ;
  assign y9522 = n40883 ;
  assign y9523 = n40887 ;
  assign y9524 = n40888 ;
  assign y9525 = ~n40891 ;
  assign y9526 = n40897 ;
  assign y9527 = n40898 ;
  assign y9528 = ~1'b0 ;
  assign y9529 = ~n40900 ;
  assign y9530 = ~n40902 ;
  assign y9531 = n40904 ;
  assign y9532 = n40914 ;
  assign y9533 = n40920 ;
  assign y9534 = n40921 ;
  assign y9535 = n40924 ;
  assign y9536 = ~n40930 ;
  assign y9537 = n40931 ;
  assign y9538 = n40934 ;
  assign y9539 = ~n40936 ;
  assign y9540 = ~n40941 ;
  assign y9541 = n40954 ;
  assign y9542 = ~n40955 ;
  assign y9543 = ~n40958 ;
  assign y9544 = ~n40961 ;
  assign y9545 = n40964 ;
  assign y9546 = n40966 ;
  assign y9547 = ~n40970 ;
  assign y9548 = n40971 ;
  assign y9549 = ~n40975 ;
  assign y9550 = n40976 ;
  assign y9551 = ~n40978 ;
  assign y9552 = ~n40980 ;
  assign y9553 = n40981 ;
  assign y9554 = n40986 ;
  assign y9555 = n40989 ;
  assign y9556 = n40990 ;
  assign y9557 = ~n40993 ;
  assign y9558 = ~n40995 ;
  assign y9559 = ~n40998 ;
  assign y9560 = ~n41004 ;
  assign y9561 = ~n41006 ;
  assign y9562 = n41012 ;
  assign y9563 = n41014 ;
  assign y9564 = ~n41016 ;
  assign y9565 = ~n41023 ;
  assign y9566 = n41026 ;
  assign y9567 = ~n41027 ;
  assign y9568 = ~n41029 ;
  assign y9569 = ~n41033 ;
  assign y9570 = n41038 ;
  assign y9571 = ~n41046 ;
  assign y9572 = ~n41052 ;
  assign y9573 = n41054 ;
  assign y9574 = n41056 ;
  assign y9575 = n41058 ;
  assign y9576 = ~n41061 ;
  assign y9577 = n41063 ;
  assign y9578 = ~n41068 ;
  assign y9579 = ~n41069 ;
  assign y9580 = ~n41073 ;
  assign y9581 = n41075 ;
  assign y9582 = n41079 ;
  assign y9583 = ~n41083 ;
  assign y9584 = n41086 ;
  assign y9585 = n41089 ;
  assign y9586 = n41091 ;
  assign y9587 = ~n41093 ;
  assign y9588 = ~n41095 ;
  assign y9589 = n41098 ;
  assign y9590 = ~n41100 ;
  assign y9591 = ~n41110 ;
  assign y9592 = ~n41115 ;
  assign y9593 = n41117 ;
  assign y9594 = n41120 ;
  assign y9595 = ~n41127 ;
  assign y9596 = n41129 ;
  assign y9597 = ~n41134 ;
  assign y9598 = n41137 ;
  assign y9599 = n41142 ;
  assign y9600 = n41143 ;
  assign y9601 = n41150 ;
  assign y9602 = ~n41153 ;
  assign y9603 = ~n41158 ;
  assign y9604 = ~n41160 ;
  assign y9605 = n41165 ;
  assign y9606 = ~n41166 ;
  assign y9607 = n41170 ;
  assign y9608 = ~n41171 ;
  assign y9609 = ~1'b0 ;
  assign y9610 = ~n41176 ;
  assign y9611 = n41177 ;
  assign y9612 = n41180 ;
  assign y9613 = n41183 ;
  assign y9614 = n41187 ;
  assign y9615 = ~n41198 ;
  assign y9616 = n41199 ;
  assign y9617 = n41200 ;
  assign y9618 = n41201 ;
  assign y9619 = ~n41203 ;
  assign y9620 = ~n41204 ;
  assign y9621 = ~n41206 ;
  assign y9622 = ~n41214 ;
  assign y9623 = ~n41219 ;
  assign y9624 = ~n41221 ;
  assign y9625 = ~n41227 ;
  assign y9626 = ~n41231 ;
  assign y9627 = ~n41233 ;
  assign y9628 = n41235 ;
  assign y9629 = n41236 ;
  assign y9630 = ~n41237 ;
  assign y9631 = ~n41238 ;
  assign y9632 = n41239 ;
  assign y9633 = ~n41242 ;
  assign y9634 = ~n41244 ;
  assign y9635 = n41245 ;
  assign y9636 = ~n41246 ;
  assign y9637 = ~n41252 ;
  assign y9638 = ~n41253 ;
  assign y9639 = ~n41256 ;
  assign y9640 = ~n41257 ;
  assign y9641 = n41259 ;
  assign y9642 = ~n41260 ;
  assign y9643 = n41262 ;
  assign y9644 = ~n41263 ;
  assign y9645 = n41264 ;
  assign y9646 = n41265 ;
  assign y9647 = ~n41270 ;
  assign y9648 = n41272 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = n41274 ;
  assign y9651 = ~n41275 ;
  assign y9652 = ~n41279 ;
  assign y9653 = ~n41280 ;
  assign y9654 = n41286 ;
  assign y9655 = n41287 ;
  assign y9656 = ~n41289 ;
  assign y9657 = ~n41294 ;
  assign y9658 = ~n41297 ;
  assign y9659 = n41299 ;
  assign y9660 = n41300 ;
  assign y9661 = ~n41303 ;
  assign y9662 = n41304 ;
  assign y9663 = n41306 ;
  assign y9664 = ~n41307 ;
  assign y9665 = n41309 ;
  assign y9666 = ~n41312 ;
  assign y9667 = ~n41314 ;
  assign y9668 = ~n41316 ;
  assign y9669 = ~n41317 ;
  assign y9670 = n41318 ;
  assign y9671 = ~n41324 ;
  assign y9672 = n41325 ;
  assign y9673 = ~n41329 ;
  assign y9674 = ~n41331 ;
  assign y9675 = ~n41333 ;
  assign y9676 = ~n41335 ;
  assign y9677 = n41342 ;
  assign y9678 = ~n41345 ;
  assign y9679 = ~n41349 ;
  assign y9680 = n41351 ;
  assign y9681 = n41353 ;
  assign y9682 = ~n41355 ;
  assign y9683 = n41356 ;
  assign y9684 = n41357 ;
  assign y9685 = n41358 ;
  assign y9686 = n41359 ;
  assign y9687 = n41363 ;
  assign y9688 = n41365 ;
  assign y9689 = n41366 ;
  assign y9690 = n41368 ;
  assign y9691 = ~n41369 ;
  assign y9692 = n41372 ;
  assign y9693 = ~n41375 ;
  assign y9694 = n41376 ;
  assign y9695 = n41378 ;
  assign y9696 = ~n41381 ;
  assign y9697 = n41384 ;
  assign y9698 = ~1'b0 ;
  assign y9699 = n41392 ;
  assign y9700 = ~n41393 ;
  assign y9701 = ~n41394 ;
  assign y9702 = ~n41395 ;
  assign y9703 = ~n41401 ;
  assign y9704 = ~n41403 ;
  assign y9705 = n41404 ;
  assign y9706 = ~n41405 ;
  assign y9707 = n41410 ;
  assign y9708 = n41414 ;
  assign y9709 = ~n41415 ;
  assign y9710 = ~n41418 ;
  assign y9711 = ~n41420 ;
  assign y9712 = ~n41427 ;
  assign y9713 = n41429 ;
  assign y9714 = ~n41431 ;
  assign y9715 = ~n41433 ;
  assign y9716 = n41434 ;
  assign y9717 = ~n41437 ;
  assign y9718 = n41439 ;
  assign y9719 = ~n41441 ;
  assign y9720 = n41442 ;
  assign y9721 = ~n41443 ;
  assign y9722 = ~n41445 ;
  assign y9723 = ~n41452 ;
  assign y9724 = n41457 ;
  assign y9725 = n41462 ;
  assign y9726 = n41467 ;
  assign y9727 = n41469 ;
  assign y9728 = ~n41470 ;
  assign y9729 = n41471 ;
  assign y9730 = ~n41477 ;
  assign y9731 = ~n41479 ;
  assign y9732 = ~n41481 ;
  assign y9733 = ~n41483 ;
  assign y9734 = ~n41491 ;
  assign y9735 = ~n41492 ;
  assign y9736 = n41494 ;
  assign y9737 = ~n41497 ;
  assign y9738 = ~n41498 ;
  assign y9739 = ~n41499 ;
  assign y9740 = ~n41505 ;
  assign y9741 = ~n41511 ;
  assign y9742 = ~n41513 ;
  assign y9743 = ~1'b0 ;
  assign y9744 = ~n41514 ;
  assign y9745 = n41517 ;
  assign y9746 = n41518 ;
  assign y9747 = ~n41522 ;
  assign y9748 = n41525 ;
  assign y9749 = n41528 ;
  assign y9750 = ~n41530 ;
  assign y9751 = n41532 ;
  assign y9752 = ~n41534 ;
  assign y9753 = ~n41535 ;
  assign y9754 = n41539 ;
  assign y9755 = n41540 ;
  assign y9756 = ~n41541 ;
  assign y9757 = n41545 ;
  assign y9758 = ~1'b0 ;
  assign y9759 = ~n41547 ;
  assign y9760 = n41548 ;
  assign y9761 = ~n41549 ;
  assign y9762 = ~n41551 ;
  assign y9763 = ~1'b0 ;
  assign y9764 = n41558 ;
  assign y9765 = n41561 ;
  assign y9766 = ~n41562 ;
  assign y9767 = ~n41563 ;
  assign y9768 = ~1'b0 ;
  assign y9769 = n41567 ;
  assign y9770 = ~n41568 ;
  assign y9771 = n41569 ;
  assign y9772 = n41571 ;
  assign y9773 = n41573 ;
  assign y9774 = ~n41578 ;
  assign y9775 = ~n41582 ;
  assign y9776 = ~n41587 ;
  assign y9777 = n41588 ;
  assign y9778 = n41591 ;
  assign y9779 = ~n41592 ;
  assign y9780 = n41598 ;
  assign y9781 = ~n41600 ;
  assign y9782 = ~n41606 ;
  assign y9783 = n41608 ;
  assign y9784 = n41610 ;
  assign y9785 = ~n41613 ;
  assign y9786 = n41617 ;
  assign y9787 = n41619 ;
  assign y9788 = ~n41621 ;
  assign y9789 = ~n41622 ;
  assign y9790 = n41624 ;
  assign y9791 = n41628 ;
  assign y9792 = n41630 ;
  assign y9793 = n41631 ;
  assign y9794 = n41632 ;
  assign y9795 = ~n41633 ;
  assign y9796 = ~1'b0 ;
  assign y9797 = ~n41635 ;
  assign y9798 = n41641 ;
  assign y9799 = n41643 ;
  assign y9800 = n41650 ;
  assign y9801 = ~n41651 ;
  assign y9802 = ~n41655 ;
  assign y9803 = n41656 ;
  assign y9804 = ~n41657 ;
  assign y9805 = n41659 ;
  assign y9806 = ~n41664 ;
  assign y9807 = ~n41665 ;
  assign y9808 = ~n41667 ;
  assign y9809 = n41669 ;
  assign y9810 = ~n41671 ;
  assign y9811 = ~n41673 ;
  assign y9812 = n41674 ;
  assign y9813 = n41675 ;
  assign y9814 = n41678 ;
  assign y9815 = ~n41679 ;
  assign y9816 = ~n41685 ;
  assign y9817 = n41687 ;
  assign y9818 = n41690 ;
  assign y9819 = ~n41692 ;
  assign y9820 = n41694 ;
  assign y9821 = ~n41697 ;
  assign y9822 = ~n41698 ;
  assign y9823 = ~n41699 ;
  assign y9824 = ~n41700 ;
  assign y9825 = n41701 ;
  assign y9826 = n41703 ;
  assign y9827 = n41704 ;
  assign y9828 = ~n41706 ;
  assign y9829 = n41707 ;
  assign y9830 = ~n41716 ;
  assign y9831 = ~n41717 ;
  assign y9832 = n41719 ;
  assign y9833 = n41725 ;
  assign y9834 = ~n41726 ;
  assign y9835 = ~n41727 ;
  assign y9836 = ~n41729 ;
  assign y9837 = ~1'b0 ;
  assign y9838 = n41734 ;
  assign y9839 = n41740 ;
  assign y9840 = n41741 ;
  assign y9841 = n41744 ;
  assign y9842 = n41745 ;
  assign y9843 = n41747 ;
  assign y9844 = n41748 ;
  assign y9845 = n41753 ;
  assign y9846 = ~n41754 ;
  assign y9847 = n41755 ;
  assign y9848 = ~n41758 ;
  assign y9849 = n41761 ;
  assign y9850 = ~n41764 ;
  assign y9851 = n41769 ;
  assign y9852 = n41772 ;
  assign y9853 = ~n41775 ;
  assign y9854 = n41779 ;
  assign y9855 = n41782 ;
  assign y9856 = ~n41784 ;
  assign y9857 = n41786 ;
  assign y9858 = ~n41789 ;
  assign y9859 = ~1'b0 ;
  assign y9860 = ~n41790 ;
  assign y9861 = ~1'b0 ;
  assign y9862 = n41792 ;
  assign y9863 = n41793 ;
  assign y9864 = ~n41794 ;
  assign y9865 = ~1'b0 ;
  assign y9866 = ~n41796 ;
  assign y9867 = n41798 ;
  assign y9868 = n41799 ;
  assign y9869 = ~n41804 ;
  assign y9870 = ~n41806 ;
  assign y9871 = ~n41807 ;
  assign y9872 = ~n41812 ;
  assign y9873 = ~n41815 ;
  assign y9874 = ~n41817 ;
  assign y9875 = n41818 ;
  assign y9876 = ~n41819 ;
  assign y9877 = n41824 ;
  assign y9878 = n41825 ;
  assign y9879 = n41829 ;
  assign y9880 = ~1'b0 ;
  assign y9881 = ~1'b0 ;
  assign y9882 = ~n41830 ;
  assign y9883 = n41831 ;
  assign y9884 = n41835 ;
  assign y9885 = n41837 ;
  assign y9886 = n41839 ;
  assign y9887 = n41840 ;
  assign y9888 = ~n41841 ;
  assign y9889 = ~n41845 ;
  assign y9890 = n41848 ;
  assign y9891 = ~n41849 ;
  assign y9892 = ~n41851 ;
  assign y9893 = n41852 ;
  assign y9894 = ~n41855 ;
  assign y9895 = ~n41857 ;
  assign y9896 = n41861 ;
  assign y9897 = ~n41868 ;
  assign y9898 = n41869 ;
  assign y9899 = n41870 ;
  assign y9900 = ~n41873 ;
  assign y9901 = ~n41874 ;
  assign y9902 = n41878 ;
  assign y9903 = n41879 ;
  assign y9904 = ~n41881 ;
  assign y9905 = n41885 ;
  assign y9906 = ~n41887 ;
  assign y9907 = n41889 ;
  assign y9908 = ~n41891 ;
  assign y9909 = ~n41893 ;
  assign y9910 = n41899 ;
  assign y9911 = n41901 ;
  assign y9912 = n41902 ;
  assign y9913 = n41903 ;
  assign y9914 = ~1'b0 ;
  assign y9915 = n41904 ;
  assign y9916 = ~n41906 ;
  assign y9917 = ~n41908 ;
  assign y9918 = n41909 ;
  assign y9919 = ~n41910 ;
  assign y9920 = ~n41911 ;
  assign y9921 = ~n41913 ;
  assign y9922 = ~n41917 ;
  assign y9923 = ~n41918 ;
  assign y9924 = n41926 ;
  assign y9925 = ~n41929 ;
  assign y9926 = n41931 ;
  assign y9927 = ~n41932 ;
  assign y9928 = n41935 ;
  assign y9929 = ~n41942 ;
  assign y9930 = ~n41944 ;
  assign y9931 = ~n41949 ;
  assign y9932 = n41951 ;
  assign y9933 = ~n41952 ;
  assign y9934 = n41958 ;
  assign y9935 = ~n41969 ;
  assign y9936 = ~n41974 ;
  assign y9937 = ~n41982 ;
  assign y9938 = n41983 ;
  assign y9939 = ~n41986 ;
  assign y9940 = ~n41991 ;
  assign y9941 = ~n41993 ;
  assign y9942 = n41998 ;
  assign y9943 = n42000 ;
  assign y9944 = ~n42001 ;
  assign y9945 = ~n42004 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = n42007 ;
  assign y9948 = n42011 ;
  assign y9949 = n42012 ;
  assign y9950 = ~n42013 ;
  assign y9951 = n42015 ;
  assign y9952 = ~n42018 ;
  assign y9953 = ~n42019 ;
  assign y9954 = n42021 ;
  assign y9955 = ~n42026 ;
  assign y9956 = n42030 ;
  assign y9957 = ~n42034 ;
  assign y9958 = n42039 ;
  assign y9959 = n42040 ;
  assign y9960 = n42042 ;
  assign y9961 = ~1'b0 ;
  assign y9962 = ~n42047 ;
  assign y9963 = ~n42051 ;
  assign y9964 = ~n42053 ;
  assign y9965 = ~n42055 ;
  assign y9966 = ~n42057 ;
  assign y9967 = n42058 ;
  assign y9968 = n42060 ;
  assign y9969 = ~n42064 ;
  assign y9970 = ~n42068 ;
  assign y9971 = n42071 ;
  assign y9972 = ~n42072 ;
  assign y9973 = n42073 ;
  assign y9974 = ~n42079 ;
  assign y9975 = ~n42081 ;
  assign y9976 = n42082 ;
  assign y9977 = ~n42084 ;
  assign y9978 = n42085 ;
  assign y9979 = n42087 ;
  assign y9980 = n42088 ;
  assign y9981 = n42091 ;
  assign y9982 = ~n42093 ;
  assign y9983 = ~1'b0 ;
  assign y9984 = n42094 ;
  assign y9985 = ~n42095 ;
  assign y9986 = ~n42096 ;
  assign y9987 = ~n42097 ;
  assign y9988 = ~n42102 ;
  assign y9989 = ~n42103 ;
  assign y9990 = ~1'b0 ;
  assign y9991 = ~n42104 ;
  assign y9992 = ~n42106 ;
  assign y9993 = ~n42107 ;
  assign y9994 = n42109 ;
  assign y9995 = n42110 ;
  assign y9996 = n42111 ;
  assign y9997 = ~n42112 ;
  assign y9998 = ~1'b0 ;
  assign y9999 = n42116 ;
  assign y10000 = ~n42120 ;
  assign y10001 = n42121 ;
  assign y10002 = n42124 ;
  assign y10003 = n42128 ;
  assign y10004 = ~n42129 ;
  assign y10005 = ~n42138 ;
  assign y10006 = ~1'b0 ;
  assign y10007 = ~n42139 ;
  assign y10008 = ~n42142 ;
  assign y10009 = n42144 ;
  assign y10010 = n42146 ;
  assign y10011 = ~n42151 ;
  assign y10012 = ~n42156 ;
  assign y10013 = n42157 ;
  assign y10014 = n42160 ;
  assign y10015 = ~n42164 ;
  assign y10016 = ~n42171 ;
  assign y10017 = ~n42176 ;
  assign y10018 = n42177 ;
  assign y10019 = ~n42179 ;
  assign y10020 = n42185 ;
  assign y10021 = n42187 ;
  assign y10022 = ~n42189 ;
  assign y10023 = n42192 ;
  assign y10024 = ~n42193 ;
  assign y10025 = n42195 ;
  assign y10026 = ~1'b0 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = ~n42196 ;
  assign y10029 = n42197 ;
  assign y10030 = n42198 ;
  assign y10031 = ~n42199 ;
  assign y10032 = ~n42200 ;
  assign y10033 = ~n42201 ;
  assign y10034 = ~n42203 ;
  assign y10035 = ~n42204 ;
  assign y10036 = ~n42205 ;
  assign y10037 = ~n42206 ;
  assign y10038 = n42208 ;
  assign y10039 = n42210 ;
  assign y10040 = ~n42211 ;
  assign y10041 = n42212 ;
  assign y10042 = n42213 ;
  assign y10043 = ~n42215 ;
  assign y10044 = ~n42217 ;
  assign y10045 = ~n42223 ;
  assign y10046 = ~n42224 ;
  assign y10047 = n42227 ;
  assign y10048 = ~n42234 ;
  assign y10049 = ~n42238 ;
  assign y10050 = n42239 ;
  assign y10051 = ~n42241 ;
  assign y10052 = n42246 ;
  assign y10053 = ~1'b0 ;
  assign y10054 = ~1'b0 ;
  assign y10055 = ~n42247 ;
  assign y10056 = n42248 ;
  assign y10057 = ~n42250 ;
  assign y10058 = n42252 ;
  assign y10059 = ~n42255 ;
  assign y10060 = n42260 ;
  assign y10061 = ~n42271 ;
  assign y10062 = ~1'b0 ;
  assign y10063 = ~n42273 ;
  assign y10064 = ~n42277 ;
  assign y10065 = n42278 ;
  assign y10066 = n42280 ;
  assign y10067 = ~n42285 ;
  assign y10068 = ~n42287 ;
  assign y10069 = n42289 ;
  assign y10070 = ~n42292 ;
  assign y10071 = ~n42294 ;
  assign y10072 = ~n42298 ;
  assign y10073 = n42301 ;
  assign y10074 = ~n42302 ;
  assign y10075 = ~n42303 ;
  assign y10076 = ~n42304 ;
  assign y10077 = n42307 ;
  assign y10078 = n42309 ;
  assign y10079 = n42315 ;
  assign y10080 = ~n42319 ;
  assign y10081 = ~n42321 ;
  assign y10082 = 1'b0 ;
  assign y10083 = ~n42322 ;
  assign y10084 = ~n42331 ;
  assign y10085 = ~n42332 ;
  assign y10086 = ~n42334 ;
  assign y10087 = n42336 ;
  assign y10088 = n42342 ;
  assign y10089 = ~n42349 ;
  assign y10090 = n42350 ;
  assign y10091 = ~n42352 ;
  assign y10092 = n42353 ;
  assign y10093 = ~n42354 ;
  assign y10094 = n42359 ;
  assign y10095 = n42363 ;
  assign y10096 = ~n42370 ;
  assign y10097 = ~n42371 ;
  assign y10098 = ~n42375 ;
  assign y10099 = ~n42380 ;
  assign y10100 = ~1'b0 ;
  assign y10101 = ~n42381 ;
  assign y10102 = n42385 ;
  assign y10103 = ~n42388 ;
  assign y10104 = n42389 ;
  assign y10105 = ~n42390 ;
  assign y10106 = ~n42393 ;
  assign y10107 = ~n42396 ;
  assign y10108 = ~n42399 ;
  assign y10109 = n42401 ;
  assign y10110 = ~n42405 ;
  assign y10111 = n42407 ;
  assign y10112 = n42408 ;
  assign y10113 = n42418 ;
  assign y10114 = ~n42419 ;
  assign y10115 = ~n42421 ;
  assign y10116 = n42422 ;
  assign y10117 = n42426 ;
  assign y10118 = ~n42433 ;
  assign y10119 = n42438 ;
  assign y10120 = ~n42439 ;
  assign y10121 = n42440 ;
  assign y10122 = n42442 ;
  assign y10123 = ~n42443 ;
  assign y10124 = ~n42446 ;
  assign y10125 = n42448 ;
  assign y10126 = n42451 ;
  assign y10127 = ~n19361 ;
  assign y10128 = n42452 ;
  assign y10129 = n42454 ;
  assign y10130 = n42455 ;
  assign y10131 = ~n42457 ;
  assign y10132 = ~n42460 ;
  assign y10133 = ~n42462 ;
  assign y10134 = ~n42463 ;
  assign y10135 = ~n42464 ;
  assign y10136 = ~n42466 ;
  assign y10137 = ~n42470 ;
  assign y10138 = ~n42472 ;
  assign y10139 = n42474 ;
  assign y10140 = ~n42476 ;
  assign y10141 = ~n42480 ;
  assign y10142 = ~n42481 ;
  assign y10143 = n42482 ;
  assign y10144 = ~n42485 ;
  assign y10145 = ~n42486 ;
  assign y10146 = n42487 ;
  assign y10147 = n42489 ;
  assign y10148 = n42493 ;
  assign y10149 = n42497 ;
  assign y10150 = n42501 ;
  assign y10151 = ~n42504 ;
  assign y10152 = n42507 ;
  assign y10153 = n42508 ;
  assign y10154 = n42511 ;
  assign y10155 = n42513 ;
  assign y10156 = n42517 ;
  assign y10157 = n42519 ;
  assign y10158 = n42522 ;
  assign y10159 = ~n42525 ;
  assign y10160 = n42527 ;
  assign y10161 = ~n42528 ;
  assign y10162 = ~n42530 ;
  assign y10163 = ~n42531 ;
  assign y10164 = ~n42535 ;
  assign y10165 = n42536 ;
  assign y10166 = n42539 ;
  assign y10167 = ~n42540 ;
  assign y10168 = n42545 ;
  assign y10169 = ~n42546 ;
  assign y10170 = ~n42547 ;
  assign y10171 = n42548 ;
  assign y10172 = n42549 ;
  assign y10173 = ~n42553 ;
  assign y10174 = n42555 ;
  assign y10175 = n42562 ;
  assign y10176 = n42564 ;
  assign y10177 = ~n42568 ;
  assign y10178 = n42569 ;
  assign y10179 = n42571 ;
  assign y10180 = n42572 ;
  assign y10181 = n42573 ;
  assign y10182 = n42574 ;
  assign y10183 = n42575 ;
  assign y10184 = ~n42578 ;
  assign y10185 = ~1'b0 ;
  assign y10186 = ~n42588 ;
  assign y10187 = ~n42591 ;
  assign y10188 = n42594 ;
  assign y10189 = ~n42595 ;
  assign y10190 = n42598 ;
  assign y10191 = ~n42600 ;
  assign y10192 = ~n42601 ;
  assign y10193 = n42604 ;
  assign y10194 = n42607 ;
  assign y10195 = ~n42609 ;
  assign y10196 = ~n42612 ;
  assign y10197 = ~n42613 ;
  assign y10198 = ~n42615 ;
  assign y10199 = n42617 ;
  assign y10200 = ~n42619 ;
  assign y10201 = ~n42622 ;
  assign y10202 = n42623 ;
  assign y10203 = ~n42626 ;
  assign y10204 = n42627 ;
  assign y10205 = n42629 ;
  assign y10206 = ~n42631 ;
  assign y10207 = n42633 ;
  assign y10208 = ~n42637 ;
  assign y10209 = ~n42642 ;
  assign y10210 = ~n42643 ;
  assign y10211 = ~n42645 ;
  assign y10212 = ~n42650 ;
  assign y10213 = ~n42651 ;
  assign y10214 = ~n42653 ;
  assign y10215 = ~n42655 ;
  assign y10216 = ~n42658 ;
  assign y10217 = n42660 ;
  assign y10218 = n42663 ;
  assign y10219 = ~n42665 ;
  assign y10220 = n42666 ;
  assign y10221 = n42667 ;
  assign y10222 = n42669 ;
  assign y10223 = ~n42670 ;
  assign y10224 = ~n42675 ;
  assign y10225 = n42676 ;
  assign y10226 = ~1'b0 ;
  assign y10227 = ~1'b0 ;
  assign y10228 = ~n42678 ;
  assign y10229 = n42679 ;
  assign y10230 = ~n42680 ;
  assign y10231 = ~n42688 ;
  assign y10232 = n42691 ;
  assign y10233 = ~n42693 ;
  assign y10234 = ~1'b0 ;
  assign y10235 = n42700 ;
  assign y10236 = ~n42701 ;
  assign y10237 = n42702 ;
  assign y10238 = n42703 ;
  assign y10239 = n42705 ;
  assign y10240 = n42709 ;
  assign y10241 = ~n42710 ;
  assign y10242 = ~n42720 ;
  assign y10243 = n42722 ;
  assign y10244 = ~n42724 ;
  assign y10245 = n42726 ;
  assign y10246 = n42727 ;
  assign y10247 = ~n42730 ;
  assign y10248 = ~n42731 ;
  assign y10249 = ~n42732 ;
  assign y10250 = n42737 ;
  assign y10251 = n42739 ;
  assign y10252 = ~n42740 ;
  assign y10253 = ~n42744 ;
  assign y10254 = ~n42745 ;
  assign y10255 = n42747 ;
  assign y10256 = ~n42748 ;
  assign y10257 = n42751 ;
  assign y10258 = n42752 ;
  assign y10259 = n42753 ;
  assign y10260 = n42756 ;
  assign y10261 = ~n42763 ;
  assign y10262 = n42764 ;
  assign y10263 = n42769 ;
  assign y10264 = ~n42774 ;
  assign y10265 = n42775 ;
  assign y10266 = ~n42777 ;
  assign y10267 = n42779 ;
  assign y10268 = n42780 ;
  assign y10269 = n42782 ;
  assign y10270 = ~n42785 ;
  assign y10271 = n42786 ;
  assign y10272 = ~n42793 ;
  assign y10273 = ~n42798 ;
  assign y10274 = ~n42804 ;
  assign y10275 = ~1'b0 ;
  assign y10276 = ~1'b0 ;
  assign y10277 = ~n42806 ;
  assign y10278 = n42808 ;
  assign y10279 = n42814 ;
  assign y10280 = ~n42815 ;
  assign y10281 = n42816 ;
  assign y10282 = n42818 ;
  assign y10283 = n42819 ;
  assign y10284 = ~n42820 ;
  assign y10285 = n42826 ;
  assign y10286 = ~n42827 ;
  assign y10287 = n42831 ;
  assign y10288 = ~n42832 ;
  assign y10289 = ~n42837 ;
  assign y10290 = n42838 ;
  assign y10291 = ~n42839 ;
  assign y10292 = ~n42843 ;
  assign y10293 = ~n5308 ;
  assign y10294 = n42845 ;
  assign y10295 = ~n42849 ;
  assign y10296 = n42853 ;
  assign y10297 = n42861 ;
  assign y10298 = ~n42865 ;
  assign y10299 = ~n42870 ;
  assign y10300 = n42873 ;
  assign y10301 = ~n42876 ;
  assign y10302 = n42878 ;
  assign y10303 = ~n42882 ;
  assign y10304 = n42886 ;
  assign y10305 = ~1'b0 ;
  assign y10306 = ~1'b0 ;
  assign y10307 = ~n42893 ;
  assign y10308 = ~n42894 ;
  assign y10309 = ~n42895 ;
  assign y10310 = n42897 ;
  assign y10311 = ~n42900 ;
  assign y10312 = ~n42901 ;
  assign y10313 = ~n42902 ;
  assign y10314 = n42906 ;
  assign y10315 = ~n42908 ;
  assign y10316 = ~n42912 ;
  assign y10317 = ~n42913 ;
  assign y10318 = ~n42922 ;
  assign y10319 = n42923 ;
  assign y10320 = ~1'b0 ;
  assign y10321 = n42925 ;
  assign y10322 = n42926 ;
  assign y10323 = n42930 ;
  assign y10324 = ~n42938 ;
  assign y10325 = ~1'b0 ;
  assign y10326 = ~n42944 ;
  assign y10327 = ~n42945 ;
  assign y10328 = n42949 ;
  assign y10329 = n42950 ;
  assign y10330 = ~n42952 ;
  assign y10331 = n42957 ;
  assign y10332 = ~n42959 ;
  assign y10333 = n42961 ;
  assign y10334 = n42962 ;
  assign y10335 = ~n42965 ;
  assign y10336 = ~n42968 ;
  assign y10337 = n42969 ;
  assign y10338 = ~n42971 ;
  assign y10339 = n42973 ;
  assign y10340 = ~n42977 ;
  assign y10341 = ~n42979 ;
  assign y10342 = ~n42982 ;
  assign y10343 = ~n42984 ;
  assign y10344 = ~n42989 ;
  assign y10345 = n42993 ;
  assign y10346 = n42998 ;
  assign y10347 = ~n43001 ;
  assign y10348 = ~n43002 ;
  assign y10349 = ~n43003 ;
  assign y10350 = n43008 ;
  assign y10351 = ~n43012 ;
  assign y10352 = n43018 ;
  assign y10353 = ~n43021 ;
  assign y10354 = n43022 ;
  assign y10355 = n43027 ;
  assign y10356 = n43030 ;
  assign y10357 = n43032 ;
  assign y10358 = n43034 ;
  assign y10359 = ~n43036 ;
  assign y10360 = n43039 ;
  assign y10361 = n43041 ;
  assign y10362 = n43043 ;
  assign y10363 = n43045 ;
  assign y10364 = ~n43046 ;
  assign y10365 = n43047 ;
  assign y10366 = n43053 ;
  assign y10367 = n43054 ;
  assign y10368 = ~n43057 ;
  assign y10369 = ~n43066 ;
  assign y10370 = ~n19777 ;
  assign y10371 = ~n43068 ;
  assign y10372 = ~n43070 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = ~n43073 ;
  assign y10375 = ~n43079 ;
  assign y10376 = ~n43083 ;
  assign y10377 = n43084 ;
  assign y10378 = ~n43086 ;
  assign y10379 = n43087 ;
  assign y10380 = ~n43092 ;
  assign y10381 = n43095 ;
  assign y10382 = ~n43099 ;
  assign y10383 = ~n43102 ;
  assign y10384 = n43105 ;
  assign y10385 = ~n43106 ;
  assign y10386 = n43110 ;
  assign y10387 = n43111 ;
  assign y10388 = n43114 ;
  assign y10389 = n43116 ;
  assign y10390 = ~n43118 ;
  assign y10391 = ~n43119 ;
  assign y10392 = ~1'b0 ;
  assign y10393 = n43120 ;
  assign y10394 = n43121 ;
  assign y10395 = n43122 ;
  assign y10396 = n43124 ;
  assign y10397 = ~n43127 ;
  assign y10398 = n43128 ;
  assign y10399 = ~n43130 ;
  assign y10400 = ~n43131 ;
  assign y10401 = ~n43134 ;
  assign y10402 = ~n43135 ;
  assign y10403 = ~n43136 ;
  assign y10404 = n43138 ;
  assign y10405 = ~n43143 ;
  assign y10406 = n43144 ;
  assign y10407 = ~n43145 ;
  assign y10408 = ~n43148 ;
  assign y10409 = ~n43149 ;
  assign y10410 = ~n43150 ;
  assign y10411 = n43152 ;
  assign y10412 = ~n43158 ;
  assign y10413 = n43163 ;
  assign y10414 = ~n43165 ;
  assign y10415 = n43166 ;
  assign y10416 = ~n43174 ;
  assign y10417 = n43175 ;
  assign y10418 = n43178 ;
  assign y10419 = ~n43181 ;
  assign y10420 = ~n43182 ;
  assign y10421 = ~n43184 ;
  assign y10422 = ~n43187 ;
  assign y10423 = n43189 ;
  assign y10424 = ~n43192 ;
  assign y10425 = n43194 ;
  assign y10426 = n43195 ;
  assign y10427 = ~n43199 ;
  assign y10428 = n43200 ;
  assign y10429 = n43204 ;
  assign y10430 = ~n43209 ;
  assign y10431 = n43214 ;
  assign y10432 = n43216 ;
  assign y10433 = ~n43219 ;
  assign y10434 = n43220 ;
  assign y10435 = ~n43223 ;
  assign y10436 = n43224 ;
  assign y10437 = ~n43226 ;
  assign y10438 = ~n43227 ;
  assign y10439 = ~n43230 ;
  assign y10440 = ~n43232 ;
  assign y10441 = ~n43233 ;
  assign y10442 = n43237 ;
  assign y10443 = ~n43239 ;
  assign y10444 = n43241 ;
  assign y10445 = ~n43244 ;
  assign y10446 = ~n43245 ;
  assign y10447 = ~n43248 ;
  assign y10448 = ~n43251 ;
  assign y10449 = n43254 ;
  assign y10450 = n43257 ;
  assign y10451 = ~n43261 ;
  assign y10452 = n43263 ;
  assign y10453 = ~n43265 ;
  assign y10454 = n43266 ;
  assign y10455 = ~n43272 ;
  assign y10456 = n43280 ;
  assign y10457 = ~n43281 ;
  assign y10458 = n43283 ;
  assign y10459 = n43286 ;
  assign y10460 = ~1'b0 ;
  assign y10461 = n43291 ;
  assign y10462 = ~n43293 ;
  assign y10463 = ~n43294 ;
  assign y10464 = n43296 ;
  assign y10465 = ~n43299 ;
  assign y10466 = ~n43300 ;
  assign y10467 = n43301 ;
  assign y10468 = ~1'b0 ;
  assign y10469 = ~n43309 ;
  assign y10470 = ~n43311 ;
  assign y10471 = n43313 ;
  assign y10472 = n43317 ;
  assign y10473 = ~n43320 ;
  assign y10474 = n43321 ;
  assign y10475 = ~n43325 ;
  assign y10476 = n43328 ;
  assign y10477 = ~1'b0 ;
  assign y10478 = ~n43330 ;
  assign y10479 = n43331 ;
  assign y10480 = n43335 ;
  assign y10481 = n43338 ;
  assign y10482 = n43339 ;
  assign y10483 = n43342 ;
  assign y10484 = n43346 ;
  assign y10485 = n43347 ;
  assign y10486 = ~n43349 ;
  assign y10487 = ~1'b0 ;
  assign y10488 = n43350 ;
  assign y10489 = n43351 ;
  assign y10490 = ~n43353 ;
  assign y10491 = n43355 ;
  assign y10492 = ~n43361 ;
  assign y10493 = ~n43362 ;
  assign y10494 = ~n43365 ;
  assign y10495 = n43368 ;
  assign y10496 = ~n43377 ;
  assign y10497 = ~n43379 ;
  assign y10498 = n43384 ;
  assign y10499 = ~n43386 ;
  assign y10500 = ~n43389 ;
  assign y10501 = ~n43390 ;
  assign y10502 = ~n43395 ;
  assign y10503 = n43396 ;
  assign y10504 = n43405 ;
  assign y10505 = ~n43407 ;
  assign y10506 = n43409 ;
  assign y10507 = ~n43412 ;
  assign y10508 = ~n43417 ;
  assign y10509 = ~n43420 ;
  assign y10510 = n43422 ;
  assign y10511 = ~n43423 ;
  assign y10512 = n43425 ;
  assign y10513 = ~n43430 ;
  assign y10514 = ~n43433 ;
  assign y10515 = ~n43436 ;
  assign y10516 = ~n43439 ;
  assign y10517 = n43444 ;
  assign y10518 = ~n43447 ;
  assign y10519 = ~1'b0 ;
  assign y10520 = n43449 ;
  assign y10521 = n43450 ;
  assign y10522 = n43451 ;
  assign y10523 = n43452 ;
  assign y10524 = n43456 ;
  assign y10525 = ~n43459 ;
  assign y10526 = n43460 ;
  assign y10527 = n43466 ;
  assign y10528 = ~n43467 ;
  assign y10529 = n43476 ;
  assign y10530 = ~n43478 ;
  assign y10531 = ~n43480 ;
  assign y10532 = n43482 ;
  assign y10533 = ~n43483 ;
  assign y10534 = n43489 ;
  assign y10535 = ~n43492 ;
  assign y10536 = ~n43494 ;
  assign y10537 = ~n43499 ;
  assign y10538 = n43500 ;
  assign y10539 = n43501 ;
  assign y10540 = n43502 ;
  assign y10541 = n43505 ;
  assign y10542 = ~1'b0 ;
  assign y10543 = n43506 ;
  assign y10544 = n43508 ;
  assign y10545 = ~n43510 ;
  assign y10546 = ~n43512 ;
  assign y10547 = ~n43515 ;
  assign y10548 = n43516 ;
  assign y10549 = n43517 ;
  assign y10550 = n43520 ;
  assign y10551 = ~n43527 ;
  assign y10552 = ~n43528 ;
  assign y10553 = ~n43529 ;
  assign y10554 = n43530 ;
  assign y10555 = ~n43532 ;
  assign y10556 = n43535 ;
  assign y10557 = n43536 ;
  assign y10558 = ~n43537 ;
  assign y10559 = ~1'b0 ;
  assign y10560 = n43544 ;
  assign y10561 = n43545 ;
  assign y10562 = n43547 ;
  assign y10563 = n43550 ;
  assign y10564 = ~n43553 ;
  assign y10565 = ~1'b0 ;
  assign y10566 = ~1'b0 ;
  assign y10567 = ~n43556 ;
  assign y10568 = ~n43560 ;
  assign y10569 = ~n43562 ;
  assign y10570 = n43565 ;
  assign y10571 = ~n43567 ;
  assign y10572 = ~n43572 ;
  assign y10573 = n43574 ;
  assign y10574 = n43575 ;
  assign y10575 = ~n43576 ;
  assign y10576 = n43582 ;
  assign y10577 = ~n43585 ;
  assign y10578 = n43587 ;
  assign y10579 = n43589 ;
  assign y10580 = n43590 ;
  assign y10581 = ~n43591 ;
  assign y10582 = ~1'b0 ;
  assign y10583 = n43592 ;
  assign y10584 = ~n43593 ;
  assign y10585 = ~n43594 ;
  assign y10586 = n43595 ;
  assign y10587 = ~n43598 ;
  assign y10588 = n43601 ;
  assign y10589 = ~n43603 ;
  assign y10590 = ~n43605 ;
  assign y10591 = n43606 ;
  assign y10592 = n43613 ;
  assign y10593 = ~n43617 ;
  assign y10594 = ~n43620 ;
  assign y10595 = n43624 ;
  assign y10596 = n43626 ;
  assign y10597 = ~n43628 ;
  assign y10598 = ~n43629 ;
  assign y10599 = n43631 ;
  assign y10600 = ~n43633 ;
  assign y10601 = n43634 ;
  assign y10602 = ~n43635 ;
  assign y10603 = n43638 ;
  assign y10604 = ~n43640 ;
  assign y10605 = ~n43644 ;
  assign y10606 = ~n43645 ;
  assign y10607 = ~n43646 ;
  assign y10608 = ~n43648 ;
  assign y10609 = n43651 ;
  assign y10610 = ~n43653 ;
  assign y10611 = n43656 ;
  assign y10612 = n43658 ;
  assign y10613 = n43663 ;
  assign y10614 = ~n43664 ;
  assign y10615 = n43665 ;
  assign y10616 = n43667 ;
  assign y10617 = n43671 ;
  assign y10618 = n43676 ;
  assign y10619 = ~n43680 ;
  assign y10620 = n43683 ;
  assign y10621 = n43689 ;
  assign y10622 = ~n43693 ;
  assign y10623 = ~n43698 ;
  assign y10624 = n43699 ;
  assign y10625 = n43701 ;
  assign y10626 = ~n43703 ;
  assign y10627 = ~n43704 ;
  assign y10628 = n43706 ;
  assign y10629 = ~n43714 ;
  assign y10630 = n43717 ;
  assign y10631 = n43718 ;
  assign y10632 = ~n43722 ;
  assign y10633 = ~n43727 ;
  assign y10634 = ~n43728 ;
  assign y10635 = ~n43731 ;
  assign y10636 = n43733 ;
  assign y10637 = ~n43734 ;
  assign y10638 = ~n43735 ;
  assign y10639 = n43741 ;
  assign y10640 = ~n43747 ;
  assign y10641 = ~n43748 ;
  assign y10642 = n43753 ;
  assign y10643 = ~n43757 ;
  assign y10644 = ~n43761 ;
  assign y10645 = n43767 ;
  assign y10646 = ~n43769 ;
  assign y10647 = ~n43776 ;
  assign y10648 = n43779 ;
  assign y10649 = n43782 ;
  assign y10650 = ~1'b0 ;
  assign y10651 = n43784 ;
  assign y10652 = ~n43791 ;
  assign y10653 = n43792 ;
  assign y10654 = ~n43793 ;
  assign y10655 = ~n43796 ;
  assign y10656 = n43797 ;
  assign y10657 = ~n43805 ;
  assign y10658 = ~n43807 ;
  assign y10659 = n43809 ;
  assign y10660 = ~n43819 ;
  assign y10661 = n43820 ;
  assign y10662 = ~n43822 ;
  assign y10663 = n43831 ;
  assign y10664 = n43832 ;
  assign y10665 = ~n43833 ;
  assign y10666 = n43838 ;
  assign y10667 = ~n43840 ;
  assign y10668 = n43843 ;
  assign y10669 = n43844 ;
  assign y10670 = ~n43846 ;
  assign y10671 = n43847 ;
  assign y10672 = n43849 ;
  assign y10673 = n43850 ;
  assign y10674 = ~n43853 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = ~n43859 ;
  assign y10677 = n43862 ;
  assign y10678 = ~n43863 ;
  assign y10679 = n43865 ;
  assign y10680 = ~n43867 ;
  assign y10681 = n43868 ;
  assign y10682 = n43870 ;
  assign y10683 = ~n43872 ;
  assign y10684 = n43873 ;
  assign y10685 = ~n43874 ;
  assign y10686 = ~n43878 ;
  assign y10687 = ~n43879 ;
  assign y10688 = ~n43882 ;
  assign y10689 = ~n43884 ;
  assign y10690 = n43886 ;
  assign y10691 = ~n43889 ;
  assign y10692 = n43890 ;
  assign y10693 = n43893 ;
  assign y10694 = ~n43899 ;
  assign y10695 = ~n43901 ;
  assign y10696 = n43902 ;
  assign y10697 = ~n43903 ;
  assign y10698 = n43907 ;
  assign y10699 = ~n43910 ;
  assign y10700 = ~n43911 ;
  assign y10701 = n43912 ;
  assign y10702 = ~n43913 ;
  assign y10703 = ~n43914 ;
  assign y10704 = n43915 ;
  assign y10705 = ~n43916 ;
  assign y10706 = ~n43917 ;
  assign y10707 = n43919 ;
  assign y10708 = ~n43920 ;
  assign y10709 = ~n43922 ;
  assign y10710 = ~n43923 ;
  assign y10711 = n43924 ;
  assign y10712 = ~n43927 ;
  assign y10713 = ~n43930 ;
  assign y10714 = n43931 ;
  assign y10715 = n43934 ;
  assign y10716 = ~n43941 ;
  assign y10717 = n43944 ;
  assign y10718 = ~n43945 ;
  assign y10719 = ~n43949 ;
  assign y10720 = n43951 ;
  assign y10721 = n43953 ;
  assign y10722 = n43958 ;
  assign y10723 = ~1'b0 ;
  assign y10724 = ~n43960 ;
  assign y10725 = ~n43961 ;
  assign y10726 = ~n43962 ;
  assign y10727 = n43965 ;
  assign y10728 = ~n43966 ;
  assign y10729 = n43969 ;
  assign y10730 = ~n43971 ;
  assign y10731 = ~n43973 ;
  assign y10732 = ~n43975 ;
  assign y10733 = ~n43979 ;
  assign y10734 = ~n43980 ;
  assign y10735 = ~n43983 ;
  assign y10736 = ~1'b0 ;
  assign y10737 = n43985 ;
  assign y10738 = ~n43988 ;
  assign y10739 = n43990 ;
  assign y10740 = n43992 ;
  assign y10741 = ~n43995 ;
  assign y10742 = ~n44000 ;
  assign y10743 = n44002 ;
  assign y10744 = ~n44005 ;
  assign y10745 = n44006 ;
  assign y10746 = n44007 ;
  assign y10747 = ~1'b0 ;
  assign y10748 = ~n44008 ;
  assign y10749 = n44009 ;
  assign y10750 = ~n44010 ;
  assign y10751 = n44018 ;
  assign y10752 = n44022 ;
  assign y10753 = ~n44027 ;
  assign y10754 = n44030 ;
  assign y10755 = ~n44033 ;
  assign y10756 = ~n44035 ;
  assign y10757 = ~1'b0 ;
  assign y10758 = ~n44038 ;
  assign y10759 = n44039 ;
  assign y10760 = n44042 ;
  assign y10761 = ~n44045 ;
  assign y10762 = n44046 ;
  assign y10763 = n44047 ;
  assign y10764 = n44049 ;
  assign y10765 = n44051 ;
  assign y10766 = ~n44052 ;
  assign y10767 = n44055 ;
  assign y10768 = ~n44056 ;
  assign y10769 = n44058 ;
  assign y10770 = n19752 ;
  assign y10771 = n44062 ;
  assign y10772 = ~n44064 ;
  assign y10773 = n44065 ;
  assign y10774 = ~n44067 ;
  assign y10775 = ~n44069 ;
  assign y10776 = n44076 ;
  assign y10777 = ~n44078 ;
  assign y10778 = n44080 ;
  assign y10779 = n44084 ;
  assign y10780 = ~n44085 ;
  assign y10781 = n44086 ;
  assign y10782 = ~n44087 ;
  assign y10783 = ~n44088 ;
  assign y10784 = ~n44089 ;
  assign y10785 = n44091 ;
  assign y10786 = n44093 ;
  assign y10787 = n44096 ;
  assign y10788 = n44099 ;
  assign y10789 = n5884 ;
  assign y10790 = ~n44102 ;
  assign y10791 = ~n44106 ;
  assign y10792 = ~n44112 ;
  assign y10793 = n44115 ;
  assign y10794 = n44118 ;
  assign y10795 = ~n44119 ;
  assign y10796 = ~1'b0 ;
  assign y10797 = ~n44122 ;
  assign y10798 = n44125 ;
  assign y10799 = n44126 ;
  assign y10800 = n44129 ;
  assign y10801 = n44130 ;
  assign y10802 = ~n44132 ;
  assign y10803 = ~n44136 ;
  assign y10804 = n44137 ;
  assign y10805 = n44138 ;
  assign y10806 = ~n44139 ;
  assign y10807 = n44142 ;
  assign y10808 = n44144 ;
  assign y10809 = ~n44146 ;
  assign y10810 = ~n44150 ;
  assign y10811 = n44152 ;
  assign y10812 = ~n44155 ;
  assign y10813 = ~n44160 ;
  assign y10814 = n44161 ;
  assign y10815 = ~n44163 ;
  assign y10816 = n44166 ;
  assign y10817 = ~n44169 ;
  assign y10818 = n44170 ;
  assign y10819 = ~n44172 ;
  assign y10820 = ~1'b0 ;
  assign y10821 = n44175 ;
  assign y10822 = n44176 ;
  assign y10823 = n44178 ;
  assign y10824 = n44180 ;
  assign y10825 = ~n44181 ;
  assign y10826 = n44182 ;
  assign y10827 = ~n44188 ;
  assign y10828 = ~n44191 ;
  assign y10829 = ~n44196 ;
  assign y10830 = ~n44200 ;
  assign y10831 = n44201 ;
  assign y10832 = ~n44204 ;
  assign y10833 = n44206 ;
  assign y10834 = ~1'b0 ;
  assign y10835 = n44208 ;
  assign y10836 = n44214 ;
  assign y10837 = ~n44215 ;
  assign y10838 = n44217 ;
  assign y10839 = ~n44219 ;
  assign y10840 = ~n44224 ;
  assign y10841 = ~n44226 ;
  assign y10842 = n44228 ;
  assign y10843 = ~n44230 ;
  assign y10844 = ~n44233 ;
  assign y10845 = ~n44234 ;
  assign y10846 = ~n44237 ;
  assign y10847 = ~n44238 ;
  assign y10848 = ~n44242 ;
  assign y10849 = n44243 ;
  assign y10850 = ~n44247 ;
  assign y10851 = ~n44254 ;
  assign y10852 = n44259 ;
  assign y10853 = n44263 ;
  assign y10854 = n44264 ;
  assign y10855 = n44266 ;
  assign y10856 = ~n44267 ;
  assign y10857 = ~n44273 ;
  assign y10858 = n44274 ;
  assign y10859 = n44279 ;
  assign y10860 = ~n44281 ;
  assign y10861 = ~n44285 ;
  assign y10862 = n44291 ;
  assign y10863 = ~n44292 ;
  assign y10864 = ~n44293 ;
  assign y10865 = ~n44294 ;
  assign y10866 = n44299 ;
  assign y10867 = ~n44300 ;
  assign y10868 = ~n44302 ;
  assign y10869 = ~1'b0 ;
  assign y10870 = ~n44304 ;
  assign y10871 = ~n44306 ;
  assign y10872 = ~n44310 ;
  assign y10873 = ~n44315 ;
  assign y10874 = n44317 ;
  assign y10875 = ~n44319 ;
  assign y10876 = n44321 ;
  assign y10877 = ~n44330 ;
  assign y10878 = ~n44331 ;
  assign y10879 = ~n44333 ;
  assign y10880 = ~n44337 ;
  assign y10881 = n44341 ;
  assign y10882 = n44342 ;
  assign y10883 = n44343 ;
  assign y10884 = ~n44344 ;
  assign y10885 = ~n44345 ;
  assign y10886 = n44349 ;
  assign y10887 = n44351 ;
  assign y10888 = n44353 ;
  assign y10889 = n44354 ;
  assign y10890 = ~n44356 ;
  assign y10891 = ~n44358 ;
  assign y10892 = n44360 ;
  assign y10893 = n44361 ;
  assign y10894 = ~n44363 ;
  assign y10895 = n44370 ;
  assign y10896 = n44371 ;
  assign y10897 = ~n44372 ;
  assign y10898 = ~n44373 ;
  assign y10899 = n44377 ;
  assign y10900 = n44380 ;
  assign y10901 = n44381 ;
  assign y10902 = n44384 ;
  assign y10903 = ~1'b0 ;
  assign y10904 = n44385 ;
  assign y10905 = ~n44386 ;
  assign y10906 = n44388 ;
  assign y10907 = ~n44390 ;
  assign y10908 = n44392 ;
  assign y10909 = n44393 ;
  assign y10910 = ~n44398 ;
  assign y10911 = n44400 ;
  assign y10912 = ~n44403 ;
  assign y10913 = ~n44407 ;
  assign y10914 = n44408 ;
  assign y10915 = ~n44410 ;
  assign y10916 = n44413 ;
  assign y10917 = ~n44416 ;
  assign y10918 = ~n44419 ;
  assign y10919 = ~n44421 ;
  assign y10920 = ~n44423 ;
  assign y10921 = ~n44424 ;
  assign y10922 = ~n44426 ;
  assign y10923 = ~n44427 ;
  assign y10924 = n44431 ;
  assign y10925 = n44434 ;
  assign y10926 = n44435 ;
  assign y10927 = n44436 ;
  assign y10928 = n44438 ;
  assign y10929 = n44444 ;
  assign y10930 = ~n44445 ;
  assign y10931 = ~n44447 ;
  assign y10932 = n44453 ;
  assign y10933 = ~n44454 ;
  assign y10934 = n44456 ;
  assign y10935 = ~n44459 ;
  assign y10936 = n44461 ;
  assign y10937 = ~n44462 ;
  assign y10938 = n44466 ;
  assign y10939 = n44470 ;
  assign y10940 = ~n44473 ;
  assign y10941 = ~n44475 ;
  assign y10942 = ~n44476 ;
  assign y10943 = n44481 ;
  assign y10944 = n44484 ;
  assign y10945 = n44486 ;
  assign y10946 = n44490 ;
  assign y10947 = ~n44493 ;
  assign y10948 = n44500 ;
  assign y10949 = ~n44508 ;
  assign y10950 = n44513 ;
  assign y10951 = n44514 ;
  assign y10952 = ~n44516 ;
  assign y10953 = ~n44518 ;
  assign y10954 = ~n44519 ;
  assign y10955 = n44520 ;
  assign y10956 = ~n44522 ;
  assign y10957 = n44524 ;
  assign y10958 = ~n44529 ;
  assign y10959 = ~n44530 ;
  assign y10960 = ~n44536 ;
  assign y10961 = ~1'b0 ;
  assign y10962 = ~n44538 ;
  assign y10963 = ~n44540 ;
  assign y10964 = n44545 ;
  assign y10965 = n44546 ;
  assign y10966 = n44549 ;
  assign y10967 = n44550 ;
  assign y10968 = ~n44553 ;
  assign y10969 = ~n44555 ;
  assign y10970 = n44556 ;
  assign y10971 = n44558 ;
  assign y10972 = ~n44560 ;
  assign y10973 = ~n44562 ;
  assign y10974 = ~n44563 ;
  assign y10975 = ~n44564 ;
  assign y10976 = ~n44566 ;
  assign y10977 = ~n44570 ;
  assign y10978 = ~n44573 ;
  assign y10979 = ~1'b0 ;
  assign y10980 = n44577 ;
  assign y10981 = ~n44581 ;
  assign y10982 = n44582 ;
  assign y10983 = n44583 ;
  assign y10984 = n44584 ;
  assign y10985 = n44590 ;
  assign y10986 = ~n44591 ;
  assign y10987 = ~n44592 ;
  assign y10988 = ~n44595 ;
  assign y10989 = ~n44601 ;
  assign y10990 = n44607 ;
  assign y10991 = ~n44609 ;
  assign y10992 = n44611 ;
  assign y10993 = ~n44615 ;
  assign y10994 = n44622 ;
  assign y10995 = ~n44623 ;
  assign y10996 = ~n44626 ;
  assign y10997 = n44627 ;
  assign y10998 = ~n44629 ;
  assign y10999 = ~1'b0 ;
  assign y11000 = ~n44630 ;
  assign y11001 = n44632 ;
  assign y11002 = n44634 ;
  assign y11003 = ~n44638 ;
  assign y11004 = ~n44643 ;
  assign y11005 = n44644 ;
  assign y11006 = n44645 ;
  assign y11007 = ~1'b0 ;
  assign y11008 = ~1'b0 ;
  assign y11009 = n44646 ;
  assign y11010 = n44651 ;
  assign y11011 = n44653 ;
  assign y11012 = ~n44655 ;
  assign y11013 = ~n44658 ;
  assign y11014 = ~n44662 ;
  assign y11015 = n44663 ;
  assign y11016 = ~n44664 ;
  assign y11017 = n44668 ;
  assign y11018 = ~n44672 ;
  assign y11019 = ~n44673 ;
  assign y11020 = n44674 ;
  assign y11021 = ~n44675 ;
  assign y11022 = n44677 ;
  assign y11023 = n44680 ;
  assign y11024 = ~n44681 ;
  assign y11025 = ~n44689 ;
  assign y11026 = n44690 ;
  assign y11027 = ~n44695 ;
  assign y11028 = n44700 ;
  assign y11029 = ~n44701 ;
  assign y11030 = ~n44702 ;
  assign y11031 = ~n44703 ;
  assign y11032 = ~n44704 ;
  assign y11033 = n44710 ;
  assign y11034 = ~n44713 ;
  assign y11035 = n44715 ;
  assign y11036 = n44720 ;
  assign y11037 = ~n44722 ;
  assign y11038 = ~n44723 ;
  assign y11039 = ~n44727 ;
  assign y11040 = ~n44729 ;
  assign y11041 = n44735 ;
  assign y11042 = n44736 ;
  assign y11043 = ~n44741 ;
  assign y11044 = ~n44743 ;
  assign y11045 = ~n44744 ;
  assign y11046 = n44747 ;
  assign y11047 = n44750 ;
  assign y11048 = ~n44752 ;
  assign y11049 = ~1'b0 ;
  assign y11050 = n44754 ;
  assign y11051 = ~n44760 ;
  assign y11052 = ~n44761 ;
  assign y11053 = n44767 ;
  assign y11054 = n44769 ;
  assign y11055 = n44770 ;
  assign y11056 = ~1'b0 ;
  assign y11057 = n44781 ;
  assign y11058 = ~n44782 ;
  assign y11059 = ~n44783 ;
  assign y11060 = n44788 ;
  assign y11061 = n44789 ;
  assign y11062 = n44792 ;
  assign y11063 = ~n44794 ;
  assign y11064 = ~n44797 ;
  assign y11065 = ~n44799 ;
  assign y11066 = ~n44803 ;
  assign y11067 = ~n44805 ;
  assign y11068 = ~n44806 ;
  assign y11069 = ~n44808 ;
  assign y11070 = ~n44811 ;
  assign y11071 = ~n44812 ;
  assign y11072 = ~n44815 ;
  assign y11073 = ~n44818 ;
  assign y11074 = ~1'b0 ;
  assign y11075 = n44823 ;
  assign y11076 = ~n44828 ;
  assign y11077 = n44829 ;
  assign y11078 = ~n44835 ;
  assign y11079 = n44840 ;
  assign y11080 = ~n44841 ;
  assign y11081 = ~1'b0 ;
  assign y11082 = n44843 ;
  assign y11083 = ~n44847 ;
  assign y11084 = ~n44849 ;
  assign y11085 = n44850 ;
  assign y11086 = ~n44852 ;
  assign y11087 = ~1'b0 ;
  assign y11088 = n44856 ;
  assign y11089 = n6132 ;
  assign y11090 = n44862 ;
  assign y11091 = n44865 ;
  assign y11092 = n44872 ;
  assign y11093 = ~n44874 ;
  assign y11094 = n44876 ;
  assign y11095 = ~n44878 ;
  assign y11096 = n44879 ;
  assign y11097 = ~n44880 ;
  assign y11098 = ~n44884 ;
  assign y11099 = n44887 ;
  assign y11100 = n44894 ;
  assign y11101 = ~n44898 ;
  assign y11102 = ~n44903 ;
  assign y11103 = ~n44904 ;
  assign y11104 = ~n44906 ;
  assign y11105 = n44908 ;
  assign y11106 = ~n44912 ;
  assign y11107 = ~n44916 ;
  assign y11108 = ~n44918 ;
  assign y11109 = ~n44920 ;
  assign y11110 = ~n44923 ;
  assign y11111 = ~n44925 ;
  assign y11112 = n44926 ;
  assign y11113 = n44929 ;
  assign y11114 = ~n44933 ;
  assign y11115 = ~n44934 ;
  assign y11116 = n44939 ;
  assign y11117 = ~n44940 ;
  assign y11118 = ~n44943 ;
  assign y11119 = n44946 ;
  assign y11120 = ~n44950 ;
  assign y11121 = n44951 ;
  assign y11122 = ~n44959 ;
  assign y11123 = ~n44961 ;
  assign y11124 = ~n44964 ;
  assign y11125 = ~n44966 ;
  assign y11126 = n44969 ;
  assign y11127 = n44970 ;
  assign y11128 = n44974 ;
  assign y11129 = ~n44979 ;
  assign y11130 = ~n44980 ;
  assign y11131 = ~n44981 ;
  assign y11132 = ~n44982 ;
  assign y11133 = n44987 ;
  assign y11134 = n44988 ;
  assign y11135 = ~n44991 ;
  assign y11136 = n44994 ;
  assign y11137 = n44995 ;
  assign y11138 = ~1'b0 ;
  assign y11139 = n45005 ;
  assign y11140 = n45006 ;
  assign y11141 = ~n45012 ;
  assign y11142 = ~n45017 ;
  assign y11143 = n45022 ;
  assign y11144 = ~n45032 ;
  assign y11145 = n45041 ;
  assign y11146 = n45043 ;
  assign y11147 = ~n45048 ;
  assign y11148 = ~n45049 ;
  assign y11149 = ~n45050 ;
  assign y11150 = ~n45058 ;
  assign y11151 = n45061 ;
  assign y11152 = ~n45064 ;
  assign y11153 = n45067 ;
  assign y11154 = n45069 ;
  assign y11155 = n45071 ;
  assign y11156 = ~n45080 ;
  assign y11157 = ~n45082 ;
  assign y11158 = ~n45085 ;
  assign y11159 = n45087 ;
  assign y11160 = ~n45090 ;
  assign y11161 = n45091 ;
  assign y11162 = n45093 ;
  assign y11163 = n45094 ;
  assign y11164 = n45102 ;
  assign y11165 = n45105 ;
  assign y11166 = n45107 ;
  assign y11167 = n45109 ;
  assign y11168 = ~n45114 ;
  assign y11169 = ~n45116 ;
  assign y11170 = ~n45119 ;
  assign y11171 = ~n45122 ;
  assign y11172 = ~n45124 ;
  assign y11173 = n45129 ;
  assign y11174 = n45131 ;
  assign y11175 = ~n45132 ;
  assign y11176 = ~n45135 ;
  assign y11177 = n45136 ;
  assign y11178 = n45146 ;
  assign y11179 = n45149 ;
  assign y11180 = ~n45154 ;
  assign y11181 = n45155 ;
  assign y11182 = n45161 ;
  assign y11183 = ~n45164 ;
  assign y11184 = ~n45167 ;
  assign y11185 = ~n45172 ;
  assign y11186 = ~n45174 ;
  assign y11187 = n45175 ;
  assign y11188 = n45176 ;
  assign y11189 = n45177 ;
  assign y11190 = ~n45181 ;
  assign y11191 = ~n45183 ;
  assign y11192 = ~n45185 ;
  assign y11193 = ~n45188 ;
  assign y11194 = n45189 ;
  assign y11195 = n45191 ;
  assign y11196 = ~n45193 ;
  assign y11197 = n45198 ;
  assign y11198 = ~n45201 ;
  assign y11199 = n45207 ;
  assign y11200 = n45208 ;
  assign y11201 = ~n45209 ;
  assign y11202 = ~n45212 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = n45217 ;
  assign y11205 = ~n45218 ;
  assign y11206 = ~n45219 ;
  assign y11207 = ~n45221 ;
  assign y11208 = ~n45222 ;
  assign y11209 = ~n45225 ;
  assign y11210 = ~n45226 ;
  assign y11211 = n45227 ;
  assign y11212 = n45228 ;
  assign y11213 = n45230 ;
  assign y11214 = ~n45231 ;
  assign y11215 = n45233 ;
  assign y11216 = n45240 ;
  assign y11217 = ~n45241 ;
  assign y11218 = n45243 ;
  assign y11219 = ~n45247 ;
  assign y11220 = n45250 ;
  assign y11221 = n45251 ;
  assign y11222 = ~n45252 ;
  assign y11223 = n45254 ;
  assign y11224 = n45255 ;
  assign y11225 = n45256 ;
  assign y11226 = n45258 ;
  assign y11227 = n45260 ;
  assign y11228 = n45261 ;
  assign y11229 = ~n45264 ;
  assign y11230 = n45266 ;
  assign y11231 = ~n45275 ;
  assign y11232 = ~n45284 ;
  assign y11233 = n45289 ;
  assign y11234 = ~n45292 ;
  assign y11235 = ~n45295 ;
  assign y11236 = ~n45296 ;
  assign y11237 = ~n45298 ;
  assign y11238 = ~n45299 ;
  assign y11239 = ~n45304 ;
  assign y11240 = ~n45306 ;
  assign y11241 = ~n45307 ;
  assign y11242 = ~n45309 ;
  assign y11243 = n45313 ;
  assign y11244 = n45315 ;
  assign y11245 = n45316 ;
  assign y11246 = ~n45322 ;
  assign y11247 = ~n45323 ;
  assign y11248 = n45324 ;
  assign y11249 = n45326 ;
  assign y11250 = ~n45329 ;
  assign y11251 = ~n45330 ;
  assign y11252 = ~n45335 ;
  assign y11253 = n45336 ;
  assign y11254 = ~n45339 ;
  assign y11255 = n45340 ;
  assign y11256 = ~n45342 ;
  assign y11257 = n45348 ;
  assign y11258 = ~n45350 ;
  assign y11259 = ~n45352 ;
  assign y11260 = ~n45355 ;
  assign y11261 = ~n45360 ;
  assign y11262 = ~n45361 ;
  assign y11263 = n45363 ;
  assign y11264 = ~n45364 ;
  assign y11265 = n45365 ;
  assign y11266 = n45366 ;
  assign y11267 = ~n45372 ;
  assign y11268 = ~n45377 ;
  assign y11269 = ~n45381 ;
  assign y11270 = n45383 ;
  assign y11271 = n45385 ;
  assign y11272 = ~n45390 ;
  assign y11273 = n45392 ;
  assign y11274 = n45395 ;
  assign y11275 = ~n45398 ;
  assign y11276 = ~n45402 ;
  assign y11277 = ~n45407 ;
  assign y11278 = ~n45408 ;
  assign y11279 = ~n45409 ;
  assign y11280 = n45411 ;
  assign y11281 = ~n45415 ;
  assign y11282 = ~n45416 ;
  assign y11283 = ~n45418 ;
  assign y11284 = ~n45422 ;
  assign y11285 = ~n45423 ;
  assign y11286 = ~n45425 ;
  assign y11287 = n45428 ;
  assign y11288 = ~n45429 ;
  assign y11289 = ~n45434 ;
  assign y11290 = n45441 ;
  assign y11291 = n45443 ;
  assign y11292 = ~n45446 ;
  assign y11293 = n45449 ;
  assign y11294 = ~n45452 ;
  assign y11295 = n45454 ;
  assign y11296 = n45455 ;
  assign y11297 = ~n45456 ;
  assign y11298 = ~n45462 ;
  assign y11299 = ~n45463 ;
  assign y11300 = n45466 ;
  assign y11301 = ~n45469 ;
  assign y11302 = ~n45471 ;
  assign y11303 = n45472 ;
  assign y11304 = ~n45476 ;
  assign y11305 = ~n45477 ;
  assign y11306 = n45479 ;
  assign y11307 = ~n45480 ;
  assign y11308 = ~n45484 ;
  assign y11309 = ~n45486 ;
  assign y11310 = ~n45489 ;
  assign y11311 = ~n45491 ;
  assign y11312 = n45492 ;
  assign y11313 = ~n45506 ;
  assign y11314 = n45507 ;
  assign y11315 = ~n45510 ;
  assign y11316 = ~n45512 ;
  assign y11317 = ~n45514 ;
  assign y11318 = ~n45522 ;
  assign y11319 = n45523 ;
  assign y11320 = ~n45525 ;
  assign y11321 = ~n45526 ;
  assign y11322 = ~n45527 ;
  assign y11323 = ~n45530 ;
  assign y11324 = ~n45532 ;
  assign y11325 = ~n45535 ;
  assign y11326 = n45536 ;
  assign y11327 = ~n45538 ;
  assign y11328 = ~n45541 ;
  assign y11329 = n45545 ;
  assign y11330 = n45552 ;
  assign y11331 = n45554 ;
  assign y11332 = ~n45559 ;
  assign y11333 = n45561 ;
  assign y11334 = n45564 ;
  assign y11335 = ~1'b0 ;
  assign y11336 = ~n45566 ;
  assign y11337 = n45570 ;
  assign y11338 = n45573 ;
  assign y11339 = ~n45576 ;
  assign y11340 = n45578 ;
  assign y11341 = ~n45581 ;
  assign y11342 = ~n45586 ;
  assign y11343 = ~n45591 ;
  assign y11344 = n45593 ;
  assign y11345 = ~1'b0 ;
  assign y11346 = n45596 ;
  assign y11347 = n45603 ;
  assign y11348 = ~n45605 ;
  assign y11349 = ~n45606 ;
  assign y11350 = n45610 ;
  assign y11351 = n45612 ;
  assign y11352 = ~n45614 ;
  assign y11353 = n45621 ;
  assign y11354 = n45623 ;
  assign y11355 = ~n45625 ;
  assign y11356 = ~n45632 ;
  assign y11357 = n45633 ;
  assign y11358 = ~n45637 ;
  assign y11359 = n45638 ;
  assign y11360 = ~n45644 ;
  assign y11361 = n45646 ;
  assign y11362 = ~n45647 ;
  assign y11363 = ~1'b0 ;
  assign y11364 = ~n45652 ;
  assign y11365 = ~n45654 ;
  assign y11366 = ~n31960 ;
  assign y11367 = n45655 ;
  assign y11368 = ~n45659 ;
  assign y11369 = n45660 ;
  assign y11370 = n45661 ;
  assign y11371 = ~1'b0 ;
  assign y11372 = ~n45667 ;
  assign y11373 = ~n45670 ;
  assign y11374 = ~n45676 ;
  assign y11375 = n45680 ;
  assign y11376 = n45681 ;
  assign y11377 = n45682 ;
  assign y11378 = ~n45683 ;
  assign y11379 = n45684 ;
  assign y11380 = n45686 ;
  assign y11381 = ~n45689 ;
  assign y11382 = ~n45691 ;
  assign y11383 = n45693 ;
  assign y11384 = ~n45701 ;
  assign y11385 = ~n45708 ;
  assign y11386 = n45714 ;
  assign y11387 = ~n45718 ;
  assign y11388 = ~1'b0 ;
  assign y11389 = ~1'b0 ;
  assign y11390 = ~n45720 ;
  assign y11391 = ~n45722 ;
  assign y11392 = n45726 ;
  assign y11393 = ~n45728 ;
  assign y11394 = ~n45736 ;
  assign y11395 = n45737 ;
  assign y11396 = n45739 ;
  assign y11397 = ~n45742 ;
  assign y11398 = n45747 ;
  assign y11399 = ~n45748 ;
  assign y11400 = n45754 ;
  assign y11401 = ~n45755 ;
  assign y11402 = ~n45756 ;
  assign y11403 = ~n45758 ;
  assign y11404 = ~n45760 ;
  assign y11405 = n45763 ;
  assign y11406 = ~n45765 ;
  assign y11407 = ~n45770 ;
  assign y11408 = n45775 ;
  assign y11409 = n45780 ;
  assign y11410 = n45783 ;
  assign y11411 = ~n45784 ;
  assign y11412 = ~n45786 ;
  assign y11413 = n45787 ;
  assign y11414 = ~n45788 ;
  assign y11415 = n45792 ;
  assign y11416 = ~n45793 ;
  assign y11417 = ~n45794 ;
  assign y11418 = n45797 ;
  assign y11419 = ~n45798 ;
  assign y11420 = n45802 ;
  assign y11421 = n45806 ;
  assign y11422 = n45809 ;
  assign y11423 = n45810 ;
  assign y11424 = ~1'b0 ;
  assign y11425 = ~n45815 ;
  assign y11426 = ~n45816 ;
  assign y11427 = n45817 ;
  assign y11428 = n45818 ;
  assign y11429 = ~n45821 ;
  assign y11430 = ~n45826 ;
  assign y11431 = n45827 ;
  assign y11432 = ~n45829 ;
  assign y11433 = ~n45832 ;
  assign y11434 = ~n45834 ;
  assign y11435 = ~n45835 ;
  assign y11436 = ~n45836 ;
  assign y11437 = n45837 ;
  assign y11438 = n45841 ;
  assign y11439 = n45842 ;
  assign y11440 = n45844 ;
  assign y11441 = ~n45849 ;
  assign y11442 = ~n45850 ;
  assign y11443 = ~n45860 ;
  assign y11444 = ~n45863 ;
  assign y11445 = n45867 ;
  assign y11446 = ~n45873 ;
  assign y11447 = n45874 ;
  assign y11448 = ~n45879 ;
  assign y11449 = ~1'b0 ;
  assign y11450 = ~n45883 ;
  assign y11451 = n45884 ;
  assign y11452 = n45892 ;
  assign y11453 = ~n45895 ;
  assign y11454 = n45900 ;
  assign y11455 = ~n45902 ;
  assign y11456 = n45903 ;
  assign y11457 = n45904 ;
  assign y11458 = n45908 ;
  assign y11459 = n45909 ;
  assign y11460 = ~n45910 ;
  assign y11461 = n45913 ;
  assign y11462 = ~n45916 ;
  assign y11463 = n45918 ;
  assign y11464 = n45922 ;
  assign y11465 = ~n45923 ;
  assign y11466 = n45929 ;
  assign y11467 = ~n45935 ;
  assign y11468 = ~n45942 ;
  assign y11469 = ~n45943 ;
  assign y11470 = ~1'b0 ;
  assign y11471 = ~n45944 ;
  assign y11472 = ~n45945 ;
  assign y11473 = ~n45946 ;
  assign y11474 = ~n45949 ;
  assign y11475 = ~n45951 ;
  assign y11476 = ~n45952 ;
  assign y11477 = ~n45954 ;
  assign y11478 = n45957 ;
  assign y11479 = ~n45962 ;
  assign y11480 = n45965 ;
  assign y11481 = n45966 ;
  assign y11482 = n45970 ;
  assign y11483 = n45971 ;
  assign y11484 = n45973 ;
  assign y11485 = n45979 ;
  assign y11486 = n45981 ;
  assign y11487 = ~n45982 ;
  assign y11488 = n45984 ;
  assign y11489 = ~n45987 ;
  assign y11490 = n45993 ;
  assign y11491 = ~n45994 ;
  assign y11492 = ~n45998 ;
  assign y11493 = n46002 ;
  assign y11494 = n46004 ;
  assign y11495 = ~n46005 ;
  assign y11496 = n46012 ;
  assign y11497 = ~1'b0 ;
  assign y11498 = ~n46013 ;
  assign y11499 = n46014 ;
  assign y11500 = n46015 ;
  assign y11501 = n46018 ;
  assign y11502 = n46019 ;
  assign y11503 = ~n46024 ;
  assign y11504 = n46025 ;
  assign y11505 = ~n46026 ;
  assign y11506 = n46027 ;
  assign y11507 = ~n46032 ;
  assign y11508 = ~n46036 ;
  assign y11509 = ~n46037 ;
  assign y11510 = ~n46042 ;
  assign y11511 = ~n46044 ;
  assign y11512 = n46049 ;
  assign y11513 = n46050 ;
  assign y11514 = n46051 ;
  assign y11515 = ~n46056 ;
  assign y11516 = n46057 ;
  assign y11517 = n46058 ;
  assign y11518 = n46061 ;
  assign y11519 = ~n46062 ;
  assign y11520 = ~n46063 ;
  assign y11521 = n46066 ;
  assign y11522 = ~1'b0 ;
  assign y11523 = n46069 ;
  assign y11524 = ~n46075 ;
  assign y11525 = ~n46077 ;
  assign y11526 = n46079 ;
  assign y11527 = n46085 ;
  assign y11528 = n46088 ;
  assign y11529 = ~n46097 ;
  assign y11530 = n46098 ;
  assign y11531 = ~n46099 ;
  assign y11532 = n46101 ;
  assign y11533 = n46105 ;
  assign y11534 = n46106 ;
  assign y11535 = n46108 ;
  assign y11536 = ~n46109 ;
  assign y11537 = ~n46111 ;
  assign y11538 = n46114 ;
  assign y11539 = ~n46117 ;
  assign y11540 = n46120 ;
  assign y11541 = n46121 ;
  assign y11542 = ~n46124 ;
  assign y11543 = n46134 ;
  assign y11544 = ~n46139 ;
  assign y11545 = ~n46146 ;
  assign y11546 = ~1'b0 ;
  assign y11547 = ~1'b0 ;
  assign y11548 = n46147 ;
  assign y11549 = n46148 ;
  assign y11550 = n46150 ;
  assign y11551 = n46151 ;
  assign y11552 = n46154 ;
  assign y11553 = n46155 ;
  assign y11554 = n46160 ;
  assign y11555 = n46163 ;
  assign y11556 = ~n46164 ;
  assign y11557 = ~n46165 ;
  assign y11558 = ~n46166 ;
  assign y11559 = n46168 ;
  assign y11560 = ~n46175 ;
  assign y11561 = n46178 ;
  assign y11562 = ~n46180 ;
  assign y11563 = n46182 ;
  assign y11564 = n46188 ;
  assign y11565 = n46190 ;
  assign y11566 = ~n46192 ;
  assign y11567 = n46193 ;
  assign y11568 = n46195 ;
  assign y11569 = n46198 ;
  assign y11570 = n46200 ;
  assign y11571 = n46201 ;
  assign y11572 = n46203 ;
  assign y11573 = ~n46204 ;
  assign y11574 = ~n46207 ;
  assign y11575 = n46209 ;
  assign y11576 = ~n46217 ;
  assign y11577 = ~n46224 ;
  assign y11578 = ~n46225 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = n46226 ;
  assign y11581 = ~n46232 ;
  assign y11582 = ~n46236 ;
  assign y11583 = ~n46244 ;
  assign y11584 = n46245 ;
  assign y11585 = ~n46247 ;
  assign y11586 = ~n46249 ;
  assign y11587 = n46253 ;
  assign y11588 = ~n46258 ;
  assign y11589 = n46260 ;
  assign y11590 = n46268 ;
  assign y11591 = ~n46270 ;
  assign y11592 = n46273 ;
  assign y11593 = ~n11249 ;
  assign y11594 = ~n46275 ;
  assign y11595 = n46280 ;
  assign y11596 = ~n46281 ;
  assign y11597 = n46284 ;
  assign y11598 = ~n46285 ;
  assign y11599 = ~n46286 ;
  assign y11600 = ~n46287 ;
  assign y11601 = ~n46288 ;
  assign y11602 = n46291 ;
  assign y11603 = ~n46294 ;
  assign y11604 = ~n46298 ;
  assign y11605 = n46301 ;
  assign y11606 = n46302 ;
  assign y11607 = n46305 ;
  assign y11608 = n46306 ;
  assign y11609 = n46307 ;
  assign y11610 = ~n46311 ;
  assign y11611 = n46312 ;
  assign y11612 = ~n46313 ;
  assign y11613 = n46314 ;
  assign y11614 = n46317 ;
  assign y11615 = n46322 ;
  assign y11616 = ~n46324 ;
  assign y11617 = ~n46326 ;
  assign y11618 = ~n46329 ;
  assign y11619 = n46332 ;
  assign y11620 = n46337 ;
  assign y11621 = n46339 ;
  assign y11622 = n46340 ;
  assign y11623 = ~1'b0 ;
  assign y11624 = ~1'b0 ;
  assign y11625 = ~n46341 ;
  assign y11626 = ~n46343 ;
  assign y11627 = ~n46347 ;
  assign y11628 = ~n46353 ;
  assign y11629 = n46358 ;
  assign y11630 = ~n46362 ;
  assign y11631 = ~n46365 ;
  assign y11632 = n46367 ;
  assign y11633 = n46368 ;
  assign y11634 = ~n46369 ;
  assign y11635 = n46370 ;
  assign y11636 = ~n46372 ;
  assign y11637 = n46379 ;
  assign y11638 = n46383 ;
  assign y11639 = ~1'b0 ;
  assign y11640 = ~n46385 ;
  assign y11641 = ~n46386 ;
  assign y11642 = ~n46387 ;
  assign y11643 = n46388 ;
  assign y11644 = n46393 ;
  assign y11645 = n46394 ;
  assign y11646 = n46396 ;
  assign y11647 = ~1'b0 ;
  assign y11648 = n46399 ;
  assign y11649 = n46401 ;
  assign y11650 = ~n46403 ;
  assign y11651 = n46405 ;
  assign y11652 = n46406 ;
  assign y11653 = ~n46407 ;
  assign y11654 = n46408 ;
  assign y11655 = n46409 ;
  assign y11656 = ~n46410 ;
  assign y11657 = n46412 ;
  assign y11658 = n46415 ;
  assign y11659 = n46421 ;
  assign y11660 = ~n46422 ;
  assign y11661 = n46423 ;
  assign y11662 = ~n46429 ;
  assign y11663 = n46435 ;
  assign y11664 = n46437 ;
  assign y11665 = n46438 ;
  assign y11666 = n46441 ;
  assign y11667 = n46443 ;
  assign y11668 = ~n46445 ;
  assign y11669 = ~n46450 ;
  assign y11670 = n46452 ;
  assign y11671 = ~n46454 ;
  assign y11672 = ~n46458 ;
  assign y11673 = n46463 ;
  assign y11674 = n46467 ;
  assign y11675 = ~n46470 ;
  assign y11676 = ~n46477 ;
  assign y11677 = ~1'b0 ;
  assign y11678 = ~n46478 ;
  assign y11679 = ~n46480 ;
  assign y11680 = n46481 ;
  assign y11681 = n46482 ;
  assign y11682 = ~n46485 ;
  assign y11683 = n46494 ;
  assign y11684 = ~n46497 ;
  assign y11685 = ~n46498 ;
  assign y11686 = ~n46499 ;
  assign y11687 = ~n46508 ;
  assign y11688 = ~n46510 ;
  assign y11689 = n46515 ;
  assign y11690 = n46517 ;
  assign y11691 = ~n46519 ;
  assign y11692 = n46520 ;
  assign y11693 = ~n46521 ;
  assign y11694 = n46522 ;
  assign y11695 = ~n46525 ;
  assign y11696 = n46527 ;
  assign y11697 = ~n46529 ;
  assign y11698 = n46530 ;
  assign y11699 = n46531 ;
  assign y11700 = n46535 ;
  assign y11701 = n46536 ;
  assign y11702 = ~n46537 ;
  assign y11703 = n46540 ;
  assign y11704 = n46547 ;
  assign y11705 = n46549 ;
  assign y11706 = ~n46553 ;
  assign y11707 = n46555 ;
  assign y11708 = n46559 ;
  assign y11709 = ~n46560 ;
  assign y11710 = n46563 ;
  assign y11711 = ~n46564 ;
  assign y11712 = ~n46565 ;
  assign y11713 = ~n46570 ;
  assign y11714 = ~n46573 ;
  assign y11715 = ~n46574 ;
  assign y11716 = n46575 ;
  assign y11717 = ~n46576 ;
  assign y11718 = ~n46578 ;
  assign y11719 = n46579 ;
  assign y11720 = ~n46581 ;
  assign y11721 = n46587 ;
  assign y11722 = ~n46588 ;
  assign y11723 = n46595 ;
  assign y11724 = ~n46596 ;
  assign y11725 = n46597 ;
  assign y11726 = n46600 ;
  assign y11727 = n46603 ;
  assign y11728 = ~n46606 ;
  assign y11729 = ~n46607 ;
  assign y11730 = ~n46611 ;
  assign y11731 = ~n46614 ;
  assign y11732 = n46616 ;
  assign y11733 = n46618 ;
  assign y11734 = n46621 ;
  assign y11735 = ~n46623 ;
  assign y11736 = ~n46626 ;
  assign y11737 = n46627 ;
  assign y11738 = n46631 ;
  assign y11739 = n46637 ;
  assign y11740 = ~n46640 ;
  assign y11741 = ~n46645 ;
  assign y11742 = n46648 ;
  assign y11743 = ~n46651 ;
  assign y11744 = ~n46652 ;
  assign y11745 = ~n46654 ;
  assign y11746 = n46656 ;
  assign y11747 = n46658 ;
  assign y11748 = ~n46663 ;
  assign y11749 = ~n46665 ;
  assign y11750 = ~1'b0 ;
  assign y11751 = n46669 ;
  assign y11752 = n46670 ;
  assign y11753 = ~n46674 ;
  assign y11754 = ~n46675 ;
  assign y11755 = n46678 ;
  assign y11756 = ~n46679 ;
  assign y11757 = n46682 ;
  assign y11758 = ~1'b0 ;
  assign y11759 = n46686 ;
  assign y11760 = n46690 ;
  assign y11761 = n46691 ;
  assign y11762 = ~n46696 ;
  assign y11763 = ~n46702 ;
  assign y11764 = n46704 ;
  assign y11765 = n46708 ;
  assign y11766 = ~n46709 ;
  assign y11767 = n46714 ;
  assign y11768 = n46715 ;
  assign y11769 = ~n46717 ;
  assign y11770 = ~n46718 ;
  assign y11771 = ~n46720 ;
  assign y11772 = n46722 ;
  assign y11773 = ~n46727 ;
  assign y11774 = ~n46729 ;
  assign y11775 = n46731 ;
  assign y11776 = ~n46732 ;
  assign y11777 = n46734 ;
  assign y11778 = n46737 ;
  assign y11779 = ~n46738 ;
  assign y11780 = n46740 ;
  assign y11781 = ~1'b0 ;
  assign y11782 = n46742 ;
  assign y11783 = ~n46746 ;
  assign y11784 = n46747 ;
  assign y11785 = ~n46748 ;
  assign y11786 = n46751 ;
  assign y11787 = n46757 ;
  assign y11788 = n46760 ;
  assign y11789 = ~n46764 ;
  assign y11790 = ~n46766 ;
  assign y11791 = ~n46772 ;
  assign y11792 = ~n46776 ;
  assign y11793 = ~n46778 ;
  assign y11794 = n46779 ;
  assign y11795 = ~n46782 ;
  assign y11796 = n46784 ;
  assign y11797 = n46786 ;
  assign y11798 = n46789 ;
  assign y11799 = ~n46791 ;
  assign y11800 = ~n46792 ;
  assign y11801 = ~n46795 ;
  assign y11802 = n46797 ;
  assign y11803 = n46800 ;
  assign y11804 = ~n46801 ;
  assign y11805 = ~n46804 ;
  assign y11806 = ~n46805 ;
  assign y11807 = ~n46806 ;
  assign y11808 = n46809 ;
  assign y11809 = ~n46811 ;
  assign y11810 = n46813 ;
  assign y11811 = ~n46814 ;
  assign y11812 = n46815 ;
  assign y11813 = ~n46822 ;
  assign y11814 = ~n46823 ;
  assign y11815 = n46825 ;
  assign y11816 = n46831 ;
  assign y11817 = n46835 ;
  assign y11818 = n46841 ;
  assign y11819 = ~1'b0 ;
  assign y11820 = ~n46846 ;
  assign y11821 = n46852 ;
  assign y11822 = ~n46854 ;
  assign y11823 = ~n46855 ;
  assign y11824 = n46858 ;
  assign y11825 = ~n46861 ;
  assign y11826 = n46862 ;
  assign y11827 = ~n46865 ;
  assign y11828 = ~n46868 ;
  assign y11829 = ~n46873 ;
  assign y11830 = n46878 ;
  assign y11831 = n46879 ;
  assign y11832 = ~n46880 ;
  assign y11833 = ~n46882 ;
  assign y11834 = ~n46885 ;
  assign y11835 = ~n46887 ;
  assign y11836 = n46889 ;
  assign y11837 = n46890 ;
  assign y11838 = ~n46894 ;
  assign y11839 = n46898 ;
  assign y11840 = ~n46901 ;
  assign y11841 = n46908 ;
  assign y11842 = ~1'b0 ;
  assign y11843 = n46912 ;
  assign y11844 = n46913 ;
  assign y11845 = ~n46915 ;
  assign y11846 = ~n46917 ;
  assign y11847 = ~n46918 ;
  assign y11848 = ~1'b0 ;
  assign y11849 = ~n46922 ;
  assign y11850 = ~n46927 ;
  assign y11851 = ~n46929 ;
  assign y11852 = n46930 ;
  assign y11853 = ~n46931 ;
  assign y11854 = n46939 ;
  assign y11855 = ~n46941 ;
  assign y11856 = ~n46944 ;
  assign y11857 = ~n46946 ;
  assign y11858 = n46950 ;
  assign y11859 = ~n46955 ;
  assign y11860 = n46958 ;
  assign y11861 = n46959 ;
  assign y11862 = ~n46963 ;
  assign y11863 = n46964 ;
  assign y11864 = ~n46965 ;
  assign y11865 = ~n46966 ;
  assign y11866 = ~n46969 ;
  assign y11867 = ~n46970 ;
  assign y11868 = n46972 ;
  assign y11869 = n46980 ;
  assign y11870 = n46981 ;
  assign y11871 = ~n46985 ;
  assign y11872 = ~n46986 ;
  assign y11873 = ~n46987 ;
  assign y11874 = n46989 ;
  assign y11875 = ~n46990 ;
  assign y11876 = n43037 ;
  assign y11877 = ~n46994 ;
  assign y11878 = ~n47000 ;
  assign y11879 = n47003 ;
  assign y11880 = ~n47006 ;
  assign y11881 = ~n47008 ;
  assign y11882 = ~n47010 ;
  assign y11883 = n47011 ;
  assign y11884 = n47013 ;
  assign y11885 = ~n47015 ;
  assign y11886 = n47019 ;
  assign y11887 = n47024 ;
  assign y11888 = ~n47026 ;
  assign y11889 = ~n47027 ;
  assign y11890 = ~n47028 ;
  assign y11891 = ~n47029 ;
  assign y11892 = ~1'b0 ;
  assign y11893 = ~n47031 ;
  assign y11894 = n47035 ;
  assign y11895 = ~n47037 ;
  assign y11896 = n47040 ;
  assign y11897 = n47041 ;
  assign y11898 = n47043 ;
  assign y11899 = n47044 ;
  assign y11900 = n47045 ;
  assign y11901 = n47047 ;
  assign y11902 = n47050 ;
  assign y11903 = n47052 ;
  assign y11904 = n47053 ;
  assign y11905 = n47054 ;
  assign y11906 = ~n47056 ;
  assign y11907 = n47059 ;
  assign y11908 = n47063 ;
  assign y11909 = ~n47065 ;
  assign y11910 = ~n22215 ;
  assign y11911 = ~n47066 ;
  assign y11912 = ~1'b0 ;
  assign y11913 = n47069 ;
  assign y11914 = ~n47074 ;
  assign y11915 = ~n47078 ;
  assign y11916 = n47080 ;
  assign y11917 = ~n47081 ;
  assign y11918 = n47082 ;
  assign y11919 = ~n47086 ;
  assign y11920 = ~n47092 ;
  assign y11921 = ~n47095 ;
  assign y11922 = ~n47098 ;
  assign y11923 = n47100 ;
  assign y11924 = n47102 ;
  assign y11925 = ~n47103 ;
  assign y11926 = n47105 ;
  assign y11927 = n47107 ;
  assign y11928 = n47109 ;
  assign y11929 = ~n47113 ;
  assign y11930 = ~n47114 ;
  assign y11931 = ~n47117 ;
  assign y11932 = ~n47118 ;
  assign y11933 = n47120 ;
  assign y11934 = ~n47121 ;
  assign y11935 = n47122 ;
  assign y11936 = n47123 ;
  assign y11937 = n47133 ;
  assign y11938 = n47140 ;
  assign y11939 = n47141 ;
  assign y11940 = n47143 ;
  assign y11941 = n47145 ;
  assign y11942 = ~n47151 ;
  assign y11943 = ~n47152 ;
  assign y11944 = n47154 ;
  assign y11945 = ~n47155 ;
  assign y11946 = ~n47159 ;
  assign y11947 = n47164 ;
  assign y11948 = n47166 ;
  assign y11949 = ~n47169 ;
  assign y11950 = n47172 ;
  assign y11951 = n47173 ;
  assign y11952 = ~n47176 ;
  assign y11953 = n47177 ;
  assign y11954 = ~n47179 ;
  assign y11955 = ~1'b0 ;
  assign y11956 = ~n47180 ;
  assign y11957 = ~n47181 ;
  assign y11958 = ~n47182 ;
  assign y11959 = ~n47186 ;
  assign y11960 = ~n47187 ;
  assign y11961 = ~n47190 ;
  assign y11962 = n47193 ;
  assign y11963 = ~n47195 ;
  assign y11964 = ~1'b0 ;
  assign y11965 = n47197 ;
  assign y11966 = ~n47200 ;
  assign y11967 = n47202 ;
  assign y11968 = n47204 ;
  assign y11969 = n47205 ;
  assign y11970 = n47206 ;
  assign y11971 = n47211 ;
  assign y11972 = ~1'b0 ;
  assign y11973 = n47215 ;
  assign y11974 = ~n47219 ;
  assign y11975 = n47223 ;
  assign y11976 = n47225 ;
  assign y11977 = n47226 ;
  assign y11978 = ~n47229 ;
  assign y11979 = n47231 ;
  assign y11980 = n47232 ;
  assign y11981 = ~n47235 ;
  assign y11982 = ~1'b0 ;
  assign y11983 = ~n47237 ;
  assign y11984 = ~n47239 ;
  assign y11985 = ~n47242 ;
  assign y11986 = n47246 ;
  assign y11987 = n47247 ;
  assign y11988 = ~n47248 ;
  assign y11989 = ~n47251 ;
  assign y11990 = ~n47252 ;
  assign y11991 = ~n47254 ;
  assign y11992 = ~1'b0 ;
  assign y11993 = ~n47258 ;
  assign y11994 = ~n47262 ;
  assign y11995 = n47265 ;
  assign y11996 = ~n47268 ;
  assign y11997 = ~n47269 ;
  assign y11998 = n47270 ;
  assign y11999 = n47273 ;
  assign y12000 = n47277 ;
  assign y12001 = n47281 ;
  assign y12002 = ~n47284 ;
  assign y12003 = ~n47288 ;
  assign y12004 = ~n47289 ;
  assign y12005 = n47291 ;
  assign y12006 = n47294 ;
  assign y12007 = ~n47296 ;
  assign y12008 = n47298 ;
  assign y12009 = ~n47300 ;
  assign y12010 = n47301 ;
  assign y12011 = n47302 ;
  assign y12012 = ~n47304 ;
  assign y12013 = n47305 ;
  assign y12014 = n47314 ;
  assign y12015 = n47315 ;
  assign y12016 = ~n47316 ;
  assign y12017 = n47319 ;
  assign y12018 = n47322 ;
  assign y12019 = n47324 ;
  assign y12020 = n47325 ;
  assign y12021 = ~n47326 ;
  assign y12022 = n47327 ;
  assign y12023 = ~n47329 ;
  assign y12024 = n47331 ;
  assign y12025 = n47332 ;
  assign y12026 = ~n47334 ;
  assign y12027 = ~n47339 ;
  assign y12028 = n47340 ;
  assign y12029 = n47346 ;
  assign y12030 = ~n47351 ;
  assign y12031 = n47353 ;
  assign y12032 = ~n47354 ;
  assign y12033 = ~n47356 ;
  assign y12034 = ~n47359 ;
  assign y12035 = n47360 ;
  assign y12036 = n47362 ;
  assign y12037 = ~n47365 ;
  assign y12038 = n47366 ;
  assign y12039 = n47371 ;
  assign y12040 = n47374 ;
  assign y12041 = ~n47376 ;
  assign y12042 = n47380 ;
  assign y12043 = n47383 ;
  assign y12044 = ~n47389 ;
  assign y12045 = n47391 ;
  assign y12046 = ~n47394 ;
  assign y12047 = n47397 ;
  assign y12048 = n47401 ;
  assign y12049 = n47403 ;
  assign y12050 = ~n47407 ;
  assign y12051 = n47408 ;
  assign y12052 = n47409 ;
  assign y12053 = ~n47412 ;
  assign y12054 = n47415 ;
  assign y12055 = ~n47416 ;
  assign y12056 = n47418 ;
  assign y12057 = ~n47423 ;
  assign y12058 = n47427 ;
  assign y12059 = ~n47429 ;
  assign y12060 = n47430 ;
  assign y12061 = ~n47431 ;
  assign y12062 = ~n47435 ;
  assign y12063 = n47441 ;
  assign y12064 = n47446 ;
  assign y12065 = ~n47450 ;
  assign y12066 = ~1'b0 ;
  assign y12067 = ~n47453 ;
  assign y12068 = ~n47458 ;
  assign y12069 = ~n47460 ;
  assign y12070 = n47461 ;
  assign y12071 = n47462 ;
  assign y12072 = n47467 ;
  assign y12073 = n47468 ;
  assign y12074 = ~n47469 ;
  assign y12075 = ~n47471 ;
  assign y12076 = n47472 ;
  assign y12077 = ~n47473 ;
  assign y12078 = n47475 ;
  assign y12079 = n47477 ;
  assign y12080 = n47478 ;
  assign y12081 = n47479 ;
  assign y12082 = ~n47480 ;
  assign y12083 = ~n47482 ;
  assign y12084 = ~n47484 ;
  assign y12085 = n47485 ;
  assign y12086 = ~n47486 ;
  assign y12087 = ~n47492 ;
  assign y12088 = ~n47495 ;
  assign y12089 = n47496 ;
  assign y12090 = n47500 ;
  assign y12091 = ~n47501 ;
  assign y12092 = n47502 ;
  assign y12093 = ~n47505 ;
  assign y12094 = n47508 ;
  assign y12095 = n47510 ;
  assign y12096 = ~n47511 ;
  assign y12097 = n47512 ;
  assign y12098 = ~n47513 ;
  assign y12099 = ~n47514 ;
  assign y12100 = ~n47515 ;
  assign y12101 = ~n47518 ;
  assign y12102 = ~n47520 ;
  assign y12103 = n47522 ;
  assign y12104 = ~n47525 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = n47528 ;
  assign y12107 = n47531 ;
  assign y12108 = ~n47532 ;
  assign y12109 = ~n47540 ;
  assign y12110 = ~n47544 ;
  assign y12111 = ~n47545 ;
  assign y12112 = ~1'b0 ;
  assign y12113 = n47548 ;
  assign y12114 = n47550 ;
  assign y12115 = ~n47554 ;
  assign y12116 = n47558 ;
  assign y12117 = n47560 ;
  assign y12118 = n47562 ;
  assign y12119 = ~n47566 ;
  assign y12120 = n47572 ;
  assign y12121 = ~n47574 ;
  assign y12122 = ~n47576 ;
  assign y12123 = ~n47577 ;
  assign y12124 = n47578 ;
  assign y12125 = n47579 ;
  assign y12126 = n47581 ;
  assign y12127 = ~n47582 ;
  assign y12128 = n47584 ;
  assign y12129 = ~n47585 ;
  assign y12130 = ~1'b0 ;
  assign y12131 = ~n47586 ;
  assign y12132 = n47587 ;
  assign y12133 = n47589 ;
  assign y12134 = ~n47591 ;
  assign y12135 = n47593 ;
  assign y12136 = n47596 ;
  assign y12137 = n47603 ;
  assign y12138 = ~n47606 ;
  assign y12139 = ~n47607 ;
  assign y12140 = n47612 ;
  assign y12141 = n47614 ;
  assign y12142 = ~n47615 ;
  assign y12143 = n47619 ;
  assign y12144 = ~n47629 ;
  assign y12145 = ~n47630 ;
  assign y12146 = ~n47631 ;
  assign y12147 = ~n47632 ;
  assign y12148 = ~n47640 ;
  assign y12149 = n47645 ;
  assign y12150 = n47646 ;
  assign y12151 = ~n47648 ;
  assign y12152 = n47650 ;
  assign y12153 = ~n47651 ;
  assign y12154 = n47652 ;
  assign y12155 = ~n47654 ;
  assign y12156 = n47656 ;
  assign y12157 = n47664 ;
  assign y12158 = n47669 ;
  assign y12159 = ~n47671 ;
  assign y12160 = n47673 ;
  assign y12161 = n47676 ;
  assign y12162 = n47677 ;
  assign y12163 = ~n47678 ;
  assign y12164 = n47679 ;
  assign y12165 = ~n47682 ;
  assign y12166 = n47683 ;
  assign y12167 = n47688 ;
  assign y12168 = n47694 ;
  assign y12169 = ~n47702 ;
  assign y12170 = ~n47703 ;
  assign y12171 = n47704 ;
  assign y12172 = ~n47705 ;
  assign y12173 = n47706 ;
  assign y12174 = ~n47708 ;
  assign y12175 = n47709 ;
  assign y12176 = ~n47715 ;
  assign y12177 = n47716 ;
  assign y12178 = n47717 ;
  assign y12179 = ~n47718 ;
  assign y12180 = n47725 ;
  assign y12181 = ~n47727 ;
  assign y12182 = ~1'b0 ;
  assign y12183 = ~n47729 ;
  assign y12184 = n47732 ;
  assign y12185 = n47737 ;
  assign y12186 = ~n47745 ;
  assign y12187 = ~n47746 ;
  assign y12188 = n47748 ;
  assign y12189 = n47749 ;
  assign y12190 = n47753 ;
  assign y12191 = ~n47755 ;
  assign y12192 = n47762 ;
  assign y12193 = n47763 ;
  assign y12194 = ~n47764 ;
  assign y12195 = ~n47766 ;
  assign y12196 = n47769 ;
  assign y12197 = ~n47770 ;
  assign y12198 = n47773 ;
  assign y12199 = ~n47774 ;
  assign y12200 = n47776 ;
  assign y12201 = ~n47780 ;
  assign y12202 = ~n47781 ;
  assign y12203 = ~n47783 ;
  assign y12204 = ~n47786 ;
  assign y12205 = n47789 ;
  assign y12206 = n47792 ;
  assign y12207 = n47794 ;
  assign y12208 = ~1'b0 ;
  assign y12209 = ~n47795 ;
  assign y12210 = ~n47798 ;
  assign y12211 = n47799 ;
  assign y12212 = n47802 ;
  assign y12213 = n47803 ;
  assign y12214 = ~n47806 ;
  assign y12215 = ~n47808 ;
  assign y12216 = n47809 ;
  assign y12217 = ~n47810 ;
  assign y12218 = ~1'b0 ;
  assign y12219 = ~n47813 ;
  assign y12220 = ~n47815 ;
  assign y12221 = ~n47817 ;
  assign y12222 = ~n47818 ;
  assign y12223 = n47821 ;
  assign y12224 = ~n47827 ;
  assign y12225 = n47828 ;
  assign y12226 = ~1'b0 ;
  assign y12227 = n47830 ;
  assign y12228 = n47834 ;
  assign y12229 = ~n47835 ;
  assign y12230 = n47836 ;
  assign y12231 = ~n47837 ;
  assign y12232 = ~n47838 ;
  assign y12233 = ~n47839 ;
  assign y12234 = n47843 ;
  assign y12235 = ~n47844 ;
  assign y12236 = ~n47848 ;
  assign y12237 = ~n47850 ;
  assign y12238 = n47854 ;
  assign y12239 = ~n47856 ;
  assign y12240 = ~1'b0 ;
  assign y12241 = ~n47858 ;
  assign y12242 = n47859 ;
  assign y12243 = n47862 ;
  assign y12244 = n47863 ;
  assign y12245 = ~n47868 ;
  assign y12246 = n47871 ;
  assign y12247 = ~n47872 ;
  assign y12248 = ~n47875 ;
  assign y12249 = ~n47878 ;
  assign y12250 = ~1'b0 ;
  assign y12251 = n47881 ;
  assign y12252 = n47886 ;
  assign y12253 = n47892 ;
  assign y12254 = ~n47893 ;
  assign y12255 = ~n47898 ;
  assign y12256 = n47901 ;
  assign y12257 = ~n47903 ;
  assign y12258 = n47906 ;
  assign y12259 = ~n47907 ;
  assign y12260 = n47909 ;
  assign y12261 = n47911 ;
  assign y12262 = n47912 ;
  assign y12263 = n47914 ;
  assign y12264 = ~n47927 ;
  assign y12265 = n47930 ;
  assign y12266 = n47934 ;
  assign y12267 = n47936 ;
  assign y12268 = n47938 ;
  assign y12269 = ~n47943 ;
  assign y12270 = ~n47950 ;
  assign y12271 = ~n47951 ;
  assign y12272 = ~n47953 ;
  assign y12273 = n47954 ;
  assign y12274 = ~n47956 ;
  assign y12275 = ~n47957 ;
  assign y12276 = ~n47959 ;
  assign y12277 = n47962 ;
  assign y12278 = ~n47968 ;
  assign y12279 = ~n47972 ;
  assign y12280 = n47976 ;
  assign y12281 = ~n47977 ;
  assign y12282 = n47979 ;
  assign y12283 = n47981 ;
  assign y12284 = ~n47986 ;
  assign y12285 = n47990 ;
  assign y12286 = ~n47994 ;
  assign y12287 = n47996 ;
  assign y12288 = ~n47998 ;
  assign y12289 = ~n48003 ;
  assign y12290 = n48004 ;
  assign y12291 = n48007 ;
  assign y12292 = n48011 ;
  assign y12293 = n48017 ;
  assign y12294 = n48024 ;
  assign y12295 = ~n48027 ;
  assign y12296 = ~n48028 ;
  assign y12297 = ~n48033 ;
  assign y12298 = ~n48036 ;
  assign y12299 = ~n48039 ;
  assign y12300 = n48046 ;
  assign y12301 = n48048 ;
  assign y12302 = ~n48051 ;
  assign y12303 = n48054 ;
  assign y12304 = n48058 ;
  assign y12305 = ~n48061 ;
  assign y12306 = ~n48062 ;
  assign y12307 = n48064 ;
  assign y12308 = n48066 ;
  assign y12309 = ~n48068 ;
  assign y12310 = n48071 ;
  assign y12311 = n48072 ;
  assign y12312 = ~1'b0 ;
  assign y12313 = ~1'b0 ;
  assign y12314 = ~n48075 ;
  assign y12315 = ~n48076 ;
  assign y12316 = ~n48077 ;
  assign y12317 = n48080 ;
  assign y12318 = ~n48083 ;
  assign y12319 = n48086 ;
  assign y12320 = n48087 ;
  assign y12321 = ~n48091 ;
  assign y12322 = ~n48097 ;
  assign y12323 = n48104 ;
  assign y12324 = n48107 ;
  assign y12325 = ~n48111 ;
  assign y12326 = n48115 ;
  assign y12327 = ~n48116 ;
  assign y12328 = n48117 ;
  assign y12329 = ~n48118 ;
  assign y12330 = ~1'b0 ;
  assign y12331 = ~n48120 ;
  assign y12332 = ~n48126 ;
  assign y12333 = ~n48129 ;
  assign y12334 = ~n48130 ;
  assign y12335 = n48131 ;
  assign y12336 = n48135 ;
  assign y12337 = ~n48138 ;
  assign y12338 = ~n48141 ;
  assign y12339 = ~n48146 ;
  assign y12340 = ~1'b0 ;
  assign y12341 = ~n48147 ;
  assign y12342 = n48153 ;
  assign y12343 = ~n48156 ;
  assign y12344 = n48160 ;
  assign y12345 = n48161 ;
  assign y12346 = n48164 ;
  assign y12347 = ~n48168 ;
  assign y12348 = n48172 ;
  assign y12349 = n48174 ;
  assign y12350 = ~1'b0 ;
  assign y12351 = n48178 ;
  assign y12352 = ~n48179 ;
  assign y12353 = n48180 ;
  assign y12354 = n48182 ;
  assign y12355 = n48183 ;
  assign y12356 = n48184 ;
  assign y12357 = n48185 ;
  assign y12358 = n48188 ;
  assign y12359 = n48190 ;
  assign y12360 = ~n48192 ;
  assign y12361 = n48194 ;
  assign y12362 = ~n48196 ;
  assign y12363 = n48198 ;
  assign y12364 = n48199 ;
  assign y12365 = n48200 ;
  assign y12366 = ~n48203 ;
  assign y12367 = n48207 ;
  assign y12368 = n48211 ;
  assign y12369 = n48216 ;
  assign y12370 = ~n48220 ;
  assign y12371 = n48225 ;
  assign y12372 = n48226 ;
  assign y12373 = ~n48230 ;
  assign y12374 = ~n48235 ;
  assign y12375 = ~1'b0 ;
  assign y12376 = n48236 ;
  assign y12377 = n48243 ;
  assign y12378 = n48244 ;
  assign y12379 = n48246 ;
  assign y12380 = ~n48247 ;
  assign y12381 = ~n48253 ;
  assign y12382 = ~n48255 ;
  assign y12383 = n48256 ;
  assign y12384 = ~n48258 ;
  assign y12385 = ~1'b0 ;
  assign y12386 = ~1'b0 ;
  assign y12387 = ~n48260 ;
  assign y12388 = n48264 ;
  assign y12389 = ~n48265 ;
  assign y12390 = n48266 ;
  assign y12391 = ~n48272 ;
  assign y12392 = ~n48273 ;
  assign y12393 = ~n48274 ;
  assign y12394 = ~1'b0 ;
  assign y12395 = n48275 ;
  assign y12396 = ~n48276 ;
  assign y12397 = ~n48279 ;
  assign y12398 = ~n48284 ;
  assign y12399 = n48288 ;
  assign y12400 = ~n48293 ;
  assign y12401 = ~n48294 ;
  assign y12402 = ~n48296 ;
  assign y12403 = n48298 ;
  assign y12404 = n48300 ;
  assign y12405 = n48304 ;
  assign y12406 = ~n48307 ;
  assign y12407 = ~n48309 ;
  assign y12408 = n48310 ;
  assign y12409 = ~n48311 ;
  assign y12410 = ~n48313 ;
  assign y12411 = ~n48315 ;
  assign y12412 = n48317 ;
  assign y12413 = ~n48320 ;
  assign y12414 = ~n48325 ;
  assign y12415 = ~n48327 ;
  assign y12416 = ~n48328 ;
  assign y12417 = ~n48334 ;
  assign y12418 = ~n48338 ;
  assign y12419 = ~n48341 ;
  assign y12420 = ~n48345 ;
  assign y12421 = ~n48346 ;
  assign y12422 = n48350 ;
  assign y12423 = n48351 ;
  assign y12424 = n48355 ;
  assign y12425 = n48356 ;
  assign y12426 = n48357 ;
  assign y12427 = ~n48365 ;
  assign y12428 = n48368 ;
  assign y12429 = ~n48369 ;
  assign y12430 = ~n48374 ;
  assign y12431 = n48375 ;
  assign y12432 = ~n48378 ;
  assign y12433 = n48379 ;
  assign y12434 = ~n48380 ;
  assign y12435 = n48381 ;
  assign y12436 = ~n48382 ;
  assign y12437 = n48383 ;
  assign y12438 = ~n48386 ;
  assign y12439 = ~n48387 ;
  assign y12440 = n48389 ;
  assign y12441 = ~n48397 ;
  assign y12442 = ~n48405 ;
  assign y12443 = ~n48406 ;
  assign y12444 = n48409 ;
  assign y12445 = n48412 ;
  assign y12446 = n48414 ;
  assign y12447 = n48417 ;
  assign y12448 = n48419 ;
  assign y12449 = ~n48421 ;
  assign y12450 = ~n48428 ;
  assign y12451 = ~n48432 ;
  assign y12452 = n48433 ;
  assign y12453 = ~n48435 ;
  assign y12454 = n48437 ;
  assign y12455 = ~n48441 ;
  assign y12456 = ~n48443 ;
  assign y12457 = n48448 ;
  assign y12458 = ~1'b0 ;
  assign y12459 = ~n48449 ;
  assign y12460 = ~n48452 ;
  assign y12461 = n48453 ;
  assign y12462 = n48459 ;
  assign y12463 = n48460 ;
  assign y12464 = ~n48461 ;
  assign y12465 = ~n48462 ;
  assign y12466 = ~n48464 ;
  assign y12467 = ~n48465 ;
  assign y12468 = ~n48466 ;
  assign y12469 = ~n48468 ;
  assign y12470 = ~n48469 ;
  assign y12471 = ~n48471 ;
  assign y12472 = ~n48473 ;
  assign y12473 = n48475 ;
  assign y12474 = ~n48478 ;
  assign y12475 = ~n48481 ;
  assign y12476 = n48482 ;
  assign y12477 = n48484 ;
  assign y12478 = ~n48489 ;
  assign y12479 = ~1'b0 ;
  assign y12480 = ~n48494 ;
  assign y12481 = n48495 ;
  assign y12482 = ~n48496 ;
  assign y12483 = ~n48497 ;
  assign y12484 = n48498 ;
  assign y12485 = ~n48499 ;
  assign y12486 = ~1'b0 ;
  assign y12487 = ~n48500 ;
  assign y12488 = ~n48503 ;
  assign y12489 = n48505 ;
  assign y12490 = ~n48507 ;
  assign y12491 = ~n48509 ;
  assign y12492 = ~n48510 ;
  assign y12493 = ~n48511 ;
  assign y12494 = ~n48514 ;
  assign y12495 = n48518 ;
  assign y12496 = ~1'b0 ;
  assign y12497 = ~n48527 ;
  assign y12498 = n48528 ;
  assign y12499 = ~n48529 ;
  assign y12500 = ~n48535 ;
  assign y12501 = ~n48536 ;
  assign y12502 = ~n48539 ;
  assign y12503 = n48541 ;
  assign y12504 = ~1'b0 ;
  assign y12505 = ~n48546 ;
  assign y12506 = n48547 ;
  assign y12507 = ~n48548 ;
  assign y12508 = ~n48549 ;
  assign y12509 = ~n48550 ;
  assign y12510 = ~n48556 ;
  assign y12511 = n48557 ;
  assign y12512 = ~n48558 ;
  assign y12513 = ~1'b0 ;
  assign y12514 = ~n48560 ;
  assign y12515 = ~n48564 ;
  assign y12516 = n48566 ;
  assign y12517 = n48569 ;
  assign y12518 = n48570 ;
  assign y12519 = n48579 ;
  assign y12520 = n48583 ;
  assign y12521 = n48584 ;
  assign y12522 = ~1'b0 ;
  assign y12523 = n48591 ;
  assign y12524 = n48595 ;
  assign y12525 = n48598 ;
  assign y12526 = n48599 ;
  assign y12527 = ~n48600 ;
  assign y12528 = ~n48601 ;
  assign y12529 = ~n48605 ;
  assign y12530 = n48607 ;
  assign y12531 = ~n48608 ;
  assign y12532 = n48610 ;
  assign y12533 = ~n48612 ;
  assign y12534 = n48613 ;
  assign y12535 = ~n48615 ;
  assign y12536 = n48616 ;
  assign y12537 = ~n48617 ;
  assign y12538 = n48619 ;
  assign y12539 = n48621 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = ~n48622 ;
  assign y12542 = n48624 ;
  assign y12543 = n48626 ;
  assign y12544 = n48627 ;
  assign y12545 = n48629 ;
  assign y12546 = n48630 ;
  assign y12547 = n48632 ;
  assign y12548 = n48638 ;
  assign y12549 = ~n48639 ;
  assign y12550 = ~1'b0 ;
  assign y12551 = ~n48641 ;
  assign y12552 = ~n48645 ;
  assign y12553 = ~n48646 ;
  assign y12554 = n48648 ;
  assign y12555 = n48651 ;
  assign y12556 = n48653 ;
  assign y12557 = ~n48658 ;
  assign y12558 = n48660 ;
  assign y12559 = ~n48662 ;
  assign y12560 = ~n48671 ;
  assign y12561 = ~n48675 ;
  assign y12562 = ~n48676 ;
  assign y12563 = n48679 ;
  assign y12564 = ~n48681 ;
  assign y12565 = ~n48684 ;
  assign y12566 = n48687 ;
  assign y12567 = ~n48689 ;
  assign y12568 = ~n48693 ;
  assign y12569 = ~n48696 ;
  assign y12570 = ~n48697 ;
  assign y12571 = ~n48702 ;
  assign y12572 = n48703 ;
  assign y12573 = ~n48706 ;
  assign y12574 = ~n48707 ;
  assign y12575 = n48710 ;
  assign y12576 = ~n48711 ;
  assign y12577 = n48715 ;
  assign y12578 = ~n48717 ;
  assign y12579 = ~n48719 ;
  assign y12580 = n48725 ;
  assign y12581 = ~n48730 ;
  assign y12582 = n48731 ;
  assign y12583 = n48732 ;
  assign y12584 = ~n48734 ;
  assign y12585 = ~n48735 ;
  assign y12586 = n48738 ;
  assign y12587 = ~n48744 ;
  assign y12588 = ~n48745 ;
  assign y12589 = ~n48747 ;
  assign y12590 = ~n48748 ;
  assign y12591 = ~n48749 ;
  assign y12592 = n48754 ;
  assign y12593 = ~n48757 ;
  assign y12594 = ~n48760 ;
  assign y12595 = n48763 ;
  assign y12596 = ~n48765 ;
  assign y12597 = ~1'b0 ;
  assign y12598 = n48767 ;
  assign y12599 = ~n48771 ;
  assign y12600 = ~n48775 ;
  assign y12601 = n48776 ;
  assign y12602 = ~n48782 ;
  assign y12603 = n48786 ;
  assign y12604 = ~n48789 ;
  assign y12605 = n48791 ;
  assign y12606 = ~n48792 ;
  assign y12607 = n48794 ;
  assign y12608 = ~n48796 ;
  assign y12609 = ~n48800 ;
  assign y12610 = n48801 ;
  assign y12611 = ~n48802 ;
  assign y12612 = n48803 ;
  assign y12613 = n48806 ;
  assign y12614 = n48807 ;
  assign y12615 = n48810 ;
  assign y12616 = n48811 ;
  assign y12617 = n48815 ;
  assign y12618 = ~n48817 ;
  assign y12619 = ~n48820 ;
  assign y12620 = n48825 ;
  assign y12621 = ~n48829 ;
  assign y12622 = n48832 ;
  assign y12623 = ~n48835 ;
  assign y12624 = ~n48836 ;
  assign y12625 = n48840 ;
  assign y12626 = n48841 ;
  assign y12627 = n48842 ;
  assign y12628 = ~n48844 ;
  assign y12629 = n48853 ;
  assign y12630 = ~n48854 ;
  assign y12631 = n48860 ;
  assign y12632 = ~n48861 ;
  assign y12633 = n48864 ;
  assign y12634 = n48866 ;
  assign y12635 = n48867 ;
  assign y12636 = n48868 ;
  assign y12637 = ~1'b0 ;
  assign y12638 = n48873 ;
  assign y12639 = n48876 ;
  assign y12640 = ~n48877 ;
  assign y12641 = n48878 ;
  assign y12642 = ~n48884 ;
  assign y12643 = ~n48888 ;
  assign y12644 = n48890 ;
  assign y12645 = n48897 ;
  assign y12646 = ~n48898 ;
  assign y12647 = ~n48900 ;
  assign y12648 = ~n48903 ;
  assign y12649 = ~n48905 ;
  assign y12650 = ~n48906 ;
  assign y12651 = ~n48909 ;
  assign y12652 = ~n48917 ;
  assign y12653 = n48920 ;
  assign y12654 = n48924 ;
  assign y12655 = n48927 ;
  assign y12656 = n48928 ;
  assign y12657 = n48931 ;
  assign y12658 = ~n48934 ;
  assign y12659 = n48936 ;
  assign y12660 = ~n48937 ;
  assign y12661 = ~n48941 ;
  assign y12662 = ~n48942 ;
  assign y12663 = ~n48944 ;
  assign y12664 = ~n48947 ;
  assign y12665 = n48949 ;
  assign y12666 = ~n48954 ;
  assign y12667 = n48959 ;
  assign y12668 = n48960 ;
  assign y12669 = ~n48961 ;
  assign y12670 = n48963 ;
  assign y12671 = n48966 ;
  assign y12672 = n48967 ;
  assign y12673 = ~n48969 ;
  assign y12674 = n48971 ;
  assign y12675 = ~1'b0 ;
  assign y12676 = n48972 ;
  assign y12677 = n48973 ;
  assign y12678 = ~n48977 ;
  assign y12679 = ~n48980 ;
  assign y12680 = ~n48982 ;
  assign y12681 = n48987 ;
  assign y12682 = n48989 ;
  assign y12683 = n48990 ;
  assign y12684 = ~n48991 ;
  assign y12685 = n48996 ;
  assign y12686 = n48997 ;
  assign y12687 = n49002 ;
  assign y12688 = n49004 ;
  assign y12689 = ~n49006 ;
  assign y12690 = ~n49011 ;
  assign y12691 = ~n49015 ;
  assign y12692 = n49017 ;
  assign y12693 = ~n49020 ;
  assign y12694 = n49021 ;
  assign y12695 = ~n49022 ;
  assign y12696 = n49025 ;
  assign y12697 = n49029 ;
  assign y12698 = ~n49031 ;
  assign y12699 = n49032 ;
  assign y12700 = n49034 ;
  assign y12701 = n49035 ;
  assign y12702 = n49039 ;
  assign y12703 = ~n49040 ;
  assign y12704 = ~n49046 ;
  assign y12705 = n49048 ;
  assign y12706 = n49050 ;
  assign y12707 = n49055 ;
  assign y12708 = n49058 ;
  assign y12709 = ~n49061 ;
  assign y12710 = ~n37436 ;
  assign y12711 = n49064 ;
  assign y12712 = n49066 ;
  assign y12713 = ~n49068 ;
  assign y12714 = n49069 ;
  assign y12715 = ~n49072 ;
  assign y12716 = n49073 ;
  assign y12717 = n49077 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = n49081 ;
  assign y12720 = ~n49089 ;
  assign y12721 = ~n49095 ;
  assign y12722 = ~n49100 ;
  assign y12723 = n49102 ;
  assign y12724 = n49111 ;
  assign y12725 = n49115 ;
  assign y12726 = n31021 ;
  assign y12727 = ~n49121 ;
  assign y12728 = n49123 ;
  assign y12729 = n49125 ;
  assign y12730 = n49128 ;
  assign y12731 = n49131 ;
  assign y12732 = n49142 ;
  assign y12733 = n49143 ;
  assign y12734 = n49144 ;
  assign y12735 = n49145 ;
  assign y12736 = ~n49147 ;
  assign y12737 = ~n49152 ;
  assign y12738 = n49158 ;
  assign y12739 = n49160 ;
  assign y12740 = n49164 ;
  assign y12741 = n49165 ;
  assign y12742 = n49166 ;
  assign y12743 = ~n49167 ;
  assign y12744 = n49169 ;
  assign y12745 = ~n49171 ;
  assign y12746 = n49176 ;
  assign y12747 = n49177 ;
  assign y12748 = n49179 ;
  assign y12749 = ~n49183 ;
  assign y12750 = n49190 ;
  assign y12751 = n49191 ;
  assign y12752 = n49196 ;
  assign y12753 = ~n49202 ;
  assign y12754 = ~n49207 ;
  assign y12755 = ~n49210 ;
  assign y12756 = n49211 ;
  assign y12757 = n49212 ;
  assign y12758 = ~n49220 ;
  assign y12759 = ~n49222 ;
  assign y12760 = ~n49225 ;
  assign y12761 = n49229 ;
  assign y12762 = n49230 ;
  assign y12763 = ~n49232 ;
  assign y12764 = ~n49233 ;
  assign y12765 = n49234 ;
  assign y12766 = ~n49236 ;
  assign y12767 = ~n49240 ;
  assign y12768 = ~n49241 ;
  assign y12769 = n49245 ;
  assign y12770 = n49247 ;
  assign y12771 = n49249 ;
  assign y12772 = n49252 ;
  assign y12773 = n49254 ;
  assign y12774 = ~n49257 ;
  assign y12775 = ~n49259 ;
  assign y12776 = n49260 ;
  assign y12777 = n49261 ;
  assign y12778 = n49262 ;
  assign y12779 = n49267 ;
  assign y12780 = ~n49269 ;
  assign y12781 = n49271 ;
  assign y12782 = n49273 ;
  assign y12783 = ~n49276 ;
  assign y12784 = ~n49280 ;
  assign y12785 = n49282 ;
  assign y12786 = ~n49291 ;
  assign y12787 = ~n49292 ;
  assign y12788 = ~n49293 ;
  assign y12789 = ~n49294 ;
  assign y12790 = ~n49297 ;
  assign y12791 = ~n49298 ;
  assign y12792 = ~n49299 ;
  assign y12793 = ~n49301 ;
  assign y12794 = n49302 ;
  assign y12795 = n49304 ;
  assign y12796 = ~n49306 ;
  assign y12797 = n49309 ;
  assign y12798 = n49311 ;
  assign y12799 = n49312 ;
  assign y12800 = ~n49314 ;
  assign y12801 = n49319 ;
  assign y12802 = n49320 ;
  assign y12803 = n49321 ;
  assign y12804 = n49322 ;
  assign y12805 = n49327 ;
  assign y12806 = ~n49329 ;
  assign y12807 = ~n49335 ;
  assign y12808 = ~n49336 ;
  assign y12809 = n49339 ;
  assign y12810 = n49342 ;
  assign y12811 = ~n49346 ;
  assign y12812 = n49349 ;
  assign y12813 = n49351 ;
  assign y12814 = n49352 ;
  assign y12815 = ~n49355 ;
  assign y12816 = n49366 ;
  assign y12817 = n49368 ;
  assign y12818 = ~n49369 ;
  assign y12819 = n49372 ;
  assign y12820 = ~1'b0 ;
  assign y12821 = ~n49373 ;
  assign y12822 = n49375 ;
  assign y12823 = n49386 ;
  assign y12824 = n49387 ;
  assign y12825 = ~n49388 ;
  assign y12826 = n49389 ;
  assign y12827 = n49396 ;
  assign y12828 = n49402 ;
  assign y12829 = n49405 ;
  assign y12830 = ~1'b0 ;
  assign y12831 = ~n49408 ;
  assign y12832 = ~n49411 ;
  assign y12833 = n49413 ;
  assign y12834 = n49419 ;
  assign y12835 = n49420 ;
  assign y12836 = ~n49422 ;
  assign y12837 = n49423 ;
  assign y12838 = ~n49424 ;
  assign y12839 = ~n49427 ;
  assign y12840 = ~1'b0 ;
  assign y12841 = ~n49429 ;
  assign y12842 = n49431 ;
  assign y12843 = ~n49436 ;
  assign y12844 = n49440 ;
  assign y12845 = n49441 ;
  assign y12846 = ~n49442 ;
  assign y12847 = ~n49443 ;
  assign y12848 = ~n49446 ;
  assign y12849 = n49452 ;
  assign y12850 = n49454 ;
  assign y12851 = n49455 ;
  assign y12852 = n49456 ;
  assign y12853 = ~n49457 ;
  assign y12854 = ~n49459 ;
  assign y12855 = n49460 ;
  assign y12856 = ~n49462 ;
  assign y12857 = ~n49466 ;
  assign y12858 = ~n49467 ;
  assign y12859 = ~n49475 ;
  assign y12860 = n49482 ;
  assign y12861 = n49488 ;
  assign y12862 = n49490 ;
  assign y12863 = ~n49491 ;
  assign y12864 = n49493 ;
  assign y12865 = ~n49495 ;
  assign y12866 = n49497 ;
  assign y12867 = n49500 ;
  assign y12868 = n49501 ;
  assign y12869 = n49503 ;
  assign y12870 = n49506 ;
  assign y12871 = n49508 ;
  assign y12872 = n49509 ;
  assign y12873 = n49518 ;
  assign y12874 = ~n49519 ;
  assign y12875 = n49520 ;
  assign y12876 = n49522 ;
  assign y12877 = ~n49523 ;
  assign y12878 = n49524 ;
  assign y12879 = ~1'b0 ;
  assign y12880 = n49525 ;
  assign y12881 = ~n49526 ;
  assign y12882 = ~n49528 ;
  assign y12883 = n49530 ;
  assign y12884 = ~n49531 ;
  assign y12885 = ~n49533 ;
  assign y12886 = n49534 ;
  assign y12887 = n49536 ;
  assign y12888 = ~n49537 ;
  assign y12889 = ~n49541 ;
  assign y12890 = ~n49543 ;
  assign y12891 = n49544 ;
  assign y12892 = ~n49548 ;
  assign y12893 = ~n49549 ;
  assign y12894 = ~n49551 ;
  assign y12895 = n49553 ;
  assign y12896 = ~n49555 ;
  assign y12897 = ~n49556 ;
  assign y12898 = ~n49557 ;
  assign y12899 = n49559 ;
  assign y12900 = ~n49561 ;
  assign y12901 = ~1'b0 ;
  assign y12902 = ~n49562 ;
  assign y12903 = ~n49567 ;
  assign y12904 = n49573 ;
  assign y12905 = ~n49576 ;
  assign y12906 = n49577 ;
  assign y12907 = ~n49578 ;
  assign y12908 = n49582 ;
  assign y12909 = n49584 ;
  assign y12910 = ~1'b0 ;
  assign y12911 = ~n49588 ;
  assign y12912 = n49591 ;
  assign y12913 = ~n49592 ;
  assign y12914 = ~n49596 ;
  assign y12915 = n49598 ;
  assign y12916 = ~n49600 ;
  assign y12917 = n49602 ;
  assign y12918 = ~n49605 ;
  assign y12919 = ~n49608 ;
  assign y12920 = n49609 ;
  assign y12921 = n49611 ;
  assign y12922 = n49616 ;
  assign y12923 = n49618 ;
  assign y12924 = n49620 ;
  assign y12925 = n49621 ;
  assign y12926 = ~n49622 ;
  assign y12927 = n49624 ;
  assign y12928 = n49626 ;
  assign y12929 = ~n49629 ;
  assign y12930 = ~n49631 ;
  assign y12931 = ~1'b0 ;
  assign y12932 = ~n49634 ;
  assign y12933 = ~n49638 ;
  assign y12934 = ~n49639 ;
  assign y12935 = n49648 ;
  assign y12936 = n49651 ;
  assign y12937 = n49655 ;
  assign y12938 = n49656 ;
  assign y12939 = ~n49657 ;
  assign y12940 = n49663 ;
  assign y12941 = ~1'b0 ;
  assign y12942 = ~n49665 ;
  assign y12943 = ~n49666 ;
  assign y12944 = ~n49668 ;
  assign y12945 = ~n49671 ;
  assign y12946 = ~n49672 ;
  assign y12947 = ~n49674 ;
  assign y12948 = n49677 ;
  assign y12949 = ~n49680 ;
  assign y12950 = ~n49681 ;
  assign y12951 = n49683 ;
  assign y12952 = n49685 ;
  assign y12953 = n49686 ;
  assign y12954 = n49690 ;
  assign y12955 = ~n49691 ;
  assign y12956 = n49693 ;
  assign y12957 = ~n49698 ;
  assign y12958 = ~n49699 ;
  assign y12959 = ~n49706 ;
  assign y12960 = ~n49710 ;
  assign y12961 = ~n49714 ;
  assign y12962 = n49715 ;
  assign y12963 = ~n49718 ;
  assign y12964 = n49720 ;
  assign y12965 = n49721 ;
  assign y12966 = ~n49725 ;
  assign y12967 = ~n49726 ;
  assign y12968 = ~n49728 ;
  assign y12969 = n49731 ;
  assign y12970 = n49733 ;
  assign y12971 = ~1'b0 ;
  assign y12972 = n49737 ;
  assign y12973 = ~n49738 ;
  assign y12974 = ~n49742 ;
  assign y12975 = ~n49745 ;
  assign y12976 = ~n49750 ;
  assign y12977 = n49751 ;
  assign y12978 = n49753 ;
  assign y12979 = ~n49754 ;
  assign y12980 = ~n49758 ;
  assign y12981 = ~n49761 ;
  assign y12982 = ~n49762 ;
  assign y12983 = n49763 ;
  assign y12984 = n49764 ;
  assign y12985 = n49766 ;
  assign y12986 = ~n49767 ;
  assign y12987 = ~n49768 ;
  assign y12988 = ~n49769 ;
  assign y12989 = ~n49770 ;
  assign y12990 = ~n49771 ;
  assign y12991 = ~n49773 ;
  assign y12992 = ~1'b0 ;
  assign y12993 = ~n49774 ;
  assign y12994 = n49777 ;
  assign y12995 = ~n49779 ;
  assign y12996 = ~n49782 ;
  assign y12997 = ~n49784 ;
  assign y12998 = ~n49786 ;
  assign y12999 = ~n49789 ;
  assign y13000 = n49792 ;
  assign y13001 = n49793 ;
  assign y13002 = n49797 ;
  assign y13003 = ~n49799 ;
  assign y13004 = ~n49800 ;
  assign y13005 = ~n49801 ;
  assign y13006 = n49805 ;
  assign y13007 = ~n49806 ;
  assign y13008 = ~n49808 ;
  assign y13009 = n49809 ;
  assign y13010 = n49814 ;
  assign y13011 = ~n49817 ;
  assign y13012 = n49819 ;
  assign y13013 = ~n49824 ;
  assign y13014 = n49827 ;
  assign y13015 = ~n49832 ;
  assign y13016 = n49834 ;
  assign y13017 = ~n49836 ;
  assign y13018 = n49842 ;
  assign y13019 = n49843 ;
  assign y13020 = n49844 ;
  assign y13021 = ~1'b0 ;
  assign y13022 = ~1'b0 ;
  assign y13023 = n49845 ;
  assign y13024 = ~n49848 ;
  assign y13025 = n49851 ;
  assign y13026 = ~n49852 ;
  assign y13027 = ~n49854 ;
  assign y13028 = n49855 ;
  assign y13029 = ~n49856 ;
  assign y13030 = ~n49858 ;
  assign y13031 = n49859 ;
  assign y13032 = ~1'b0 ;
  assign y13033 = ~n49861 ;
  assign y13034 = ~n49863 ;
  assign y13035 = n49871 ;
  assign y13036 = ~n49872 ;
  assign y13037 = n49873 ;
  assign y13038 = n49874 ;
  assign y13039 = n49876 ;
  assign y13040 = ~n49879 ;
  assign y13041 = n49882 ;
  assign y13042 = ~1'b0 ;
  assign y13043 = ~n49885 ;
  assign y13044 = ~n49887 ;
  assign y13045 = ~n49890 ;
  assign y13046 = ~n49892 ;
  assign y13047 = ~n49893 ;
  assign y13048 = n49898 ;
  assign y13049 = n49901 ;
  assign y13050 = ~n49902 ;
  assign y13051 = n49915 ;
  assign y13052 = n49917 ;
  assign y13053 = n49922 ;
  assign y13054 = ~n49923 ;
  assign y13055 = ~n49926 ;
  assign y13056 = n49929 ;
  assign y13057 = n49930 ;
  assign y13058 = ~n49936 ;
  assign y13059 = n49940 ;
  assign y13060 = ~n49942 ;
  assign y13061 = ~n49946 ;
  assign y13062 = ~n49948 ;
  assign y13063 = n49949 ;
  assign y13064 = n49950 ;
  assign y13065 = n49951 ;
  assign y13066 = n49954 ;
  assign y13067 = ~n49955 ;
  assign y13068 = ~n49956 ;
  assign y13069 = n49958 ;
  assign y13070 = ~n49959 ;
  assign y13071 = ~n49963 ;
  assign y13072 = n49967 ;
  assign y13073 = ~1'b0 ;
  assign y13074 = n49969 ;
  assign y13075 = n49970 ;
  assign y13076 = n49972 ;
  assign y13077 = n49973 ;
  assign y13078 = n49974 ;
  assign y13079 = n49976 ;
  assign y13080 = n49984 ;
  assign y13081 = n49986 ;
  assign y13082 = ~1'b0 ;
  assign y13083 = ~n49989 ;
  assign y13084 = n49991 ;
  assign y13085 = n49998 ;
  assign y13086 = n49999 ;
  assign y13087 = ~n50000 ;
  assign y13088 = n50001 ;
  assign y13089 = n50003 ;
  assign y13090 = n50005 ;
  assign y13091 = ~n50006 ;
  assign y13092 = ~n50008 ;
  assign y13093 = n50015 ;
  assign y13094 = n50016 ;
  assign y13095 = n50018 ;
  assign y13096 = ~n50020 ;
  assign y13097 = n50028 ;
  assign y13098 = n50034 ;
  assign y13099 = ~n50036 ;
  assign y13100 = n50038 ;
  assign y13101 = ~n50040 ;
  assign y13102 = n50043 ;
  assign y13103 = ~n50045 ;
  assign y13104 = n31417 ;
  assign y13105 = ~n50046 ;
  assign y13106 = n50047 ;
  assign y13107 = ~n50051 ;
  assign y13108 = ~n50052 ;
  assign y13109 = ~n50055 ;
  assign y13110 = n50057 ;
  assign y13111 = ~1'b0 ;
  assign y13112 = n50060 ;
  assign y13113 = n50062 ;
  assign y13114 = n50065 ;
  assign y13115 = ~n50066 ;
  assign y13116 = n50070 ;
  assign y13117 = ~n50071 ;
  assign y13118 = ~n50073 ;
  assign y13119 = n50078 ;
  assign y13120 = n50081 ;
  assign y13121 = ~n50082 ;
  assign y13122 = ~n50084 ;
  assign y13123 = ~n50086 ;
  assign y13124 = ~n50087 ;
  assign y13125 = n50088 ;
  assign y13126 = n50089 ;
  assign y13127 = ~n50095 ;
  assign y13128 = ~n50097 ;
  assign y13129 = ~n50099 ;
  assign y13130 = ~n50100 ;
  assign y13131 = ~n50102 ;
  assign y13132 = n50108 ;
  assign y13133 = ~n50110 ;
  assign y13134 = n50117 ;
  assign y13135 = n50119 ;
  assign y13136 = ~n50120 ;
  assign y13137 = n50121 ;
  assign y13138 = n50122 ;
  assign y13139 = ~n50123 ;
  assign y13140 = ~n50126 ;
  assign y13141 = ~n50129 ;
  assign y13142 = ~n50132 ;
  assign y13143 = n50133 ;
  assign y13144 = ~n50136 ;
  assign y13145 = ~n50137 ;
  assign y13146 = ~n50144 ;
  assign y13147 = ~n50148 ;
  assign y13148 = ~n50151 ;
  assign y13149 = ~n50158 ;
  assign y13150 = ~n50160 ;
  assign y13151 = n50161 ;
  assign y13152 = ~n50163 ;
  assign y13153 = ~n50164 ;
  assign y13154 = n50166 ;
  assign y13155 = ~n50168 ;
  assign y13156 = ~n50172 ;
  assign y13157 = ~n50176 ;
  assign y13158 = n50177 ;
  assign y13159 = ~n50182 ;
  assign y13160 = ~1'b0 ;
  assign y13161 = ~n50183 ;
  assign y13162 = ~n50188 ;
  assign y13163 = ~n50190 ;
  assign y13164 = n50192 ;
  assign y13165 = n50193 ;
  assign y13166 = ~n50194 ;
  assign y13167 = n50197 ;
  assign y13168 = ~n50202 ;
  assign y13169 = ~1'b0 ;
  assign y13170 = ~n50203 ;
  assign y13171 = ~n50204 ;
  assign y13172 = ~n50205 ;
  assign y13173 = n50207 ;
  assign y13174 = n50208 ;
  assign y13175 = n50209 ;
  assign y13176 = n50210 ;
  assign y13177 = n50214 ;
  assign y13178 = n50218 ;
  assign y13179 = ~n50219 ;
  assign y13180 = n50223 ;
  assign y13181 = ~n50228 ;
  assign y13182 = n50231 ;
  assign y13183 = n50233 ;
  assign y13184 = ~n50238 ;
  assign y13185 = ~n50239 ;
  assign y13186 = n50241 ;
  assign y13187 = n50246 ;
  assign y13188 = n50249 ;
  assign y13189 = n50250 ;
  assign y13190 = n50251 ;
  assign y13191 = ~n50254 ;
  assign y13192 = n50261 ;
  assign y13193 = ~n50262 ;
  assign y13194 = n50266 ;
  assign y13195 = n50267 ;
  assign y13196 = ~n50269 ;
  assign y13197 = ~n50271 ;
  assign y13198 = ~n50273 ;
  assign y13199 = ~n50274 ;
  assign y13200 = ~n50275 ;
  assign y13201 = ~n50276 ;
  assign y13202 = n50280 ;
  assign y13203 = n50284 ;
  assign y13204 = ~1'b0 ;
  assign y13205 = n50286 ;
  assign y13206 = ~n50289 ;
  assign y13207 = n50290 ;
  assign y13208 = ~n50291 ;
  assign y13209 = n50295 ;
  assign y13210 = ~n50296 ;
  assign y13211 = n50297 ;
  assign y13212 = n50299 ;
  assign y13213 = ~n50301 ;
  assign y13214 = ~n50302 ;
  assign y13215 = n50303 ;
  assign y13216 = n50305 ;
  assign y13217 = n50310 ;
  assign y13218 = n50311 ;
  assign y13219 = n50313 ;
  assign y13220 = ~n50314 ;
  assign y13221 = n50317 ;
  assign y13222 = n50318 ;
  assign y13223 = ~1'b0 ;
  assign y13224 = n50320 ;
  assign y13225 = n50323 ;
  assign y13226 = n50324 ;
  assign y13227 = n50328 ;
  assign y13228 = ~n50330 ;
  assign y13229 = ~n50331 ;
  assign y13230 = n50335 ;
  assign y13231 = n50337 ;
  assign y13232 = n50339 ;
  assign y13233 = n50341 ;
  assign y13234 = n50344 ;
  assign y13235 = ~1'b0 ;
  assign y13236 = ~n50346 ;
  assign y13237 = n50347 ;
  assign y13238 = n50348 ;
  assign y13239 = ~n50351 ;
  assign y13240 = ~n50353 ;
  assign y13241 = ~n50358 ;
  assign y13242 = ~n50360 ;
  assign y13243 = ~1'b0 ;
  assign y13244 = n50362 ;
  assign y13245 = ~n50364 ;
  assign y13246 = ~n50365 ;
  assign y13247 = ~n50367 ;
  assign y13248 = n50368 ;
  assign y13249 = n50369 ;
  assign y13250 = ~n50372 ;
  assign y13251 = ~n50375 ;
  assign y13252 = n50377 ;
  assign y13253 = n50380 ;
  assign y13254 = n50381 ;
  assign y13255 = ~n50384 ;
  assign y13256 = ~n50386 ;
  assign y13257 = n50390 ;
  assign y13258 = ~n50392 ;
  assign y13259 = ~n50393 ;
  assign y13260 = n50394 ;
  assign y13261 = ~n50396 ;
  assign y13262 = ~n50398 ;
  assign y13263 = n50402 ;
  assign y13264 = ~n50404 ;
  assign y13265 = ~n50407 ;
  assign y13266 = ~n50408 ;
  assign y13267 = n50410 ;
  assign y13268 = ~n50413 ;
  assign y13269 = ~1'b0 ;
  assign y13270 = n50415 ;
  assign y13271 = ~n50422 ;
  assign y13272 = n50423 ;
  assign y13273 = ~n50424 ;
  assign y13274 = n50425 ;
  assign y13275 = ~n50426 ;
  assign y13276 = ~n50430 ;
  assign y13277 = n50435 ;
  assign y13278 = ~n50440 ;
  assign y13279 = n50449 ;
  assign y13280 = ~n50451 ;
  assign y13281 = ~n50453 ;
  assign y13282 = ~n50455 ;
  assign y13283 = n50456 ;
  assign y13284 = n50458 ;
  assign y13285 = ~n50461 ;
  assign y13286 = n50462 ;
  assign y13287 = n50464 ;
  assign y13288 = n50465 ;
  assign y13289 = n50466 ;
  assign y13290 = 1'b0 ;
  assign y13291 = n50468 ;
  assign y13292 = n50469 ;
  assign y13293 = ~n50470 ;
  assign y13294 = ~n50471 ;
  assign y13295 = ~n50472 ;
  assign y13296 = n50476 ;
  assign y13297 = n50478 ;
  assign y13298 = ~n50479 ;
  assign y13299 = ~n50481 ;
  assign y13300 = n50485 ;
  assign y13301 = n50487 ;
  assign y13302 = n50488 ;
  assign y13303 = ~n50491 ;
  assign y13304 = ~n50496 ;
  assign y13305 = n50497 ;
  assign y13306 = n50500 ;
  assign y13307 = n28841 ;
  assign y13308 = n50502 ;
  assign y13309 = ~n50504 ;
  assign y13310 = ~1'b0 ;
  assign y13311 = ~n50506 ;
  assign y13312 = n50507 ;
  assign y13313 = n50509 ;
  assign y13314 = n50511 ;
  assign y13315 = ~n50513 ;
  assign y13316 = n50514 ;
  assign y13317 = ~n50516 ;
  assign y13318 = n50517 ;
  assign y13319 = ~n50530 ;
  assign y13320 = ~n50536 ;
  assign y13321 = n50538 ;
  assign y13322 = ~n50542 ;
  assign y13323 = n50543 ;
  assign y13324 = n50544 ;
  assign y13325 = ~n50545 ;
  assign y13326 = ~n50546 ;
  assign y13327 = n50547 ;
  assign y13328 = n50549 ;
  assign y13329 = ~n50550 ;
  assign y13330 = ~n50553 ;
  assign y13331 = ~n50556 ;
  assign y13332 = ~n50565 ;
  assign y13333 = n50567 ;
  assign y13334 = ~n50568 ;
  assign y13335 = n50570 ;
  assign y13336 = n50571 ;
  assign y13337 = n50572 ;
  assign y13338 = ~n50573 ;
  assign y13339 = ~n50575 ;
  assign y13340 = ~1'b0 ;
  assign y13341 = ~1'b0 ;
  assign y13342 = ~n50576 ;
  assign y13343 = ~n50580 ;
  assign y13344 = n50583 ;
  assign y13345 = ~n50588 ;
  assign y13346 = ~n50589 ;
  assign y13347 = ~n50591 ;
  assign y13348 = n50595 ;
  assign y13349 = n50597 ;
  assign y13350 = ~n50599 ;
  assign y13351 = ~n50600 ;
  assign y13352 = ~n50602 ;
  assign y13353 = n50603 ;
  assign y13354 = ~n50604 ;
  assign y13355 = ~n50609 ;
  assign y13356 = ~n50611 ;
  assign y13357 = ~n50614 ;
  assign y13358 = n50615 ;
  assign y13359 = n50617 ;
  assign y13360 = n50619 ;
  assign y13361 = ~n50620 ;
  assign y13362 = ~n50623 ;
  assign y13363 = n50627 ;
  assign y13364 = ~n50633 ;
  assign y13365 = n50635 ;
  assign y13366 = n50636 ;
  assign y13367 = n50638 ;
  assign y13368 = ~n50642 ;
  assign y13369 = n50643 ;
  assign y13370 = ~n50648 ;
  assign y13371 = ~n50657 ;
  assign y13372 = ~n50658 ;
  assign y13373 = ~n50659 ;
  assign y13374 = ~n50663 ;
  assign y13375 = n50666 ;
  assign y13376 = n50669 ;
  assign y13377 = ~1'b0 ;
  assign y13378 = ~n50670 ;
  assign y13379 = n50675 ;
  assign y13380 = n50677 ;
  assign y13381 = ~n50681 ;
  assign y13382 = n50682 ;
  assign y13383 = n50683 ;
  assign y13384 = ~1'b0 ;
  assign y13385 = ~n50685 ;
  assign y13386 = n50691 ;
  assign y13387 = n50692 ;
  assign y13388 = n50697 ;
  assign y13389 = n50698 ;
  assign y13390 = ~n50700 ;
  assign y13391 = ~n50704 ;
  assign y13392 = n50705 ;
  assign y13393 = ~1'b0 ;
  assign y13394 = ~n50712 ;
  assign y13395 = ~n50713 ;
  assign y13396 = n50714 ;
  assign y13397 = ~n50720 ;
  assign y13398 = ~n50722 ;
  assign y13399 = ~n50726 ;
  assign y13400 = ~n50727 ;
  assign y13401 = n50728 ;
  assign y13402 = n50729 ;
  assign y13403 = ~n50734 ;
  assign y13404 = ~1'b0 ;
  assign y13405 = n50735 ;
  assign y13406 = ~n50737 ;
  assign y13407 = n50740 ;
  assign y13408 = ~n50742 ;
  assign y13409 = n50743 ;
  assign y13410 = n50746 ;
  assign y13411 = n50748 ;
  assign y13412 = ~n50753 ;
  assign y13413 = n50757 ;
  assign y13414 = n50758 ;
  assign y13415 = ~1'b0 ;
  assign y13416 = ~1'b0 ;
  assign y13417 = n50759 ;
  assign y13418 = n50761 ;
  assign y13419 = n50766 ;
  assign y13420 = n50767 ;
  assign y13421 = ~n50773 ;
  assign y13422 = ~n50774 ;
  assign y13423 = ~n50780 ;
  assign y13424 = n50781 ;
  assign y13425 = ~n50785 ;
  assign y13426 = ~n50787 ;
  assign y13427 = n50789 ;
  assign y13428 = n50790 ;
  assign y13429 = n50792 ;
  assign y13430 = ~n50796 ;
  assign y13431 = n50800 ;
  assign y13432 = n50803 ;
  assign y13433 = ~n50807 ;
  assign y13434 = ~n50808 ;
  assign y13435 = ~n50812 ;
  assign y13436 = n50814 ;
  assign y13437 = ~n50816 ;
  assign y13438 = ~n50818 ;
  assign y13439 = n50820 ;
  assign y13440 = n50822 ;
  assign y13441 = n50827 ;
  assign y13442 = n50828 ;
  assign y13443 = n50829 ;
  assign y13444 = ~n50833 ;
  assign y13445 = ~n50834 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = ~n50836 ;
  assign y13448 = ~n50837 ;
  assign y13449 = n50838 ;
  assign y13450 = ~n50841 ;
  assign y13451 = n50842 ;
  assign y13452 = ~n50843 ;
  assign y13453 = n50845 ;
  assign y13454 = n50846 ;
  assign y13455 = ~1'b0 ;
  assign y13456 = ~n50848 ;
  assign y13457 = ~n50850 ;
  assign y13458 = ~n50851 ;
  assign y13459 = ~n50855 ;
  assign y13460 = n50856 ;
  assign y13461 = ~n50859 ;
  assign y13462 = ~n50860 ;
  assign y13463 = n50861 ;
  assign y13464 = ~n50863 ;
  assign y13465 = ~1'b0 ;
  assign y13466 = ~1'b0 ;
  assign y13467 = n50867 ;
  assign y13468 = n50871 ;
  assign y13469 = n50872 ;
  assign y13470 = n50874 ;
  assign y13471 = ~n50879 ;
  assign y13472 = ~n50881 ;
  assign y13473 = ~n50883 ;
  assign y13474 = n50884 ;
  assign y13475 = n50886 ;
  assign y13476 = ~n50887 ;
  assign y13477 = n50888 ;
  assign y13478 = ~n50892 ;
  assign y13479 = ~n50893 ;
  assign y13480 = ~n50894 ;
  assign y13481 = n50901 ;
  assign y13482 = n50902 ;
  assign y13483 = ~n50905 ;
  assign y13484 = ~n50908 ;
  assign y13485 = ~n50910 ;
  assign y13486 = n50914 ;
  assign y13487 = ~n50917 ;
  assign y13488 = n50918 ;
  assign y13489 = ~n50921 ;
  assign y13490 = n26093 ;
  assign y13491 = ~n50924 ;
  assign y13492 = ~n50925 ;
  assign y13493 = n50928 ;
  assign y13494 = n50931 ;
  assign y13495 = ~n50937 ;
  assign y13496 = n50939 ;
  assign y13497 = n50941 ;
  assign y13498 = ~n50942 ;
  assign y13499 = ~n50945 ;
  assign y13500 = n50949 ;
  assign y13501 = n50950 ;
  assign y13502 = n50951 ;
  assign y13503 = n50954 ;
  assign y13504 = n50958 ;
  assign y13505 = ~n50960 ;
  assign y13506 = n50962 ;
  assign y13507 = ~n50965 ;
  assign y13508 = n50968 ;
  assign y13509 = n50969 ;
  assign y13510 = n50971 ;
  assign y13511 = ~n50978 ;
  assign y13512 = n50979 ;
  assign y13513 = ~1'b0 ;
  assign y13514 = ~n50981 ;
  assign y13515 = n50982 ;
  assign y13516 = ~n50985 ;
  assign y13517 = ~n50986 ;
  assign y13518 = n50990 ;
  assign y13519 = n50993 ;
  assign y13520 = ~n50994 ;
  assign y13521 = n50995 ;
  assign y13522 = n51001 ;
  assign y13523 = n51005 ;
  assign y13524 = ~n51009 ;
  assign y13525 = n51012 ;
  assign y13526 = ~n51014 ;
  assign y13527 = n51016 ;
  assign y13528 = ~n51017 ;
  assign y13529 = n51021 ;
  assign y13530 = ~n51022 ;
  assign y13531 = n51024 ;
  assign y13532 = n51026 ;
  assign y13533 = ~n51027 ;
  assign y13534 = ~n51029 ;
  assign y13535 = n51033 ;
  assign y13536 = n51035 ;
  assign y13537 = n51036 ;
  assign y13538 = ~n51038 ;
  assign y13539 = ~n51040 ;
  assign y13540 = n51045 ;
  assign y13541 = n51049 ;
  assign y13542 = ~n51053 ;
  assign y13543 = n51057 ;
  assign y13544 = ~n51058 ;
  assign y13545 = n51061 ;
  assign y13546 = ~n51063 ;
  assign y13547 = ~n51064 ;
  assign y13548 = n51070 ;
  assign y13549 = ~n51072 ;
  assign y13550 = n51074 ;
  assign y13551 = ~n51079 ;
  assign y13552 = n51080 ;
  assign y13553 = n51082 ;
  assign y13554 = ~n51084 ;
  assign y13555 = n51086 ;
  assign y13556 = n51090 ;
  assign y13557 = ~n51092 ;
  assign y13558 = n51094 ;
  assign y13559 = ~n51095 ;
  assign y13560 = ~n51102 ;
  assign y13561 = n51103 ;
  assign y13562 = n51104 ;
  assign y13563 = ~n51106 ;
  assign y13564 = n51109 ;
  assign y13565 = ~n51111 ;
  assign y13566 = ~n51113 ;
  assign y13567 = n51116 ;
  assign y13568 = ~n51122 ;
  assign y13569 = n51129 ;
  assign y13570 = ~n51130 ;
  assign y13571 = ~n51136 ;
  assign y13572 = ~n51138 ;
  assign y13573 = ~n51140 ;
  assign y13574 = n51141 ;
  assign y13575 = ~n51143 ;
  assign y13576 = n51145 ;
  assign y13577 = n51153 ;
  assign y13578 = ~n51155 ;
  assign y13579 = ~n51156 ;
  assign y13580 = n51162 ;
  assign y13581 = n51166 ;
  assign y13582 = ~n51167 ;
  assign y13583 = ~n51168 ;
  assign y13584 = ~n51169 ;
  assign y13585 = n51170 ;
  assign y13586 = n51172 ;
  assign y13587 = ~n51174 ;
  assign y13588 = n51175 ;
  assign y13589 = ~n51176 ;
  assign y13590 = n51182 ;
  assign y13591 = ~n51185 ;
  assign y13592 = ~n51187 ;
  assign y13593 = ~n51192 ;
  assign y13594 = n51195 ;
  assign y13595 = n51198 ;
  assign y13596 = ~n51201 ;
  assign y13597 = n51202 ;
  assign y13598 = n51203 ;
  assign y13599 = n51206 ;
  assign y13600 = ~n51207 ;
  assign y13601 = ~n51210 ;
  assign y13602 = n51211 ;
  assign y13603 = ~n51214 ;
  assign y13604 = ~n51215 ;
  assign y13605 = ~n51218 ;
  assign y13606 = ~1'b0 ;
  assign y13607 = ~n51222 ;
  assign y13608 = n51226 ;
  assign y13609 = ~1'b0 ;
  assign y13610 = n51228 ;
  assign y13611 = ~n51230 ;
  assign y13612 = ~n51231 ;
  assign y13613 = n51232 ;
  assign y13614 = ~n51235 ;
  assign y13615 = ~n51236 ;
  assign y13616 = ~n51237 ;
  assign y13617 = ~1'b0 ;
  assign y13618 = ~1'b0 ;
  assign y13619 = ~n51238 ;
  assign y13620 = ~n51241 ;
  assign y13621 = n51242 ;
  assign y13622 = ~n51243 ;
  assign y13623 = n51244 ;
  assign y13624 = n51245 ;
  assign y13625 = ~n51248 ;
  assign y13626 = ~1'b0 ;
  assign y13627 = n51249 ;
  assign y13628 = n51251 ;
  assign y13629 = n51254 ;
  assign y13630 = ~n51255 ;
  assign y13631 = ~n51256 ;
  assign y13632 = ~n51258 ;
  assign y13633 = n51259 ;
  assign y13634 = n51261 ;
  assign y13635 = n51262 ;
  assign y13636 = n51264 ;
  assign y13637 = ~1'b0 ;
  assign y13638 = ~n51268 ;
  assign y13639 = n51269 ;
  assign y13640 = ~n51271 ;
  assign y13641 = n51272 ;
  assign y13642 = n51278 ;
  assign y13643 = n51279 ;
  assign y13644 = ~n51280 ;
  assign y13645 = n51282 ;
  assign y13646 = ~n51286 ;
  assign y13647 = ~1'b0 ;
  assign y13648 = n51287 ;
  assign y13649 = ~n51288 ;
  assign y13650 = n51289 ;
  assign y13651 = ~n51291 ;
  assign y13652 = ~n51292 ;
  assign y13653 = n51293 ;
  assign y13654 = n51295 ;
  assign y13655 = ~n51296 ;
  assign y13656 = n51298 ;
  assign y13657 = ~n51299 ;
  assign y13658 = n51303 ;
  assign y13659 = n51304 ;
  assign y13660 = ~n51305 ;
  assign y13661 = n51315 ;
  assign y13662 = ~n51317 ;
  assign y13663 = n51319 ;
  assign y13664 = ~n51322 ;
  assign y13665 = ~n51323 ;
  assign y13666 = ~1'b0 ;
  assign y13667 = n51324 ;
  assign y13668 = n51329 ;
  assign y13669 = ~n51332 ;
  assign y13670 = ~n51337 ;
  assign y13671 = ~n51339 ;
  assign y13672 = n51341 ;
  assign y13673 = ~n51343 ;
  assign y13674 = n51344 ;
  assign y13675 = ~n51345 ;
  assign y13676 = ~n51350 ;
  assign y13677 = n51353 ;
  assign y13678 = ~n51356 ;
  assign y13679 = n51357 ;
  assign y13680 = ~n51358 ;
  assign y13681 = n51361 ;
  assign y13682 = ~n51366 ;
  assign y13683 = n51367 ;
  assign y13684 = n51368 ;
  assign y13685 = n51370 ;
  assign y13686 = n51373 ;
  assign y13687 = n51375 ;
  assign y13688 = n51376 ;
  assign y13689 = n51380 ;
  assign y13690 = ~n51384 ;
  assign y13691 = n51386 ;
  assign y13692 = n51388 ;
  assign y13693 = n51391 ;
  assign y13694 = n51392 ;
  assign y13695 = ~n51395 ;
  assign y13696 = ~n51396 ;
  assign y13697 = n51397 ;
  assign y13698 = n51399 ;
  assign y13699 = ~n51401 ;
  assign y13700 = ~n51404 ;
  assign y13701 = n51406 ;
  assign y13702 = n51407 ;
  assign y13703 = ~n51410 ;
  assign y13704 = n51412 ;
  assign y13705 = n51416 ;
  assign y13706 = ~n51418 ;
  assign y13707 = n51419 ;
  assign y13708 = n51421 ;
  assign y13709 = n51425 ;
  assign y13710 = n51427 ;
  assign y13711 = ~n51429 ;
  assign y13712 = n51430 ;
  assign y13713 = ~n51433 ;
  assign y13714 = n51439 ;
  assign y13715 = ~n51440 ;
  assign y13716 = n51441 ;
  assign y13717 = ~n51442 ;
  assign y13718 = ~n51444 ;
  assign y13719 = ~n51449 ;
  assign y13720 = n51452 ;
  assign y13721 = ~n51454 ;
  assign y13722 = n51457 ;
  assign y13723 = n51459 ;
  assign y13724 = n51461 ;
  assign y13725 = n51463 ;
  assign y13726 = ~n51464 ;
  assign y13727 = ~n51465 ;
  assign y13728 = ~n51466 ;
  assign y13729 = n51467 ;
  assign y13730 = n51470 ;
  assign y13731 = n51471 ;
  assign y13732 = ~1'b0 ;
  assign y13733 = ~n51473 ;
  assign y13734 = n51476 ;
  assign y13735 = ~n51478 ;
  assign y13736 = n51480 ;
  assign y13737 = n51481 ;
  assign y13738 = ~n51482 ;
  assign y13739 = ~n51484 ;
  assign y13740 = n51486 ;
  assign y13741 = ~n51491 ;
  assign y13742 = ~1'b0 ;
  assign y13743 = n51493 ;
  assign y13744 = ~n51494 ;
  assign y13745 = n51495 ;
  assign y13746 = ~n51496 ;
  assign y13747 = n51497 ;
  assign y13748 = n51502 ;
  assign y13749 = n51503 ;
  assign y13750 = ~n51505 ;
  assign y13751 = n51507 ;
  assign y13752 = ~n51509 ;
  assign y13753 = n51511 ;
  assign y13754 = n51516 ;
  assign y13755 = n51519 ;
  assign y13756 = n51524 ;
  assign y13757 = ~n51526 ;
  assign y13758 = n51528 ;
  assign y13759 = ~n51529 ;
  assign y13760 = n51534 ;
  assign y13761 = ~n51535 ;
  assign y13762 = n51541 ;
  assign y13763 = ~n51545 ;
  assign y13764 = ~n51548 ;
  assign y13765 = n51551 ;
  assign y13766 = ~n51552 ;
  assign y13767 = n51554 ;
  assign y13768 = n51566 ;
  assign y13769 = ~n51567 ;
  assign y13770 = ~n51571 ;
  assign y13771 = n51573 ;
  assign y13772 = n51574 ;
  assign y13773 = n51579 ;
  assign y13774 = ~n51583 ;
  assign y13775 = ~n51586 ;
  assign y13776 = ~n51589 ;
  assign y13777 = n51590 ;
  assign y13778 = ~n51591 ;
  assign y13779 = n51592 ;
  assign y13780 = n51594 ;
  assign y13781 = ~n51598 ;
  assign y13782 = ~n51600 ;
  assign y13783 = ~n51604 ;
  assign y13784 = ~n51615 ;
  assign y13785 = n51616 ;
  assign y13786 = n51618 ;
  assign y13787 = ~n51621 ;
  assign y13788 = n51622 ;
  assign y13789 = ~n51623 ;
  assign y13790 = ~n51624 ;
  assign y13791 = n51625 ;
  assign y13792 = ~n51628 ;
  assign y13793 = n51635 ;
  assign y13794 = n51638 ;
  assign y13795 = n51640 ;
  assign y13796 = n51641 ;
  assign y13797 = n51642 ;
  assign y13798 = ~n51643 ;
  assign y13799 = ~n51644 ;
  assign y13800 = ~n51645 ;
  assign y13801 = ~n51649 ;
  assign y13802 = ~n51650 ;
  assign y13803 = ~n51652 ;
  assign y13804 = ~n51654 ;
  assign y13805 = ~n51656 ;
  assign y13806 = n51657 ;
  assign y13807 = n51659 ;
  assign y13808 = ~n51661 ;
  assign y13809 = n51662 ;
  assign y13810 = n51663 ;
  assign y13811 = n51667 ;
  assign y13812 = ~n51670 ;
  assign y13813 = ~1'b0 ;
  assign y13814 = n51671 ;
  assign y13815 = n51672 ;
  assign y13816 = ~n51674 ;
  assign y13817 = n51676 ;
  assign y13818 = ~n51684 ;
  assign y13819 = ~n51685 ;
  assign y13820 = n51688 ;
  assign y13821 = ~n51690 ;
  assign y13822 = ~1'b0 ;
  assign y13823 = ~n51694 ;
  assign y13824 = ~n51698 ;
  assign y13825 = ~n51699 ;
  assign y13826 = n51703 ;
  assign y13827 = n51704 ;
  assign y13828 = ~n51705 ;
  assign y13829 = ~n51706 ;
  assign y13830 = n51707 ;
  assign y13831 = n51708 ;
  assign y13832 = n51712 ;
  assign y13833 = n51714 ;
  assign y13834 = ~n51715 ;
  assign y13835 = n51716 ;
  assign y13836 = n51718 ;
  assign y13837 = n51721 ;
  assign y13838 = n51724 ;
  assign y13839 = n51729 ;
  assign y13840 = ~n51730 ;
  assign y13841 = ~n51732 ;
  assign y13842 = ~n51735 ;
  assign y13843 = n51738 ;
  assign y13844 = ~n51740 ;
  assign y13845 = ~n51746 ;
  assign y13846 = ~n51747 ;
  assign y13847 = n51751 ;
  assign y13848 = ~n51752 ;
  assign y13849 = n51756 ;
  assign y13850 = n51757 ;
  assign y13851 = ~n51764 ;
  assign y13852 = ~n51768 ;
  assign y13853 = ~1'b0 ;
  assign y13854 = ~n51769 ;
  assign y13855 = n51772 ;
  assign y13856 = ~n51776 ;
  assign y13857 = ~n51777 ;
  assign y13858 = ~n51780 ;
  assign y13859 = ~n51781 ;
  assign y13860 = n51783 ;
  assign y13861 = n51784 ;
  assign y13862 = n51787 ;
  assign y13863 = ~n51789 ;
  assign y13864 = ~n51792 ;
  assign y13865 = n51794 ;
  assign y13866 = ~n51795 ;
  assign y13867 = ~n51796 ;
  assign y13868 = n51798 ;
  assign y13869 = n51801 ;
  assign y13870 = ~n51802 ;
  assign y13871 = ~n51805 ;
  assign y13872 = ~1'b0 ;
  assign y13873 = ~n51810 ;
  assign y13874 = n51813 ;
  assign y13875 = n51815 ;
  assign y13876 = n51816 ;
  assign y13877 = n51819 ;
  assign y13878 = ~n51823 ;
  assign y13879 = n51824 ;
  assign y13880 = ~1'b0 ;
  assign y13881 = ~n51829 ;
  assign y13882 = ~n51830 ;
  assign y13883 = ~n51831 ;
  assign y13884 = ~n51838 ;
  assign y13885 = n51841 ;
  assign y13886 = n51844 ;
  assign y13887 = ~n51845 ;
  assign y13888 = ~n51847 ;
  assign y13889 = ~1'b0 ;
  assign y13890 = n51849 ;
  assign y13891 = n51852 ;
  assign y13892 = ~n51853 ;
  assign y13893 = n51855 ;
  assign y13894 = ~n51856 ;
  assign y13895 = n51857 ;
  assign y13896 = ~n51861 ;
  assign y13897 = n51864 ;
  assign y13898 = n51867 ;
  assign y13899 = ~1'b0 ;
  assign y13900 = ~n51869 ;
  assign y13901 = n51873 ;
  assign y13902 = n51877 ;
  assign y13903 = ~n51884 ;
  assign y13904 = ~n51885 ;
  assign y13905 = n51886 ;
  assign y13906 = ~n51888 ;
  assign y13907 = ~1'b0 ;
  assign y13908 = ~n51889 ;
  assign y13909 = n51896 ;
  assign y13910 = ~n51897 ;
  assign y13911 = ~n51900 ;
  assign y13912 = n51903 ;
  assign y13913 = n51905 ;
  assign y13914 = ~n51907 ;
  assign y13915 = ~n51908 ;
  assign y13916 = n51915 ;
  assign y13917 = ~1'b0 ;
  assign y13918 = ~n51917 ;
  assign y13919 = n51918 ;
  assign y13920 = n51922 ;
  assign y13921 = ~n51924 ;
  assign y13922 = ~n51931 ;
  assign y13923 = ~n51941 ;
  assign y13924 = ~n51942 ;
  assign y13925 = n51946 ;
  assign y13926 = n51947 ;
  assign y13927 = ~1'b0 ;
  assign y13928 = n51951 ;
  assign y13929 = ~n51952 ;
  assign y13930 = n51956 ;
  assign y13931 = ~n51957 ;
  assign y13932 = ~n51960 ;
  assign y13933 = ~n51961 ;
  assign y13934 = ~n51962 ;
  assign y13935 = ~n51967 ;
  assign y13936 = ~n51972 ;
  assign y13937 = ~n51973 ;
  assign y13938 = ~1'b0 ;
  assign y13939 = ~n51978 ;
  assign y13940 = ~n51979 ;
  assign y13941 = n51982 ;
  assign y13942 = n51984 ;
  assign y13943 = n51986 ;
  assign y13944 = n51987 ;
  assign y13945 = n51993 ;
  assign y13946 = n51995 ;
  assign y13947 = ~n51996 ;
  assign y13948 = ~1'b0 ;
  assign y13949 = ~n51997 ;
  assign y13950 = n51999 ;
  assign y13951 = ~n52000 ;
  assign y13952 = ~n52001 ;
  assign y13953 = n52009 ;
  assign y13954 = n52010 ;
  assign y13955 = n52013 ;
  assign y13956 = ~n52014 ;
  assign y13957 = ~1'b0 ;
  assign y13958 = ~n52016 ;
  assign y13959 = ~n52019 ;
  assign y13960 = n52020 ;
  assign y13961 = ~n52022 ;
  assign y13962 = n52027 ;
  assign y13963 = ~n52028 ;
  assign y13964 = n52032 ;
  assign y13965 = ~n52034 ;
  assign y13966 = ~n52039 ;
  assign y13967 = ~1'b0 ;
  assign y13968 = n52041 ;
  assign y13969 = ~n52042 ;
  assign y13970 = n52046 ;
  assign y13971 = n52047 ;
  assign y13972 = ~n52048 ;
  assign y13973 = n52049 ;
  assign y13974 = ~n52052 ;
  assign y13975 = ~n52058 ;
  assign y13976 = ~n52061 ;
  assign y13977 = ~n52063 ;
  assign y13978 = ~n52070 ;
  assign y13979 = n52072 ;
  assign y13980 = n52073 ;
  assign y13981 = n52074 ;
  assign y13982 = n52079 ;
  assign y13983 = n52083 ;
  assign y13984 = ~n52085 ;
  assign y13985 = n52087 ;
  assign y13986 = n52088 ;
  assign y13987 = ~n52090 ;
  assign y13988 = ~n52092 ;
  assign y13989 = ~n52093 ;
  assign y13990 = n52096 ;
  assign y13991 = n52099 ;
  assign y13992 = ~n52100 ;
  assign y13993 = n52101 ;
  assign y13994 = ~n52102 ;
  assign y13995 = n52105 ;
  assign y13996 = ~n52110 ;
  assign y13997 = ~n52111 ;
  assign y13998 = ~1'b0 ;
  assign y13999 = ~1'b0 ;
  assign y14000 = ~n52114 ;
  assign y14001 = ~n52115 ;
  assign y14002 = ~n52117 ;
  assign y14003 = n52118 ;
  assign y14004 = ~n52120 ;
  assign y14005 = n52121 ;
  assign y14006 = ~n52127 ;
  assign y14007 = n52128 ;
  assign y14008 = n52129 ;
  assign y14009 = n52131 ;
  assign y14010 = n52133 ;
  assign y14011 = n52134 ;
  assign y14012 = ~n52135 ;
  assign y14013 = n52137 ;
  assign y14014 = n52143 ;
  assign y14015 = ~n52144 ;
  assign y14016 = ~n52145 ;
  assign y14017 = n52146 ;
  assign y14018 = ~n52149 ;
  assign y14019 = ~1'b0 ;
  assign y14020 = n52151 ;
  assign y14021 = n52153 ;
  assign y14022 = n52154 ;
  assign y14023 = ~n52155 ;
  assign y14024 = n52156 ;
  assign y14025 = n52159 ;
  assign y14026 = n52161 ;
  assign y14027 = n52162 ;
  assign y14028 = n52163 ;
  assign y14029 = n52166 ;
  assign y14030 = ~n52171 ;
  assign y14031 = ~n52172 ;
  assign y14032 = n52173 ;
  assign y14033 = ~n52179 ;
  assign y14034 = n52182 ;
  assign y14035 = ~n52185 ;
  assign y14036 = ~n52186 ;
  assign y14037 = n52188 ;
  assign y14038 = n52189 ;
  assign y14039 = ~n52192 ;
  assign y14040 = ~n52198 ;
  assign y14041 = ~1'b0 ;
  assign y14042 = n52199 ;
  assign y14043 = ~n52201 ;
  assign y14044 = ~n52203 ;
  assign y14045 = ~n52207 ;
  assign y14046 = n52213 ;
  assign y14047 = n52215 ;
  assign y14048 = n52217 ;
  assign y14049 = ~1'b0 ;
  assign y14050 = ~n52224 ;
  assign y14051 = ~n52226 ;
  assign y14052 = n52228 ;
  assign y14053 = ~n52229 ;
  assign y14054 = n52230 ;
  assign y14055 = ~n52231 ;
  assign y14056 = n52232 ;
  assign y14057 = ~n52236 ;
  assign y14058 = n52237 ;
  assign y14059 = n52241 ;
  assign y14060 = ~n52243 ;
  assign y14061 = ~1'b0 ;
  assign y14062 = ~n52250 ;
  assign y14063 = ~n52254 ;
  assign y14064 = ~n52255 ;
  assign y14065 = ~n52258 ;
  assign y14066 = n52260 ;
  assign y14067 = ~n52268 ;
  assign y14068 = ~n52272 ;
  assign y14069 = ~n52274 ;
  assign y14070 = ~n52276 ;
  assign y14071 = ~1'b0 ;
  assign y14072 = ~n52278 ;
  assign y14073 = n52279 ;
  assign y14074 = n52281 ;
  assign y14075 = n52284 ;
  assign y14076 = ~n52288 ;
  assign y14077 = n52289 ;
  assign y14078 = ~n52290 ;
  assign y14079 = n52292 ;
  assign y14080 = ~n52298 ;
  assign y14081 = ~n52304 ;
  assign y14082 = ~n52306 ;
  assign y14083 = n52307 ;
  assign y14084 = ~n52312 ;
  assign y14085 = n52315 ;
  assign y14086 = n52316 ;
  assign y14087 = ~n52317 ;
  assign y14088 = ~n52319 ;
  assign y14089 = n52320 ;
  assign y14090 = n52327 ;
  assign y14091 = ~n52329 ;
  assign y14092 = n52331 ;
  assign y14093 = n52332 ;
  assign y14094 = ~n52334 ;
  assign y14095 = n52337 ;
  assign y14096 = n52340 ;
  assign y14097 = ~n52342 ;
  assign y14098 = n52343 ;
  assign y14099 = ~n52344 ;
  assign y14100 = ~n52345 ;
  assign y14101 = ~n52347 ;
  assign y14102 = ~n52348 ;
  assign y14103 = ~n52350 ;
  assign y14104 = ~n52356 ;
  assign y14105 = ~n52358 ;
  assign y14106 = n52365 ;
  assign y14107 = n52367 ;
  assign y14108 = n52369 ;
  assign y14109 = ~n52372 ;
  assign y14110 = n52376 ;
  assign y14111 = n52379 ;
  assign y14112 = n52380 ;
  assign y14113 = ~n52387 ;
  assign y14114 = n52392 ;
  assign y14115 = ~n52394 ;
  assign y14116 = ~n52400 ;
  assign y14117 = ~1'b0 ;
  assign y14118 = n52402 ;
  assign y14119 = n52403 ;
  assign y14120 = ~n52405 ;
  assign y14121 = n52408 ;
  assign y14122 = n52411 ;
  assign y14123 = n52419 ;
  assign y14124 = ~n52422 ;
  assign y14125 = n52426 ;
  assign y14126 = ~1'b0 ;
  assign y14127 = n52431 ;
  assign y14128 = n52433 ;
  assign y14129 = ~n52434 ;
  assign y14130 = ~n52436 ;
  assign y14131 = ~n52438 ;
  assign y14132 = ~n52444 ;
  assign y14133 = ~n52450 ;
  assign y14134 = n52457 ;
  assign y14135 = ~n52459 ;
  assign y14136 = ~n52463 ;
  assign y14137 = n52466 ;
  assign y14138 = n52467 ;
  assign y14139 = ~n52471 ;
  assign y14140 = n52473 ;
  assign y14141 = ~n52474 ;
  assign y14142 = ~n52476 ;
  assign y14143 = n52477 ;
  assign y14144 = n52480 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = ~n52484 ;
  assign y14147 = ~n52485 ;
  assign y14148 = ~n52489 ;
  assign y14149 = n52490 ;
  assign y14150 = n52491 ;
  assign y14151 = n52494 ;
  assign y14152 = ~n52496 ;
  assign y14153 = ~n52501 ;
  assign y14154 = ~n52502 ;
  assign y14155 = n52507 ;
  assign y14156 = ~n52511 ;
  assign y14157 = ~n52514 ;
  assign y14158 = ~n52515 ;
  assign y14159 = n52517 ;
  assign y14160 = ~n52519 ;
  assign y14161 = n52522 ;
  assign y14162 = ~n52525 ;
  assign y14163 = ~n52526 ;
  assign y14164 = ~n52528 ;
  assign y14165 = ~n52529 ;
  assign y14166 = n52531 ;
  assign y14167 = ~1'b0 ;
  assign y14168 = ~n52535 ;
  assign y14169 = ~n52537 ;
  assign y14170 = n52538 ;
  assign y14171 = ~n52540 ;
  assign y14172 = ~n52541 ;
  assign y14173 = n52542 ;
  assign y14174 = ~n52543 ;
  assign y14175 = n52549 ;
  assign y14176 = n52551 ;
  assign y14177 = ~1'b0 ;
  assign y14178 = ~n52554 ;
  assign y14179 = ~n52556 ;
  assign y14180 = n52561 ;
  assign y14181 = ~n52564 ;
  assign y14182 = n52565 ;
  assign y14183 = ~n52566 ;
  assign y14184 = ~n52569 ;
  assign y14185 = n52571 ;
  assign y14186 = ~1'b0 ;
  assign y14187 = ~1'b0 ;
  assign y14188 = n17040 ;
  assign y14189 = ~n52576 ;
  assign y14190 = ~n52579 ;
  assign y14191 = ~n52583 ;
  assign y14192 = ~n52585 ;
  assign y14193 = n52587 ;
  assign y14194 = ~n52588 ;
  assign y14195 = n52591 ;
  assign y14196 = ~n52602 ;
  assign y14197 = ~n52605 ;
  assign y14198 = n52607 ;
  assign y14199 = ~n52608 ;
  assign y14200 = ~n52612 ;
  assign y14201 = n52613 ;
  assign y14202 = n52617 ;
  assign y14203 = ~n52618 ;
  assign y14204 = n52623 ;
  assign y14205 = ~1'b0 ;
  assign y14206 = n52627 ;
  assign y14207 = ~n52629 ;
  assign y14208 = n52631 ;
  assign y14209 = ~n52632 ;
  assign y14210 = ~n52635 ;
  assign y14211 = ~n52638 ;
  assign y14212 = ~n52642 ;
  assign y14213 = n52643 ;
  assign y14214 = n52645 ;
  assign y14215 = n52648 ;
  assign y14216 = ~n52652 ;
  assign y14217 = ~1'b0 ;
  assign y14218 = n52656 ;
  assign y14219 = ~n52660 ;
  assign y14220 = n52663 ;
  assign y14221 = n52666 ;
  assign y14222 = ~n52668 ;
  assign y14223 = ~n52670 ;
  assign y14224 = n52672 ;
  assign y14225 = ~n52674 ;
  assign y14226 = ~n52676 ;
  assign y14227 = ~n52678 ;
  assign y14228 = n52680 ;
  assign y14229 = n52681 ;
  assign y14230 = ~n52682 ;
  assign y14231 = n52684 ;
  assign y14232 = ~n52685 ;
  assign y14233 = ~n52690 ;
  assign y14234 = ~n52692 ;
  assign y14235 = ~n52695 ;
  assign y14236 = ~n52697 ;
  assign y14237 = n52703 ;
  assign y14238 = ~n52708 ;
  assign y14239 = ~n52709 ;
  assign y14240 = ~n52715 ;
  assign y14241 = n52716 ;
  assign y14242 = n52717 ;
  assign y14243 = ~n52718 ;
  assign y14244 = ~n52720 ;
  assign y14245 = n52721 ;
  assign y14246 = n52722 ;
  assign y14247 = ~n52725 ;
  assign y14248 = n52726 ;
  assign y14249 = n52729 ;
  assign y14250 = n52730 ;
  assign y14251 = ~n52731 ;
  assign y14252 = ~n52738 ;
  assign y14253 = ~n52739 ;
  assign y14254 = n52740 ;
  assign y14255 = ~n52741 ;
  assign y14256 = n52742 ;
  assign y14257 = ~n52748 ;
  assign y14258 = ~1'b0 ;
  assign y14259 = n52752 ;
  assign y14260 = n52753 ;
  assign y14261 = n52757 ;
  assign y14262 = n52758 ;
  assign y14263 = ~n52759 ;
  assign y14264 = n52760 ;
  assign y14265 = ~n52761 ;
  assign y14266 = n52762 ;
  assign y14267 = ~n52763 ;
  assign y14268 = n52767 ;
  assign y14269 = ~n52772 ;
  assign y14270 = ~n52774 ;
  assign y14271 = n52776 ;
  assign y14272 = n52783 ;
  assign y14273 = ~n52784 ;
  assign y14274 = n52785 ;
  assign y14275 = n52789 ;
  assign y14276 = ~n52790 ;
  assign y14277 = n52792 ;
  assign y14278 = n52793 ;
  assign y14279 = n52795 ;
  assign y14280 = n52797 ;
  assign y14281 = n52800 ;
  assign y14282 = ~n52803 ;
  assign y14283 = ~n52804 ;
  assign y14284 = ~n52807 ;
  assign y14285 = n52812 ;
  assign y14286 = ~n52813 ;
  assign y14287 = n52814 ;
  assign y14288 = n52815 ;
  assign y14289 = n52818 ;
  assign y14290 = n52820 ;
  assign y14291 = ~n52822 ;
  assign y14292 = n52827 ;
  assign y14293 = n52828 ;
  assign y14294 = ~n52830 ;
  assign y14295 = ~n52834 ;
  assign y14296 = ~n52835 ;
  assign y14297 = n52838 ;
  assign y14298 = n52844 ;
  assign y14299 = n52850 ;
  assign y14300 = ~n52852 ;
  assign y14301 = ~n52854 ;
  assign y14302 = ~n52856 ;
  assign y14303 = ~n52858 ;
  assign y14304 = ~n52860 ;
  assign y14305 = n52862 ;
  assign y14306 = n52863 ;
  assign y14307 = n52864 ;
  assign y14308 = n52865 ;
  assign y14309 = n52868 ;
  assign y14310 = n52870 ;
  assign y14311 = n52871 ;
  assign y14312 = n52875 ;
  assign y14313 = n52879 ;
  assign y14314 = ~n52882 ;
  assign y14315 = n52884 ;
  assign y14316 = ~n52886 ;
  assign y14317 = n52893 ;
  assign y14318 = n52896 ;
  assign y14319 = ~n52897 ;
  assign y14320 = n52899 ;
  assign y14321 = n52900 ;
  assign y14322 = ~n52902 ;
  assign y14323 = ~n52904 ;
  assign y14324 = n52907 ;
  assign y14325 = ~n52915 ;
  assign y14326 = ~n52917 ;
  assign y14327 = n52919 ;
  assign y14328 = ~n52920 ;
  assign y14329 = n52923 ;
  assign y14330 = n52926 ;
  assign y14331 = n52929 ;
  assign y14332 = ~n52932 ;
  assign y14333 = n52933 ;
  assign y14334 = ~1'b0 ;
  assign y14335 = ~1'b0 ;
  assign y14336 = ~n52935 ;
  assign y14337 = n52938 ;
  assign y14338 = ~n52941 ;
  assign y14339 = ~n52943 ;
  assign y14340 = ~n52944 ;
  assign y14341 = ~n52948 ;
  assign y14342 = ~n52950 ;
  assign y14343 = n52951 ;
  assign y14344 = ~n52952 ;
  assign y14345 = n52954 ;
  assign y14346 = n52955 ;
  assign y14347 = n52957 ;
  assign y14348 = ~n52960 ;
  assign y14349 = n52961 ;
  assign y14350 = n52963 ;
  assign y14351 = n52964 ;
  assign y14352 = n52966 ;
  assign y14353 = ~n52967 ;
  assign y14354 = n52971 ;
  assign y14355 = n52973 ;
  assign y14356 = n52976 ;
  assign y14357 = n52977 ;
  assign y14358 = n52979 ;
  assign y14359 = ~n52981 ;
  assign y14360 = ~n52982 ;
  assign y14361 = ~n52983 ;
  assign y14362 = ~n52985 ;
  assign y14363 = ~n52992 ;
  assign y14364 = n52993 ;
  assign y14365 = n52994 ;
  assign y14366 = ~n52996 ;
  assign y14367 = ~n53001 ;
  assign y14368 = n53003 ;
  assign y14369 = ~n53004 ;
  assign y14370 = n53006 ;
  assign y14371 = n53007 ;
  assign y14372 = n53008 ;
  assign y14373 = n53009 ;
  assign y14374 = n53010 ;
  assign y14375 = ~n53011 ;
  assign y14376 = n53013 ;
  assign y14377 = ~n53016 ;
  assign y14378 = n53017 ;
  assign y14379 = ~n53019 ;
  assign y14380 = ~n53023 ;
  assign y14381 = ~n53025 ;
  assign y14382 = ~n53028 ;
  assign y14383 = ~n53031 ;
  assign y14384 = ~n53033 ;
  assign y14385 = ~n53035 ;
  assign y14386 = n53038 ;
  assign y14387 = ~1'b0 ;
  assign y14388 = ~1'b0 ;
  assign y14389 = n53040 ;
  assign y14390 = ~n53043 ;
  assign y14391 = n53051 ;
  assign y14392 = n53052 ;
  assign y14393 = n53057 ;
  assign y14394 = ~n53058 ;
  assign y14395 = ~n53061 ;
  assign y14396 = n53063 ;
  assign y14397 = ~1'b0 ;
  assign y14398 = ~n53065 ;
  assign y14399 = n53066 ;
  assign y14400 = n53068 ;
  assign y14401 = n53070 ;
  assign y14402 = n53072 ;
  assign y14403 = n53074 ;
  assign y14404 = ~n53078 ;
  assign y14405 = ~n53081 ;
  assign y14406 = n53087 ;
  assign y14407 = ~1'b0 ;
  assign y14408 = ~n53088 ;
  assign y14409 = ~n53091 ;
  assign y14410 = ~n53092 ;
  assign y14411 = n53094 ;
  assign y14412 = ~n53097 ;
  assign y14413 = n53098 ;
  assign y14414 = ~n53100 ;
  assign y14415 = ~n53104 ;
  assign y14416 = n53107 ;
  assign y14417 = n53109 ;
  assign y14418 = n53110 ;
  assign y14419 = n53116 ;
  assign y14420 = ~n53120 ;
  assign y14421 = n53122 ;
  assign y14422 = ~n53127 ;
  assign y14423 = ~n53131 ;
  assign y14424 = ~n53132 ;
  assign y14425 = ~n53136 ;
  assign y14426 = n53139 ;
  assign y14427 = n53141 ;
  assign y14428 = ~n53143 ;
  assign y14429 = n53144 ;
  assign y14430 = ~n53146 ;
  assign y14431 = ~n53150 ;
  assign y14432 = ~n53156 ;
  assign y14433 = n53158 ;
  assign y14434 = ~n53159 ;
  assign y14435 = n53161 ;
  assign y14436 = ~n53163 ;
  assign y14437 = n53165 ;
  assign y14438 = ~n53167 ;
  assign y14439 = ~n53171 ;
  assign y14440 = n53173 ;
  assign y14441 = ~n53178 ;
  assign y14442 = ~n53183 ;
  assign y14443 = n53186 ;
  assign y14444 = ~n53191 ;
  assign y14445 = n53193 ;
  assign y14446 = n53196 ;
  assign y14447 = ~n53204 ;
  assign y14448 = ~n53206 ;
  assign y14449 = n53207 ;
  assign y14450 = n53210 ;
  assign y14451 = ~n53213 ;
  assign y14452 = ~n53217 ;
  assign y14453 = ~n53218 ;
  assign y14454 = ~n53219 ;
  assign y14455 = n53220 ;
  assign y14456 = ~n53221 ;
  assign y14457 = ~1'b0 ;
  assign y14458 = ~n53226 ;
  assign y14459 = ~n53227 ;
  assign y14460 = ~n53230 ;
  assign y14461 = n53232 ;
  assign y14462 = ~n53241 ;
  assign y14463 = n53242 ;
  assign y14464 = ~n53243 ;
  assign y14465 = n53247 ;
  assign y14466 = n53253 ;
  assign y14467 = ~n53255 ;
  assign y14468 = ~1'b0 ;
  assign y14469 = n53258 ;
  assign y14470 = n53261 ;
  assign y14471 = n53264 ;
  assign y14472 = ~n53268 ;
  assign y14473 = ~n53270 ;
  assign y14474 = ~n53271 ;
  assign y14475 = n53276 ;
  assign y14476 = ~n53277 ;
  assign y14477 = ~n53279 ;
  assign y14478 = ~1'b0 ;
  assign y14479 = n53282 ;
  assign y14480 = ~n53283 ;
  assign y14481 = ~n53286 ;
  assign y14482 = ~n53290 ;
  assign y14483 = ~n53292 ;
  assign y14484 = n53296 ;
  assign y14485 = ~n53297 ;
  assign y14486 = n53299 ;
  assign y14487 = ~n53303 ;
  assign y14488 = ~n53305 ;
  assign y14489 = ~n53308 ;
  assign y14490 = n53309 ;
  assign y14491 = ~n53314 ;
  assign y14492 = ~n53317 ;
  assign y14493 = n53320 ;
  assign y14494 = ~n53321 ;
  assign y14495 = ~n53322 ;
  assign y14496 = ~n53324 ;
  assign y14497 = n53327 ;
  assign y14498 = ~n53330 ;
  assign y14499 = ~n53332 ;
  assign y14500 = n53334 ;
  assign y14501 = ~n53335 ;
  assign y14502 = n53336 ;
  assign y14503 = n53347 ;
  assign y14504 = ~n53348 ;
  assign y14505 = n53349 ;
  assign y14506 = ~n53351 ;
  assign y14507 = ~1'b0 ;
  assign y14508 = ~n53354 ;
  assign y14509 = n53356 ;
  assign y14510 = n53357 ;
  assign y14511 = n53358 ;
  assign y14512 = ~n53359 ;
  assign y14513 = ~n53361 ;
  assign y14514 = n53365 ;
  assign y14515 = ~n53367 ;
  assign y14516 = n53368 ;
  assign y14517 = ~n53371 ;
  assign y14518 = ~1'b0 ;
  assign y14519 = n53375 ;
  assign y14520 = n53377 ;
  assign y14521 = ~n53378 ;
  assign y14522 = n53379 ;
  assign y14523 = ~n53380 ;
  assign y14524 = ~n53381 ;
  assign y14525 = n53385 ;
  assign y14526 = ~n53386 ;
  assign y14527 = ~n53388 ;
  assign y14528 = ~1'b0 ;
  assign y14529 = n53389 ;
  assign y14530 = n53390 ;
  assign y14531 = ~n53391 ;
  assign y14532 = ~n53392 ;
  assign y14533 = ~n53395 ;
  assign y14534 = ~n53398 ;
  assign y14535 = n53400 ;
  assign y14536 = ~n53401 ;
  assign y14537 = ~n53404 ;
  assign y14538 = ~n53405 ;
  assign y14539 = ~n53409 ;
  assign y14540 = ~n53413 ;
  assign y14541 = n53414 ;
  assign y14542 = n53416 ;
  assign y14543 = ~n53420 ;
  assign y14544 = ~n53422 ;
  assign y14545 = ~n53423 ;
  assign y14546 = n53428 ;
  assign y14547 = ~n53436 ;
  assign y14548 = n53437 ;
  assign y14549 = n53440 ;
  assign y14550 = n53441 ;
  assign y14551 = ~n53443 ;
  assign y14552 = n53444 ;
  assign y14553 = ~n53446 ;
  assign y14554 = ~n53448 ;
  assign y14555 = n53449 ;
  assign y14556 = n53450 ;
  assign y14557 = n53454 ;
  assign y14558 = ~n53455 ;
  assign y14559 = n53458 ;
  assign y14560 = ~1'b0 ;
  assign y14561 = ~n53459 ;
  assign y14562 = ~n53464 ;
  assign y14563 = n53465 ;
  assign y14564 = ~n53468 ;
  assign y14565 = ~n53470 ;
  assign y14566 = n53472 ;
  assign y14567 = ~n53473 ;
  assign y14568 = n53474 ;
  assign y14569 = n53476 ;
  assign y14570 = ~1'b0 ;
  assign y14571 = n53480 ;
  assign y14572 = n53481 ;
  assign y14573 = ~n53482 ;
  assign y14574 = n53486 ;
  assign y14575 = ~n53488 ;
  assign y14576 = n53489 ;
  assign y14577 = n53492 ;
  assign y14578 = n53494 ;
  assign y14579 = ~n53495 ;
  assign y14580 = n53498 ;
  assign y14581 = ~n53500 ;
  assign y14582 = ~n53501 ;
  assign y14583 = ~n53502 ;
  assign y14584 = n53505 ;
  assign y14585 = n53506 ;
  assign y14586 = n53507 ;
  assign y14587 = ~n53510 ;
  assign y14588 = ~n53516 ;
  assign y14589 = ~n53519 ;
  assign y14590 = ~n53521 ;
  assign y14591 = ~n53525 ;
  assign y14592 = ~n53526 ;
  assign y14593 = n53527 ;
  assign y14594 = ~n53528 ;
  assign y14595 = ~n53530 ;
  assign y14596 = n53531 ;
  assign y14597 = ~n53532 ;
  assign y14598 = n53533 ;
  assign y14599 = ~n53534 ;
  assign y14600 = n53536 ;
  assign y14601 = n53539 ;
  assign y14602 = ~n53543 ;
  assign y14603 = n53544 ;
  assign y14604 = n53546 ;
  assign y14605 = ~n53547 ;
  assign y14606 = ~n53548 ;
  assign y14607 = n53549 ;
  assign y14608 = ~n53550 ;
  assign y14609 = n53551 ;
  assign y14610 = n53553 ;
  assign y14611 = ~1'b0 ;
  assign y14612 = n53556 ;
  assign y14613 = n53559 ;
  assign y14614 = ~n53566 ;
  assign y14615 = n53575 ;
  assign y14616 = ~n53577 ;
  assign y14617 = n53585 ;
  assign y14618 = n53587 ;
  assign y14619 = ~n53590 ;
  assign y14620 = ~n53601 ;
  assign y14621 = ~n53603 ;
  assign y14622 = n53604 ;
  assign y14623 = ~n53607 ;
  assign y14624 = n53608 ;
  assign y14625 = ~n53610 ;
  assign y14626 = n53614 ;
  assign y14627 = ~n53618 ;
  assign y14628 = ~n53625 ;
  assign y14629 = ~n53628 ;
  assign y14630 = n53629 ;
  assign y14631 = ~n53631 ;
  assign y14632 = ~1'b0 ;
  assign y14633 = n53634 ;
  assign y14634 = n53635 ;
  assign y14635 = n53637 ;
  assign y14636 = ~n53646 ;
  assign y14637 = n53647 ;
  assign y14638 = ~n53649 ;
  assign y14639 = n53653 ;
  assign y14640 = n53654 ;
  assign y14641 = ~n53655 ;
  assign y14642 = n53657 ;
  assign y14643 = ~1'b0 ;
  assign y14644 = n53658 ;
  assign y14645 = n53660 ;
  assign y14646 = n53663 ;
  assign y14647 = n53664 ;
  assign y14648 = ~n53666 ;
  assign y14649 = n53669 ;
  assign y14650 = n53670 ;
  assign y14651 = n53671 ;
  assign y14652 = ~n53672 ;
  assign y14653 = ~n53675 ;
  assign y14654 = ~n53680 ;
  assign y14655 = n53685 ;
  assign y14656 = ~n53692 ;
  assign y14657 = ~n53693 ;
  assign y14658 = n53694 ;
  assign y14659 = ~n53698 ;
  assign y14660 = n53699 ;
  assign y14661 = ~n53700 ;
  assign y14662 = ~n53701 ;
  assign y14663 = ~n53706 ;
  assign y14664 = n53708 ;
  assign y14665 = ~n53713 ;
  assign y14666 = n53715 ;
  assign y14667 = n53719 ;
  assign y14668 = ~n53725 ;
  assign y14669 = ~n53727 ;
  assign y14670 = n53728 ;
  assign y14671 = n53732 ;
  assign y14672 = n53735 ;
  assign y14673 = ~n53736 ;
  assign y14674 = ~n53739 ;
  assign y14675 = ~1'b0 ;
  assign y14676 = ~n53748 ;
  assign y14677 = ~n53749 ;
  assign y14678 = n53750 ;
  assign y14679 = ~n53752 ;
  assign y14680 = n53754 ;
  assign y14681 = n53755 ;
  assign y14682 = n53758 ;
  assign y14683 = n53766 ;
  assign y14684 = n53769 ;
  assign y14685 = n53770 ;
  assign y14686 = ~1'b0 ;
  assign y14687 = n53772 ;
  assign y14688 = n53773 ;
  assign y14689 = n53776 ;
  assign y14690 = n53777 ;
  assign y14691 = ~n53778 ;
  assign y14692 = ~n53779 ;
  assign y14693 = ~n53781 ;
  assign y14694 = n53784 ;
  assign y14695 = ~1'b0 ;
  assign y14696 = n53786 ;
  assign y14697 = ~n53791 ;
  assign y14698 = ~n53792 ;
  assign y14699 = ~n53795 ;
  assign y14700 = ~n53797 ;
  assign y14701 = ~n53799 ;
  assign y14702 = ~n53807 ;
  assign y14703 = ~n53810 ;
  assign y14704 = ~n53811 ;
  assign y14705 = ~n53812 ;
  assign y14706 = n53813 ;
  assign y14707 = ~n53815 ;
  assign y14708 = ~n53819 ;
  assign y14709 = n53822 ;
  assign y14710 = ~n53825 ;
  assign y14711 = n53826 ;
  assign y14712 = n53828 ;
  assign y14713 = ~n53830 ;
  assign y14714 = n53831 ;
  assign y14715 = ~n53834 ;
  assign y14716 = ~1'b0 ;
  assign y14717 = n53837 ;
  assign y14718 = ~n53838 ;
  assign y14719 = n53842 ;
  assign y14720 = ~n53851 ;
  assign y14721 = ~n53854 ;
  assign y14722 = n53858 ;
  assign y14723 = ~n53859 ;
  assign y14724 = ~n53860 ;
  assign y14725 = n53861 ;
  assign y14726 = n53862 ;
  assign y14727 = ~n53864 ;
  assign y14728 = ~n53868 ;
  assign y14729 = n53878 ;
  assign y14730 = ~n53879 ;
  assign y14731 = n53882 ;
  assign y14732 = ~n53890 ;
  assign y14733 = ~n53891 ;
  assign y14734 = n53894 ;
  assign y14735 = ~n53896 ;
  assign y14736 = n53898 ;
  assign y14737 = n53902 ;
  assign y14738 = ~1'b0 ;
  assign y14739 = ~n53903 ;
  assign y14740 = ~n53909 ;
  assign y14741 = n53911 ;
  assign y14742 = n53912 ;
  assign y14743 = ~n53914 ;
  assign y14744 = ~n53916 ;
  assign y14745 = n53919 ;
  assign y14746 = n53920 ;
  assign y14747 = n53922 ;
  assign y14748 = ~n53924 ;
  assign y14749 = ~1'b0 ;
  assign y14750 = ~n53926 ;
  assign y14751 = n53930 ;
  assign y14752 = ~n53932 ;
  assign y14753 = ~n53934 ;
  assign y14754 = ~n53937 ;
  assign y14755 = ~n53938 ;
  assign y14756 = ~n53941 ;
  assign y14757 = ~n53944 ;
  assign y14758 = ~1'b0 ;
  assign y14759 = n53946 ;
  assign y14760 = ~n53947 ;
  assign y14761 = ~n53950 ;
  assign y14762 = n53952 ;
  assign y14763 = ~n53953 ;
  assign y14764 = n53958 ;
  assign y14765 = ~n53959 ;
  assign y14766 = n53961 ;
  assign y14767 = n53962 ;
  assign y14768 = n53964 ;
  assign y14769 = n53966 ;
  assign y14770 = ~n53968 ;
  assign y14771 = ~n53970 ;
  assign y14772 = n53974 ;
  assign y14773 = n53977 ;
  assign y14774 = n53978 ;
  assign y14775 = n53980 ;
  assign y14776 = ~n53981 ;
  assign y14777 = n53984 ;
  assign y14778 = n53986 ;
  assign y14779 = n53989 ;
  assign y14780 = n53992 ;
  assign y14781 = ~n53993 ;
  assign y14782 = ~n53996 ;
  assign y14783 = ~n54000 ;
  assign y14784 = ~n54004 ;
  assign y14785 = n54005 ;
  assign y14786 = ~n54011 ;
  assign y14787 = ~n54013 ;
  assign y14788 = n54014 ;
  assign y14789 = n54015 ;
  assign y14790 = ~n54019 ;
  assign y14791 = ~n54021 ;
  assign y14792 = ~n54023 ;
  assign y14793 = ~n54024 ;
  assign y14794 = n54030 ;
  assign y14795 = n54031 ;
  assign y14796 = n54035 ;
  assign y14797 = n54037 ;
  assign y14798 = ~n54040 ;
  assign y14799 = n54041 ;
  assign y14800 = n54042 ;
  assign y14801 = ~n54044 ;
  assign y14802 = n54048 ;
  assign y14803 = ~n54051 ;
  assign y14804 = n54052 ;
  assign y14805 = n11875 ;
  assign y14806 = n18998 ;
  assign y14807 = ~n54053 ;
  assign y14808 = ~n54055 ;
  assign y14809 = n54058 ;
  assign y14810 = n54060 ;
  assign y14811 = ~n54061 ;
  assign y14812 = ~n54063 ;
  assign y14813 = n54066 ;
  assign y14814 = n54067 ;
  assign y14815 = ~n54069 ;
  assign y14816 = ~n54070 ;
  assign y14817 = n54072 ;
  assign y14818 = n54074 ;
  assign y14819 = n54078 ;
  assign y14820 = ~n54080 ;
  assign y14821 = ~1'b0 ;
  assign y14822 = n54084 ;
  assign y14823 = ~n54085 ;
  assign y14824 = ~n54087 ;
  assign y14825 = ~n54090 ;
  assign y14826 = ~n54091 ;
  assign y14827 = ~n54093 ;
  assign y14828 = n54094 ;
  assign y14829 = ~n54096 ;
  assign y14830 = n54097 ;
  assign y14831 = n54101 ;
  assign y14832 = n54104 ;
  assign y14833 = n54105 ;
  assign y14834 = n54106 ;
  assign y14835 = ~n54108 ;
  assign y14836 = n54113 ;
  assign y14837 = ~n54114 ;
  assign y14838 = ~n54115 ;
  assign y14839 = n54116 ;
  assign y14840 = n54117 ;
  assign y14841 = ~n54119 ;
  assign y14842 = ~1'b0 ;
  assign y14843 = ~n54123 ;
  assign y14844 = n54127 ;
  assign y14845 = n54128 ;
  assign y14846 = ~n54129 ;
  assign y14847 = n54130 ;
  assign y14848 = ~n54132 ;
  assign y14849 = n54133 ;
  assign y14850 = n54137 ;
  assign y14851 = n54142 ;
  assign y14852 = ~n54144 ;
  assign y14853 = ~n54146 ;
  assign y14854 = n54147 ;
  assign y14855 = n54151 ;
  assign y14856 = ~n54153 ;
  assign y14857 = n54160 ;
  assign y14858 = ~n54166 ;
  assign y14859 = n54167 ;
  assign y14860 = ~n54168 ;
  assign y14861 = ~n54169 ;
  assign y14862 = n54170 ;
  assign y14863 = ~n54172 ;
  assign y14864 = n54174 ;
  assign y14865 = n54178 ;
  assign y14866 = n54181 ;
  assign y14867 = ~n54184 ;
  assign y14868 = n54185 ;
  assign y14869 = n54187 ;
  assign y14870 = ~n54188 ;
  assign y14871 = ~n54189 ;
  assign y14872 = n54191 ;
  assign y14873 = ~n54192 ;
  assign y14874 = n54194 ;
  assign y14875 = n54198 ;
  assign y14876 = ~n54199 ;
  assign y14877 = ~n54200 ;
  assign y14878 = ~n54203 ;
  assign y14879 = ~n54206 ;
  assign y14880 = ~n54214 ;
  assign y14881 = ~n54218 ;
  assign y14882 = ~n54219 ;
  assign y14883 = ~n54222 ;
  assign y14884 = n54223 ;
  assign y14885 = ~n54227 ;
  assign y14886 = ~1'b0 ;
  assign y14887 = n54229 ;
  assign y14888 = ~n54238 ;
  assign y14889 = ~n54239 ;
  assign y14890 = n54245 ;
  assign y14891 = ~n54250 ;
  assign y14892 = ~n54251 ;
  assign y14893 = ~n54252 ;
  assign y14894 = ~n54253 ;
  assign y14895 = ~n54254 ;
  assign y14896 = n54255 ;
  assign y14897 = ~1'b0 ;
  assign y14898 = n54258 ;
  assign y14899 = ~n54260 ;
  assign y14900 = n54262 ;
  assign y14901 = n54265 ;
  assign y14902 = n54268 ;
  assign y14903 = ~n54269 ;
  assign y14904 = n54271 ;
  assign y14905 = n54273 ;
  assign y14906 = ~n54276 ;
  assign y14907 = ~1'b0 ;
  assign y14908 = ~1'b0 ;
  assign y14909 = n54278 ;
  assign y14910 = ~n54279 ;
  assign y14911 = n54280 ;
  assign y14912 = ~n54281 ;
  assign y14913 = n54282 ;
  assign y14914 = ~n54283 ;
  assign y14915 = n54285 ;
  assign y14916 = ~n54286 ;
  assign y14917 = ~n54288 ;
  assign y14918 = n54290 ;
  assign y14919 = ~n54291 ;
  assign y14920 = n54296 ;
  assign y14921 = ~n54297 ;
  assign y14922 = n54300 ;
  assign y14923 = ~n54302 ;
  assign y14924 = n54305 ;
  assign y14925 = n54306 ;
  assign y14926 = ~n54310 ;
  assign y14927 = ~n54313 ;
  assign y14928 = ~n54314 ;
  assign y14929 = n54316 ;
  assign y14930 = ~1'b0 ;
  assign y14931 = n54317 ;
  assign y14932 = n54318 ;
  assign y14933 = ~n54321 ;
  assign y14934 = ~n54322 ;
  assign y14935 = ~n54323 ;
  assign y14936 = ~n54324 ;
  assign y14937 = n54325 ;
  assign y14938 = ~n54326 ;
  assign y14939 = ~n54328 ;
  assign y14940 = ~1'b0 ;
  assign y14941 = ~1'b0 ;
  assign y14942 = n54331 ;
  assign y14943 = ~n54332 ;
  assign y14944 = ~n54333 ;
  assign y14945 = ~n54335 ;
  assign y14946 = ~n54343 ;
  assign y14947 = ~n54345 ;
  assign y14948 = ~n54348 ;
  assign y14949 = ~n54349 ;
  assign y14950 = ~n54351 ;
  assign y14951 = n54353 ;
  assign y14952 = n54355 ;
  assign y14953 = ~n54365 ;
  assign y14954 = n54366 ;
  assign y14955 = n54367 ;
  assign y14956 = n54368 ;
  assign y14957 = ~n54371 ;
  assign y14958 = n54375 ;
  assign y14959 = n54378 ;
  assign y14960 = n54380 ;
  assign y14961 = n54382 ;
  assign y14962 = ~1'b0 ;
  assign y14963 = ~n54387 ;
  assign y14964 = ~n54388 ;
  assign y14965 = ~n54390 ;
  assign y14966 = ~n54392 ;
  assign y14967 = n54397 ;
  assign y14968 = n54400 ;
  assign y14969 = n54401 ;
  assign y14970 = ~n54402 ;
  assign y14971 = ~n54404 ;
  assign y14972 = ~n54405 ;
  assign y14973 = ~1'b0 ;
  assign y14974 = ~n54407 ;
  assign y14975 = ~n54408 ;
  assign y14976 = ~n54409 ;
  assign y14977 = ~n54410 ;
  assign y14978 = ~n54413 ;
  assign y14979 = ~n54417 ;
  assign y14980 = ~n54418 ;
  assign y14981 = ~n54419 ;
  assign y14982 = n54420 ;
  assign y14983 = n54425 ;
  assign y14984 = n54428 ;
  assign y14985 = ~1'b0 ;
  assign y14986 = n54429 ;
  assign y14987 = n54435 ;
  assign y14988 = n54436 ;
  assign y14989 = ~n54437 ;
  assign y14990 = n54441 ;
  assign y14991 = n54443 ;
  assign y14992 = n54444 ;
  assign y14993 = ~n54446 ;
  assign y14994 = n54447 ;
  assign y14995 = ~n54449 ;
  assign y14996 = ~1'b0 ;
  assign y14997 = n54453 ;
  assign y14998 = n54455 ;
  assign y14999 = n54456 ;
  assign y15000 = ~n54459 ;
  assign y15001 = ~n54460 ;
  assign y15002 = ~n54462 ;
  assign y15003 = n54465 ;
  assign y15004 = n54466 ;
  assign y15005 = n54468 ;
  assign y15006 = ~1'b0 ;
  assign y15007 = ~1'b0 ;
  assign y15008 = n54470 ;
  assign y15009 = ~n54471 ;
  assign y15010 = ~n54472 ;
  assign y15011 = n54473 ;
  assign y15012 = ~n54477 ;
  assign y15013 = n54479 ;
  assign y15014 = n54482 ;
  assign y15015 = n54483 ;
  assign y15016 = n54484 ;
  assign y15017 = n54486 ;
  assign y15018 = ~1'b0 ;
  assign y15019 = ~n54493 ;
  assign y15020 = ~n54494 ;
  assign y15021 = ~n54495 ;
  assign y15022 = ~n54496 ;
  assign y15023 = n54497 ;
  assign y15024 = n54499 ;
  assign y15025 = ~n54500 ;
  assign y15026 = ~n54502 ;
  assign y15027 = n54506 ;
  assign y15028 = ~1'b0 ;
  assign y15029 = n54510 ;
  assign y15030 = ~n54511 ;
  assign y15031 = ~n54512 ;
  assign y15032 = ~n54515 ;
  assign y15033 = n54519 ;
  assign y15034 = ~n54521 ;
  assign y15035 = ~n54523 ;
  assign y15036 = n54525 ;
  assign y15037 = ~n54526 ;
  assign y15038 = ~n54527 ;
  assign y15039 = n54529 ;
  assign y15040 = n54535 ;
  assign y15041 = ~n54537 ;
  assign y15042 = ~n54541 ;
  assign y15043 = ~n54544 ;
  assign y15044 = ~n54549 ;
  assign y15045 = ~n54550 ;
  assign y15046 = ~n54554 ;
  assign y15047 = n54557 ;
  assign y15048 = ~n54558 ;
  assign y15049 = n54559 ;
  assign y15050 = ~n54561 ;
  assign y15051 = ~1'b0 ;
  assign y15052 = n54568 ;
  assign y15053 = ~n54569 ;
  assign y15054 = n54571 ;
  assign y15055 = n54573 ;
  assign y15056 = ~n54574 ;
  assign y15057 = n54575 ;
  assign y15058 = ~n9287 ;
  assign y15059 = ~n54576 ;
  assign y15060 = n54578 ;
  assign y15061 = ~1'b0 ;
  assign y15062 = ~1'b0 ;
  assign y15063 = n54581 ;
  assign y15064 = n54584 ;
  assign y15065 = ~n54585 ;
  assign y15066 = n54587 ;
  assign y15067 = n54588 ;
  assign y15068 = n54595 ;
  assign y15069 = ~n54597 ;
  assign y15070 = n54598 ;
  assign y15071 = ~n54601 ;
  assign y15072 = n54604 ;
  assign y15073 = ~1'b0 ;
  assign y15074 = ~n54605 ;
  assign y15075 = n54609 ;
  assign y15076 = ~n54612 ;
  assign y15077 = ~n54619 ;
  assign y15078 = ~n54623 ;
  assign y15079 = ~n54624 ;
  assign y15080 = ~n54626 ;
  assign y15081 = n54627 ;
  assign y15082 = n54628 ;
  assign y15083 = ~n54632 ;
  assign y15084 = ~n54634 ;
  assign y15085 = ~n54635 ;
  assign y15086 = n54636 ;
  assign y15087 = n54639 ;
  assign y15088 = ~n54640 ;
  assign y15089 = n54641 ;
  assign y15090 = n54642 ;
  assign y15091 = ~n54649 ;
  assign y15092 = n54650 ;
  assign y15093 = ~n54651 ;
  assign y15094 = ~n54652 ;
  assign y15095 = ~n54654 ;
  assign y15096 = ~n54655 ;
  assign y15097 = n54656 ;
  assign y15098 = n54658 ;
  assign y15099 = ~n54660 ;
  assign y15100 = ~n54661 ;
  assign y15101 = ~n54662 ;
  assign y15102 = n54666 ;
  assign y15103 = n54671 ;
  assign y15104 = n54672 ;
  assign y15105 = ~n54677 ;
  assign y15106 = ~n54679 ;
  assign y15107 = ~n54681 ;
  assign y15108 = ~n54685 ;
  assign y15109 = n54690 ;
  assign y15110 = ~n54692 ;
  assign y15111 = n54697 ;
  assign y15112 = n54698 ;
  assign y15113 = ~n54700 ;
  assign y15114 = ~n54705 ;
  assign y15115 = n54708 ;
  assign y15116 = ~n54713 ;
  assign y15117 = ~n54718 ;
  assign y15118 = ~n54719 ;
  assign y15119 = n54720 ;
  assign y15120 = n54724 ;
  assign y15121 = ~n54725 ;
  assign y15122 = ~n54728 ;
  assign y15123 = ~n54729 ;
  assign y15124 = n54735 ;
  assign y15125 = n54736 ;
  assign y15126 = ~n54740 ;
  assign y15127 = ~n54744 ;
  assign y15128 = ~1'b0 ;
  assign y15129 = n54747 ;
  assign y15130 = ~n54751 ;
  assign y15131 = n54753 ;
  assign y15132 = ~n54757 ;
  assign y15133 = n54759 ;
  assign y15134 = ~n54764 ;
  assign y15135 = n54769 ;
  assign y15136 = ~n54780 ;
  assign y15137 = ~n54783 ;
  assign y15138 = ~1'b0 ;
  assign y15139 = ~n54785 ;
  assign y15140 = ~n54788 ;
  assign y15141 = ~n54789 ;
  assign y15142 = n54791 ;
  assign y15143 = n54792 ;
  assign y15144 = ~n54797 ;
  assign y15145 = n54800 ;
  assign y15146 = ~n54804 ;
  assign y15147 = n54805 ;
  assign y15148 = ~n54807 ;
  assign y15149 = ~1'b0 ;
  assign y15150 = ~1'b0 ;
  assign y15151 = n54811 ;
  assign y15152 = n54812 ;
  assign y15153 = n54813 ;
  assign y15154 = n54815 ;
  assign y15155 = ~n54816 ;
  assign y15156 = n54819 ;
  assign y15157 = ~n54820 ;
  assign y15158 = ~n54823 ;
  assign y15159 = n54826 ;
  assign y15160 = n54828 ;
  assign y15161 = n54829 ;
  assign y15162 = ~n54831 ;
  assign y15163 = ~n54832 ;
  assign y15164 = n54837 ;
  assign y15165 = ~n54838 ;
  assign y15166 = ~n54843 ;
  assign y15167 = ~n54845 ;
  assign y15168 = ~n54846 ;
  assign y15169 = n54847 ;
  assign y15170 = n54850 ;
  assign y15171 = ~n54852 ;
  assign y15172 = n54853 ;
  assign y15173 = ~n54855 ;
  assign y15174 = ~n54858 ;
  assign y15175 = n54859 ;
  assign y15176 = n54860 ;
  assign y15177 = ~n54863 ;
  assign y15178 = ~n54865 ;
  assign y15179 = n54866 ;
  assign y15180 = n54867 ;
  assign y15181 = ~n54869 ;
  assign y15182 = n54871 ;
  assign y15183 = n54880 ;
  assign y15184 = ~n54883 ;
  assign y15185 = n54886 ;
  assign y15186 = ~n54889 ;
  assign y15187 = n54890 ;
  assign y15188 = n54891 ;
  assign y15189 = n54896 ;
  assign y15190 = n54900 ;
  assign y15191 = ~1'b0 ;
  assign y15192 = ~n54902 ;
  assign y15193 = ~n54904 ;
  assign y15194 = ~n54910 ;
  assign y15195 = ~n54913 ;
  assign y15196 = n54919 ;
  assign y15197 = n54920 ;
  assign y15198 = n54922 ;
  assign y15199 = n54924 ;
  assign y15200 = n54925 ;
  assign y15201 = ~n54929 ;
  assign y15202 = ~n54931 ;
  assign y15203 = ~n54932 ;
  assign y15204 = ~n54936 ;
  assign y15205 = ~n54938 ;
  assign y15206 = ~n54939 ;
  assign y15207 = ~n54940 ;
  assign y15208 = n54944 ;
  assign y15209 = n54950 ;
  assign y15210 = ~n54951 ;
  assign y15211 = n54953 ;
  assign y15212 = n54955 ;
  assign y15213 = n54961 ;
  assign y15214 = ~n54962 ;
  assign y15215 = n54965 ;
  assign y15216 = ~n54966 ;
  assign y15217 = n54967 ;
  assign y15218 = ~n54971 ;
  assign y15219 = n54972 ;
  assign y15220 = ~n54974 ;
  assign y15221 = ~n54977 ;
  assign y15222 = ~n54979 ;
  assign y15223 = n54980 ;
  assign y15224 = n54982 ;
  assign y15225 = n54984 ;
  assign y15226 = n54991 ;
  assign y15227 = n54993 ;
  assign y15228 = n54994 ;
  assign y15229 = ~n54995 ;
  assign y15230 = n54998 ;
  assign y15231 = ~n55001 ;
  assign y15232 = n55003 ;
  assign y15233 = n55005 ;
  assign y15234 = ~1'b0 ;
  assign y15235 = ~1'b0 ;
  assign y15236 = n55011 ;
  assign y15237 = ~n55014 ;
  assign y15238 = ~n55015 ;
  assign y15239 = n55018 ;
  assign y15240 = ~n55022 ;
  assign y15241 = ~n55026 ;
  assign y15242 = ~n55029 ;
  assign y15243 = n55030 ;
  assign y15244 = n55031 ;
  assign y15245 = ~n55036 ;
  assign y15246 = ~1'b0 ;
  assign y15247 = n55038 ;
  assign y15248 = ~n55039 ;
  assign y15249 = ~n55040 ;
  assign y15250 = ~n55043 ;
  assign y15251 = ~n55044 ;
  assign y15252 = n55047 ;
  assign y15253 = n55052 ;
  assign y15254 = ~n55057 ;
  assign y15255 = ~n55058 ;
  assign y15256 = ~n55060 ;
  assign y15257 = n55063 ;
  assign y15258 = ~n55067 ;
  assign y15259 = n55068 ;
  assign y15260 = n55069 ;
  assign y15261 = ~n55071 ;
  assign y15262 = n55072 ;
  assign y15263 = n55075 ;
  assign y15264 = n55080 ;
  assign y15265 = n55082 ;
  assign y15266 = ~n55090 ;
  assign y15267 = n55092 ;
  assign y15268 = ~1'b0 ;
  assign y15269 = ~n55093 ;
  assign y15270 = n55095 ;
  assign y15271 = ~n55096 ;
  assign y15272 = n55098 ;
  assign y15273 = n55099 ;
  assign y15274 = n55100 ;
  assign y15275 = n55101 ;
  assign y15276 = ~n55102 ;
  assign y15277 = n55104 ;
  assign y15278 = n55106 ;
  assign y15279 = n55113 ;
  assign y15280 = ~n55116 ;
  assign y15281 = ~n55117 ;
  assign y15282 = n55118 ;
  assign y15283 = n55119 ;
  assign y15284 = n55122 ;
  assign y15285 = ~n55124 ;
  assign y15286 = ~n55126 ;
  assign y15287 = n55127 ;
  assign y15288 = ~n55128 ;
  assign y15289 = ~n55130 ;
  assign y15290 = ~1'b0 ;
  assign y15291 = n55133 ;
  assign y15292 = ~n55134 ;
  assign y15293 = ~n55135 ;
  assign y15294 = n55136 ;
  assign y15295 = ~n55146 ;
  assign y15296 = ~n55148 ;
  assign y15297 = ~n55149 ;
  assign y15298 = n55155 ;
  assign y15299 = ~n55157 ;
  assign y15300 = ~1'b0 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = n55158 ;
  assign y15303 = n55159 ;
  assign y15304 = n55160 ;
  assign y15305 = ~n55162 ;
  assign y15306 = ~n55163 ;
  assign y15307 = n55164 ;
  assign y15308 = ~n55169 ;
  assign y15309 = ~n55170 ;
  assign y15310 = n55171 ;
  assign y15311 = n55173 ;
  assign y15312 = ~n55177 ;
  assign y15313 = ~n55178 ;
  assign y15314 = ~n55182 ;
  assign y15315 = ~n55183 ;
  assign y15316 = n55185 ;
  assign y15317 = n55190 ;
  assign y15318 = ~n55191 ;
  assign y15319 = n55192 ;
  assign y15320 = ~n55199 ;
  assign y15321 = ~n55200 ;
  assign y15322 = n55201 ;
  assign y15323 = ~1'b0 ;
  assign y15324 = ~n55202 ;
  assign y15325 = ~n55203 ;
  assign y15326 = n55204 ;
  assign y15327 = n55208 ;
  assign y15328 = n55209 ;
  assign y15329 = ~n55210 ;
  assign y15330 = n55215 ;
  assign y15331 = ~n55216 ;
  assign y15332 = n55217 ;
  assign y15333 = ~1'b0 ;
  assign y15334 = n55219 ;
  assign y15335 = n55220 ;
  assign y15336 = ~n55221 ;
  assign y15337 = ~n55223 ;
  assign y15338 = ~n55225 ;
  assign y15339 = ~n55226 ;
  assign y15340 = n55227 ;
  assign y15341 = ~n55228 ;
  assign y15342 = n55229 ;
  assign y15343 = n55230 ;
  assign y15344 = n55231 ;
  assign y15345 = n55233 ;
  assign y15346 = ~n55236 ;
  assign y15347 = ~n55238 ;
  assign y15348 = ~n55239 ;
  assign y15349 = n55240 ;
  assign y15350 = ~n55243 ;
  assign y15351 = ~n55244 ;
  assign y15352 = n55247 ;
  assign y15353 = ~n55251 ;
  assign y15354 = ~n55254 ;
  assign y15355 = ~1'b0 ;
  assign y15356 = ~n55257 ;
  assign y15357 = n55259 ;
  assign y15358 = n55260 ;
  assign y15359 = ~n55261 ;
  assign y15360 = ~n55263 ;
  assign y15361 = ~n55266 ;
  assign y15362 = n55267 ;
  assign y15363 = n55268 ;
  assign y15364 = n55273 ;
  assign y15365 = n55276 ;
  assign y15366 = ~1'b0 ;
  assign y15367 = ~n55279 ;
  assign y15368 = n55280 ;
  assign y15369 = ~n55282 ;
  assign y15370 = ~n55283 ;
  assign y15371 = n55284 ;
  assign y15372 = ~n55285 ;
  assign y15373 = ~n55286 ;
  assign y15374 = n55288 ;
  assign y15375 = n55289 ;
  assign y15376 = ~n55292 ;
  assign y15377 = n55293 ;
  assign y15378 = ~n55295 ;
  assign y15379 = n55296 ;
  assign y15380 = n55297 ;
  assign y15381 = ~n55307 ;
  assign y15382 = n55312 ;
  assign y15383 = n55316 ;
  assign y15384 = ~n55320 ;
  assign y15385 = n55321 ;
  assign y15386 = ~n55324 ;
  assign y15387 = ~n55326 ;
  assign y15388 = n55330 ;
  assign y15389 = ~1'b0 ;
  assign y15390 = ~n55331 ;
  assign y15391 = ~n55332 ;
  assign y15392 = n55333 ;
  assign y15393 = ~n55334 ;
  assign y15394 = ~1'b0 ;
  assign y15395 = n55338 ;
  assign y15396 = ~n55342 ;
  assign y15397 = n55343 ;
  assign y15398 = ~n55345 ;
  assign y15399 = ~n55348 ;
  assign y15400 = ~1'b0 ;
  assign y15401 = ~n55349 ;
  assign y15402 = ~n55351 ;
  assign y15403 = n55357 ;
  assign y15404 = n55358 ;
  assign y15405 = n55362 ;
  assign y15406 = ~n55363 ;
  assign y15407 = n55365 ;
  assign y15408 = n55368 ;
endmodule
