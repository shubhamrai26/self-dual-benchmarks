module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1362 , n1363 , n1364 ;
  assign n11 = ~x3 & ~x5 ;
  assign n12 = ~x1 & x9 ;
  assign n13 = ~x0 & x9 ;
  assign n14 = x1 & ~n13 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = n11 & n15 ;
  assign n17 = x0 & ~x9 ;
  assign n18 = ~x1 & ~n17 ;
  assign n19 = x1 & ~x9 ;
  assign n20 = ~x7 & ~n19 ;
  assign n21 = ~n18 & n20 ;
  assign n22 = ~n16 & ~n21 ;
  assign n23 = ~x2 & ~n22 ;
  assign n24 = ~x2 & ~x5 ;
  assign n25 = ~x0 & ~n24 ;
  assign n26 = x1 & x2 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = ~x9 & ~n27 ;
  assign n29 = ~x2 & ~x3 ;
  assign n30 = x9 & ~n29 ;
  assign n31 = x0 & x3 ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~x1 & ~n32 ;
  assign n34 = x1 & ~x3 ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~n28 & n35 ;
  assign n37 = ~x7 & ~n36 ;
  assign n38 = ~n23 & ~n37 ;
  assign n39 = ~x8 & ~n38 ;
  assign n40 = x7 & x8 ;
  assign n41 = ~x5 & n40 ;
  assign n42 = ~x7 & x9 ;
  assign n43 = ~n41 & ~n42 ;
  assign n44 = x1 & ~n43 ;
  assign n45 = x1 & ~x7 ;
  assign n46 = ~x5 & ~x9 ;
  assign n47 = ~n45 & n46 ;
  assign n48 = ~n44 & ~n47 ;
  assign n49 = x0 & ~x2 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = x2 & ~x9 ;
  assign n52 = ~x0 & ~x1 ;
  assign n53 = n51 & n52 ;
  assign n54 = n41 & n53 ;
  assign n55 = ~n50 & ~n54 ;
  assign n56 = ~x3 & ~n55 ;
  assign n57 = ~n39 & ~n56 ;
  assign n58 = ~x6 & ~n57 ;
  assign n59 = ~x0 & ~x2 ;
  assign n60 = n12 & n59 ;
  assign n61 = ~x5 & ~n60 ;
  assign n62 = x6 & ~n61 ;
  assign n63 = ~x0 & ~x9 ;
  assign n64 = x0 & x9 ;
  assign n65 = ~n63 & ~n64 ;
  assign n66 = x1 & ~n65 ;
  assign n67 = x2 & n66 ;
  assign n68 = x5 & n67 ;
  assign n69 = ~n62 & ~n68 ;
  assign n70 = x8 & ~n69 ;
  assign n71 = ~x1 & ~n13 ;
  assign n72 = ~x8 & ~n71 ;
  assign n73 = ~x1 & x2 ;
  assign n74 = n17 & n73 ;
  assign n75 = ~n72 & ~n74 ;
  assign n76 = ~x5 & ~n75 ;
  assign n77 = ~n70 & ~n76 ;
  assign n78 = x3 & ~n77 ;
  assign n79 = ~x2 & ~n17 ;
  assign n80 = x6 & ~n79 ;
  assign n81 = n29 & n66 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = x5 & ~n82 ;
  assign n84 = x2 & x9 ;
  assign n85 = ~x2 & n19 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = ~x0 & ~x3 ;
  assign n88 = ~n86 & n87 ;
  assign n89 = x6 & n88 ;
  assign n90 = ~n83 & ~n89 ;
  assign n91 = x8 & ~n90 ;
  assign n92 = x2 & ~x3 ;
  assign n93 = n12 & n92 ;
  assign n94 = x1 & ~x8 ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = ~x0 & ~n95 ;
  assign n97 = ~x1 & ~x9 ;
  assign n98 = ~x2 & x6 ;
  assign n99 = x3 & ~n98 ;
  assign n100 = n97 & ~n99 ;
  assign n101 = ~n84 & ~n100 ;
  assign n102 = ~x8 & ~n101 ;
  assign n103 = ~n96 & ~n102 ;
  assign n104 = ~x5 & ~n103 ;
  assign n105 = ~x0 & n29 ;
  assign n106 = ~x8 & n97 ;
  assign n107 = n105 & n106 ;
  assign n108 = ~n104 & ~n107 ;
  assign n109 = ~n91 & n108 ;
  assign n110 = ~n78 & n109 ;
  assign n111 = ~x7 & ~n110 ;
  assign n112 = ~n58 & ~n111 ;
  assign n113 = ~x4 & ~n112 ;
  assign n114 = ~x8 & ~x9 ;
  assign n115 = ~x6 & n114 ;
  assign n116 = x4 & x8 ;
  assign n117 = x6 & n116 ;
  assign n118 = ~n115 & ~n117 ;
  assign n119 = x5 & ~n118 ;
  assign n120 = x6 & ~x9 ;
  assign n121 = x4 & x9 ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = x5 & x6 ;
  assign n124 = ~n122 & ~n123 ;
  assign n125 = ~x8 & n124 ;
  assign n126 = ~n119 & ~n125 ;
  assign n127 = ~x7 & ~n126 ;
  assign n128 = ~x1 & ~x3 ;
  assign n129 = ~x2 & n128 ;
  assign n130 = n127 & n129 ;
  assign n131 = ~x0 & n130 ;
  assign n132 = ~n113 & ~n131 ;
  assign n245 = ~n132 & x10 ;
  assign n133 = x3 & x5 ;
  assign n134 = ~n18 & ~n19 ;
  assign n135 = n133 & n134 ;
  assign n136 = x7 & ~n12 ;
  assign n137 = ~n14 & n136 ;
  assign n138 = ~n135 & ~n137 ;
  assign n139 = x2 & ~n138 ;
  assign n140 = x2 & x5 ;
  assign n141 = x0 & ~n140 ;
  assign n142 = ~x1 & ~x2 ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = x9 & ~n143 ;
  assign n145 = x2 & x3 ;
  assign n146 = ~x9 & ~n145 ;
  assign n147 = ~n87 & ~n146 ;
  assign n148 = x1 & ~n147 ;
  assign n149 = ~x1 & x3 ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = ~n144 & n150 ;
  assign n152 = x7 & ~n151 ;
  assign n153 = ~n139 & ~n152 ;
  assign n154 = x8 & ~n153 ;
  assign n155 = ~x7 & ~x8 ;
  assign n156 = x5 & n155 ;
  assign n157 = x7 & ~x9 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = ~x1 & ~n158 ;
  assign n160 = ~x1 & x7 ;
  assign n161 = x5 & x9 ;
  assign n162 = ~n160 & n161 ;
  assign n163 = ~n159 & ~n162 ;
  assign n164 = ~x0 & x2 ;
  assign n165 = ~n163 & n164 ;
  assign n166 = ~x2 & x9 ;
  assign n167 = x0 & x1 ;
  assign n168 = n166 & n167 ;
  assign n169 = n156 & n168 ;
  assign n170 = ~n165 & ~n169 ;
  assign n171 = x3 & ~n170 ;
  assign n172 = ~n154 & ~n171 ;
  assign n173 = x6 & ~n172 ;
  assign n174 = x0 & x2 ;
  assign n175 = n19 & n174 ;
  assign n176 = x5 & ~n175 ;
  assign n177 = ~x6 & ~n176 ;
  assign n178 = ~x1 & ~n65 ;
  assign n179 = ~x2 & n178 ;
  assign n180 = ~x5 & n179 ;
  assign n181 = ~n177 & ~n180 ;
  assign n182 = ~x8 & ~n181 ;
  assign n183 = x1 & ~n17 ;
  assign n184 = x8 & ~n183 ;
  assign n185 = x1 & ~x2 ;
  assign n186 = n13 & n185 ;
  assign n187 = ~n184 & ~n186 ;
  assign n188 = x5 & ~n187 ;
  assign n189 = ~n182 & ~n188 ;
  assign n190 = ~x3 & ~n189 ;
  assign n191 = x2 & ~n13 ;
  assign n192 = ~x6 & ~n191 ;
  assign n193 = n145 & n178 ;
  assign n194 = ~n192 & ~n193 ;
  assign n195 = ~x5 & ~n194 ;
  assign n196 = ~x2 & ~x9 ;
  assign n197 = x2 & n12 ;
  assign n198 = ~n196 & ~n197 ;
  assign n199 = n31 & ~n198 ;
  assign n200 = ~x6 & n199 ;
  assign n201 = ~n195 & ~n200 ;
  assign n202 = ~x8 & ~n201 ;
  assign n203 = ~x2 & x3 ;
  assign n204 = n19 & n203 ;
  assign n205 = ~x1 & x8 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = x0 & ~n206 ;
  assign n208 = x1 & x9 ;
  assign n209 = x2 & ~x6 ;
  assign n210 = ~x3 & ~n209 ;
  assign n211 = n208 & ~n210 ;
  assign n212 = ~n196 & ~n211 ;
  assign n213 = x8 & ~n212 ;
  assign n214 = ~n207 & ~n213 ;
  assign n215 = x5 & ~n214 ;
  assign n216 = x0 & n145 ;
  assign n217 = x8 & n208 ;
  assign n218 = n216 & n217 ;
  assign n219 = ~n215 & ~n218 ;
  assign n220 = ~n202 & n219 ;
  assign n221 = ~n190 & n220 ;
  assign n222 = x7 & ~n221 ;
  assign n223 = ~n173 & ~n222 ;
  assign n224 = x4 & ~n223 ;
  assign n225 = x8 & x9 ;
  assign n226 = x6 & n225 ;
  assign n227 = ~x4 & ~x8 ;
  assign n228 = ~x6 & n227 ;
  assign n229 = ~n226 & ~n228 ;
  assign n230 = ~x5 & ~n229 ;
  assign n231 = ~x6 & x9 ;
  assign n232 = ~x4 & ~x9 ;
  assign n233 = ~n231 & ~n232 ;
  assign n234 = ~x5 & ~x6 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = x8 & n235 ;
  assign n237 = ~n230 & ~n236 ;
  assign n238 = x7 & ~n237 ;
  assign n239 = x1 & x3 ;
  assign n240 = x2 & n239 ;
  assign n241 = n238 & n240 ;
  assign n242 = x0 & n241 ;
  assign n243 = ~n224 & ~n242 ;
  assign n246 = n243 & ~x10 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = x0 & x8 ;
  assign n249 = n84 & n248 ;
  assign n250 = ~x2 & ~x8 ;
  assign n251 = n63 & n250 ;
  assign n252 = ~n249 & ~n251 ;
  assign n253 = x5 & ~n252 ;
  assign n254 = ~x5 & x8 ;
  assign n255 = x6 & x9 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = ~x0 & ~n256 ;
  assign n258 = x8 & n255 ;
  assign n259 = ~x8 & n46 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = ~n257 & n260 ;
  assign n262 = x2 & ~n261 ;
  assign n263 = ~n253 & ~n262 ;
  assign n264 = ~x4 & ~n263 ;
  assign n265 = x5 & ~x8 ;
  assign n266 = ~n116 & ~n265 ;
  assign n267 = ~x6 & ~n266 ;
  assign n268 = ~n121 & ~n267 ;
  assign n269 = ~n231 & ~n268 ;
  assign n270 = n59 & n269 ;
  assign n271 = ~n264 & ~n270 ;
  assign n272 = ~x1 & ~n271 ;
  assign n273 = x6 & x8 ;
  assign n274 = ~n256 & ~n273 ;
  assign n275 = x0 & n274 ;
  assign n276 = ~x0 & x5 ;
  assign n277 = ~x8 & x9 ;
  assign n278 = n276 & n277 ;
  assign n279 = ~n275 & ~n278 ;
  assign n280 = ~x2 & ~n279 ;
  assign n281 = ~x6 & ~x8 ;
  assign n282 = ~x0 & x6 ;
  assign n283 = ~x2 & ~n282 ;
  assign n284 = n254 & ~n283 ;
  assign n285 = ~n281 & ~n284 ;
  assign n286 = ~x9 & ~n285 ;
  assign n287 = ~n280 & ~n286 ;
  assign n288 = x1 & ~n287 ;
  assign n289 = ~x6 & x8 ;
  assign n290 = n51 & n289 ;
  assign n291 = ~n288 & ~n290 ;
  assign n292 = ~x4 & ~n291 ;
  assign n293 = ~n272 & ~n292 ;
  assign n294 = ~x3 & ~n293 ;
  assign n295 = x5 & n250 ;
  assign n296 = ~x3 & ~x8 ;
  assign n297 = ~n254 & ~n296 ;
  assign n298 = x0 & n297 ;
  assign n299 = ~n295 & ~n298 ;
  assign n300 = ~x1 & ~n299 ;
  assign n301 = x3 & x8 ;
  assign n302 = ~x2 & ~n301 ;
  assign n303 = ~x0 & ~n302 ;
  assign n304 = ~x2 & x8 ;
  assign n305 = x0 & n304 ;
  assign n306 = x0 & ~x5 ;
  assign n307 = ~n276 & ~n306 ;
  assign n308 = ~n305 & n307 ;
  assign n309 = x1 & ~n308 ;
  assign n310 = ~n303 & ~n309 ;
  assign n311 = ~n300 & n310 ;
  assign n312 = ~x6 & ~n311 ;
  assign n313 = ~x1 & x6 ;
  assign n314 = x2 & ~n313 ;
  assign n315 = ~x1 & ~x8 ;
  assign n316 = ~n314 & ~n315 ;
  assign n317 = x3 & n316 ;
  assign n318 = ~x0 & x8 ;
  assign n319 = ~x1 & ~x6 ;
  assign n320 = ~n167 & ~n319 ;
  assign n321 = ~n318 & n320 ;
  assign n322 = ~x2 & n321 ;
  assign n323 = ~n317 & ~n322 ;
  assign n324 = ~x5 & ~n323 ;
  assign n325 = ~n312 & ~n324 ;
  assign n326 = ~x9 & ~n325 ;
  assign n327 = x1 & x5 ;
  assign n328 = x3 & ~x8 ;
  assign n329 = n142 & n328 ;
  assign n330 = ~n327 & ~n329 ;
  assign n331 = x0 & ~n330 ;
  assign n332 = x5 & ~n29 ;
  assign n333 = x3 & n26 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = ~n331 & n334 ;
  assign n336 = x6 & ~n335 ;
  assign n337 = n265 & n333 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = x9 & ~n338 ;
  assign n340 = ~n326 & ~n339 ;
  assign n341 = ~x4 & ~n340 ;
  assign n342 = ~n294 & ~n341 ;
  assign n343 = ~x7 & ~n342 ;
  assign n344 = x2 & ~n52 ;
  assign n345 = n79 & ~n167 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = ~x8 & n346 ;
  assign n348 = n19 & n304 ;
  assign n349 = ~n347 & ~n348 ;
  assign n350 = x7 & ~n349 ;
  assign n351 = ~n53 & ~n350 ;
  assign n352 = ~x4 & ~n351 ;
  assign n353 = ~x6 & n352 ;
  assign n354 = n11 & n353 ;
  assign n355 = ~n343 & ~n354 ;
  assign n456 = ~n355 & x11 ;
  assign n356 = ~x0 & ~x8 ;
  assign n357 = n196 & n356 ;
  assign n358 = x2 & x8 ;
  assign n359 = n64 & n358 ;
  assign n360 = ~n357 & ~n359 ;
  assign n361 = ~x5 & ~n360 ;
  assign n362 = ~x6 & ~x9 ;
  assign n363 = ~n265 & ~n362 ;
  assign n364 = x0 & ~n363 ;
  assign n365 = ~x8 & n362 ;
  assign n366 = x8 & n161 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = ~n364 & n367 ;
  assign n369 = ~x2 & ~n368 ;
  assign n370 = ~n361 & ~n369 ;
  assign n371 = x4 & ~n370 ;
  assign n372 = ~n227 & ~n254 ;
  assign n373 = x6 & ~n372 ;
  assign n374 = ~n232 & ~n373 ;
  assign n375 = ~n120 & ~n374 ;
  assign n376 = n174 & n375 ;
  assign n377 = ~n371 & ~n376 ;
  assign n378 = x1 & ~n377 ;
  assign n379 = ~n281 & ~n363 ;
  assign n380 = ~x0 & n379 ;
  assign n381 = x8 & ~x9 ;
  assign n382 = n306 & n381 ;
  assign n383 = ~n380 & ~n382 ;
  assign n384 = x2 & ~n383 ;
  assign n385 = x0 & ~x6 ;
  assign n386 = x2 & ~n385 ;
  assign n387 = n265 & ~n386 ;
  assign n388 = ~n273 & ~n387 ;
  assign n389 = x9 & ~n388 ;
  assign n390 = ~n384 & ~n389 ;
  assign n391 = ~x1 & ~n390 ;
  assign n392 = x6 & ~x8 ;
  assign n393 = n166 & n392 ;
  assign n394 = ~n391 & ~n393 ;
  assign n395 = x4 & ~n394 ;
  assign n396 = ~n378 & ~n395 ;
  assign n397 = x3 & ~n396 ;
  assign n398 = ~x5 & n358 ;
  assign n399 = ~n265 & ~n301 ;
  assign n400 = ~x0 & n399 ;
  assign n401 = ~n398 & ~n400 ;
  assign n402 = x1 & ~n401 ;
  assign n403 = x2 & ~n296 ;
  assign n404 = x0 & ~n403 ;
  assign n405 = x2 & ~x8 ;
  assign n406 = ~x0 & n405 ;
  assign n407 = n307 & ~n406 ;
  assign n408 = ~x1 & ~n407 ;
  assign n409 = ~n404 & ~n408 ;
  assign n410 = ~n402 & n409 ;
  assign n411 = x6 & ~n410 ;
  assign n412 = x1 & ~x6 ;
  assign n413 = ~x2 & ~n412 ;
  assign n414 = x1 & x8 ;
  assign n415 = ~n413 & ~n414 ;
  assign n416 = ~x3 & n415 ;
  assign n417 = x0 & ~x8 ;
  assign n418 = x1 & x6 ;
  assign n419 = ~n52 & ~n418 ;
  assign n420 = ~n417 & n419 ;
  assign n421 = x2 & n420 ;
  assign n422 = ~n416 & ~n421 ;
  assign n423 = x5 & ~n422 ;
  assign n424 = ~n411 & ~n423 ;
  assign n425 = x9 & ~n424 ;
  assign n426 = ~x1 & ~x5 ;
  assign n427 = ~x3 & x8 ;
  assign n428 = n26 & n427 ;
  assign n429 = ~n426 & ~n428 ;
  assign n430 = ~x0 & ~n429 ;
  assign n431 = ~x5 & ~n145 ;
  assign n432 = ~x3 & n142 ;
  assign n433 = ~n431 & ~n432 ;
  assign n434 = ~n430 & n433 ;
  assign n435 = ~x6 & ~n434 ;
  assign n436 = n254 & n432 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = ~x9 & ~n437 ;
  assign n439 = ~n425 & ~n438 ;
  assign n440 = x4 & ~n439 ;
  assign n441 = ~n397 & ~n440 ;
  assign n442 = x7 & ~n441 ;
  assign n443 = ~x2 & ~n167 ;
  assign n444 = ~n52 & n191 ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = x8 & n445 ;
  assign n447 = n12 & n405 ;
  assign n448 = ~n446 & ~n447 ;
  assign n449 = ~x7 & ~n448 ;
  assign n450 = ~n168 & ~n449 ;
  assign n451 = x4 & ~n450 ;
  assign n452 = x6 & n451 ;
  assign n453 = n133 & n452 ;
  assign n454 = ~n442 & ~n453 ;
  assign n457 = n454 & ~x11 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = ~x3 & x9 ;
  assign n460 = ~n34 & ~n277 ;
  assign n461 = ~n459 & ~n460 ;
  assign n462 = ~x6 & n461 ;
  assign n463 = x3 & ~n304 ;
  assign n464 = x5 & ~n463 ;
  assign n465 = x2 & ~x5 ;
  assign n466 = x3 & ~n465 ;
  assign n467 = x8 & ~n466 ;
  assign n468 = ~n464 & ~n467 ;
  assign n469 = x1 & ~n468 ;
  assign n470 = ~x5 & x6 ;
  assign n471 = ~x8 & n470 ;
  assign n472 = n128 & n471 ;
  assign n473 = ~n469 & ~n472 ;
  assign n474 = ~x9 & ~n473 ;
  assign n475 = ~x1 & ~n302 ;
  assign n476 = x2 & ~n289 ;
  assign n477 = ~n475 & ~n476 ;
  assign n478 = x5 & ~n477 ;
  assign n479 = x6 & ~n414 ;
  assign n480 = ~x9 & ~n479 ;
  assign n481 = ~x2 & ~n480 ;
  assign n482 = ~x1 & n277 ;
  assign n483 = ~n481 & ~n482 ;
  assign n484 = x3 & ~n483 ;
  assign n485 = x1 & n459 ;
  assign n486 = n392 & n485 ;
  assign n487 = ~n484 & ~n486 ;
  assign n488 = ~n478 & n487 ;
  assign n489 = ~n474 & n488 ;
  assign n490 = ~n462 & n489 ;
  assign n491 = ~x4 & ~n490 ;
  assign n492 = ~n281 & ~n381 ;
  assign n493 = ~x5 & n492 ;
  assign n494 = ~x3 & x4 ;
  assign n495 = ~x1 & n494 ;
  assign n496 = ~n493 & n495 ;
  assign n497 = ~x2 & n496 ;
  assign n498 = ~n491 & ~n497 ;
  assign n499 = ~x0 & ~n498 ;
  assign n500 = x8 & n64 ;
  assign n501 = ~n114 & ~n500 ;
  assign n502 = x5 & ~n501 ;
  assign n503 = ~x5 & n84 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = x1 & ~n504 ;
  assign n506 = ~n277 & ~n381 ;
  assign n507 = ~n97 & n506 ;
  assign n508 = x2 & ~n507 ;
  assign n509 = ~n505 & ~n508 ;
  assign n510 = ~x3 & ~n509 ;
  assign n511 = x5 & ~n149 ;
  assign n512 = ~x2 & n114 ;
  assign n513 = ~n511 & n512 ;
  assign n514 = n30 & n205 ;
  assign n515 = ~n513 & ~n514 ;
  assign n516 = x0 & ~n515 ;
  assign n517 = ~n510 & ~n516 ;
  assign n518 = ~x6 & ~n517 ;
  assign n519 = x2 & n208 ;
  assign n520 = ~n205 & ~n519 ;
  assign n521 = x6 & ~n520 ;
  assign n522 = x8 & ~n51 ;
  assign n523 = x2 & n114 ;
  assign n524 = ~n522 & ~n523 ;
  assign n525 = ~n521 & n524 ;
  assign n526 = x3 & ~n525 ;
  assign n527 = x6 & ~n12 ;
  assign n528 = ~n19 & ~n527 ;
  assign n529 = x8 & ~n528 ;
  assign n530 = ~n97 & ~n208 ;
  assign n531 = n296 & ~n530 ;
  assign n532 = ~n529 & ~n531 ;
  assign n533 = ~x2 & ~n532 ;
  assign n534 = ~n526 & ~n533 ;
  assign n535 = n306 & ~n534 ;
  assign n536 = ~n518 & ~n535 ;
  assign n537 = ~x4 & ~n536 ;
  assign n538 = ~n499 & ~n537 ;
  assign n539 = ~x7 & ~n538 ;
  assign n540 = n40 & n64 ;
  assign n541 = ~n63 & ~n540 ;
  assign n542 = x1 & ~n541 ;
  assign n543 = n17 & n315 ;
  assign n544 = ~n542 & ~n543 ;
  assign n545 = ~x4 & ~n544 ;
  assign n546 = n29 & n545 ;
  assign n547 = n234 & n546 ;
  assign n548 = ~n539 & ~n547 ;
  assign n638 = ~n548 & x12 ;
  assign n549 = x3 & ~x9 ;
  assign n550 = ~n149 & ~n381 ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = x6 & n551 ;
  assign n553 = ~x3 & ~n405 ;
  assign n554 = ~x5 & ~n553 ;
  assign n555 = ~x2 & x5 ;
  assign n556 = ~x3 & ~n555 ;
  assign n557 = ~x8 & ~n556 ;
  assign n558 = ~n554 & ~n557 ;
  assign n559 = ~x1 & ~n558 ;
  assign n560 = x5 & ~x6 ;
  assign n561 = x8 & n560 ;
  assign n562 = n239 & n561 ;
  assign n563 = ~n559 & ~n562 ;
  assign n564 = x9 & ~n563 ;
  assign n565 = x1 & ~n403 ;
  assign n566 = ~x2 & ~n392 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = ~x5 & ~n567 ;
  assign n569 = ~x6 & ~n315 ;
  assign n570 = x9 & ~n569 ;
  assign n571 = x2 & ~n570 ;
  assign n572 = x1 & n381 ;
  assign n573 = ~n571 & ~n572 ;
  assign n574 = ~x3 & ~n573 ;
  assign n575 = ~x1 & n549 ;
  assign n576 = n289 & n575 ;
  assign n577 = ~n574 & ~n576 ;
  assign n578 = ~n568 & n577 ;
  assign n579 = ~n564 & n578 ;
  assign n580 = ~n552 & n579 ;
  assign n581 = x4 & ~n580 ;
  assign n582 = ~n273 & ~n277 ;
  assign n583 = x5 & n582 ;
  assign n584 = x3 & ~x4 ;
  assign n585 = x1 & n584 ;
  assign n586 = ~n583 & n585 ;
  assign n587 = x2 & n586 ;
  assign n588 = ~n581 & ~n587 ;
  assign n589 = x0 & ~n588 ;
  assign n590 = ~x8 & n63 ;
  assign n591 = ~n225 & ~n590 ;
  assign n592 = ~x5 & ~n591 ;
  assign n593 = x5 & n196 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~x1 & ~n594 ;
  assign n596 = ~n208 & n506 ;
  assign n597 = ~x2 & ~n596 ;
  assign n598 = ~n595 & ~n597 ;
  assign n599 = x3 & ~n598 ;
  assign n600 = ~x5 & ~n34 ;
  assign n601 = x2 & n225 ;
  assign n602 = ~n600 & n601 ;
  assign n603 = n94 & n146 ;
  assign n604 = ~n602 & ~n603 ;
  assign n605 = ~x0 & ~n604 ;
  assign n606 = ~n599 & ~n605 ;
  assign n607 = x6 & ~n606 ;
  assign n608 = ~x2 & n97 ;
  assign n609 = ~n94 & ~n608 ;
  assign n610 = ~x6 & ~n609 ;
  assign n611 = ~x8 & ~n166 ;
  assign n612 = ~x2 & n225 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = ~n610 & n613 ;
  assign n615 = ~x3 & ~n614 ;
  assign n616 = ~x6 & ~n19 ;
  assign n617 = ~n12 & ~n616 ;
  assign n618 = ~x8 & ~n617 ;
  assign n619 = n301 & ~n530 ;
  assign n620 = ~n618 & ~n619 ;
  assign n621 = x2 & ~n620 ;
  assign n622 = ~n615 & ~n621 ;
  assign n623 = n276 & ~n622 ;
  assign n624 = ~n607 & ~n623 ;
  assign n625 = x4 & ~n624 ;
  assign n626 = ~n589 & ~n625 ;
  assign n627 = x7 & ~n626 ;
  assign n628 = n63 & n155 ;
  assign n629 = ~n64 & ~n628 ;
  assign n630 = ~x1 & ~n629 ;
  assign n631 = n13 & n414 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = x4 & ~n632 ;
  assign n634 = n145 & n633 ;
  assign n635 = n123 & n634 ;
  assign n636 = ~n627 & ~n635 ;
  assign n639 = n636 & ~x12 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = x3 & ~n231 ;
  assign n642 = x2 & x6 ;
  assign n643 = ~n641 & ~n642 ;
  assign n644 = ~x4 & ~n643 ;
  assign n645 = n225 & n234 ;
  assign n646 = ~n123 & ~n645 ;
  assign n647 = ~x2 & n494 ;
  assign n648 = ~n646 & n647 ;
  assign n649 = ~n644 & ~n648 ;
  assign n650 = ~x1 & ~n649 ;
  assign n651 = x5 & x8 ;
  assign n652 = n231 & n651 ;
  assign n653 = ~n259 & ~n652 ;
  assign n654 = x2 & ~n653 ;
  assign n655 = x5 & ~n289 ;
  assign n656 = x3 & ~n655 ;
  assign n657 = ~n471 & ~n656 ;
  assign n658 = ~n654 & n657 ;
  assign n659 = x1 & ~n658 ;
  assign n660 = x2 & n470 ;
  assign n661 = ~n659 & ~n660 ;
  assign n662 = ~x4 & ~n661 ;
  assign n663 = ~n650 & ~n662 ;
  assign n664 = ~x0 & ~n663 ;
  assign n665 = x2 & ~n297 ;
  assign n666 = ~x2 & n651 ;
  assign n667 = ~n665 & ~n666 ;
  assign n668 = ~x9 & ~n667 ;
  assign n669 = ~x8 & n161 ;
  assign n670 = ~x3 & ~n669 ;
  assign n671 = ~x2 & ~n670 ;
  assign n672 = ~x6 & ~n328 ;
  assign n673 = x3 & ~x5 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~n671 & ~n674 ;
  assign n676 = ~n668 & n675 ;
  assign n677 = x1 & ~n676 ;
  assign n678 = ~x3 & n470 ;
  assign n679 = n295 & n319 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = ~x9 & ~n680 ;
  assign n682 = ~n677 & ~n681 ;
  assign n683 = x0 & ~n682 ;
  assign n684 = ~n29 & n470 ;
  assign n685 = x3 & ~x6 ;
  assign n686 = x2 & n685 ;
  assign n687 = ~n684 & ~n686 ;
  assign n688 = x9 & ~n687 ;
  assign n689 = ~x9 & n470 ;
  assign n690 = ~n685 & ~n689 ;
  assign n691 = ~x8 & ~n690 ;
  assign n692 = ~n688 & ~n691 ;
  assign n693 = ~x1 & ~n692 ;
  assign n694 = ~n46 & ~n281 ;
  assign n695 = ~x2 & ~n694 ;
  assign n696 = ~x6 & ~n161 ;
  assign n697 = ~n208 & ~n651 ;
  assign n698 = n696 & ~n697 ;
  assign n699 = ~n695 & ~n698 ;
  assign n700 = x3 & ~n699 ;
  assign n701 = n470 & n572 ;
  assign n702 = ~n700 & ~n701 ;
  assign n703 = ~n693 & n702 ;
  assign n704 = ~n683 & n703 ;
  assign n705 = ~x4 & ~n704 ;
  assign n706 = ~n664 & ~n705 ;
  assign n707 = ~x7 & ~n706 ;
  assign n776 = n707 & x13 ;
  assign n708 = ~x3 & ~n120 ;
  assign n709 = ~x2 & ~x6 ;
  assign n710 = ~n708 & ~n709 ;
  assign n711 = x4 & ~n710 ;
  assign n712 = n114 & n123 ;
  assign n713 = ~n234 & ~n712 ;
  assign n714 = x2 & n584 ;
  assign n715 = ~n713 & n714 ;
  assign n716 = ~n711 & ~n715 ;
  assign n717 = x1 & ~n716 ;
  assign n718 = ~x5 & ~x8 ;
  assign n719 = n120 & n718 ;
  assign n720 = ~n366 & ~n719 ;
  assign n721 = ~x2 & ~n720 ;
  assign n722 = ~x5 & ~n392 ;
  assign n723 = ~x3 & ~n722 ;
  assign n724 = ~n561 & ~n723 ;
  assign n725 = ~n721 & n724 ;
  assign n726 = ~x1 & ~n725 ;
  assign n727 = ~x2 & n560 ;
  assign n728 = ~n726 & ~n727 ;
  assign n729 = x4 & ~n728 ;
  assign n730 = ~n717 & ~n729 ;
  assign n731 = x0 & ~n730 ;
  assign n732 = ~x2 & ~n399 ;
  assign n733 = x2 & n718 ;
  assign n734 = ~n732 & ~n733 ;
  assign n735 = x9 & ~n734 ;
  assign n736 = x8 & n46 ;
  assign n737 = x3 & ~n736 ;
  assign n738 = x2 & ~n737 ;
  assign n739 = x6 & ~n427 ;
  assign n740 = ~x3 & x5 ;
  assign n741 = ~n739 & ~n740 ;
  assign n742 = ~n738 & ~n741 ;
  assign n743 = ~n735 & n742 ;
  assign n744 = ~x1 & ~n743 ;
  assign n745 = x3 & n560 ;
  assign n746 = n398 & n418 ;
  assign n747 = ~n745 & ~n746 ;
  assign n748 = x9 & ~n747 ;
  assign n749 = ~n744 & ~n748 ;
  assign n750 = ~x0 & ~n749 ;
  assign n751 = ~n145 & n560 ;
  assign n752 = ~x3 & x6 ;
  assign n753 = ~x2 & n752 ;
  assign n754 = ~n751 & ~n753 ;
  assign n755 = ~x9 & ~n754 ;
  assign n756 = x9 & n560 ;
  assign n757 = ~n752 & ~n756 ;
  assign n758 = x8 & ~n757 ;
  assign n759 = ~n755 & ~n758 ;
  assign n760 = x1 & ~n759 ;
  assign n761 = ~n161 & ~n273 ;
  assign n762 = x2 & ~n761 ;
  assign n763 = x6 & ~n46 ;
  assign n764 = ~n97 & ~n718 ;
  assign n765 = n763 & ~n764 ;
  assign n766 = ~n762 & ~n765 ;
  assign n767 = ~x3 & ~n766 ;
  assign n768 = n482 & n560 ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~n760 & n769 ;
  assign n771 = ~n750 & n770 ;
  assign n772 = x4 & ~n771 ;
  assign n773 = ~n731 & ~n772 ;
  assign n774 = x7 & ~n773 ;
  assign n777 = ~n774 & ~x13 ;
  assign n778 = ~n776 & ~n777 ;
  assign n779 = ~x4 & n344 ;
  assign n780 = ~n494 & ~n584 ;
  assign n781 = ~x0 & n142 ;
  assign n782 = ~n780 & n781 ;
  assign n783 = ~n779 & ~n782 ;
  assign n784 = ~x7 & ~n783 ;
  assign n785 = n123 & n784 ;
  assign n793 = n785 & x14 ;
  assign n786 = x4 & n443 ;
  assign n787 = x0 & n26 ;
  assign n788 = ~n780 & n787 ;
  assign n789 = ~n786 & ~n788 ;
  assign n790 = x7 & ~n789 ;
  assign n791 = n234 & n790 ;
  assign n794 = ~n791 & ~x14 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = n52 & n647 ;
  assign n797 = n584 & ~n781 ;
  assign n798 = ~n796 & ~n797 ;
  assign n799 = ~x7 & ~n798 ;
  assign n800 = n123 & n799 ;
  assign n807 = n800 & x15 ;
  assign n801 = n167 & n714 ;
  assign n802 = n494 & ~n787 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = x7 & ~n803 ;
  assign n805 = n234 & n804 ;
  assign n808 = ~n805 & ~x15 ;
  assign n809 = ~n807 & ~n808 ;
  assign n810 = x2 & ~n426 ;
  assign n811 = ~x9 & ~n810 ;
  assign n812 = ~x6 & n811 ;
  assign n813 = x5 & n208 ;
  assign n814 = ~n812 & ~n813 ;
  assign n815 = x0 & ~n814 ;
  assign n816 = ~x0 & ~n46 ;
  assign n817 = x2 & n816 ;
  assign n818 = ~n815 & ~n817 ;
  assign n819 = x8 & ~n818 ;
  assign n820 = x2 & n13 ;
  assign n821 = ~n106 & ~n820 ;
  assign n822 = x5 & ~n821 ;
  assign n823 = ~n819 & ~n822 ;
  assign n824 = ~n114 & ~n225 ;
  assign n825 = x6 & ~n824 ;
  assign n826 = ~n51 & ~n166 ;
  assign n827 = n825 & n826 ;
  assign n828 = n823 & ~n827 ;
  assign n829 = ~x7 & ~n828 ;
  assign n830 = x8 & ~n157 ;
  assign n831 = n73 & ~n830 ;
  assign n832 = ~n85 & ~n831 ;
  assign n833 = ~x0 & ~n832 ;
  assign n834 = n208 & n248 ;
  assign n835 = ~n114 & ~n834 ;
  assign n836 = x7 & ~n835 ;
  assign n837 = ~x2 & n836 ;
  assign n838 = ~n833 & ~n837 ;
  assign n839 = n234 & ~n838 ;
  assign n840 = ~n829 & ~n839 ;
  assign n841 = ~x3 & ~n840 ;
  assign n842 = ~n106 & ~n208 ;
  assign n843 = x0 & ~n842 ;
  assign n844 = x2 & n19 ;
  assign n845 = ~n843 & ~n844 ;
  assign n846 = ~x0 & ~x6 ;
  assign n847 = ~n315 & n530 ;
  assign n848 = n846 & n847 ;
  assign n849 = n845 & ~n848 ;
  assign n850 = ~x5 & ~n849 ;
  assign n851 = ~x8 & n167 ;
  assign n852 = x0 & n273 ;
  assign n853 = ~n94 & ~n852 ;
  assign n854 = ~x2 & ~n853 ;
  assign n855 = ~n851 & ~n854 ;
  assign n856 = x9 & ~n855 ;
  assign n857 = ~n306 & ~n356 ;
  assign n858 = n19 & n857 ;
  assign n859 = ~n856 & ~n858 ;
  assign n860 = ~n850 & n859 ;
  assign n861 = x3 & ~n860 ;
  assign n862 = ~n65 & n555 ;
  assign n863 = ~x6 & ~n465 ;
  assign n864 = n13 & ~n863 ;
  assign n865 = ~n862 & ~n864 ;
  assign n866 = ~x8 & ~n865 ;
  assign n867 = x2 & ~n114 ;
  assign n868 = ~n500 & ~n867 ;
  assign n869 = x6 & ~n868 ;
  assign n870 = ~n866 & ~n869 ;
  assign n871 = x1 & ~n870 ;
  assign n872 = ~x8 & ~n846 ;
  assign n873 = ~n306 & ~n872 ;
  assign n874 = ~x9 & ~n873 ;
  assign n875 = ~x2 & n874 ;
  assign n876 = n13 & n358 ;
  assign n877 = ~n875 & ~n876 ;
  assign n878 = ~x1 & ~n877 ;
  assign n879 = ~n871 & ~n878 ;
  assign n880 = ~n861 & n879 ;
  assign n881 = ~x7 & ~n880 ;
  assign n882 = ~n841 & ~n881 ;
  assign n883 = ~x4 & ~n882 ;
  assign n884 = ~x1 & x4 ;
  assign n885 = n105 & n884 ;
  assign n886 = ~n123 & ~n885 ;
  assign n887 = ~x7 & ~n886 ;
  assign n888 = ~n883 & ~n887 ;
  assign n967 = n888 & x16 ;
  assign n889 = ~x2 & ~n327 ;
  assign n890 = x9 & ~n889 ;
  assign n891 = x6 & n890 ;
  assign n892 = ~x5 & n97 ;
  assign n893 = ~n891 & ~n892 ;
  assign n894 = ~x0 & ~n893 ;
  assign n895 = x0 & ~n161 ;
  assign n896 = ~x2 & n895 ;
  assign n897 = ~n894 & ~n896 ;
  assign n898 = ~x8 & ~n897 ;
  assign n899 = ~x2 & n17 ;
  assign n900 = ~n217 & ~n899 ;
  assign n901 = ~x5 & ~n900 ;
  assign n902 = ~n898 & ~n901 ;
  assign n903 = ~x6 & ~n824 ;
  assign n904 = n826 & n903 ;
  assign n905 = n902 & ~n904 ;
  assign n906 = x7 & ~n905 ;
  assign n907 = ~x8 & ~n42 ;
  assign n908 = n185 & ~n907 ;
  assign n909 = ~n197 & ~n908 ;
  assign n910 = x0 & ~n909 ;
  assign n911 = n97 & n356 ;
  assign n912 = ~n225 & ~n911 ;
  assign n913 = ~x7 & ~n912 ;
  assign n914 = x2 & n913 ;
  assign n915 = ~n910 & ~n914 ;
  assign n916 = n123 & ~n915 ;
  assign n917 = ~n906 & ~n916 ;
  assign n918 = x3 & ~n917 ;
  assign n919 = ~n97 & ~n217 ;
  assign n920 = ~x0 & ~n919 ;
  assign n921 = ~x2 & n12 ;
  assign n922 = ~n920 & ~n921 ;
  assign n923 = x0 & x6 ;
  assign n924 = ~n414 & n530 ;
  assign n925 = n923 & n924 ;
  assign n926 = n922 & ~n925 ;
  assign n927 = x5 & ~n926 ;
  assign n928 = x8 & n52 ;
  assign n929 = ~x0 & n281 ;
  assign n930 = ~n205 & ~n929 ;
  assign n931 = x2 & ~n930 ;
  assign n932 = ~n928 & ~n931 ;
  assign n933 = ~x9 & ~n932 ;
  assign n934 = ~n248 & ~n276 ;
  assign n935 = n12 & n934 ;
  assign n936 = ~n933 & ~n935 ;
  assign n937 = ~n927 & n936 ;
  assign n938 = ~x3 & ~n937 ;
  assign n939 = ~n65 & n465 ;
  assign n940 = x6 & ~n555 ;
  assign n941 = n17 & ~n940 ;
  assign n942 = ~n939 & ~n941 ;
  assign n943 = x8 & ~n942 ;
  assign n944 = ~x2 & ~n225 ;
  assign n945 = ~n590 & ~n944 ;
  assign n946 = ~x6 & ~n945 ;
  assign n947 = ~n943 & ~n946 ;
  assign n948 = ~x1 & ~n947 ;
  assign n949 = x8 & ~n923 ;
  assign n950 = ~n276 & ~n949 ;
  assign n951 = x9 & ~n950 ;
  assign n952 = x2 & n951 ;
  assign n953 = n17 & n250 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = x1 & ~n954 ;
  assign n956 = ~n948 & ~n955 ;
  assign n957 = ~n938 & n956 ;
  assign n958 = x7 & ~n957 ;
  assign n959 = ~n918 & ~n958 ;
  assign n960 = x4 & ~n959 ;
  assign n961 = x1 & ~x4 ;
  assign n962 = n216 & n961 ;
  assign n963 = ~n234 & ~n962 ;
  assign n964 = x7 & ~n963 ;
  assign n965 = ~n960 & ~n964 ;
  assign n968 = ~n965 & ~x16 ;
  assign n969 = ~n967 & ~n968 ;
  assign n970 = ~n255 & ~n427 ;
  assign n971 = x0 & ~n970 ;
  assign n972 = n318 & n685 ;
  assign n973 = ~n392 & ~n972 ;
  assign n974 = x9 & ~n973 ;
  assign n975 = ~x9 & n273 ;
  assign n976 = ~n974 & ~n975 ;
  assign n977 = ~n971 & n976 ;
  assign n978 = ~x2 & ~n977 ;
  assign n979 = ~x3 & n225 ;
  assign n980 = x3 & ~n225 ;
  assign n981 = ~n248 & ~n980 ;
  assign n982 = ~x6 & ~n981 ;
  assign n983 = ~n979 & ~n982 ;
  assign n984 = x2 & ~n983 ;
  assign n985 = ~x3 & n115 ;
  assign n986 = ~n984 & ~n985 ;
  assign n987 = ~n978 & n986 ;
  assign n988 = x1 & ~n987 ;
  assign n989 = ~n63 & ~n277 ;
  assign n990 = ~x6 & ~n989 ;
  assign n991 = ~x2 & n990 ;
  assign n992 = ~x0 & n825 ;
  assign n993 = ~n991 & ~n992 ;
  assign n994 = x3 & ~n993 ;
  assign n995 = ~x0 & n250 ;
  assign n996 = ~n852 & ~n995 ;
  assign n997 = ~x9 & ~n996 ;
  assign n998 = ~x6 & ~n296 ;
  assign n999 = n867 & ~n998 ;
  assign n1000 = ~n997 & ~n999 ;
  assign n1001 = ~n994 & n1000 ;
  assign n1002 = ~x1 & ~n1001 ;
  assign n1003 = ~x9 & n392 ;
  assign n1004 = n203 & n1003 ;
  assign n1005 = ~n1002 & ~n1004 ;
  assign n1006 = ~n988 & n1005 ;
  assign n1007 = ~x5 & ~n1006 ;
  assign n1008 = x0 & ~n826 ;
  assign n1009 = x5 & ~x9 ;
  assign n1010 = ~x0 & n1009 ;
  assign n1011 = ~n1008 & ~n1010 ;
  assign n1012 = x8 & ~n1011 ;
  assign n1013 = n84 & n265 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = ~x3 & ~n1014 ;
  assign n1016 = ~n51 & ~n133 ;
  assign n1017 = ~x0 & ~n1016 ;
  assign n1018 = x3 & n555 ;
  assign n1019 = ~n1017 & ~n1018 ;
  assign n1020 = ~x8 & ~n1019 ;
  assign n1021 = n203 & n1009 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = ~n1015 & n1022 ;
  assign n1024 = x1 & ~n1023 ;
  assign n1025 = ~x2 & ~n31 ;
  assign n1026 = ~n824 & ~n1025 ;
  assign n1027 = ~n145 & ~n1026 ;
  assign n1028 = x5 & ~n1027 ;
  assign n1029 = n31 & n523 ;
  assign n1030 = ~n1028 & ~n1029 ;
  assign n1031 = ~x1 & ~n1030 ;
  assign n1032 = n145 & n366 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = ~n1024 & n1033 ;
  assign n1035 = ~x6 & ~n1034 ;
  assign n1036 = ~n1007 & ~n1035 ;
  assign n1037 = ~x7 & ~n1036 ;
  assign n1038 = x2 & ~n506 ;
  assign n1039 = ~x0 & n1038 ;
  assign n1040 = ~x9 & n40 ;
  assign n1041 = n49 & n1040 ;
  assign n1042 = ~n1039 & ~n1041 ;
  assign n1043 = n319 & ~n1042 ;
  assign n1044 = n11 & n1043 ;
  assign n1045 = ~n1037 & ~n1044 ;
  assign n1046 = ~x4 & ~n1045 ;
  assign n1047 = n24 & n87 ;
  assign n1048 = x4 & ~x7 ;
  assign n1049 = n319 & n1048 ;
  assign n1050 = n1047 & n1049 ;
  assign n1051 = ~n1046 & ~n1050 ;
  assign n1135 = n1051 & x17 ;
  assign n1052 = ~n328 & ~n362 ;
  assign n1053 = ~x0 & ~n1052 ;
  assign n1054 = n417 & n752 ;
  assign n1055 = ~n289 & ~n1054 ;
  assign n1056 = ~x9 & ~n1055 ;
  assign n1057 = x9 & n281 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = ~n1053 & n1058 ;
  assign n1060 = x2 & ~n1059 ;
  assign n1061 = x3 & n114 ;
  assign n1062 = ~x3 & ~n114 ;
  assign n1063 = ~n356 & ~n1062 ;
  assign n1064 = x6 & ~n1063 ;
  assign n1065 = ~n1061 & ~n1064 ;
  assign n1066 = ~x2 & ~n1065 ;
  assign n1067 = x3 & n226 ;
  assign n1068 = ~n1066 & ~n1067 ;
  assign n1069 = ~n1060 & n1068 ;
  assign n1070 = ~x1 & ~n1069 ;
  assign n1071 = ~n64 & ~n381 ;
  assign n1072 = x6 & ~n1071 ;
  assign n1073 = x2 & n1072 ;
  assign n1074 = x0 & n903 ;
  assign n1075 = ~n1073 & ~n1074 ;
  assign n1076 = ~x3 & ~n1075 ;
  assign n1077 = x0 & n358 ;
  assign n1078 = ~n929 & ~n1077 ;
  assign n1079 = x9 & ~n1078 ;
  assign n1080 = x6 & ~n301 ;
  assign n1081 = n944 & ~n1080 ;
  assign n1082 = ~n1079 & ~n1081 ;
  assign n1083 = ~n1076 & n1082 ;
  assign n1084 = x1 & ~n1083 ;
  assign n1085 = x9 & n289 ;
  assign n1086 = n92 & n1085 ;
  assign n1087 = ~n1084 & ~n1086 ;
  assign n1088 = ~n1070 & n1087 ;
  assign n1089 = x5 & ~n1088 ;
  assign n1090 = ~x0 & ~n826 ;
  assign n1091 = ~x5 & x9 ;
  assign n1092 = x0 & n1091 ;
  assign n1093 = ~n1090 & ~n1092 ;
  assign n1094 = ~x8 & ~n1093 ;
  assign n1095 = n196 & n254 ;
  assign n1096 = ~n1094 & ~n1095 ;
  assign n1097 = x3 & ~n1096 ;
  assign n1098 = ~n11 & ~n166 ;
  assign n1099 = x0 & ~n1098 ;
  assign n1100 = ~x3 & n465 ;
  assign n1101 = ~n1099 & ~n1100 ;
  assign n1102 = x8 & ~n1101 ;
  assign n1103 = n92 & n1091 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1105 = ~n1097 & n1104 ;
  assign n1106 = ~x1 & ~n1105 ;
  assign n1107 = x2 & ~n87 ;
  assign n1108 = ~n824 & ~n1107 ;
  assign n1109 = ~n29 & ~n1108 ;
  assign n1110 = ~x5 & ~n1109 ;
  assign n1111 = n87 & n612 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1113 = x1 & ~n1112 ;
  assign n1114 = n29 & n259 ;
  assign n1115 = ~n1113 & ~n1114 ;
  assign n1116 = ~n1106 & n1115 ;
  assign n1117 = x6 & ~n1116 ;
  assign n1118 = ~n1089 & ~n1117 ;
  assign n1119 = x7 & ~n1118 ;
  assign n1120 = ~x2 & ~n506 ;
  assign n1121 = x0 & n1120 ;
  assign n1122 = x9 & n155 ;
  assign n1123 = n164 & n1122 ;
  assign n1124 = ~n1121 & ~n1123 ;
  assign n1125 = n418 & ~n1124 ;
  assign n1126 = n133 & n1125 ;
  assign n1127 = ~n1119 & ~n1126 ;
  assign n1128 = x4 & ~n1127 ;
  assign n1129 = n31 & n140 ;
  assign n1130 = ~x4 & x7 ;
  assign n1131 = n418 & n1130 ;
  assign n1132 = n1129 & n1131 ;
  assign n1133 = ~n1128 & ~n1132 ;
  assign n1136 = ~n1133 & ~x17 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = n142 & n1009 ;
  assign n1139 = ~n485 & ~n1138 ;
  assign n1140 = ~x0 & ~n1139 ;
  assign n1141 = ~x1 & x5 ;
  assign n1142 = ~n11 & ~n1141 ;
  assign n1143 = ~n97 & ~n459 ;
  assign n1144 = ~n1142 & n1143 ;
  assign n1145 = ~x2 & n1144 ;
  assign n1146 = ~n426 & n530 ;
  assign n1147 = n92 & ~n1146 ;
  assign n1148 = ~n1145 & ~n1147 ;
  assign n1149 = ~n1140 & n1148 ;
  assign n1150 = ~x8 & ~n1149 ;
  assign n1151 = ~n87 & ~n1142 ;
  assign n1152 = ~x2 & n1151 ;
  assign n1153 = n128 & n306 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = x8 & ~n1154 ;
  assign n1156 = ~x5 & ~n318 ;
  assign n1157 = ~n133 & ~n1156 ;
  assign n1158 = n26 & n1157 ;
  assign n1159 = ~n1155 & ~n1158 ;
  assign n1160 = ~x9 & ~n1159 ;
  assign n1161 = ~n133 & ~n465 ;
  assign n1162 = ~n463 & ~n1161 ;
  assign n1163 = x1 & n1162 ;
  assign n1164 = n149 & ~n276 ;
  assign n1165 = n304 & n1164 ;
  assign n1166 = ~n1163 & ~n1165 ;
  assign n1167 = x9 & ~n1166 ;
  assign n1168 = ~n1160 & ~n1167 ;
  assign n1169 = ~n1150 & n1168 ;
  assign n1170 = ~x6 & ~n1169 ;
  assign n1171 = ~x1 & ~n114 ;
  assign n1172 = x2 & ~n1171 ;
  assign n1173 = ~n527 & ~n1172 ;
  assign n1174 = x0 & ~n1173 ;
  assign n1175 = ~x6 & ~n94 ;
  assign n1176 = x2 & ~n1175 ;
  assign n1177 = x8 & ~n19 ;
  assign n1178 = n527 & ~n1177 ;
  assign n1179 = ~n1176 & ~n1178 ;
  assign n1180 = ~n1174 & n1179 ;
  assign n1181 = n673 & ~n1180 ;
  assign n1182 = ~n1170 & ~n1181 ;
  assign n1183 = ~x7 & ~n1182 ;
  assign n1184 = ~n250 & ~n358 ;
  assign n1185 = ~x0 & ~n1184 ;
  assign n1186 = ~n305 & ~n1185 ;
  assign n1187 = ~x9 & ~n1186 ;
  assign n1188 = n84 & n356 ;
  assign n1189 = ~n1187 & ~n1188 ;
  assign n1190 = ~x1 & ~n1189 ;
  assign n1191 = n208 & n995 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1193 = n11 & ~n1192 ;
  assign n1194 = ~x6 & n1193 ;
  assign n1195 = ~n1183 & ~n1194 ;
  assign n1196 = ~x4 & ~n1195 ;
  assign n1197 = n11 & n1048 ;
  assign n1198 = n781 & n1197 ;
  assign n1199 = ~n1196 & ~n1198 ;
  assign n1262 = n1199 & x18 ;
  assign n1200 = n26 & n1091 ;
  assign n1201 = ~n575 & ~n1200 ;
  assign n1202 = x0 & ~n1201 ;
  assign n1203 = x1 & ~x5 ;
  assign n1204 = ~n133 & ~n1203 ;
  assign n1205 = ~n208 & ~n549 ;
  assign n1206 = ~n1204 & n1205 ;
  assign n1207 = x2 & n1206 ;
  assign n1208 = ~n327 & n530 ;
  assign n1209 = n203 & ~n1208 ;
  assign n1210 = ~n1207 & ~n1209 ;
  assign n1211 = ~n1202 & n1210 ;
  assign n1212 = x8 & ~n1211 ;
  assign n1213 = ~n31 & ~n1204 ;
  assign n1214 = x2 & n1213 ;
  assign n1215 = n239 & n276 ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = ~x8 & ~n1216 ;
  assign n1218 = x5 & ~n417 ;
  assign n1219 = ~n11 & ~n1218 ;
  assign n1220 = n142 & n1219 ;
  assign n1221 = ~n1217 & ~n1220 ;
  assign n1222 = x9 & ~n1221 ;
  assign n1223 = ~n11 & ~n555 ;
  assign n1224 = ~n553 & ~n1223 ;
  assign n1225 = ~x1 & n1224 ;
  assign n1226 = n34 & ~n306 ;
  assign n1227 = n405 & n1226 ;
  assign n1228 = ~n1225 & ~n1227 ;
  assign n1229 = ~x9 & ~n1228 ;
  assign n1230 = ~n1222 & ~n1229 ;
  assign n1231 = ~n1212 & n1230 ;
  assign n1232 = x6 & ~n1231 ;
  assign n1233 = x1 & ~n225 ;
  assign n1234 = ~x2 & ~n1233 ;
  assign n1235 = ~n616 & ~n1234 ;
  assign n1236 = ~x0 & ~n1235 ;
  assign n1237 = x6 & ~n205 ;
  assign n1238 = ~x2 & ~n1237 ;
  assign n1239 = ~x8 & ~n12 ;
  assign n1240 = n616 & ~n1239 ;
  assign n1241 = ~n1238 & ~n1240 ;
  assign n1242 = ~n1236 & n1241 ;
  assign n1243 = n740 & ~n1242 ;
  assign n1244 = ~n1232 & ~n1243 ;
  assign n1245 = x7 & ~n1244 ;
  assign n1246 = x0 & ~n1184 ;
  assign n1247 = ~n406 & ~n1246 ;
  assign n1248 = x9 & ~n1247 ;
  assign n1249 = n196 & n248 ;
  assign n1250 = ~n1248 & ~n1249 ;
  assign n1251 = x1 & ~n1250 ;
  assign n1252 = n97 & n1077 ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = n133 & ~n1253 ;
  assign n1255 = x6 & n1254 ;
  assign n1256 = ~n1245 & ~n1255 ;
  assign n1257 = x4 & ~n1256 ;
  assign n1258 = n133 & n1130 ;
  assign n1259 = n787 & n1258 ;
  assign n1260 = ~n1257 & ~n1259 ;
  assign n1263 = ~n1260 & ~x18 ;
  assign n1264 = ~n1262 & ~n1263 ;
  assign n1265 = x4 & ~n129 ;
  assign n1266 = n306 & n686 ;
  assign n1267 = ~x7 & ~n1266 ;
  assign n1268 = ~n1171 & ~n1267 ;
  assign n1269 = ~x7 & ~n129 ;
  assign n1270 = x0 & ~n1269 ;
  assign n1271 = x7 & ~n92 ;
  assign n1272 = ~x3 & ~n46 ;
  assign n1273 = x3 & ~n255 ;
  assign n1274 = n318 & ~n1273 ;
  assign n1275 = ~n1272 & ~n1274 ;
  assign n1276 = ~x2 & ~n1275 ;
  assign n1277 = ~n225 & n686 ;
  assign n1278 = ~x5 & n1277 ;
  assign n1279 = ~x6 & ~n366 ;
  assign n1280 = ~x3 & ~n1279 ;
  assign n1281 = ~n1278 & ~n1280 ;
  assign n1282 = ~n1276 & n1281 ;
  assign n1283 = x1 & ~n1282 ;
  assign n1284 = n318 & ~n696 ;
  assign n1285 = ~n255 & ~n1284 ;
  assign n1286 = x3 & ~n1285 ;
  assign n1287 = x4 & ~n234 ;
  assign n1288 = ~x3 & ~n1287 ;
  assign n1289 = ~n1286 & ~n1288 ;
  assign n1290 = ~x2 & ~n1289 ;
  assign n1291 = ~x8 & ~n161 ;
  assign n1292 = n1272 & ~n1291 ;
  assign n1293 = x2 & n1292 ;
  assign n1294 = ~n1290 & ~n1293 ;
  assign n1295 = ~x1 & ~n1294 ;
  assign n1296 = ~x5 & ~n92 ;
  assign n1297 = x6 & ~n1296 ;
  assign n1298 = ~n1295 & ~n1297 ;
  assign n1299 = ~n1283 & n1298 ;
  assign n1300 = ~n1271 & n1299 ;
  assign n1301 = ~n1270 & n1300 ;
  assign n1302 = ~n1268 & n1301 ;
  assign n1303 = ~n1265 & n1302 ;
  assign n1344 = n1303 & x19 ;
  assign n1304 = ~x4 & ~n240 ;
  assign n1305 = n276 & n753 ;
  assign n1306 = x7 & ~n1305 ;
  assign n1307 = ~n1233 & ~n1306 ;
  assign n1308 = x7 & ~n240 ;
  assign n1309 = ~x0 & ~n1308 ;
  assign n1310 = ~x7 & ~n203 ;
  assign n1311 = x3 & ~n161 ;
  assign n1312 = ~x3 & ~n362 ;
  assign n1313 = n417 & ~n1312 ;
  assign n1314 = ~n1311 & ~n1313 ;
  assign n1315 = x2 & ~n1314 ;
  assign n1316 = ~n114 & n753 ;
  assign n1317 = x5 & n1316 ;
  assign n1318 = x6 & ~n259 ;
  assign n1319 = x3 & ~n1318 ;
  assign n1320 = ~n1317 & ~n1319 ;
  assign n1321 = ~n1315 & n1320 ;
  assign n1322 = ~x1 & ~n1321 ;
  assign n1323 = n417 & ~n763 ;
  assign n1324 = ~n362 & ~n1323 ;
  assign n1325 = ~x3 & ~n1324 ;
  assign n1326 = ~x4 & ~n123 ;
  assign n1327 = x3 & ~n1326 ;
  assign n1328 = ~n1325 & ~n1327 ;
  assign n1329 = x2 & ~n1328 ;
  assign n1330 = x8 & ~n46 ;
  assign n1331 = n1311 & ~n1330 ;
  assign n1332 = ~x2 & n1331 ;
  assign n1333 = ~n1329 & ~n1332 ;
  assign n1334 = x1 & ~n1333 ;
  assign n1335 = x5 & ~n203 ;
  assign n1336 = ~x6 & ~n1335 ;
  assign n1337 = ~n1334 & ~n1336 ;
  assign n1338 = ~n1322 & n1337 ;
  assign n1339 = ~n1310 & n1338 ;
  assign n1340 = ~n1309 & n1339 ;
  assign n1341 = ~n1307 & n1340 ;
  assign n1342 = ~n1304 & n1341 ;
  assign n1345 = ~n1342 & ~x19 ;
  assign n1346 = ~n1344 & ~n1345 ;
  assign n1347 = ~x8 & ~n18 ;
  assign n1348 = ~n14 & ~n1347 ;
  assign n1349 = n584 & ~n1348 ;
  assign n1350 = x2 & n1349 ;
  assign n1351 = ~n796 & ~n1350 ;
  assign n1352 = ~x7 & ~n1351 ;
  assign n1353 = n234 & n1352 ;
  assign n1362 = n1353 & x20 ;
  assign n1354 = x8 & ~n14 ;
  assign n1355 = ~n18 & ~n1354 ;
  assign n1356 = n494 & ~n1355 ;
  assign n1357 = ~x2 & n1356 ;
  assign n1358 = ~n801 & ~n1357 ;
  assign n1359 = x7 & ~n1358 ;
  assign n1360 = n123 & n1359 ;
  assign n1363 = ~n1360 & ~x20 ;
  assign n1364 = ~n1362 & ~n1363 ;
  assign y0 = ~n247 ;
  assign y1 = ~n458 ;
  assign y2 = ~n640 ;
  assign y3 = ~n778 ;
  assign y4 = ~n795 ;
  assign y5 = ~n809 ;
  assign y6 = ~n969 ;
  assign y7 = ~n1137 ;
  assign y8 = ~n1264 ;
  assign y9 = ~n1346 ;
  assign y10 = ~n1364 ;
endmodule
