module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 , y10320 , y10321 , y10322 , y10323 , y10324 , y10325 , y10326 , y10327 , y10328 , y10329 , y10330 , y10331 , y10332 , y10333 , y10334 , y10335 , y10336 , y10337 , y10338 , y10339 , y10340 , y10341 , y10342 , y10343 , y10344 , y10345 , y10346 , y10347 , y10348 , y10349 , y10350 , y10351 , y10352 , y10353 , y10354 , y10355 , y10356 , y10357 , y10358 , y10359 , y10360 , y10361 , y10362 , y10363 , y10364 , y10365 , y10366 , y10367 , y10368 , y10369 , y10370 , y10371 , y10372 , y10373 , y10374 , y10375 , y10376 , y10377 , y10378 , y10379 , y10380 , y10381 , y10382 , y10383 , y10384 , y10385 , y10386 , y10387 , y10388 , y10389 , y10390 , y10391 , y10392 , y10393 , y10394 , y10395 , y10396 , y10397 , y10398 , y10399 , y10400 , y10401 , y10402 , y10403 , y10404 , y10405 , y10406 , y10407 , y10408 , y10409 , y10410 , y10411 , y10412 , y10413 , y10414 , y10415 , y10416 , y10417 , y10418 , y10419 , y10420 , y10421 , y10422 , y10423 , y10424 , y10425 , y10426 , y10427 , y10428 , y10429 , y10430 , y10431 , y10432 , y10433 , y10434 , y10435 , y10436 , y10437 , y10438 , y10439 , y10440 , y10441 , y10442 , y10443 , y10444 , y10445 , y10446 , y10447 , y10448 , y10449 , y10450 , y10451 , y10452 , y10453 , y10454 , y10455 , y10456 , y10457 , y10458 , y10459 , y10460 , y10461 , y10462 , y10463 , y10464 , y10465 , y10466 , y10467 , y10468 , y10469 , y10470 , y10471 , y10472 , y10473 , y10474 , y10475 , y10476 , y10477 , y10478 , y10479 , y10480 , y10481 , y10482 , y10483 , y10484 , y10485 , y10486 , y10487 , y10488 , y10489 , y10490 , y10491 , y10492 , y10493 , y10494 , y10495 , y10496 , y10497 , y10498 , y10499 , y10500 , y10501 , y10502 , y10503 , y10504 , y10505 , y10506 , y10507 , y10508 , y10509 , y10510 , y10511 , y10512 , y10513 , y10514 , y10515 , y10516 , y10517 , y10518 , y10519 , y10520 , y10521 , y10522 , y10523 , y10524 , y10525 , y10526 , y10527 , y10528 , y10529 , y10530 , y10531 , y10532 , y10533 , y10534 , y10535 , y10536 , y10537 , y10538 , y10539 , y10540 , y10541 , y10542 , y10543 , y10544 , y10545 , y10546 , y10547 , y10548 , y10549 , y10550 , y10551 , y10552 , y10553 , y10554 , y10555 , y10556 , y10557 , y10558 , y10559 , y10560 , y10561 , y10562 , y10563 , y10564 , y10565 , y10566 , y10567 , y10568 , y10569 , y10570 , y10571 , y10572 , y10573 , y10574 , y10575 , y10576 , y10577 , y10578 , y10579 , y10580 , y10581 , y10582 , y10583 , y10584 , y10585 , y10586 , y10587 , y10588 , y10589 , y10590 , y10591 , y10592 , y10593 , y10594 , y10595 , y10596 , y10597 , y10598 , y10599 , y10600 , y10601 , y10602 , y10603 , y10604 , y10605 , y10606 , y10607 , y10608 , y10609 , y10610 , y10611 , y10612 , y10613 , y10614 , y10615 , y10616 , y10617 , y10618 , y10619 , y10620 , y10621 , y10622 , y10623 , y10624 , y10625 , y10626 , y10627 , y10628 , y10629 , y10630 , y10631 , y10632 , y10633 , y10634 , y10635 , y10636 , y10637 , y10638 , y10639 , y10640 , y10641 , y10642 , y10643 , y10644 , y10645 , y10646 , y10647 , y10648 , y10649 , y10650 , y10651 , y10652 , y10653 , y10654 , y10655 , y10656 , y10657 , y10658 , y10659 , y10660 , y10661 , y10662 , y10663 , y10664 , y10665 , y10666 , y10667 , y10668 , y10669 , y10670 , y10671 , y10672 , y10673 , y10674 , y10675 , y10676 , y10677 , y10678 , y10679 , y10680 , y10681 , y10682 , y10683 , y10684 , y10685 , y10686 , y10687 , y10688 , y10689 , y10690 , y10691 , y10692 , y10693 , y10694 , y10695 , y10696 , y10697 , y10698 , y10699 , y10700 , y10701 , y10702 , y10703 , y10704 , y10705 , y10706 , y10707 , y10708 , y10709 , y10710 , y10711 , y10712 , y10713 , y10714 , y10715 , y10716 , y10717 , y10718 , y10719 , y10720 , y10721 , y10722 , y10723 , y10724 , y10725 , y10726 , y10727 , y10728 , y10729 , y10730 , y10731 , y10732 , y10733 , y10734 , y10735 , y10736 , y10737 , y10738 , y10739 , y10740 , y10741 , y10742 , y10743 , y10744 , y10745 , y10746 , y10747 , y10748 , y10749 , y10750 , y10751 , y10752 , y10753 , y10754 , y10755 , y10756 , y10757 , y10758 , y10759 , y10760 , y10761 , y10762 , y10763 , y10764 , y10765 , y10766 , y10767 , y10768 , y10769 , y10770 , y10771 , y10772 , y10773 , y10774 , y10775 , y10776 , y10777 , y10778 , y10779 , y10780 , y10781 , y10782 , y10783 , y10784 , y10785 , y10786 , y10787 , y10788 , y10789 , y10790 , y10791 , y10792 , y10793 , y10794 , y10795 , y10796 , y10797 , y10798 , y10799 , y10800 , y10801 , y10802 , y10803 , y10804 , y10805 , y10806 , y10807 , y10808 , y10809 , y10810 , y10811 , y10812 , y10813 , y10814 , y10815 , y10816 , y10817 , y10818 , y10819 , y10820 , y10821 , y10822 , y10823 , y10824 , y10825 , y10826 , y10827 , y10828 , y10829 , y10830 , y10831 , y10832 , y10833 , y10834 , y10835 , y10836 , y10837 , y10838 , y10839 , y10840 , y10841 , y10842 , y10843 , y10844 , y10845 , y10846 , y10847 , y10848 , y10849 , y10850 , y10851 , y10852 , y10853 , y10854 , y10855 , y10856 , y10857 , y10858 , y10859 , y10860 , y10861 , y10862 , y10863 , y10864 , y10865 , y10866 , y10867 , y10868 , y10869 , y10870 , y10871 , y10872 , y10873 , y10874 , y10875 , y10876 , y10877 , y10878 , y10879 , y10880 , y10881 , y10882 , y10883 , y10884 , y10885 , y10886 , y10887 , y10888 , y10889 , y10890 , y10891 , y10892 , y10893 , y10894 , y10895 , y10896 , y10897 , y10898 , y10899 , y10900 , y10901 , y10902 , y10903 , y10904 , y10905 , y10906 , y10907 , y10908 , y10909 , y10910 , y10911 , y10912 , y10913 , y10914 , y10915 , y10916 , y10917 , y10918 , y10919 , y10920 , y10921 , y10922 , y10923 , y10924 , y10925 , y10926 , y10927 , y10928 , y10929 , y10930 , y10931 , y10932 , y10933 , y10934 , y10935 , y10936 , y10937 , y10938 , y10939 , y10940 , y10941 , y10942 , y10943 , y10944 , y10945 , y10946 , y10947 , y10948 , y10949 , y10950 , y10951 , y10952 , y10953 , y10954 , y10955 , y10956 , y10957 , y10958 , y10959 , y10960 , y10961 , y10962 , y10963 , y10964 , y10965 , y10966 , y10967 , y10968 , y10969 , y10970 , y10971 , y10972 , y10973 , y10974 , y10975 , y10976 , y10977 , y10978 , y10979 , y10980 , y10981 , y10982 , y10983 , y10984 , y10985 , y10986 , y10987 , y10988 , y10989 , y10990 , y10991 , y10992 , y10993 , y10994 , y10995 , y10996 , y10997 , y10998 , y10999 , y11000 , y11001 , y11002 , y11003 , y11004 , y11005 , y11006 , y11007 , y11008 , y11009 , y11010 , y11011 , y11012 , y11013 , y11014 , y11015 , y11016 , y11017 , y11018 , y11019 , y11020 , y11021 , y11022 , y11023 , y11024 , y11025 , y11026 , y11027 , y11028 , y11029 , y11030 , y11031 , y11032 , y11033 , y11034 , y11035 , y11036 , y11037 , y11038 , y11039 , y11040 , y11041 , y11042 , y11043 , y11044 , y11045 , y11046 , y11047 , y11048 , y11049 , y11050 , y11051 , y11052 , y11053 , y11054 , y11055 , y11056 , y11057 , y11058 , y11059 , y11060 , y11061 , y11062 , y11063 , y11064 , y11065 , y11066 , y11067 , y11068 , y11069 , y11070 , y11071 , y11072 , y11073 , y11074 , y11075 , y11076 , y11077 , y11078 , y11079 , y11080 , y11081 , y11082 , y11083 , y11084 , y11085 , y11086 , y11087 , y11088 , y11089 , y11090 , y11091 , y11092 , y11093 , y11094 , y11095 , y11096 , y11097 , y11098 , y11099 , y11100 , y11101 , y11102 , y11103 , y11104 , y11105 , y11106 , y11107 , y11108 , y11109 , y11110 , y11111 , y11112 , y11113 , y11114 , y11115 , y11116 , y11117 , y11118 , y11119 , y11120 , y11121 , y11122 , y11123 , y11124 , y11125 , y11126 , y11127 , y11128 , y11129 , y11130 , y11131 , y11132 , y11133 , y11134 , y11135 , y11136 , y11137 , y11138 , y11139 , y11140 , y11141 , y11142 , y11143 , y11144 , y11145 , y11146 , y11147 , y11148 , y11149 , y11150 , y11151 , y11152 , y11153 , y11154 , y11155 , y11156 , y11157 , y11158 , y11159 , y11160 , y11161 , y11162 , y11163 , y11164 , y11165 , y11166 , y11167 , y11168 , y11169 , y11170 , y11171 , y11172 , y11173 , y11174 , y11175 , y11176 , y11177 , y11178 , y11179 , y11180 , y11181 , y11182 , y11183 , y11184 , y11185 , y11186 , y11187 , y11188 , y11189 , y11190 , y11191 , y11192 , y11193 , y11194 , y11195 , y11196 , y11197 , y11198 , y11199 , y11200 , y11201 , y11202 , y11203 , y11204 , y11205 , y11206 , y11207 , y11208 , y11209 , y11210 , y11211 , y11212 , y11213 , y11214 , y11215 , y11216 , y11217 , y11218 , y11219 , y11220 , y11221 , y11222 , y11223 , y11224 , y11225 , y11226 , y11227 , y11228 , y11229 , y11230 , y11231 , y11232 , y11233 , y11234 , y11235 , y11236 , y11237 , y11238 , y11239 , y11240 , y11241 , y11242 , y11243 , y11244 , y11245 , y11246 , y11247 , y11248 , y11249 , y11250 , y11251 , y11252 , y11253 , y11254 , y11255 , y11256 , y11257 , y11258 , y11259 , y11260 , y11261 , y11262 , y11263 , y11264 , y11265 , y11266 , y11267 , y11268 , y11269 , y11270 , y11271 , y11272 , y11273 , y11274 , y11275 , y11276 , y11277 , y11278 , y11279 , y11280 , y11281 , y11282 , y11283 , y11284 , y11285 , y11286 , y11287 , y11288 , y11289 , y11290 , y11291 , y11292 , y11293 , y11294 , y11295 , y11296 , y11297 , y11298 , y11299 , y11300 , y11301 , y11302 , y11303 , y11304 , y11305 , y11306 , y11307 , y11308 , y11309 , y11310 , y11311 , y11312 , y11313 , y11314 , y11315 , y11316 , y11317 , y11318 , y11319 , y11320 , y11321 , y11322 , y11323 , y11324 , y11325 , y11326 , y11327 , y11328 , y11329 , y11330 , y11331 , y11332 , y11333 , y11334 , y11335 , y11336 , y11337 , y11338 , y11339 , y11340 , y11341 , y11342 , y11343 , y11344 , y11345 , y11346 , y11347 , y11348 , y11349 , y11350 , y11351 , y11352 , y11353 , y11354 , y11355 , y11356 , y11357 , y11358 , y11359 , y11360 , y11361 , y11362 , y11363 , y11364 , y11365 , y11366 , y11367 , y11368 , y11369 , y11370 , y11371 , y11372 , y11373 , y11374 , y11375 , y11376 , y11377 , y11378 , y11379 , y11380 , y11381 , y11382 , y11383 , y11384 , y11385 , y11386 , y11387 , y11388 , y11389 , y11390 , y11391 , y11392 , y11393 , y11394 , y11395 , y11396 , y11397 , y11398 , y11399 , y11400 , y11401 , y11402 , y11403 , y11404 , y11405 , y11406 , y11407 , y11408 , y11409 , y11410 , y11411 , y11412 , y11413 , y11414 , y11415 , y11416 , y11417 , y11418 , y11419 , y11420 , y11421 , y11422 , y11423 , y11424 , y11425 , y11426 , y11427 , y11428 , y11429 , y11430 , y11431 , y11432 , y11433 , y11434 , y11435 , y11436 , y11437 , y11438 , y11439 , y11440 , y11441 , y11442 , y11443 , y11444 , y11445 , y11446 , y11447 , y11448 , y11449 , y11450 , y11451 , y11452 , y11453 , y11454 , y11455 , y11456 , y11457 , y11458 , y11459 , y11460 , y11461 , y11462 , y11463 , y11464 , y11465 , y11466 , y11467 , y11468 , y11469 , y11470 , y11471 , y11472 , y11473 , y11474 , y11475 , y11476 , y11477 , y11478 , y11479 , y11480 , y11481 , y11482 , y11483 , y11484 , y11485 , y11486 , y11487 , y11488 , y11489 , y11490 , y11491 , y11492 , y11493 , y11494 , y11495 , y11496 , y11497 , y11498 , y11499 , y11500 , y11501 , y11502 , y11503 , y11504 , y11505 , y11506 , y11507 , y11508 , y11509 , y11510 , y11511 , y11512 , y11513 , y11514 , y11515 , y11516 , y11517 , y11518 , y11519 , y11520 , y11521 , y11522 , y11523 , y11524 , y11525 , y11526 , y11527 , y11528 , y11529 , y11530 , y11531 , y11532 , y11533 , y11534 , y11535 , y11536 , y11537 , y11538 , y11539 , y11540 , y11541 , y11542 , y11543 , y11544 , y11545 , y11546 , y11547 , y11548 , y11549 , y11550 , y11551 , y11552 , y11553 , y11554 , y11555 , y11556 , y11557 , y11558 , y11559 , y11560 , y11561 , y11562 , y11563 , y11564 , y11565 , y11566 , y11567 , y11568 , y11569 , y11570 , y11571 , y11572 , y11573 , y11574 , y11575 , y11576 , y11577 , y11578 , y11579 , y11580 , y11581 , y11582 , y11583 , y11584 , y11585 , y11586 , y11587 , y11588 , y11589 , y11590 , y11591 , y11592 , y11593 , y11594 , y11595 , y11596 , y11597 , y11598 , y11599 , y11600 , y11601 , y11602 , y11603 , y11604 , y11605 , y11606 , y11607 , y11608 , y11609 , y11610 , y11611 , y11612 , y11613 , y11614 , y11615 , y11616 , y11617 , y11618 , y11619 , y11620 , y11621 , y11622 , y11623 , y11624 , y11625 , y11626 , y11627 , y11628 , y11629 , y11630 , y11631 , y11632 , y11633 , y11634 , y11635 , y11636 , y11637 , y11638 , y11639 , y11640 , y11641 , y11642 , y11643 , y11644 , y11645 , y11646 , y11647 , y11648 , y11649 , y11650 , y11651 , y11652 , y11653 , y11654 , y11655 , y11656 , y11657 , y11658 , y11659 , y11660 , y11661 , y11662 , y11663 , y11664 , y11665 , y11666 , y11667 , y11668 , y11669 , y11670 , y11671 , y11672 , y11673 , y11674 , y11675 , y11676 , y11677 , y11678 , y11679 , y11680 , y11681 , y11682 , y11683 , y11684 , y11685 , y11686 , y11687 , y11688 , y11689 , y11690 , y11691 , y11692 , y11693 , y11694 , y11695 , y11696 , y11697 , y11698 , y11699 , y11700 , y11701 , y11702 , y11703 , y11704 , y11705 , y11706 , y11707 , y11708 , y11709 , y11710 , y11711 , y11712 , y11713 , y11714 , y11715 , y11716 , y11717 , y11718 , y11719 , y11720 , y11721 , y11722 , y11723 , y11724 , y11725 , y11726 , y11727 , y11728 , y11729 , y11730 , y11731 , y11732 , y11733 , y11734 , y11735 , y11736 , y11737 , y11738 , y11739 , y11740 , y11741 , y11742 , y11743 , y11744 , y11745 , y11746 , y11747 , y11748 , y11749 , y11750 , y11751 , y11752 , y11753 , y11754 , y11755 , y11756 , y11757 , y11758 , y11759 , y11760 , y11761 , y11762 , y11763 , y11764 , y11765 , y11766 , y11767 , y11768 , y11769 , y11770 , y11771 , y11772 , y11773 , y11774 , y11775 , y11776 , y11777 , y11778 , y11779 , y11780 , y11781 , y11782 , y11783 , y11784 , y11785 , y11786 , y11787 , y11788 , y11789 , y11790 , y11791 , y11792 , y11793 , y11794 , y11795 , y11796 , y11797 , y11798 , y11799 , y11800 , y11801 , y11802 , y11803 , y11804 , y11805 , y11806 , y11807 , y11808 , y11809 , y11810 , y11811 , y11812 , y11813 , y11814 , y11815 , y11816 , y11817 , y11818 , y11819 , y11820 , y11821 , y11822 , y11823 , y11824 , y11825 , y11826 , y11827 , y11828 , y11829 , y11830 , y11831 , y11832 , y11833 , y11834 , y11835 , y11836 , y11837 , y11838 , y11839 , y11840 , y11841 , y11842 , y11843 , y11844 , y11845 , y11846 , y11847 , y11848 , y11849 , y11850 , y11851 , y11852 , y11853 , y11854 , y11855 , y11856 , y11857 , y11858 , y11859 , y11860 , y11861 , y11862 , y11863 , y11864 , y11865 , y11866 , y11867 , y11868 , y11869 , y11870 , y11871 , y11872 , y11873 , y11874 , y11875 , y11876 , y11877 , y11878 , y11879 , y11880 , y11881 , y11882 , y11883 , y11884 , y11885 , y11886 , y11887 , y11888 , y11889 , y11890 , y11891 , y11892 , y11893 , y11894 , y11895 , y11896 , y11897 , y11898 , y11899 , y11900 , y11901 , y11902 , y11903 , y11904 , y11905 , y11906 , y11907 , y11908 , y11909 , y11910 , y11911 , y11912 , y11913 , y11914 , y11915 , y11916 , y11917 , y11918 , y11919 , y11920 , y11921 , y11922 , y11923 , y11924 , y11925 , y11926 , y11927 , y11928 , y11929 , y11930 , y11931 , y11932 , y11933 , y11934 , y11935 , y11936 , y11937 , y11938 , y11939 , y11940 , y11941 , y11942 , y11943 , y11944 , y11945 , y11946 , y11947 , y11948 , y11949 , y11950 , y11951 , y11952 , y11953 , y11954 , y11955 , y11956 , y11957 , y11958 , y11959 , y11960 , y11961 , y11962 , y11963 , y11964 , y11965 , y11966 , y11967 , y11968 , y11969 , y11970 , y11971 , y11972 , y11973 , y11974 , y11975 , y11976 , y11977 , y11978 , y11979 , y11980 , y11981 , y11982 , y11983 , y11984 , y11985 , y11986 , y11987 , y11988 , y11989 , y11990 , y11991 , y11992 , y11993 , y11994 , y11995 , y11996 , y11997 , y11998 , y11999 , y12000 , y12001 , y12002 , y12003 , y12004 , y12005 , y12006 , y12007 , y12008 , y12009 , y12010 , y12011 , y12012 , y12013 , y12014 , y12015 , y12016 , y12017 , y12018 , y12019 , y12020 , y12021 , y12022 , y12023 , y12024 , y12025 , y12026 , y12027 , y12028 , y12029 , y12030 , y12031 , y12032 , y12033 , y12034 , y12035 , y12036 , y12037 , y12038 , y12039 , y12040 , y12041 , y12042 , y12043 , y12044 , y12045 , y12046 , y12047 , y12048 , y12049 , y12050 , y12051 , y12052 , y12053 , y12054 , y12055 , y12056 , y12057 , y12058 , y12059 , y12060 , y12061 , y12062 , y12063 , y12064 , y12065 , y12066 , y12067 , y12068 , y12069 , y12070 , y12071 , y12072 , y12073 , y12074 , y12075 , y12076 , y12077 , y12078 , y12079 , y12080 , y12081 , y12082 , y12083 , y12084 , y12085 , y12086 , y12087 , y12088 , y12089 , y12090 , y12091 , y12092 , y12093 , y12094 , y12095 , y12096 , y12097 , y12098 , y12099 , y12100 , y12101 , y12102 , y12103 , y12104 , y12105 , y12106 , y12107 , y12108 , y12109 , y12110 , y12111 , y12112 , y12113 , y12114 , y12115 , y12116 , y12117 , y12118 , y12119 , y12120 , y12121 , y12122 , y12123 , y12124 , y12125 , y12126 , y12127 , y12128 , y12129 , y12130 , y12131 , y12132 , y12133 , y12134 , y12135 , y12136 , y12137 , y12138 , y12139 , y12140 , y12141 , y12142 , y12143 , y12144 , y12145 , y12146 , y12147 , y12148 , y12149 , y12150 , y12151 , y12152 , y12153 , y12154 , y12155 , y12156 , y12157 , y12158 , y12159 , y12160 , y12161 , y12162 , y12163 , y12164 , y12165 , y12166 , y12167 , y12168 , y12169 , y12170 , y12171 , y12172 , y12173 , y12174 , y12175 , y12176 , y12177 , y12178 , y12179 , y12180 , y12181 , y12182 , y12183 , y12184 , y12185 , y12186 , y12187 , y12188 , y12189 , y12190 , y12191 , y12192 , y12193 , y12194 , y12195 , y12196 , y12197 , y12198 , y12199 , y12200 , y12201 , y12202 , y12203 , y12204 , y12205 , y12206 , y12207 , y12208 , y12209 , y12210 , y12211 , y12212 , y12213 , y12214 , y12215 , y12216 , y12217 , y12218 , y12219 , y12220 , y12221 , y12222 , y12223 , y12224 , y12225 , y12226 , y12227 , y12228 , y12229 , y12230 , y12231 , y12232 , y12233 , y12234 , y12235 , y12236 , y12237 , y12238 , y12239 , y12240 , y12241 , y12242 , y12243 , y12244 , y12245 , y12246 , y12247 , y12248 , y12249 , y12250 , y12251 , y12252 , y12253 , y12254 , y12255 , y12256 , y12257 , y12258 , y12259 , y12260 , y12261 , y12262 , y12263 , y12264 , y12265 , y12266 , y12267 , y12268 , y12269 , y12270 , y12271 , y12272 , y12273 , y12274 , y12275 , y12276 , y12277 , y12278 , y12279 , y12280 , y12281 , y12282 , y12283 , y12284 , y12285 , y12286 , y12287 , y12288 , y12289 , y12290 , y12291 , y12292 , y12293 , y12294 , y12295 , y12296 , y12297 , y12298 , y12299 , y12300 , y12301 , y12302 , y12303 , y12304 , y12305 , y12306 , y12307 , y12308 , y12309 , y12310 , y12311 , y12312 , y12313 , y12314 , y12315 , y12316 , y12317 , y12318 , y12319 , y12320 , y12321 , y12322 , y12323 , y12324 , y12325 , y12326 , y12327 , y12328 , y12329 , y12330 , y12331 , y12332 , y12333 , y12334 , y12335 , y12336 , y12337 , y12338 , y12339 , y12340 , y12341 , y12342 , y12343 , y12344 , y12345 , y12346 , y12347 , y12348 , y12349 , y12350 , y12351 , y12352 , y12353 , y12354 , y12355 , y12356 , y12357 , y12358 , y12359 , y12360 , y12361 , y12362 , y12363 , y12364 , y12365 , y12366 , y12367 , y12368 , y12369 , y12370 , y12371 , y12372 , y12373 , y12374 , y12375 , y12376 , y12377 , y12378 , y12379 , y12380 , y12381 , y12382 , y12383 , y12384 , y12385 , y12386 , y12387 , y12388 , y12389 , y12390 , y12391 , y12392 , y12393 , y12394 , y12395 , y12396 , y12397 , y12398 , y12399 , y12400 , y12401 , y12402 , y12403 , y12404 , y12405 , y12406 , y12407 , y12408 , y12409 , y12410 , y12411 , y12412 , y12413 , y12414 , y12415 , y12416 , y12417 , y12418 , y12419 , y12420 , y12421 , y12422 , y12423 , y12424 , y12425 , y12426 , y12427 , y12428 , y12429 , y12430 , y12431 , y12432 , y12433 , y12434 , y12435 , y12436 , y12437 , y12438 , y12439 , y12440 , y12441 , y12442 , y12443 , y12444 , y12445 , y12446 , y12447 , y12448 , y12449 , y12450 , y12451 , y12452 , y12453 , y12454 , y12455 , y12456 , y12457 , y12458 , y12459 , y12460 , y12461 , y12462 , y12463 , y12464 , y12465 , y12466 , y12467 , y12468 , y12469 , y12470 , y12471 , y12472 , y12473 , y12474 , y12475 , y12476 , y12477 , y12478 , y12479 , y12480 , y12481 , y12482 , y12483 , y12484 , y12485 , y12486 , y12487 , y12488 , y12489 , y12490 , y12491 , y12492 , y12493 , y12494 , y12495 , y12496 , y12497 , y12498 , y12499 , y12500 , y12501 , y12502 , y12503 , y12504 , y12505 , y12506 , y12507 , y12508 , y12509 , y12510 , y12511 , y12512 , y12513 , y12514 , y12515 , y12516 , y12517 , y12518 , y12519 , y12520 , y12521 , y12522 , y12523 , y12524 , y12525 , y12526 , y12527 , y12528 , y12529 , y12530 , y12531 , y12532 , y12533 , y12534 , y12535 , y12536 , y12537 , y12538 , y12539 , y12540 , y12541 , y12542 , y12543 , y12544 , y12545 , y12546 , y12547 , y12548 , y12549 , y12550 , y12551 , y12552 , y12553 , y12554 , y12555 , y12556 , y12557 , y12558 , y12559 , y12560 , y12561 , y12562 , y12563 , y12564 , y12565 , y12566 , y12567 , y12568 , y12569 , y12570 , y12571 , y12572 , y12573 , y12574 , y12575 , y12576 , y12577 , y12578 , y12579 , y12580 , y12581 , y12582 , y12583 , y12584 , y12585 , y12586 , y12587 , y12588 , y12589 , y12590 , y12591 , y12592 , y12593 , y12594 , y12595 , y12596 , y12597 , y12598 , y12599 , y12600 , y12601 , y12602 , y12603 , y12604 , y12605 , y12606 , y12607 , y12608 , y12609 , y12610 , y12611 , y12612 , y12613 , y12614 , y12615 , y12616 , y12617 , y12618 , y12619 , y12620 , y12621 , y12622 , y12623 , y12624 , y12625 , y12626 , y12627 , y12628 , y12629 , y12630 , y12631 , y12632 , y12633 , y12634 , y12635 , y12636 , y12637 , y12638 , y12639 , y12640 , y12641 , y12642 , y12643 , y12644 , y12645 , y12646 , y12647 , y12648 , y12649 , y12650 , y12651 , y12652 , y12653 , y12654 , y12655 , y12656 , y12657 , y12658 , y12659 , y12660 , y12661 , y12662 , y12663 , y12664 , y12665 , y12666 , y12667 , y12668 , y12669 , y12670 , y12671 , y12672 , y12673 , y12674 , y12675 , y12676 , y12677 , y12678 , y12679 , y12680 , y12681 , y12682 , y12683 , y12684 , y12685 , y12686 , y12687 , y12688 , y12689 , y12690 , y12691 , y12692 , y12693 , y12694 , y12695 , y12696 , y12697 , y12698 , y12699 , y12700 , y12701 , y12702 , y12703 , y12704 , y12705 , y12706 , y12707 , y12708 , y12709 , y12710 , y12711 , y12712 , y12713 , y12714 , y12715 , y12716 , y12717 , y12718 , y12719 , y12720 , y12721 , y12722 , y12723 , y12724 , y12725 , y12726 , y12727 , y12728 , y12729 , y12730 , y12731 , y12732 , y12733 , y12734 , y12735 , y12736 , y12737 , y12738 , y12739 , y12740 , y12741 , y12742 , y12743 , y12744 , y12745 , y12746 , y12747 , y12748 , y12749 , y12750 , y12751 , y12752 , y12753 , y12754 , y12755 , y12756 , y12757 , y12758 , y12759 , y12760 , y12761 , y12762 , y12763 , y12764 , y12765 , y12766 , y12767 , y12768 , y12769 , y12770 , y12771 , y12772 , y12773 , y12774 , y12775 , y12776 , y12777 , y12778 , y12779 , y12780 , y12781 , y12782 , y12783 , y12784 , y12785 , y12786 , y12787 , y12788 , y12789 , y12790 , y12791 , y12792 , y12793 , y12794 , y12795 , y12796 , y12797 , y12798 , y12799 , y12800 , y12801 , y12802 , y12803 , y12804 , y12805 , y12806 , y12807 , y12808 , y12809 , y12810 , y12811 , y12812 , y12813 , y12814 , y12815 , y12816 , y12817 , y12818 , y12819 , y12820 , y12821 , y12822 , y12823 , y12824 , y12825 , y12826 , y12827 , y12828 , y12829 , y12830 , y12831 , y12832 , y12833 , y12834 , y12835 , y12836 , y12837 , y12838 , y12839 , y12840 , y12841 , y12842 , y12843 , y12844 , y12845 , y12846 , y12847 , y12848 , y12849 , y12850 , y12851 , y12852 , y12853 , y12854 , y12855 , y12856 , y12857 , y12858 , y12859 , y12860 , y12861 , y12862 , y12863 , y12864 , y12865 , y12866 , y12867 , y12868 , y12869 , y12870 , y12871 , y12872 , y12873 , y12874 , y12875 , y12876 , y12877 , y12878 , y12879 , y12880 , y12881 , y12882 , y12883 , y12884 , y12885 , y12886 , y12887 , y12888 , y12889 , y12890 , y12891 , y12892 , y12893 , y12894 , y12895 , y12896 , y12897 , y12898 , y12899 , y12900 , y12901 , y12902 , y12903 , y12904 , y12905 , y12906 , y12907 , y12908 , y12909 , y12910 , y12911 , y12912 , y12913 , y12914 , y12915 , y12916 , y12917 , y12918 , y12919 , y12920 , y12921 , y12922 , y12923 , y12924 , y12925 , y12926 , y12927 , y12928 , y12929 , y12930 , y12931 , y12932 , y12933 , y12934 , y12935 , y12936 , y12937 , y12938 , y12939 , y12940 , y12941 , y12942 , y12943 , y12944 , y12945 , y12946 , y12947 , y12948 , y12949 , y12950 , y12951 , y12952 , y12953 , y12954 , y12955 , y12956 , y12957 , y12958 , y12959 , y12960 , y12961 , y12962 , y12963 , y12964 , y12965 , y12966 , y12967 , y12968 , y12969 , y12970 , y12971 , y12972 , y12973 , y12974 , y12975 , y12976 , y12977 , y12978 , y12979 , y12980 , y12981 , y12982 , y12983 , y12984 , y12985 , y12986 , y12987 , y12988 , y12989 , y12990 , y12991 , y12992 , y12993 , y12994 , y12995 , y12996 , y12997 , y12998 , y12999 , y13000 , y13001 , y13002 , y13003 , y13004 , y13005 , y13006 , y13007 , y13008 , y13009 , y13010 , y13011 , y13012 , y13013 , y13014 , y13015 , y13016 , y13017 , y13018 , y13019 , y13020 , y13021 , y13022 , y13023 , y13024 , y13025 , y13026 , y13027 , y13028 , y13029 , y13030 , y13031 , y13032 , y13033 , y13034 , y13035 , y13036 , y13037 , y13038 , y13039 , y13040 , y13041 , y13042 , y13043 , y13044 , y13045 , y13046 , y13047 , y13048 , y13049 , y13050 , y13051 , y13052 , y13053 , y13054 , y13055 , y13056 , y13057 , y13058 , y13059 , y13060 , y13061 , y13062 , y13063 , y13064 , y13065 , y13066 , y13067 , y13068 , y13069 , y13070 , y13071 , y13072 , y13073 , y13074 , y13075 , y13076 , y13077 , y13078 , y13079 , y13080 , y13081 , y13082 , y13083 , y13084 , y13085 , y13086 , y13087 , y13088 , y13089 , y13090 , y13091 , y13092 , y13093 , y13094 , y13095 , y13096 , y13097 , y13098 , y13099 , y13100 , y13101 , y13102 , y13103 , y13104 , y13105 , y13106 , y13107 , y13108 , y13109 , y13110 , y13111 , y13112 , y13113 , y13114 , y13115 , y13116 , y13117 , y13118 , y13119 , y13120 , y13121 , y13122 , y13123 , y13124 , y13125 , y13126 , y13127 , y13128 , y13129 , y13130 , y13131 , y13132 , y13133 , y13134 , y13135 , y13136 , y13137 , y13138 , y13139 , y13140 , y13141 , y13142 , y13143 , y13144 , y13145 , y13146 , y13147 , y13148 , y13149 , y13150 , y13151 , y13152 , y13153 , y13154 , y13155 , y13156 , y13157 , y13158 , y13159 , y13160 , y13161 , y13162 , y13163 , y13164 , y13165 , y13166 , y13167 , y13168 , y13169 , y13170 , y13171 , y13172 , y13173 , y13174 , y13175 , y13176 , y13177 , y13178 , y13179 , y13180 , y13181 , y13182 , y13183 , y13184 , y13185 , y13186 , y13187 , y13188 , y13189 , y13190 , y13191 , y13192 , y13193 , y13194 , y13195 , y13196 , y13197 , y13198 , y13199 , y13200 , y13201 , y13202 , y13203 , y13204 , y13205 , y13206 , y13207 , y13208 , y13209 , y13210 , y13211 , y13212 , y13213 , y13214 , y13215 , y13216 , y13217 , y13218 , y13219 , y13220 , y13221 , y13222 , y13223 , y13224 , y13225 , y13226 , y13227 , y13228 , y13229 , y13230 , y13231 , y13232 , y13233 , y13234 , y13235 , y13236 , y13237 , y13238 , y13239 , y13240 , y13241 , y13242 , y13243 , y13244 , y13245 , y13246 , y13247 , y13248 , y13249 , y13250 , y13251 , y13252 , y13253 , y13254 , y13255 , y13256 , y13257 , y13258 , y13259 , y13260 , y13261 , y13262 , y13263 , y13264 , y13265 , y13266 , y13267 , y13268 , y13269 , y13270 , y13271 , y13272 , y13273 , y13274 , y13275 , y13276 , y13277 , y13278 , y13279 , y13280 , y13281 , y13282 , y13283 , y13284 , y13285 , y13286 , y13287 , y13288 , y13289 , y13290 , y13291 , y13292 , y13293 , y13294 , y13295 , y13296 , y13297 , y13298 , y13299 , y13300 , y13301 , y13302 , y13303 , y13304 , y13305 , y13306 , y13307 , y13308 , y13309 , y13310 , y13311 , y13312 , y13313 , y13314 , y13315 , y13316 , y13317 , y13318 , y13319 , y13320 , y13321 , y13322 , y13323 , y13324 , y13325 , y13326 , y13327 , y13328 , y13329 , y13330 , y13331 , y13332 , y13333 , y13334 , y13335 , y13336 , y13337 , y13338 , y13339 , y13340 , y13341 , y13342 , y13343 , y13344 , y13345 , y13346 , y13347 , y13348 , y13349 , y13350 , y13351 , y13352 , y13353 , y13354 , y13355 , y13356 , y13357 , y13358 , y13359 , y13360 , y13361 , y13362 , y13363 , y13364 , y13365 , y13366 , y13367 , y13368 , y13369 , y13370 , y13371 , y13372 , y13373 , y13374 , y13375 , y13376 , y13377 , y13378 , y13379 , y13380 , y13381 , y13382 , y13383 , y13384 , y13385 , y13386 , y13387 , y13388 , y13389 , y13390 , y13391 , y13392 , y13393 , y13394 , y13395 , y13396 , y13397 , y13398 , y13399 , y13400 , y13401 , y13402 , y13403 , y13404 , y13405 , y13406 , y13407 , y13408 , y13409 , y13410 , y13411 , y13412 , y13413 , y13414 , y13415 , y13416 , y13417 , y13418 , y13419 , y13420 , y13421 , y13422 , y13423 , y13424 , y13425 , y13426 , y13427 , y13428 , y13429 , y13430 , y13431 , y13432 , y13433 , y13434 , y13435 , y13436 , y13437 , y13438 , y13439 , y13440 , y13441 , y13442 , y13443 , y13444 , y13445 , y13446 , y13447 , y13448 , y13449 , y13450 , y13451 , y13452 , y13453 , y13454 , y13455 , y13456 , y13457 , y13458 , y13459 , y13460 , y13461 , y13462 , y13463 , y13464 , y13465 , y13466 , y13467 , y13468 , y13469 , y13470 , y13471 , y13472 , y13473 , y13474 , y13475 , y13476 , y13477 , y13478 , y13479 , y13480 , y13481 , y13482 , y13483 , y13484 , y13485 , y13486 , y13487 , y13488 , y13489 , y13490 , y13491 , y13492 , y13493 , y13494 , y13495 , y13496 , y13497 , y13498 , y13499 , y13500 , y13501 , y13502 , y13503 , y13504 , y13505 , y13506 , y13507 , y13508 , y13509 , y13510 , y13511 , y13512 , y13513 , y13514 , y13515 , y13516 , y13517 , y13518 , y13519 , y13520 , y13521 , y13522 , y13523 , y13524 , y13525 , y13526 , y13527 , y13528 , y13529 , y13530 , y13531 , y13532 , y13533 , y13534 , y13535 , y13536 , y13537 , y13538 , y13539 , y13540 , y13541 , y13542 , y13543 , y13544 , y13545 , y13546 , y13547 , y13548 , y13549 , y13550 , y13551 , y13552 , y13553 , y13554 , y13555 , y13556 , y13557 , y13558 , y13559 , y13560 , y13561 , y13562 , y13563 , y13564 , y13565 , y13566 , y13567 , y13568 , y13569 , y13570 , y13571 , y13572 , y13573 , y13574 , y13575 , y13576 , y13577 , y13578 , y13579 , y13580 , y13581 , y13582 , y13583 , y13584 , y13585 , y13586 , y13587 , y13588 , y13589 , y13590 , y13591 , y13592 , y13593 , y13594 , y13595 , y13596 , y13597 , y13598 , y13599 , y13600 , y13601 , y13602 , y13603 , y13604 , y13605 , y13606 , y13607 , y13608 , y13609 , y13610 , y13611 , y13612 , y13613 , y13614 , y13615 , y13616 , y13617 , y13618 , y13619 , y13620 , y13621 , y13622 , y13623 , y13624 , y13625 , y13626 , y13627 , y13628 , y13629 , y13630 , y13631 , y13632 , y13633 , y13634 , y13635 , y13636 , y13637 , y13638 , y13639 , y13640 , y13641 , y13642 , y13643 , y13644 , y13645 , y13646 , y13647 , y13648 , y13649 , y13650 , y13651 , y13652 , y13653 , y13654 , y13655 , y13656 , y13657 , y13658 , y13659 , y13660 , y13661 , y13662 , y13663 , y13664 , y13665 , y13666 , y13667 , y13668 , y13669 , y13670 , y13671 , y13672 , y13673 , y13674 , y13675 , y13676 , y13677 , y13678 , y13679 , y13680 , y13681 , y13682 , y13683 , y13684 , y13685 , y13686 , y13687 , y13688 , y13689 , y13690 , y13691 , y13692 , y13693 , y13694 , y13695 , y13696 , y13697 , y13698 , y13699 , y13700 , y13701 , y13702 , y13703 , y13704 , y13705 , y13706 , y13707 , y13708 , y13709 , y13710 , y13711 , y13712 , y13713 , y13714 , y13715 , y13716 , y13717 , y13718 , y13719 , y13720 , y13721 , y13722 , y13723 , y13724 , y13725 , y13726 , y13727 , y13728 , y13729 , y13730 , y13731 , y13732 , y13733 , y13734 , y13735 , y13736 , y13737 , y13738 , y13739 , y13740 , y13741 , y13742 , y13743 , y13744 , y13745 , y13746 , y13747 , y13748 , y13749 , y13750 , y13751 , y13752 , y13753 , y13754 , y13755 , y13756 , y13757 , y13758 , y13759 , y13760 , y13761 , y13762 , y13763 , y13764 , y13765 , y13766 , y13767 , y13768 , y13769 , y13770 , y13771 , y13772 , y13773 , y13774 , y13775 , y13776 , y13777 , y13778 , y13779 , y13780 , y13781 , y13782 , y13783 , y13784 , y13785 , y13786 , y13787 , y13788 , y13789 , y13790 , y13791 , y13792 , y13793 , y13794 , y13795 , y13796 , y13797 , y13798 , y13799 , y13800 , y13801 , y13802 , y13803 , y13804 , y13805 , y13806 , y13807 , y13808 , y13809 , y13810 , y13811 , y13812 , y13813 , y13814 , y13815 , y13816 , y13817 , y13818 , y13819 , y13820 , y13821 , y13822 , y13823 , y13824 , y13825 , y13826 , y13827 , y13828 , y13829 , y13830 , y13831 , y13832 , y13833 , y13834 , y13835 , y13836 , y13837 , y13838 , y13839 , y13840 , y13841 , y13842 , y13843 , y13844 , y13845 , y13846 , y13847 , y13848 , y13849 , y13850 , y13851 , y13852 , y13853 , y13854 , y13855 , y13856 , y13857 , y13858 , y13859 , y13860 , y13861 , y13862 , y13863 , y13864 , y13865 , y13866 , y13867 , y13868 , y13869 , y13870 , y13871 , y13872 , y13873 , y13874 , y13875 , y13876 , y13877 , y13878 , y13879 , y13880 , y13881 , y13882 , y13883 , y13884 , y13885 , y13886 , y13887 , y13888 , y13889 , y13890 , y13891 , y13892 , y13893 , y13894 , y13895 , y13896 , y13897 , y13898 , y13899 , y13900 , y13901 , y13902 , y13903 , y13904 , y13905 , y13906 , y13907 , y13908 , y13909 , y13910 , y13911 , y13912 , y13913 , y13914 , y13915 , y13916 , y13917 , y13918 , y13919 , y13920 , y13921 , y13922 , y13923 , y13924 , y13925 , y13926 , y13927 , y13928 , y13929 , y13930 , y13931 , y13932 , y13933 , y13934 , y13935 , y13936 , y13937 , y13938 , y13939 , y13940 , y13941 , y13942 , y13943 , y13944 , y13945 , y13946 , y13947 , y13948 , y13949 , y13950 , y13951 , y13952 , y13953 , y13954 , y13955 , y13956 , y13957 , y13958 , y13959 , y13960 , y13961 , y13962 , y13963 , y13964 , y13965 , y13966 , y13967 , y13968 , y13969 , y13970 , y13971 , y13972 , y13973 , y13974 , y13975 , y13976 , y13977 , y13978 , y13979 , y13980 , y13981 , y13982 , y13983 , y13984 , y13985 , y13986 , y13987 , y13988 , y13989 , y13990 , y13991 , y13992 , y13993 , y13994 , y13995 , y13996 , y13997 , y13998 , y13999 , y14000 , y14001 , y14002 , y14003 , y14004 , y14005 , y14006 , y14007 , y14008 , y14009 , y14010 , y14011 , y14012 , y14013 , y14014 , y14015 , y14016 , y14017 , y14018 , y14019 , y14020 , y14021 , y14022 , y14023 , y14024 , y14025 , y14026 , y14027 , y14028 , y14029 , y14030 , y14031 , y14032 , y14033 , y14034 , y14035 , y14036 , y14037 , y14038 , y14039 , y14040 , y14041 , y14042 , y14043 , y14044 , y14045 , y14046 , y14047 , y14048 , y14049 , y14050 , y14051 , y14052 , y14053 , y14054 , y14055 , y14056 , y14057 , y14058 , y14059 , y14060 , y14061 , y14062 , y14063 , y14064 , y14065 , y14066 , y14067 , y14068 , y14069 , y14070 , y14071 , y14072 , y14073 , y14074 , y14075 , y14076 , y14077 , y14078 , y14079 , y14080 , y14081 , y14082 , y14083 , y14084 , y14085 , y14086 , y14087 , y14088 , y14089 , y14090 , y14091 , y14092 , y14093 , y14094 , y14095 , y14096 , y14097 , y14098 , y14099 , y14100 , y14101 , y14102 , y14103 , y14104 , y14105 , y14106 , y14107 , y14108 , y14109 , y14110 , y14111 , y14112 , y14113 , y14114 , y14115 , y14116 , y14117 , y14118 , y14119 , y14120 , y14121 , y14122 , y14123 , y14124 , y14125 , y14126 , y14127 , y14128 , y14129 , y14130 , y14131 , y14132 , y14133 , y14134 , y14135 , y14136 , y14137 , y14138 , y14139 , y14140 , y14141 , y14142 , y14143 , y14144 , y14145 , y14146 , y14147 , y14148 , y14149 , y14150 , y14151 , y14152 , y14153 , y14154 , y14155 , y14156 , y14157 , y14158 , y14159 , y14160 , y14161 , y14162 , y14163 , y14164 , y14165 , y14166 , y14167 , y14168 , y14169 , y14170 , y14171 , y14172 , y14173 , y14174 , y14175 , y14176 , y14177 , y14178 , y14179 , y14180 , y14181 , y14182 , y14183 , y14184 , y14185 , y14186 , y14187 , y14188 , y14189 , y14190 , y14191 , y14192 , y14193 , y14194 , y14195 , y14196 , y14197 , y14198 , y14199 , y14200 , y14201 , y14202 , y14203 , y14204 , y14205 , y14206 , y14207 , y14208 , y14209 , y14210 , y14211 , y14212 , y14213 , y14214 , y14215 , y14216 , y14217 , y14218 , y14219 , y14220 , y14221 , y14222 , y14223 , y14224 , y14225 , y14226 , y14227 , y14228 , y14229 , y14230 , y14231 , y14232 , y14233 , y14234 , y14235 , y14236 , y14237 , y14238 , y14239 , y14240 , y14241 , y14242 , y14243 , y14244 , y14245 , y14246 , y14247 , y14248 , y14249 , y14250 , y14251 , y14252 , y14253 , y14254 , y14255 , y14256 , y14257 , y14258 , y14259 , y14260 , y14261 , y14262 , y14263 , y14264 , y14265 , y14266 , y14267 , y14268 , y14269 , y14270 , y14271 , y14272 , y14273 , y14274 , y14275 , y14276 , y14277 , y14278 , y14279 , y14280 , y14281 , y14282 , y14283 , y14284 , y14285 , y14286 , y14287 , y14288 , y14289 , y14290 , y14291 , y14292 , y14293 , y14294 , y14295 , y14296 , y14297 , y14298 , y14299 , y14300 , y14301 , y14302 , y14303 , y14304 , y14305 , y14306 , y14307 , y14308 , y14309 , y14310 , y14311 , y14312 , y14313 , y14314 , y14315 , y14316 , y14317 , y14318 , y14319 , y14320 , y14321 , y14322 , y14323 , y14324 , y14325 , y14326 , y14327 , y14328 , y14329 , y14330 , y14331 , y14332 , y14333 , y14334 , y14335 , y14336 , y14337 , y14338 , y14339 , y14340 , y14341 , y14342 , y14343 , y14344 , y14345 , y14346 , y14347 , y14348 , y14349 , y14350 , y14351 , y14352 , y14353 , y14354 , y14355 , y14356 , y14357 , y14358 , y14359 , y14360 , y14361 , y14362 , y14363 , y14364 , y14365 , y14366 , y14367 , y14368 , y14369 , y14370 , y14371 , y14372 , y14373 , y14374 , y14375 , y14376 , y14377 , y14378 , y14379 , y14380 , y14381 , y14382 , y14383 , y14384 , y14385 , y14386 , y14387 , y14388 , y14389 , y14390 , y14391 , y14392 , y14393 , y14394 , y14395 , y14396 , y14397 , y14398 , y14399 , y14400 , y14401 , y14402 , y14403 , y14404 , y14405 , y14406 , y14407 , y14408 , y14409 , y14410 , y14411 , y14412 , y14413 , y14414 , y14415 , y14416 , y14417 , y14418 , y14419 , y14420 , y14421 , y14422 , y14423 , y14424 , y14425 , y14426 , y14427 , y14428 , y14429 , y14430 , y14431 , y14432 , y14433 , y14434 , y14435 , y14436 , y14437 , y14438 , y14439 , y14440 , y14441 , y14442 , y14443 , y14444 , y14445 , y14446 , y14447 , y14448 , y14449 , y14450 , y14451 , y14452 , y14453 , y14454 , y14455 , y14456 , y14457 , y14458 , y14459 , y14460 , y14461 , y14462 , y14463 , y14464 , y14465 , y14466 , y14467 , y14468 , y14469 , y14470 , y14471 , y14472 , y14473 , y14474 , y14475 , y14476 , y14477 , y14478 , y14479 , y14480 , y14481 , y14482 , y14483 , y14484 , y14485 , y14486 , y14487 , y14488 , y14489 , y14490 , y14491 , y14492 , y14493 , y14494 , y14495 , y14496 , y14497 , y14498 , y14499 , y14500 , y14501 , y14502 , y14503 , y14504 , y14505 , y14506 , y14507 , y14508 , y14509 , y14510 , y14511 , y14512 , y14513 , y14514 , y14515 , y14516 , y14517 , y14518 , y14519 , y14520 , y14521 , y14522 , y14523 , y14524 , y14525 , y14526 , y14527 , y14528 , y14529 , y14530 , y14531 , y14532 , y14533 , y14534 , y14535 , y14536 , y14537 , y14538 , y14539 , y14540 , y14541 , y14542 , y14543 , y14544 , y14545 , y14546 , y14547 , y14548 , y14549 , y14550 , y14551 , y14552 , y14553 , y14554 , y14555 , y14556 , y14557 , y14558 , y14559 , y14560 , y14561 , y14562 , y14563 , y14564 , y14565 , y14566 , y14567 , y14568 , y14569 , y14570 , y14571 , y14572 , y14573 , y14574 , y14575 , y14576 , y14577 , y14578 , y14579 , y14580 , y14581 , y14582 , y14583 , y14584 , y14585 , y14586 , y14587 , y14588 , y14589 , y14590 , y14591 , y14592 , y14593 , y14594 , y14595 , y14596 , y14597 , y14598 , y14599 , y14600 , y14601 , y14602 , y14603 , y14604 , y14605 , y14606 , y14607 , y14608 , y14609 , y14610 , y14611 , y14612 , y14613 , y14614 , y14615 , y14616 , y14617 , y14618 , y14619 , y14620 , y14621 , y14622 , y14623 , y14624 , y14625 , y14626 , y14627 , y14628 , y14629 , y14630 , y14631 , y14632 , y14633 , y14634 , y14635 , y14636 , y14637 , y14638 , y14639 , y14640 , y14641 , y14642 , y14643 , y14644 , y14645 , y14646 , y14647 , y14648 , y14649 , y14650 , y14651 , y14652 , y14653 , y14654 , y14655 , y14656 , y14657 , y14658 , y14659 , y14660 , y14661 , y14662 , y14663 , y14664 , y14665 , y14666 , y14667 , y14668 , y14669 , y14670 , y14671 , y14672 , y14673 , y14674 , y14675 , y14676 , y14677 , y14678 , y14679 , y14680 , y14681 , y14682 , y14683 , y14684 , y14685 , y14686 , y14687 , y14688 , y14689 , y14690 , y14691 , y14692 , y14693 , y14694 , y14695 , y14696 , y14697 , y14698 , y14699 , y14700 , y14701 , y14702 , y14703 , y14704 , y14705 , y14706 , y14707 , y14708 , y14709 , y14710 , y14711 , y14712 , y14713 , y14714 , y14715 , y14716 , y14717 , y14718 , y14719 , y14720 , y14721 , y14722 , y14723 , y14724 , y14725 , y14726 , y14727 , y14728 , y14729 , y14730 , y14731 , y14732 , y14733 , y14734 , y14735 , y14736 , y14737 , y14738 , y14739 , y14740 , y14741 , y14742 , y14743 , y14744 , y14745 , y14746 , y14747 , y14748 , y14749 , y14750 , y14751 , y14752 , y14753 , y14754 , y14755 , y14756 , y14757 , y14758 , y14759 , y14760 , y14761 , y14762 , y14763 , y14764 , y14765 , y14766 , y14767 , y14768 , y14769 , y14770 , y14771 , y14772 , y14773 , y14774 , y14775 , y14776 , y14777 , y14778 , y14779 , y14780 , y14781 , y14782 , y14783 , y14784 , y14785 , y14786 , y14787 , y14788 , y14789 , y14790 , y14791 , y14792 , y14793 , y14794 , y14795 , y14796 , y14797 , y14798 , y14799 , y14800 , y14801 , y14802 , y14803 , y14804 , y14805 , y14806 , y14807 , y14808 , y14809 , y14810 , y14811 , y14812 , y14813 , y14814 , y14815 , y14816 , y14817 , y14818 , y14819 , y14820 , y14821 , y14822 , y14823 , y14824 , y14825 , y14826 , y14827 , y14828 , y14829 , y14830 , y14831 , y14832 , y14833 , y14834 , y14835 , y14836 , y14837 , y14838 , y14839 , y14840 , y14841 , y14842 , y14843 , y14844 , y14845 , y14846 , y14847 , y14848 , y14849 , y14850 , y14851 , y14852 , y14853 , y14854 , y14855 , y14856 , y14857 , y14858 , y14859 , y14860 , y14861 , y14862 , y14863 , y14864 , y14865 , y14866 , y14867 , y14868 , y14869 , y14870 , y14871 , y14872 , y14873 , y14874 , y14875 , y14876 , y14877 , y14878 , y14879 , y14880 , y14881 , y14882 , y14883 , y14884 , y14885 , y14886 , y14887 , y14888 , y14889 , y14890 , y14891 , y14892 , y14893 , y14894 , y14895 , y14896 , y14897 , y14898 , y14899 , y14900 , y14901 , y14902 , y14903 , y14904 , y14905 , y14906 , y14907 , y14908 , y14909 , y14910 , y14911 , y14912 , y14913 , y14914 , y14915 , y14916 , y14917 , y14918 , y14919 , y14920 , y14921 , y14922 , y14923 , y14924 , y14925 , y14926 , y14927 , y14928 , y14929 , y14930 , y14931 , y14932 , y14933 , y14934 , y14935 , y14936 , y14937 , y14938 , y14939 , y14940 , y14941 , y14942 , y14943 , y14944 , y14945 , y14946 , y14947 , y14948 , y14949 , y14950 , y14951 , y14952 , y14953 , y14954 , y14955 , y14956 , y14957 , y14958 , y14959 , y14960 , y14961 , y14962 , y14963 , y14964 , y14965 , y14966 , y14967 , y14968 , y14969 , y14970 , y14971 , y14972 , y14973 , y14974 , y14975 , y14976 , y14977 , y14978 , y14979 , y14980 , y14981 , y14982 , y14983 , y14984 , y14985 , y14986 , y14987 , y14988 , y14989 , y14990 , y14991 , y14992 , y14993 , y14994 , y14995 , y14996 , y14997 , y14998 , y14999 , y15000 , y15001 , y15002 , y15003 , y15004 , y15005 , y15006 , y15007 , y15008 , y15009 , y15010 , y15011 , y15012 , y15013 , y15014 , y15015 , y15016 , y15017 , y15018 , y15019 , y15020 , y15021 , y15022 , y15023 , y15024 , y15025 , y15026 , y15027 , y15028 , y15029 , y15030 , y15031 , y15032 , y15033 , y15034 , y15035 , y15036 , y15037 , y15038 , y15039 , y15040 , y15041 , y15042 , y15043 , y15044 , y15045 , y15046 , y15047 , y15048 , y15049 , y15050 , y15051 , y15052 , y15053 , y15054 , y15055 , y15056 , y15057 , y15058 , y15059 , y15060 , y15061 , y15062 , y15063 , y15064 , y15065 , y15066 , y15067 , y15068 , y15069 , y15070 , y15071 , y15072 , y15073 , y15074 , y15075 , y15076 , y15077 , y15078 , y15079 , y15080 , y15081 , y15082 , y15083 , y15084 , y15085 , y15086 , y15087 , y15088 , y15089 , y15090 , y15091 , y15092 , y15093 , y15094 , y15095 , y15096 , y15097 , y15098 , y15099 , y15100 , y15101 , y15102 , y15103 , y15104 , y15105 , y15106 , y15107 , y15108 , y15109 , y15110 , y15111 , y15112 , y15113 , y15114 , y15115 , y15116 , y15117 , y15118 , y15119 , y15120 , y15121 , y15122 , y15123 , y15124 , y15125 , y15126 , y15127 , y15128 , y15129 , y15130 , y15131 , y15132 , y15133 , y15134 , y15135 , y15136 , y15137 , y15138 , y15139 , y15140 , y15141 , y15142 , y15143 , y15144 , y15145 , y15146 , y15147 , y15148 , y15149 , y15150 , y15151 , y15152 , y15153 , y15154 , y15155 , y15156 , y15157 , y15158 , y15159 , y15160 , y15161 , y15162 , y15163 , y15164 , y15165 , y15166 , y15167 , y15168 , y15169 , y15170 , y15171 , y15172 , y15173 , y15174 , y15175 , y15176 , y15177 , y15178 , y15179 , y15180 , y15181 , y15182 , y15183 , y15184 , y15185 , y15186 , y15187 , y15188 , y15189 , y15190 , y15191 , y15192 , y15193 , y15194 , y15195 , y15196 , y15197 , y15198 , y15199 , y15200 , y15201 , y15202 , y15203 , y15204 , y15205 , y15206 , y15207 , y15208 , y15209 , y15210 , y15211 , y15212 , y15213 , y15214 , y15215 , y15216 , y15217 , y15218 , y15219 , y15220 , y15221 , y15222 , y15223 , y15224 , y15225 , y15226 , y15227 , y15228 , y15229 , y15230 , y15231 , y15232 , y15233 , y15234 , y15235 , y15236 , y15237 , y15238 , y15239 , y15240 , y15241 , y15242 , y15243 , y15244 , y15245 , y15246 , y15247 , y15248 , y15249 , y15250 , y15251 , y15252 , y15253 , y15254 , y15255 , y15256 , y15257 , y15258 , y15259 , y15260 , y15261 , y15262 , y15263 , y15264 , y15265 , y15266 , y15267 , y15268 , y15269 , y15270 , y15271 , y15272 , y15273 , y15274 , y15275 , y15276 , y15277 , y15278 , y15279 , y15280 , y15281 , y15282 , y15283 , y15284 , y15285 , y15286 , y15287 , y15288 , y15289 , y15290 , y15291 , y15292 , y15293 , y15294 , y15295 , y15296 , y15297 , y15298 , y15299 , y15300 , y15301 , y15302 , y15303 , y15304 , y15305 , y15306 , y15307 , y15308 , y15309 , y15310 , y15311 , y15312 , y15313 , y15314 , y15315 , y15316 , y15317 , y15318 , y15319 , y15320 , y15321 , y15322 , y15323 , y15324 , y15325 , y15326 , y15327 , y15328 , y15329 , y15330 , y15331 , y15332 , y15333 , y15334 , y15335 , y15336 , y15337 , y15338 , y15339 , y15340 , y15341 , y15342 , y15343 , y15344 , y15345 , y15346 , y15347 , y15348 , y15349 , y15350 , y15351 , y15352 , y15353 , y15354 , y15355 , y15356 , y15357 , y15358 , y15359 , y15360 , y15361 , y15362 , y15363 , y15364 , y15365 , y15366 , y15367 , y15368 , y15369 , y15370 , y15371 , y15372 , y15373 , y15374 , y15375 , y15376 , y15377 , y15378 , y15379 , y15380 , y15381 , y15382 , y15383 , y15384 , y15385 , y15386 , y15387 , y15388 , y15389 , y15390 , y15391 , y15392 , y15393 , y15394 , y15395 , y15396 , y15397 , y15398 , y15399 , y15400 , y15401 , y15402 , y15403 , y15404 , y15405 , y15406 , y15407 , y15408 , y15409 , y15410 , y15411 , y15412 , y15413 , y15414 , y15415 , y15416 , y15417 , y15418 , y15419 , y15420 , y15421 , y15422 , y15423 , y15424 , y15425 , y15426 , y15427 , y15428 , y15429 , y15430 , y15431 , y15432 , y15433 , y15434 , y15435 , y15436 , y15437 , y15438 , y15439 , y15440 , y15441 , y15442 , y15443 , y15444 , y15445 , y15446 , y15447 , y15448 , y15449 , y15450 , y15451 , y15452 , y15453 , y15454 , y15455 , y15456 , y15457 , y15458 , y15459 , y15460 , y15461 , y15462 , y15463 , y15464 , y15465 , y15466 , y15467 , y15468 , y15469 , y15470 , y15471 , y15472 , y15473 , y15474 , y15475 , y15476 , y15477 , y15478 , y15479 , y15480 , y15481 , y15482 , y15483 , y15484 , y15485 , y15486 , y15487 , y15488 , y15489 , y15490 , y15491 , y15492 , y15493 , y15494 , y15495 , y15496 , y15497 , y15498 , y15499 , y15500 , y15501 , y15502 , y15503 , y15504 , y15505 , y15506 , y15507 , y15508 , y15509 , y15510 , y15511 , y15512 , y15513 , y15514 , y15515 , y15516 , y15517 , y15518 , y15519 , y15520 , y15521 , y15522 , y15523 , y15524 , y15525 , y15526 , y15527 , y15528 , y15529 , y15530 , y15531 , y15532 , y15533 , y15534 , y15535 , y15536 , y15537 , y15538 , y15539 , y15540 , y15541 , y15542 , y15543 , y15544 , y15545 , y15546 , y15547 , y15548 , y15549 , y15550 , y15551 , y15552 , y15553 , y15554 , y15555 , y15556 , y15557 , y15558 , y15559 , y15560 , y15561 , y15562 , y15563 , y15564 , y15565 , y15566 , y15567 , y15568 , y15569 , y15570 , y15571 , y15572 , y15573 , y15574 , y15575 , y15576 , y15577 , y15578 , y15579 , y15580 , y15581 , y15582 , y15583 , y15584 , y15585 , y15586 , y15587 , y15588 , y15589 , y15590 , y15591 , y15592 , y15593 , y15594 , y15595 , y15596 , y15597 , y15598 , y15599 , y15600 , y15601 , y15602 , y15603 , y15604 , y15605 , y15606 , y15607 , y15608 , y15609 , y15610 , y15611 , y15612 , y15613 , y15614 , y15615 , y15616 , y15617 , y15618 , y15619 , y15620 , y15621 , y15622 , y15623 , y15624 , y15625 , y15626 , y15627 , y15628 , y15629 , y15630 , y15631 , y15632 , y15633 , y15634 , y15635 , y15636 , y15637 , y15638 , y15639 , y15640 , y15641 , y15642 , y15643 , y15644 , y15645 , y15646 , y15647 , y15648 , y15649 , y15650 , y15651 , y15652 , y15653 , y15654 , y15655 , y15656 , y15657 , y15658 , y15659 , y15660 , y15661 , y15662 , y15663 , y15664 , y15665 , y15666 , y15667 , y15668 , y15669 , y15670 , y15671 , y15672 , y15673 , y15674 , y15675 , y15676 , y15677 , y15678 , y15679 , y15680 , y15681 , y15682 , y15683 , y15684 , y15685 , y15686 , y15687 , y15688 , y15689 , y15690 , y15691 , y15692 , y15693 , y15694 , y15695 , y15696 , y15697 , y15698 , y15699 , y15700 , y15701 , y15702 , y15703 , y15704 , y15705 , y15706 , y15707 , y15708 , y15709 , y15710 , y15711 , y15712 , y15713 , y15714 , y15715 , y15716 , y15717 , y15718 , y15719 , y15720 , y15721 , y15722 , y15723 , y15724 , y15725 , y15726 , y15727 , y15728 , y15729 , y15730 , y15731 , y15732 , y15733 , y15734 , y15735 , y15736 , y15737 , y15738 , y15739 , y15740 , y15741 , y15742 , y15743 , y15744 , y15745 , y15746 , y15747 , y15748 , y15749 , y15750 , y15751 , y15752 , y15753 , y15754 , y15755 , y15756 , y15757 , y15758 , y15759 , y15760 , y15761 , y15762 , y15763 , y15764 , y15765 , y15766 , y15767 , y15768 , y15769 , y15770 , y15771 , y15772 , y15773 , y15774 , y15775 , y15776 , y15777 , y15778 , y15779 , y15780 , y15781 , y15782 , y15783 , y15784 , y15785 , y15786 , y15787 , y15788 , y15789 , y15790 , y15791 , y15792 , y15793 , y15794 , y15795 , y15796 , y15797 , y15798 , y15799 , y15800 , y15801 , y15802 , y15803 , y15804 , y15805 , y15806 , y15807 , y15808 , y15809 , y15810 , y15811 , y15812 , y15813 , y15814 , y15815 , y15816 , y15817 , y15818 , y15819 , y15820 , y15821 , y15822 , y15823 , y15824 , y15825 , y15826 , y15827 , y15828 , y15829 , y15830 , y15831 , y15832 , y15833 , y15834 , y15835 , y15836 , y15837 , y15838 , y15839 , y15840 , y15841 , y15842 , y15843 , y15844 , y15845 , y15846 , y15847 , y15848 , y15849 , y15850 , y15851 , y15852 , y15853 , y15854 , y15855 , y15856 , y15857 , y15858 , y15859 , y15860 , y15861 , y15862 , y15863 , y15864 , y15865 , y15866 , y15867 , y15868 , y15869 , y15870 , y15871 , y15872 , y15873 , y15874 , y15875 , y15876 , y15877 , y15878 , y15879 , y15880 , y15881 , y15882 , y15883 , y15884 , y15885 , y15886 , y15887 , y15888 , y15889 , y15890 , y15891 , y15892 , y15893 , y15894 , y15895 , y15896 , y15897 , y15898 , y15899 , y15900 , y15901 , y15902 , y15903 , y15904 , y15905 , y15906 , y15907 , y15908 , y15909 , y15910 , y15911 , y15912 , y15913 , y15914 , y15915 , y15916 , y15917 , y15918 , y15919 , y15920 , y15921 , y15922 , y15923 , y15924 , y15925 , y15926 , y15927 , y15928 , y15929 , y15930 , y15931 , y15932 , y15933 , y15934 , y15935 , y15936 , y15937 , y15938 , y15939 , y15940 , y15941 , y15942 , y15943 , y15944 , y15945 , y15946 , y15947 , y15948 , y15949 , y15950 , y15951 , y15952 , y15953 , y15954 , y15955 , y15956 , y15957 , y15958 , y15959 , y15960 , y15961 , y15962 , y15963 , y15964 , y15965 , y15966 , y15967 , y15968 , y15969 , y15970 , y15971 , y15972 , y15973 , y15974 , y15975 , y15976 , y15977 , y15978 , y15979 , y15980 , y15981 , y15982 , y15983 , y15984 , y15985 , y15986 , y15987 , y15988 , y15989 , y15990 , y15991 , y15992 , y15993 , y15994 , y15995 , y15996 , y15997 , y15998 , y15999 , y16000 , y16001 , y16002 , y16003 , y16004 , y16005 , y16006 , y16007 , y16008 , y16009 , y16010 , y16011 , y16012 , y16013 , y16014 , y16015 , y16016 , y16017 , y16018 , y16019 , y16020 , y16021 , y16022 , y16023 , y16024 , y16025 , y16026 , y16027 , y16028 , y16029 , y16030 , y16031 , y16032 , y16033 , y16034 , y16035 , y16036 , y16037 , y16038 , y16039 , y16040 , y16041 , y16042 , y16043 , y16044 , y16045 , y16046 , y16047 , y16048 , y16049 , y16050 , y16051 , y16052 , y16053 , y16054 , y16055 , y16056 , y16057 , y16058 , y16059 , y16060 , y16061 , y16062 , y16063 , y16064 , y16065 , y16066 , y16067 , y16068 , y16069 , y16070 , y16071 , y16072 , y16073 , y16074 , y16075 , y16076 , y16077 , y16078 , y16079 , y16080 , y16081 , y16082 , y16083 , y16084 , y16085 , y16086 , y16087 , y16088 , y16089 , y16090 , y16091 , y16092 , y16093 , y16094 , y16095 , y16096 , y16097 , y16098 , y16099 , y16100 , y16101 , y16102 , y16103 , y16104 , y16105 , y16106 , y16107 , y16108 , y16109 , y16110 , y16111 , y16112 , y16113 , y16114 , y16115 , y16116 , y16117 , y16118 , y16119 , y16120 , y16121 , y16122 , y16123 , y16124 , y16125 , y16126 , y16127 , y16128 , y16129 , y16130 , y16131 , y16132 , y16133 , y16134 , y16135 , y16136 , y16137 , y16138 , y16139 , y16140 , y16141 , y16142 , y16143 , y16144 , y16145 , y16146 , y16147 , y16148 , y16149 , y16150 , y16151 , y16152 , y16153 , y16154 , y16155 , y16156 , y16157 , y16158 , y16159 , y16160 , y16161 , y16162 , y16163 , y16164 , y16165 , y16166 , y16167 , y16168 , y16169 , y16170 , y16171 , y16172 , y16173 , y16174 , y16175 , y16176 , y16177 , y16178 , y16179 , y16180 , y16181 , y16182 , y16183 , y16184 , y16185 , y16186 , y16187 , y16188 , y16189 , y16190 , y16191 , y16192 , y16193 , y16194 , y16195 , y16196 , y16197 , y16198 , y16199 , y16200 , y16201 , y16202 , y16203 , y16204 , y16205 , y16206 , y16207 , y16208 , y16209 , y16210 , y16211 , y16212 , y16213 , y16214 , y16215 , y16216 , y16217 , y16218 , y16219 , y16220 , y16221 , y16222 , y16223 , y16224 , y16225 , y16226 , y16227 , y16228 , y16229 , y16230 , y16231 , y16232 , y16233 , y16234 , y16235 , y16236 , y16237 , y16238 , y16239 , y16240 , y16241 , y16242 , y16243 , y16244 , y16245 , y16246 , y16247 , y16248 , y16249 , y16250 , y16251 , y16252 , y16253 , y16254 , y16255 , y16256 , y16257 , y16258 , y16259 , y16260 , y16261 , y16262 , y16263 , y16264 , y16265 , y16266 , y16267 , y16268 , y16269 , y16270 , y16271 , y16272 , y16273 , y16274 , y16275 , y16276 , y16277 , y16278 , y16279 , y16280 , y16281 , y16282 , y16283 , y16284 , y16285 , y16286 , y16287 , y16288 , y16289 , y16290 , y16291 , y16292 , y16293 , y16294 , y16295 , y16296 , y16297 , y16298 , y16299 , y16300 , y16301 , y16302 , y16303 , y16304 , y16305 , y16306 , y16307 , y16308 , y16309 , y16310 , y16311 , y16312 , y16313 , y16314 , y16315 , y16316 , y16317 , y16318 , y16319 , y16320 , y16321 , y16322 , y16323 , y16324 , y16325 , y16326 , y16327 , y16328 , y16329 , y16330 , y16331 , y16332 , y16333 , y16334 , y16335 , y16336 , y16337 , y16338 , y16339 , y16340 , y16341 , y16342 , y16343 , y16344 , y16345 , y16346 , y16347 , y16348 , y16349 , y16350 , y16351 , y16352 , y16353 , y16354 , y16355 , y16356 , y16357 , y16358 , y16359 , y16360 , y16361 , y16362 , y16363 , y16364 , y16365 , y16366 , y16367 , y16368 , y16369 , y16370 , y16371 , y16372 , y16373 , y16374 , y16375 , y16376 , y16377 , y16378 , y16379 , y16380 , y16381 , y16382 , y16383 , y16384 , y16385 , y16386 , y16387 , y16388 , y16389 , y16390 , y16391 , y16392 , y16393 , y16394 , y16395 , y16396 , y16397 , y16398 , y16399 , y16400 , y16401 , y16402 , y16403 , y16404 , y16405 , y16406 , y16407 , y16408 , y16409 , y16410 , y16411 , y16412 , y16413 , y16414 , y16415 , y16416 , y16417 , y16418 , y16419 , y16420 , y16421 , y16422 , y16423 , y16424 , y16425 , y16426 , y16427 , y16428 , y16429 , y16430 , y16431 , y16432 , y16433 , y16434 , y16435 , y16436 , y16437 , y16438 , y16439 , y16440 , y16441 , y16442 , y16443 , y16444 , y16445 , y16446 , y16447 , y16448 , y16449 , y16450 , y16451 , y16452 , y16453 , y16454 , y16455 , y16456 , y16457 , y16458 , y16459 , y16460 , y16461 , y16462 , y16463 , y16464 , y16465 , y16466 , y16467 , y16468 , y16469 , y16470 , y16471 , y16472 , y16473 , y16474 , y16475 , y16476 , y16477 , y16478 , y16479 , y16480 , y16481 , y16482 , y16483 , y16484 , y16485 , y16486 , y16487 , y16488 , y16489 , y16490 , y16491 , y16492 , y16493 , y16494 , y16495 , y16496 , y16497 , y16498 , y16499 , y16500 , y16501 , y16502 , y16503 , y16504 , y16505 , y16506 , y16507 , y16508 , y16509 , y16510 , y16511 , y16512 , y16513 , y16514 , y16515 , y16516 , y16517 , y16518 , y16519 , y16520 , y16521 , y16522 , y16523 , y16524 , y16525 , y16526 , y16527 , y16528 , y16529 , y16530 , y16531 , y16532 , y16533 , y16534 , y16535 , y16536 , y16537 , y16538 , y16539 , y16540 , y16541 , y16542 , y16543 , y16544 , y16545 , y16546 , y16547 , y16548 , y16549 , y16550 , y16551 , y16552 , y16553 , y16554 , y16555 , y16556 , y16557 , y16558 , y16559 , y16560 , y16561 , y16562 , y16563 , y16564 , y16565 , y16566 , y16567 , y16568 , y16569 , y16570 , y16571 , y16572 , y16573 , y16574 , y16575 , y16576 , y16577 , y16578 , y16579 , y16580 , y16581 , y16582 , y16583 , y16584 , y16585 , y16586 , y16587 , y16588 , y16589 , y16590 , y16591 , y16592 , y16593 , y16594 , y16595 , y16596 , y16597 , y16598 , y16599 , y16600 , y16601 , y16602 , y16603 , y16604 , y16605 , y16606 , y16607 , y16608 , y16609 , y16610 , y16611 , y16612 , y16613 , y16614 , y16615 , y16616 , y16617 , y16618 , y16619 , y16620 , y16621 , y16622 , y16623 , y16624 , y16625 , y16626 , y16627 , y16628 , y16629 , y16630 , y16631 , y16632 , y16633 , y16634 , y16635 , y16636 , y16637 , y16638 , y16639 , y16640 , y16641 , y16642 , y16643 , y16644 , y16645 , y16646 , y16647 , y16648 , y16649 , y16650 , y16651 , y16652 , y16653 , y16654 , y16655 , y16656 , y16657 , y16658 , y16659 , y16660 , y16661 , y16662 , y16663 , y16664 , y16665 , y16666 , y16667 , y16668 , y16669 , y16670 , y16671 , y16672 , y16673 , y16674 , y16675 , y16676 , y16677 , y16678 , y16679 , y16680 , y16681 , y16682 , y16683 , y16684 , y16685 , y16686 , y16687 , y16688 , y16689 , y16690 , y16691 , y16692 , y16693 , y16694 , y16695 , y16696 , y16697 , y16698 , y16699 , y16700 , y16701 , y16702 , y16703 , y16704 , y16705 , y16706 , y16707 , y16708 , y16709 , y16710 , y16711 , y16712 , y16713 , y16714 , y16715 , y16716 , y16717 , y16718 , y16719 , y16720 , y16721 , y16722 , y16723 , y16724 , y16725 , y16726 , y16727 , y16728 , y16729 , y16730 , y16731 , y16732 , y16733 , y16734 , y16735 , y16736 , y16737 , y16738 , y16739 , y16740 , y16741 , y16742 , y16743 , y16744 , y16745 , y16746 , y16747 , y16748 , y16749 , y16750 , y16751 , y16752 , y16753 , y16754 , y16755 , y16756 , y16757 , y16758 , y16759 , y16760 , y16761 , y16762 , y16763 , y16764 , y16765 , y16766 , y16767 , y16768 , y16769 , y16770 , y16771 , y16772 , y16773 , y16774 , y16775 , y16776 , y16777 , y16778 , y16779 , y16780 , y16781 , y16782 , y16783 , y16784 , y16785 , y16786 , y16787 , y16788 , y16789 , y16790 , y16791 , y16792 , y16793 , y16794 , y16795 , y16796 , y16797 , y16798 , y16799 , y16800 , y16801 , y16802 , y16803 , y16804 , y16805 , y16806 , y16807 , y16808 , y16809 , y16810 , y16811 , y16812 , y16813 , y16814 , y16815 , y16816 , y16817 , y16818 , y16819 , y16820 , y16821 , y16822 , y16823 , y16824 , y16825 , y16826 , y16827 , y16828 , y16829 , y16830 , y16831 , y16832 , y16833 , y16834 , y16835 , y16836 , y16837 , y16838 , y16839 , y16840 , y16841 , y16842 , y16843 , y16844 , y16845 , y16846 , y16847 , y16848 , y16849 , y16850 , y16851 , y16852 , y16853 , y16854 , y16855 , y16856 , y16857 , y16858 , y16859 , y16860 , y16861 , y16862 , y16863 , y16864 , y16865 , y16866 , y16867 , y16868 , y16869 , y16870 , y16871 , y16872 , y16873 , y16874 , y16875 , y16876 , y16877 , y16878 , y16879 , y16880 , y16881 , y16882 , y16883 , y16884 , y16885 , y16886 , y16887 , y16888 , y16889 , y16890 , y16891 , y16892 , y16893 , y16894 , y16895 , y16896 , y16897 , y16898 , y16899 , y16900 , y16901 , y16902 , y16903 , y16904 , y16905 , y16906 , y16907 , y16908 , y16909 , y16910 , y16911 , y16912 , y16913 , y16914 , y16915 , y16916 , y16917 , y16918 , y16919 , y16920 , y16921 , y16922 , y16923 , y16924 , y16925 , y16926 , y16927 , y16928 , y16929 , y16930 , y16931 , y16932 , y16933 , y16934 , y16935 , y16936 , y16937 , y16938 , y16939 , y16940 , y16941 , y16942 , y16943 , y16944 , y16945 , y16946 , y16947 , y16948 , y16949 , y16950 , y16951 , y16952 , y16953 , y16954 , y16955 , y16956 , y16957 , y16958 , y16959 , y16960 , y16961 , y16962 , y16963 , y16964 , y16965 , y16966 , y16967 , y16968 , y16969 , y16970 , y16971 , y16972 , y16973 , y16974 , y16975 , y16976 , y16977 , y16978 , y16979 , y16980 , y16981 , y16982 , y16983 , y16984 , y16985 , y16986 , y16987 , y16988 , y16989 , y16990 , y16991 , y16992 , y16993 , y16994 , y16995 , y16996 , y16997 , y16998 , y16999 , y17000 , y17001 , y17002 , y17003 , y17004 , y17005 , y17006 , y17007 , y17008 , y17009 , y17010 , y17011 , y17012 , y17013 , y17014 , y17015 , y17016 , y17017 , y17018 , y17019 , y17020 , y17021 , y17022 , y17023 , y17024 , y17025 , y17026 , y17027 , y17028 , y17029 , y17030 , y17031 , y17032 , y17033 , y17034 , y17035 , y17036 , y17037 , y17038 , y17039 , y17040 , y17041 , y17042 , y17043 , y17044 , y17045 , y17046 , y17047 , y17048 , y17049 , y17050 , y17051 , y17052 , y17053 , y17054 , y17055 , y17056 , y17057 , y17058 , y17059 , y17060 , y17061 , y17062 , y17063 , y17064 , y17065 , y17066 , y17067 , y17068 , y17069 , y17070 , y17071 , y17072 , y17073 , y17074 , y17075 , y17076 , y17077 , y17078 , y17079 , y17080 , y17081 , y17082 , y17083 , y17084 , y17085 , y17086 , y17087 , y17088 , y17089 , y17090 , y17091 , y17092 , y17093 , y17094 , y17095 , y17096 , y17097 , y17098 , y17099 , y17100 , y17101 , y17102 , y17103 , y17104 , y17105 , y17106 , y17107 , y17108 , y17109 , y17110 , y17111 , y17112 , y17113 , y17114 , y17115 , y17116 , y17117 , y17118 , y17119 , y17120 , y17121 , y17122 , y17123 , y17124 , y17125 , y17126 , y17127 , y17128 , y17129 , y17130 , y17131 , y17132 , y17133 , y17134 , y17135 , y17136 , y17137 , y17138 , y17139 , y17140 , y17141 , y17142 , y17143 , y17144 , y17145 , y17146 , y17147 , y17148 , y17149 , y17150 , y17151 , y17152 , y17153 , y17154 , y17155 , y17156 , y17157 , y17158 , y17159 , y17160 , y17161 , y17162 , y17163 , y17164 , y17165 , y17166 , y17167 , y17168 , y17169 , y17170 , y17171 , y17172 , y17173 , y17174 , y17175 , y17176 , y17177 , y17178 , y17179 , y17180 , y17181 , y17182 , y17183 , y17184 , y17185 , y17186 , y17187 , y17188 , y17189 , y17190 , y17191 , y17192 , y17193 , y17194 , y17195 , y17196 , y17197 , y17198 , y17199 , y17200 , y17201 , y17202 , y17203 , y17204 , y17205 , y17206 , y17207 , y17208 , y17209 , y17210 , y17211 , y17212 , y17213 , y17214 , y17215 , y17216 , y17217 , y17218 , y17219 , y17220 , y17221 , y17222 , y17223 , y17224 , y17225 , y17226 , y17227 , y17228 , y17229 , y17230 , y17231 , y17232 , y17233 , y17234 , y17235 , y17236 , y17237 , y17238 , y17239 , y17240 , y17241 , y17242 , y17243 , y17244 , y17245 , y17246 , y17247 , y17248 , y17249 , y17250 , y17251 , y17252 , y17253 , y17254 , y17255 , y17256 , y17257 , y17258 , y17259 , y17260 , y17261 , y17262 , y17263 , y17264 , y17265 , y17266 , y17267 , y17268 , y17269 , y17270 , y17271 , y17272 , y17273 , y17274 , y17275 , y17276 , y17277 , y17278 , y17279 , y17280 , y17281 , y17282 , y17283 , y17284 , y17285 , y17286 , y17287 , y17288 , y17289 , y17290 , y17291 , y17292 , y17293 , y17294 , y17295 , y17296 , y17297 , y17298 , y17299 , y17300 , y17301 , y17302 , y17303 , y17304 , y17305 , y17306 , y17307 , y17308 , y17309 , y17310 , y17311 , y17312 , y17313 , y17314 , y17315 , y17316 , y17317 , y17318 , y17319 , y17320 , y17321 , y17322 , y17323 , y17324 , y17325 , y17326 , y17327 , y17328 , y17329 , y17330 , y17331 , y17332 , y17333 , y17334 , y17335 , y17336 , y17337 , y17338 , y17339 , y17340 , y17341 , y17342 , y17343 , y17344 , y17345 , y17346 , y17347 , y17348 , y17349 , y17350 , y17351 , y17352 , y17353 , y17354 , y17355 , y17356 , y17357 , y17358 , y17359 , y17360 , y17361 , y17362 , y17363 , y17364 , y17365 , y17366 , y17367 , y17368 , y17369 , y17370 , y17371 , y17372 , y17373 , y17374 , y17375 , y17376 , y17377 , y17378 , y17379 , y17380 , y17381 , y17382 , y17383 , y17384 , y17385 , y17386 , y17387 , y17388 , y17389 , y17390 , y17391 , y17392 , y17393 , y17394 , y17395 , y17396 , y17397 , y17398 , y17399 , y17400 , y17401 , y17402 , y17403 , y17404 , y17405 , y17406 , y17407 , y17408 , y17409 , y17410 , y17411 , y17412 , y17413 , y17414 , y17415 , y17416 , y17417 , y17418 , y17419 , y17420 , y17421 , y17422 , y17423 , y17424 , y17425 , y17426 , y17427 , y17428 , y17429 , y17430 , y17431 , y17432 , y17433 , y17434 , y17435 , y17436 , y17437 , y17438 , y17439 , y17440 , y17441 , y17442 , y17443 , y17444 , y17445 , y17446 , y17447 , y17448 , y17449 , y17450 , y17451 , y17452 , y17453 , y17454 , y17455 , y17456 , y17457 , y17458 , y17459 , y17460 , y17461 , y17462 , y17463 , y17464 , y17465 , y17466 , y17467 , y17468 , y17469 , y17470 , y17471 , y17472 , y17473 , y17474 , y17475 , y17476 , y17477 , y17478 , y17479 , y17480 , y17481 , y17482 , y17483 , y17484 , y17485 , y17486 , y17487 , y17488 , y17489 , y17490 , y17491 , y17492 , y17493 , y17494 , y17495 , y17496 , y17497 , y17498 , y17499 , y17500 , y17501 , y17502 , y17503 , y17504 , y17505 , y17506 , y17507 , y17508 , y17509 , y17510 , y17511 , y17512 , y17513 , y17514 , y17515 , y17516 , y17517 , y17518 , y17519 , y17520 , y17521 , y17522 , y17523 , y17524 , y17525 , y17526 , y17527 , y17528 , y17529 , y17530 , y17531 , y17532 , y17533 , y17534 , y17535 , y17536 , y17537 , y17538 , y17539 , y17540 , y17541 , y17542 , y17543 , y17544 , y17545 , y17546 , y17547 , y17548 , y17549 , y17550 , y17551 , y17552 , y17553 , y17554 , y17555 , y17556 , y17557 , y17558 , y17559 , y17560 , y17561 , y17562 , y17563 , y17564 , y17565 , y17566 , y17567 , y17568 , y17569 , y17570 , y17571 , y17572 , y17573 , y17574 , y17575 , y17576 , y17577 , y17578 , y17579 , y17580 , y17581 , y17582 , y17583 , y17584 , y17585 , y17586 , y17587 , y17588 , y17589 , y17590 , y17591 , y17592 , y17593 , y17594 , y17595 , y17596 , y17597 , y17598 , y17599 , y17600 , y17601 , y17602 , y17603 , y17604 , y17605 , y17606 , y17607 , y17608 , y17609 , y17610 , y17611 , y17612 , y17613 , y17614 , y17615 , y17616 , y17617 , y17618 , y17619 , y17620 , y17621 , y17622 , y17623 , y17624 , y17625 , y17626 , y17627 , y17628 , y17629 , y17630 , y17631 , y17632 , y17633 , y17634 , y17635 , y17636 , y17637 , y17638 , y17639 , y17640 , y17641 , y17642 , y17643 , y17644 , y17645 , y17646 , y17647 , y17648 , y17649 , y17650 , y17651 , y17652 , y17653 , y17654 , y17655 , y17656 , y17657 , y17658 , y17659 , y17660 , y17661 , y17662 , y17663 , y17664 , y17665 , y17666 , y17667 , y17668 , y17669 , y17670 , y17671 , y17672 , y17673 , y17674 , y17675 , y17676 , y17677 , y17678 , y17679 , y17680 , y17681 , y17682 , y17683 , y17684 , y17685 , y17686 , y17687 , y17688 , y17689 , y17690 , y17691 , y17692 , y17693 , y17694 , y17695 , y17696 , y17697 , y17698 , y17699 , y17700 , y17701 , y17702 , y17703 , y17704 , y17705 , y17706 , y17707 , y17708 , y17709 , y17710 , y17711 , y17712 , y17713 , y17714 , y17715 , y17716 , y17717 , y17718 , y17719 , y17720 , y17721 , y17722 , y17723 , y17724 , y17725 , y17726 , y17727 , y17728 , y17729 , y17730 , y17731 , y17732 , y17733 , y17734 , y17735 , y17736 , y17737 , y17738 , y17739 , y17740 , y17741 , y17742 , y17743 , y17744 , y17745 , y17746 , y17747 , y17748 , y17749 , y17750 , y17751 , y17752 , y17753 , y17754 , y17755 , y17756 , y17757 , y17758 , y17759 , y17760 , y17761 , y17762 , y17763 , y17764 , y17765 , y17766 , y17767 , y17768 , y17769 , y17770 , y17771 , y17772 , y17773 , y17774 , y17775 , y17776 , y17777 , y17778 , y17779 , y17780 , y17781 , y17782 , y17783 , y17784 , y17785 , y17786 , y17787 , y17788 , y17789 , y17790 , y17791 , y17792 , y17793 , y17794 , y17795 , y17796 , y17797 , y17798 , y17799 , y17800 , y17801 , y17802 , y17803 , y17804 , y17805 , y17806 , y17807 , y17808 , y17809 , y17810 , y17811 , y17812 , y17813 , y17814 , y17815 , y17816 , y17817 , y17818 , y17819 , y17820 , y17821 , y17822 , y17823 , y17824 , y17825 , y17826 , y17827 , y17828 , y17829 , y17830 , y17831 , y17832 , y17833 , y17834 , y17835 , y17836 , y17837 , y17838 , y17839 , y17840 , y17841 , y17842 , y17843 , y17844 , y17845 , y17846 , y17847 , y17848 , y17849 , y17850 , y17851 , y17852 , y17853 , y17854 , y17855 , y17856 , y17857 , y17858 , y17859 , y17860 , y17861 , y17862 , y17863 , y17864 , y17865 , y17866 , y17867 , y17868 , y17869 , y17870 , y17871 , y17872 , y17873 , y17874 , y17875 , y17876 , y17877 , y17878 , y17879 , y17880 , y17881 , y17882 , y17883 , y17884 , y17885 , y17886 , y17887 , y17888 , y17889 , y17890 , y17891 , y17892 , y17893 , y17894 , y17895 , y17896 , y17897 , y17898 , y17899 , y17900 , y17901 , y17902 , y17903 , y17904 , y17905 , y17906 , y17907 , y17908 , y17909 , y17910 , y17911 , y17912 , y17913 , y17914 , y17915 , y17916 , y17917 , y17918 , y17919 , y17920 , y17921 , y17922 , y17923 , y17924 , y17925 , y17926 , y17927 , y17928 , y17929 , y17930 , y17931 , y17932 , y17933 , y17934 , y17935 , y17936 , y17937 , y17938 , y17939 , y17940 , y17941 , y17942 , y17943 , y17944 , y17945 , y17946 , y17947 , y17948 , y17949 , y17950 , y17951 , y17952 , y17953 , y17954 , y17955 , y17956 , y17957 , y17958 , y17959 , y17960 , y17961 , y17962 , y17963 , y17964 , y17965 , y17966 , y17967 , y17968 , y17969 , y17970 , y17971 , y17972 , y17973 , y17974 , y17975 , y17976 , y17977 , y17978 , y17979 , y17980 , y17981 , y17982 , y17983 , y17984 , y17985 , y17986 , y17987 , y17988 , y17989 , y17990 , y17991 , y17992 , y17993 , y17994 , y17995 , y17996 , y17997 , y17998 , y17999 , y18000 , y18001 , y18002 , y18003 , y18004 , y18005 , y18006 , y18007 , y18008 , y18009 , y18010 , y18011 , y18012 , y18013 , y18014 , y18015 , y18016 , y18017 , y18018 , y18019 , y18020 , y18021 , y18022 , y18023 , y18024 , y18025 , y18026 , y18027 , y18028 , y18029 , y18030 , y18031 , y18032 , y18033 , y18034 , y18035 , y18036 , y18037 , y18038 , y18039 , y18040 , y18041 , y18042 , y18043 , y18044 , y18045 , y18046 , y18047 , y18048 , y18049 , y18050 , y18051 , y18052 , y18053 , y18054 , y18055 , y18056 , y18057 , y18058 , y18059 , y18060 , y18061 , y18062 , y18063 , y18064 , y18065 , y18066 , y18067 , y18068 , y18069 , y18070 , y18071 , y18072 , y18073 , y18074 , y18075 , y18076 , y18077 , y18078 , y18079 , y18080 , y18081 , y18082 , y18083 , y18084 , y18085 , y18086 , y18087 , y18088 , y18089 , y18090 , y18091 , y18092 , y18093 , y18094 , y18095 , y18096 , y18097 , y18098 , y18099 , y18100 , y18101 , y18102 , y18103 , y18104 , y18105 , y18106 , y18107 , y18108 , y18109 , y18110 , y18111 , y18112 , y18113 , y18114 , y18115 , y18116 , y18117 , y18118 , y18119 , y18120 , y18121 , y18122 , y18123 , y18124 , y18125 , y18126 , y18127 , y18128 , y18129 , y18130 , y18131 , y18132 , y18133 , y18134 , y18135 , y18136 , y18137 , y18138 , y18139 , y18140 , y18141 , y18142 , y18143 , y18144 , y18145 , y18146 , y18147 , y18148 , y18149 , y18150 , y18151 , y18152 , y18153 , y18154 , y18155 , y18156 , y18157 , y18158 , y18159 , y18160 , y18161 , y18162 , y18163 , y18164 , y18165 , y18166 , y18167 , y18168 , y18169 , y18170 , y18171 , y18172 , y18173 , y18174 , y18175 , y18176 , y18177 , y18178 , y18179 , y18180 , y18181 , y18182 , y18183 , y18184 , y18185 , y18186 , y18187 , y18188 , y18189 , y18190 , y18191 , y18192 , y18193 , y18194 , y18195 , y18196 , y18197 , y18198 , y18199 , y18200 , y18201 , y18202 , y18203 , y18204 , y18205 , y18206 , y18207 , y18208 , y18209 , y18210 , y18211 , y18212 , y18213 , y18214 , y18215 , y18216 , y18217 , y18218 , y18219 , y18220 , y18221 , y18222 , y18223 , y18224 , y18225 , y18226 , y18227 , y18228 , y18229 , y18230 , y18231 , y18232 , y18233 , y18234 , y18235 , y18236 , y18237 , y18238 , y18239 , y18240 , y18241 , y18242 , y18243 , y18244 , y18245 , y18246 , y18247 , y18248 , y18249 , y18250 , y18251 , y18252 , y18253 , y18254 , y18255 , y18256 , y18257 , y18258 , y18259 , y18260 , y18261 , y18262 , y18263 , y18264 , y18265 , y18266 , y18267 , y18268 , y18269 , y18270 , y18271 , y18272 , y18273 , y18274 , y18275 , y18276 , y18277 , y18278 , y18279 , y18280 , y18281 , y18282 , y18283 , y18284 , y18285 , y18286 , y18287 , y18288 , y18289 , y18290 , y18291 , y18292 , y18293 , y18294 , y18295 , y18296 , y18297 , y18298 , y18299 , y18300 , y18301 , y18302 , y18303 , y18304 , y18305 , y18306 , y18307 , y18308 , y18309 , y18310 , y18311 , y18312 , y18313 , y18314 , y18315 , y18316 , y18317 , y18318 , y18319 , y18320 , y18321 , y18322 , y18323 , y18324 , y18325 , y18326 , y18327 , y18328 , y18329 , y18330 , y18331 , y18332 , y18333 , y18334 , y18335 , y18336 , y18337 , y18338 , y18339 , y18340 , y18341 , y18342 , y18343 , y18344 , y18345 , y18346 , y18347 , y18348 , y18349 , y18350 , y18351 , y18352 , y18353 , y18354 , y18355 , y18356 , y18357 , y18358 , y18359 , y18360 , y18361 , y18362 , y18363 , y18364 , y18365 , y18366 , y18367 , y18368 , y18369 , y18370 , y18371 , y18372 , y18373 , y18374 , y18375 , y18376 , y18377 , y18378 , y18379 , y18380 , y18381 , y18382 , y18383 , y18384 , y18385 , y18386 , y18387 , y18388 , y18389 , y18390 , y18391 , y18392 , y18393 , y18394 , y18395 , y18396 , y18397 , y18398 , y18399 , y18400 , y18401 , y18402 , y18403 , y18404 , y18405 , y18406 , y18407 , y18408 , y18409 , y18410 , y18411 , y18412 , y18413 , y18414 , y18415 , y18416 , y18417 , y18418 , y18419 , y18420 , y18421 , y18422 , y18423 , y18424 , y18425 , y18426 , y18427 , y18428 , y18429 , y18430 , y18431 , y18432 , y18433 , y18434 , y18435 , y18436 , y18437 , y18438 , y18439 , y18440 , y18441 , y18442 , y18443 , y18444 , y18445 , y18446 , y18447 , y18448 , y18449 , y18450 , y18451 , y18452 , y18453 , y18454 , y18455 , y18456 , y18457 , y18458 , y18459 , y18460 , y18461 , y18462 , y18463 , y18464 , y18465 , y18466 , y18467 , y18468 , y18469 , y18470 , y18471 , y18472 , y18473 , y18474 , y18475 , y18476 , y18477 , y18478 , y18479 , y18480 , y18481 , y18482 , y18483 , y18484 , y18485 , y18486 , y18487 , y18488 , y18489 , y18490 , y18491 , y18492 , y18493 , y18494 , y18495 , y18496 , y18497 , y18498 , y18499 , y18500 , y18501 , y18502 , y18503 , y18504 , y18505 , y18506 , y18507 , y18508 , y18509 , y18510 , y18511 , y18512 , y18513 , y18514 , y18515 , y18516 , y18517 , y18518 , y18519 , y18520 , y18521 , y18522 , y18523 , y18524 , y18525 , y18526 , y18527 , y18528 , y18529 , y18530 , y18531 , y18532 , y18533 , y18534 , y18535 , y18536 , y18537 , y18538 , y18539 , y18540 , y18541 , y18542 , y18543 , y18544 , y18545 , y18546 , y18547 , y18548 , y18549 , y18550 , y18551 , y18552 , y18553 , y18554 , y18555 , y18556 , y18557 , y18558 , y18559 , y18560 , y18561 , y18562 , y18563 , y18564 , y18565 , y18566 , y18567 , y18568 , y18569 , y18570 , y18571 , y18572 , y18573 , y18574 , y18575 , y18576 , y18577 , y18578 , y18579 , y18580 , y18581 , y18582 , y18583 , y18584 , y18585 , y18586 , y18587 , y18588 , y18589 , y18590 , y18591 , y18592 , y18593 , y18594 , y18595 , y18596 , y18597 , y18598 , y18599 , y18600 , y18601 , y18602 , y18603 , y18604 , y18605 , y18606 , y18607 , y18608 , y18609 , y18610 , y18611 , y18612 , y18613 , y18614 , y18615 , y18616 , y18617 , y18618 , y18619 , y18620 , y18621 , y18622 , y18623 , y18624 , y18625 , y18626 , y18627 , y18628 , y18629 , y18630 , y18631 , y18632 , y18633 , y18634 , y18635 , y18636 , y18637 , y18638 , y18639 , y18640 , y18641 , y18642 , y18643 , y18644 , y18645 , y18646 , y18647 , y18648 , y18649 , y18650 , y18651 , y18652 , y18653 , y18654 , y18655 , y18656 , y18657 , y18658 , y18659 , y18660 , y18661 , y18662 , y18663 , y18664 , y18665 , y18666 , y18667 , y18668 , y18669 , y18670 , y18671 , y18672 , y18673 , y18674 , y18675 , y18676 , y18677 , y18678 , y18679 , y18680 , y18681 , y18682 , y18683 , y18684 , y18685 , y18686 , y18687 , y18688 , y18689 , y18690 , y18691 , y18692 , y18693 , y18694 , y18695 , y18696 , y18697 , y18698 , y18699 , y18700 , y18701 , y18702 , y18703 , y18704 , y18705 , y18706 , y18707 , y18708 , y18709 , y18710 , y18711 , y18712 , y18713 , y18714 , y18715 , y18716 , y18717 , y18718 , y18719 , y18720 , y18721 , y18722 , y18723 , y18724 , y18725 , y18726 , y18727 , y18728 , y18729 , y18730 , y18731 , y18732 , y18733 , y18734 , y18735 , y18736 , y18737 , y18738 , y18739 , y18740 , y18741 , y18742 , y18743 , y18744 , y18745 , y18746 , y18747 , y18748 , y18749 , y18750 , y18751 , y18752 , y18753 , y18754 , y18755 , y18756 , y18757 , y18758 , y18759 , y18760 , y18761 , y18762 , y18763 , y18764 , y18765 , y18766 , y18767 , y18768 , y18769 , y18770 , y18771 , y18772 , y18773 , y18774 , y18775 , y18776 , y18777 , y18778 , y18779 , y18780 , y18781 , y18782 , y18783 , y18784 , y18785 , y18786 , y18787 , y18788 , y18789 , y18790 , y18791 , y18792 , y18793 , y18794 , y18795 , y18796 , y18797 , y18798 , y18799 , y18800 , y18801 , y18802 , y18803 , y18804 , y18805 , y18806 , y18807 , y18808 , y18809 , y18810 , y18811 , y18812 , y18813 , y18814 , y18815 , y18816 , y18817 , y18818 , y18819 , y18820 , y18821 , y18822 , y18823 , y18824 , y18825 , y18826 , y18827 , y18828 , y18829 , y18830 , y18831 , y18832 , y18833 , y18834 , y18835 , y18836 , y18837 , y18838 , y18839 , y18840 , y18841 , y18842 , y18843 , y18844 , y18845 , y18846 , y18847 , y18848 , y18849 , y18850 , y18851 , y18852 , y18853 , y18854 , y18855 , y18856 , y18857 , y18858 , y18859 , y18860 , y18861 , y18862 , y18863 , y18864 , y18865 , y18866 , y18867 , y18868 , y18869 , y18870 , y18871 , y18872 , y18873 , y18874 , y18875 , y18876 , y18877 , y18878 , y18879 , y18880 , y18881 , y18882 , y18883 , y18884 , y18885 , y18886 , y18887 , y18888 , y18889 , y18890 , y18891 , y18892 , y18893 , y18894 , y18895 , y18896 , y18897 , y18898 , y18899 , y18900 , y18901 , y18902 , y18903 , y18904 , y18905 , y18906 , y18907 , y18908 , y18909 , y18910 , y18911 , y18912 , y18913 , y18914 , y18915 , y18916 , y18917 , y18918 , y18919 , y18920 , y18921 , y18922 , y18923 , y18924 , y18925 , y18926 , y18927 , y18928 , y18929 , y18930 , y18931 , y18932 , y18933 , y18934 , y18935 , y18936 , y18937 , y18938 , y18939 , y18940 , y18941 , y18942 , y18943 , y18944 , y18945 , y18946 , y18947 , y18948 , y18949 , y18950 , y18951 , y18952 , y18953 , y18954 , y18955 , y18956 , y18957 , y18958 , y18959 , y18960 , y18961 , y18962 , y18963 , y18964 , y18965 , y18966 , y18967 , y18968 , y18969 , y18970 , y18971 , y18972 , y18973 , y18974 , y18975 , y18976 , y18977 , y18978 , y18979 , y18980 , y18981 , y18982 , y18983 , y18984 , y18985 , y18986 , y18987 , y18988 , y18989 , y18990 , y18991 , y18992 , y18993 , y18994 , y18995 , y18996 , y18997 , y18998 , y18999 , y19000 , y19001 , y19002 , y19003 , y19004 , y19005 , y19006 , y19007 , y19008 , y19009 , y19010 , y19011 , y19012 , y19013 , y19014 , y19015 , y19016 , y19017 , y19018 , y19019 , y19020 , y19021 , y19022 , y19023 , y19024 , y19025 , y19026 , y19027 , y19028 , y19029 , y19030 , y19031 , y19032 , y19033 , y19034 , y19035 , y19036 , y19037 , y19038 , y19039 , y19040 , y19041 , y19042 , y19043 , y19044 , y19045 , y19046 , y19047 , y19048 , y19049 , y19050 , y19051 , y19052 , y19053 , y19054 , y19055 , y19056 , y19057 , y19058 , y19059 , y19060 , y19061 , y19062 , y19063 , y19064 , y19065 , y19066 , y19067 , y19068 , y19069 , y19070 , y19071 , y19072 , y19073 , y19074 , y19075 , y19076 , y19077 , y19078 , y19079 , y19080 , y19081 , y19082 , y19083 , y19084 , y19085 , y19086 , y19087 , y19088 , y19089 , y19090 , y19091 , y19092 , y19093 , y19094 , y19095 , y19096 , y19097 , y19098 , y19099 , y19100 , y19101 , y19102 , y19103 , y19104 , y19105 , y19106 , y19107 , y19108 , y19109 , y19110 , y19111 , y19112 , y19113 , y19114 , y19115 , y19116 , y19117 , y19118 , y19119 , y19120 , y19121 , y19122 , y19123 , y19124 , y19125 , y19126 , y19127 , y19128 , y19129 , y19130 , y19131 , y19132 , y19133 , y19134 , y19135 , y19136 , y19137 , y19138 , y19139 , y19140 , y19141 , y19142 , y19143 , y19144 , y19145 , y19146 , y19147 , y19148 , y19149 , y19150 , y19151 , y19152 , y19153 , y19154 , y19155 , y19156 , y19157 , y19158 , y19159 , y19160 , y19161 , y19162 , y19163 , y19164 , y19165 , y19166 , y19167 , y19168 , y19169 , y19170 , y19171 , y19172 , y19173 , y19174 , y19175 , y19176 , y19177 , y19178 , y19179 , y19180 , y19181 , y19182 , y19183 , y19184 , y19185 , y19186 , y19187 , y19188 , y19189 , y19190 , y19191 , y19192 , y19193 , y19194 , y19195 , y19196 , y19197 , y19198 , y19199 , y19200 , y19201 , y19202 , y19203 , y19204 , y19205 , y19206 , y19207 , y19208 , y19209 , y19210 , y19211 , y19212 , y19213 , y19214 , y19215 , y19216 , y19217 , y19218 , y19219 , y19220 , y19221 , y19222 , y19223 , y19224 , y19225 , y19226 , y19227 , y19228 , y19229 , y19230 , y19231 , y19232 , y19233 , y19234 , y19235 , y19236 , y19237 , y19238 , y19239 , y19240 , y19241 , y19242 , y19243 , y19244 , y19245 , y19246 , y19247 , y19248 , y19249 , y19250 , y19251 , y19252 , y19253 , y19254 , y19255 , y19256 , y19257 , y19258 , y19259 , y19260 , y19261 , y19262 , y19263 , y19264 , y19265 , y19266 , y19267 , y19268 , y19269 , y19270 , y19271 , y19272 , y19273 , y19274 , y19275 , y19276 , y19277 , y19278 , y19279 , y19280 , y19281 , y19282 , y19283 , y19284 , y19285 , y19286 , y19287 , y19288 , y19289 , y19290 , y19291 , y19292 , y19293 , y19294 , y19295 , y19296 , y19297 , y19298 , y19299 , y19300 , y19301 , y19302 , y19303 , y19304 , y19305 , y19306 , y19307 , y19308 , y19309 , y19310 , y19311 , y19312 , y19313 , y19314 , y19315 , y19316 , y19317 , y19318 , y19319 , y19320 , y19321 , y19322 , y19323 , y19324 , y19325 , y19326 , y19327 , y19328 , y19329 , y19330 , y19331 , y19332 , y19333 , y19334 , y19335 , y19336 , y19337 , y19338 , y19339 , y19340 , y19341 , y19342 , y19343 , y19344 , y19345 , y19346 , y19347 , y19348 , y19349 , y19350 , y19351 , y19352 , y19353 , y19354 , y19355 , y19356 , y19357 , y19358 , y19359 , y19360 , y19361 , y19362 , y19363 , y19364 , y19365 , y19366 , y19367 , y19368 , y19369 , y19370 , y19371 , y19372 , y19373 , y19374 , y19375 , y19376 , y19377 , y19378 , y19379 , y19380 , y19381 , y19382 , y19383 , y19384 , y19385 , y19386 , y19387 , y19388 , y19389 , y19390 , y19391 , y19392 , y19393 , y19394 , y19395 , y19396 , y19397 , y19398 , y19399 , y19400 , y19401 , y19402 , y19403 , y19404 , y19405 , y19406 , y19407 , y19408 , y19409 , y19410 , y19411 , y19412 , y19413 , y19414 , y19415 , y19416 , y19417 , y19418 , y19419 , y19420 , y19421 , y19422 , y19423 , y19424 , y19425 , y19426 , y19427 , y19428 , y19429 , y19430 , y19431 , y19432 , y19433 , y19434 , y19435 , y19436 , y19437 , y19438 , y19439 , y19440 , y19441 , y19442 , y19443 , y19444 , y19445 , y19446 , y19447 , y19448 , y19449 , y19450 , y19451 , y19452 , y19453 , y19454 , y19455 , y19456 , y19457 , y19458 , y19459 , y19460 , y19461 , y19462 , y19463 , y19464 , y19465 , y19466 , y19467 , y19468 , y19469 , y19470 , y19471 , y19472 , y19473 , y19474 , y19475 , y19476 , y19477 , y19478 , y19479 , y19480 , y19481 , y19482 , y19483 , y19484 , y19485 , y19486 , y19487 , y19488 , y19489 , y19490 , y19491 , y19492 , y19493 , y19494 , y19495 , y19496 , y19497 , y19498 , y19499 , y19500 , y19501 , y19502 , y19503 , y19504 , y19505 , y19506 , y19507 , y19508 , y19509 , y19510 , y19511 , y19512 , y19513 , y19514 , y19515 , y19516 , y19517 , y19518 , y19519 , y19520 , y19521 , y19522 , y19523 , y19524 , y19525 , y19526 , y19527 , y19528 , y19529 , y19530 , y19531 , y19532 , y19533 , y19534 , y19535 , y19536 , y19537 , y19538 , y19539 , y19540 , y19541 , y19542 , y19543 , y19544 , y19545 , y19546 , y19547 , y19548 , y19549 , y19550 , y19551 , y19552 , y19553 , y19554 , y19555 , y19556 , y19557 , y19558 , y19559 , y19560 , y19561 , y19562 , y19563 , y19564 , y19565 , y19566 , y19567 , y19568 , y19569 , y19570 , y19571 , y19572 , y19573 , y19574 , y19575 , y19576 , y19577 , y19578 , y19579 , y19580 , y19581 , y19582 , y19583 , y19584 , y19585 , y19586 , y19587 , y19588 , y19589 , y19590 , y19591 , y19592 , y19593 , y19594 , y19595 , y19596 , y19597 , y19598 , y19599 , y19600 , y19601 , y19602 , y19603 , y19604 , y19605 , y19606 , y19607 , y19608 , y19609 , y19610 , y19611 , y19612 , y19613 , y19614 , y19615 , y19616 , y19617 , y19618 , y19619 , y19620 , y19621 , y19622 , y19623 , y19624 , y19625 , y19626 , y19627 , y19628 , y19629 , y19630 , y19631 , y19632 , y19633 , y19634 , y19635 , y19636 , y19637 , y19638 , y19639 , y19640 , y19641 , y19642 , y19643 , y19644 , y19645 , y19646 , y19647 , y19648 , y19649 , y19650 , y19651 , y19652 , y19653 , y19654 , y19655 , y19656 , y19657 , y19658 , y19659 , y19660 , y19661 , y19662 , y19663 , y19664 , y19665 , y19666 , y19667 , y19668 , y19669 , y19670 , y19671 , y19672 , y19673 , y19674 , y19675 , y19676 , y19677 , y19678 , y19679 , y19680 , y19681 , y19682 , y19683 , y19684 , y19685 , y19686 , y19687 , y19688 , y19689 , y19690 , y19691 , y19692 , y19693 , y19694 , y19695 , y19696 , y19697 , y19698 , y19699 , y19700 , y19701 , y19702 , y19703 , y19704 , y19705 , y19706 , y19707 , y19708 , y19709 , y19710 , y19711 , y19712 , y19713 , y19714 , y19715 , y19716 , y19717 , y19718 , y19719 , y19720 , y19721 , y19722 , y19723 , y19724 , y19725 , y19726 , y19727 , y19728 , y19729 , y19730 , y19731 , y19732 , y19733 , y19734 , y19735 , y19736 , y19737 , y19738 , y19739 , y19740 , y19741 , y19742 , y19743 , y19744 , y19745 , y19746 , y19747 , y19748 , y19749 , y19750 , y19751 , y19752 , y19753 , y19754 , y19755 , y19756 , y19757 , y19758 , y19759 , y19760 , y19761 , y19762 , y19763 , y19764 , y19765 , y19766 , y19767 , y19768 , y19769 , y19770 , y19771 , y19772 , y19773 , y19774 , y19775 , y19776 , y19777 , y19778 , y19779 , y19780 , y19781 , y19782 , y19783 , y19784 , y19785 , y19786 , y19787 , y19788 , y19789 , y19790 , y19791 , y19792 , y19793 , y19794 , y19795 , y19796 , y19797 , y19798 , y19799 , y19800 , y19801 , y19802 , y19803 , y19804 , y19805 , y19806 , y19807 , y19808 , y19809 , y19810 , y19811 , y19812 , y19813 , y19814 , y19815 , y19816 , y19817 , y19818 , y19819 , y19820 , y19821 , y19822 , y19823 , y19824 , y19825 , y19826 , y19827 , y19828 , y19829 , y19830 , y19831 , y19832 , y19833 , y19834 , y19835 , y19836 , y19837 , y19838 , y19839 , y19840 , y19841 , y19842 , y19843 , y19844 , y19845 , y19846 , y19847 , y19848 , y19849 , y19850 , y19851 , y19852 , y19853 , y19854 , y19855 , y19856 , y19857 , y19858 , y19859 , y19860 , y19861 , y19862 , y19863 , y19864 , y19865 , y19866 , y19867 , y19868 , y19869 , y19870 , y19871 , y19872 , y19873 , y19874 , y19875 , y19876 , y19877 , y19878 , y19879 , y19880 , y19881 , y19882 , y19883 , y19884 , y19885 , y19886 , y19887 , y19888 , y19889 , y19890 , y19891 , y19892 , y19893 , y19894 , y19895 , y19896 , y19897 , y19898 , y19899 , y19900 , y19901 , y19902 , y19903 , y19904 , y19905 , y19906 , y19907 , y19908 , y19909 , y19910 , y19911 , y19912 , y19913 , y19914 , y19915 , y19916 , y19917 , y19918 , y19919 , y19920 , y19921 , y19922 , y19923 , y19924 , y19925 , y19926 , y19927 , y19928 , y19929 , y19930 , y19931 , y19932 , y19933 , y19934 , y19935 , y19936 , y19937 , y19938 , y19939 , y19940 , y19941 , y19942 , y19943 , y19944 , y19945 , y19946 , y19947 , y19948 , y19949 , y19950 , y19951 , y19952 , y19953 , y19954 , y19955 , y19956 , y19957 , y19958 , y19959 , y19960 , y19961 , y19962 , y19963 , y19964 , y19965 , y19966 , y19967 , y19968 , y19969 , y19970 , y19971 , y19972 , y19973 , y19974 , y19975 , y19976 , y19977 , y19978 , y19979 , y19980 , y19981 , y19982 , y19983 , y19984 , y19985 , y19986 , y19987 , y19988 , y19989 , y19990 , y19991 , y19992 , y19993 , y19994 , y19995 , y19996 , y19997 , y19998 , y19999 , y20000 , y20001 , y20002 , y20003 , y20004 , y20005 , y20006 , y20007 , y20008 , y20009 , y20010 , y20011 , y20012 , y20013 , y20014 , y20015 , y20016 , y20017 , y20018 , y20019 , y20020 , y20021 , y20022 , y20023 , y20024 , y20025 , y20026 , y20027 , y20028 , y20029 , y20030 , y20031 , y20032 , y20033 , y20034 , y20035 , y20036 , y20037 , y20038 , y20039 , y20040 , y20041 , y20042 , y20043 , y20044 , y20045 , y20046 , y20047 , y20048 , y20049 , y20050 , y20051 , y20052 , y20053 , y20054 , y20055 , y20056 , y20057 , y20058 , y20059 , y20060 , y20061 , y20062 , y20063 , y20064 , y20065 , y20066 , y20067 , y20068 , y20069 , y20070 , y20071 , y20072 , y20073 , y20074 , y20075 , y20076 , y20077 , y20078 , y20079 , y20080 , y20081 , y20082 , y20083 , y20084 , y20085 , y20086 , y20087 , y20088 , y20089 , y20090 , y20091 , y20092 , y20093 , y20094 , y20095 , y20096 , y20097 , y20098 , y20099 , y20100 , y20101 , y20102 , y20103 , y20104 , y20105 , y20106 , y20107 , y20108 , y20109 , y20110 , y20111 , y20112 , y20113 , y20114 , y20115 , y20116 , y20117 , y20118 , y20119 , y20120 , y20121 , y20122 , y20123 , y20124 , y20125 , y20126 , y20127 , y20128 , y20129 , y20130 , y20131 , y20132 , y20133 , y20134 , y20135 , y20136 , y20137 , y20138 , y20139 , y20140 , y20141 , y20142 , y20143 , y20144 , y20145 , y20146 , y20147 , y20148 , y20149 , y20150 , y20151 , y20152 , y20153 , y20154 , y20155 , y20156 , y20157 , y20158 , y20159 , y20160 , y20161 , y20162 , y20163 , y20164 , y20165 , y20166 , y20167 , y20168 , y20169 , y20170 , y20171 , y20172 , y20173 , y20174 , y20175 , y20176 , y20177 , y20178 , y20179 , y20180 , y20181 , y20182 , y20183 , y20184 , y20185 , y20186 , y20187 , y20188 , y20189 , y20190 , y20191 , y20192 , y20193 , y20194 , y20195 , y20196 , y20197 , y20198 , y20199 , y20200 , y20201 , y20202 , y20203 , y20204 , y20205 , y20206 , y20207 , y20208 , y20209 , y20210 , y20211 , y20212 , y20213 , y20214 , y20215 , y20216 , y20217 , y20218 , y20219 , y20220 , y20221 , y20222 , y20223 , y20224 , y20225 , y20226 , y20227 , y20228 , y20229 , y20230 , y20231 , y20232 , y20233 , y20234 , y20235 , y20236 , y20237 , y20238 , y20239 , y20240 , y20241 , y20242 , y20243 , y20244 , y20245 , y20246 , y20247 , y20248 , y20249 , y20250 , y20251 , y20252 , y20253 , y20254 , y20255 , y20256 , y20257 , y20258 , y20259 , y20260 , y20261 , y20262 , y20263 , y20264 , y20265 , y20266 , y20267 , y20268 , y20269 , y20270 , y20271 , y20272 , y20273 , y20274 , y20275 , y20276 , y20277 , y20278 , y20279 , y20280 , y20281 , y20282 , y20283 , y20284 , y20285 , y20286 , y20287 , y20288 , y20289 , y20290 , y20291 , y20292 , y20293 , y20294 , y20295 , y20296 , y20297 , y20298 , y20299 , y20300 , y20301 , y20302 , y20303 , y20304 , y20305 , y20306 , y20307 , y20308 , y20309 , y20310 , y20311 , y20312 , y20313 , y20314 , y20315 , y20316 , y20317 , y20318 , y20319 , y20320 , y20321 , y20322 , y20323 , y20324 , y20325 , y20326 , y20327 , y20328 , y20329 , y20330 , y20331 , y20332 , y20333 , y20334 , y20335 , y20336 , y20337 , y20338 , y20339 , y20340 , y20341 , y20342 , y20343 , y20344 , y20345 , y20346 , y20347 , y20348 , y20349 , y20350 , y20351 , y20352 , y20353 , y20354 , y20355 , y20356 , y20357 , y20358 , y20359 , y20360 , y20361 , y20362 , y20363 , y20364 , y20365 , y20366 , y20367 , y20368 , y20369 , y20370 , y20371 , y20372 , y20373 , y20374 , y20375 , y20376 , y20377 , y20378 , y20379 , y20380 , y20381 , y20382 , y20383 , y20384 , y20385 , y20386 , y20387 , y20388 , y20389 , y20390 , y20391 , y20392 , y20393 , y20394 , y20395 , y20396 , y20397 , y20398 , y20399 , y20400 , y20401 , y20402 , y20403 , y20404 , y20405 , y20406 , y20407 , y20408 , y20409 , y20410 , y20411 , y20412 , y20413 , y20414 , y20415 , y20416 , y20417 , y20418 , y20419 , y20420 , y20421 , y20422 , y20423 , y20424 , y20425 , y20426 , y20427 , y20428 , y20429 , y20430 , y20431 , y20432 , y20433 , y20434 , y20435 , y20436 , y20437 , y20438 , y20439 , y20440 , y20441 , y20442 , y20443 , y20444 , y20445 , y20446 , y20447 , y20448 , y20449 , y20450 , y20451 , y20452 , y20453 , y20454 , y20455 , y20456 , y20457 , y20458 , y20459 , y20460 , y20461 , y20462 , y20463 , y20464 , y20465 , y20466 , y20467 , y20468 , y20469 , y20470 , y20471 , y20472 , y20473 , y20474 , y20475 , y20476 , y20477 , y20478 , y20479 , y20480 , y20481 , y20482 , y20483 , y20484 , y20485 , y20486 , y20487 , y20488 , y20489 , y20490 , y20491 , y20492 , y20493 , y20494 , y20495 , y20496 , y20497 , y20498 , y20499 , y20500 , y20501 , y20502 , y20503 , y20504 , y20505 , y20506 , y20507 , y20508 , y20509 , y20510 , y20511 , y20512 , y20513 , y20514 , y20515 , y20516 , y20517 , y20518 , y20519 , y20520 , y20521 , y20522 , y20523 , y20524 , y20525 , y20526 , y20527 , y20528 , y20529 , y20530 , y20531 , y20532 , y20533 , y20534 , y20535 , y20536 , y20537 , y20538 , y20539 , y20540 , y20541 , y20542 , y20543 , y20544 , y20545 , y20546 , y20547 , y20548 , y20549 , y20550 , y20551 , y20552 , y20553 , y20554 , y20555 , y20556 , y20557 , y20558 , y20559 , y20560 , y20561 , y20562 , y20563 , y20564 , y20565 , y20566 , y20567 , y20568 , y20569 , y20570 , y20571 , y20572 , y20573 , y20574 , y20575 , y20576 , y20577 , y20578 , y20579 , y20580 , y20581 , y20582 , y20583 , y20584 , y20585 , y20586 , y20587 , y20588 , y20589 , y20590 , y20591 , y20592 , y20593 , y20594 , y20595 , y20596 , y20597 , y20598 , y20599 , y20600 , y20601 , y20602 , y20603 , y20604 , y20605 , y20606 , y20607 , y20608 , y20609 , y20610 , y20611 , y20612 , y20613 , y20614 , y20615 , y20616 , y20617 , y20618 , y20619 , y20620 , y20621 , y20622 , y20623 , y20624 , y20625 , y20626 , y20627 , y20628 , y20629 , y20630 , y20631 , y20632 , y20633 , y20634 , y20635 , y20636 , y20637 , y20638 , y20639 , y20640 , y20641 , y20642 , y20643 , y20644 , y20645 , y20646 , y20647 , y20648 , y20649 , y20650 , y20651 , y20652 , y20653 , y20654 , y20655 , y20656 , y20657 , y20658 , y20659 , y20660 , y20661 , y20662 , y20663 , y20664 , y20665 , y20666 , y20667 , y20668 , y20669 , y20670 , y20671 , y20672 , y20673 , y20674 , y20675 , y20676 , y20677 , y20678 , y20679 , y20680 , y20681 , y20682 , y20683 , y20684 , y20685 , y20686 , y20687 , y20688 , y20689 , y20690 , y20691 , y20692 , y20693 , y20694 , y20695 , y20696 , y20697 , y20698 , y20699 , y20700 , y20701 , y20702 , y20703 , y20704 , y20705 , y20706 , y20707 , y20708 , y20709 , y20710 , y20711 , y20712 , y20713 , y20714 , y20715 , y20716 , y20717 , y20718 , y20719 , y20720 , y20721 , y20722 , y20723 , y20724 , y20725 , y20726 , y20727 , y20728 , y20729 , y20730 , y20731 , y20732 , y20733 , y20734 , y20735 , y20736 , y20737 , y20738 , y20739 , y20740 , y20741 , y20742 , y20743 , y20744 , y20745 , y20746 , y20747 , y20748 , y20749 , y20750 , y20751 , y20752 , y20753 , y20754 , y20755 , y20756 , y20757 , y20758 , y20759 , y20760 , y20761 , y20762 , y20763 , y20764 , y20765 , y20766 , y20767 , y20768 , y20769 , y20770 , y20771 , y20772 , y20773 , y20774 , y20775 , y20776 , y20777 , y20778 , y20779 , y20780 , y20781 , y20782 , y20783 , y20784 , y20785 , y20786 , y20787 , y20788 , y20789 , y20790 , y20791 , y20792 , y20793 , y20794 , y20795 , y20796 , y20797 , y20798 , y20799 , y20800 , y20801 , y20802 , y20803 , y20804 , y20805 , y20806 , y20807 , y20808 , y20809 , y20810 , y20811 , y20812 , y20813 , y20814 , y20815 , y20816 , y20817 , y20818 , y20819 , y20820 , y20821 , y20822 , y20823 , y20824 , y20825 , y20826 , y20827 , y20828 , y20829 , y20830 , y20831 , y20832 , y20833 , y20834 , y20835 , y20836 , y20837 , y20838 , y20839 , y20840 , y20841 , y20842 , y20843 , y20844 , y20845 , y20846 , y20847 , y20848 , y20849 , y20850 , y20851 , y20852 , y20853 , y20854 , y20855 , y20856 , y20857 , y20858 , y20859 , y20860 , y20861 , y20862 , y20863 , y20864 , y20865 , y20866 , y20867 , y20868 , y20869 , y20870 , y20871 , y20872 , y20873 , y20874 , y20875 , y20876 , y20877 , y20878 , y20879 , y20880 , y20881 , y20882 , y20883 , y20884 , y20885 , y20886 , y20887 , y20888 , y20889 , y20890 , y20891 , y20892 , y20893 , y20894 , y20895 , y20896 , y20897 , y20898 , y20899 , y20900 , y20901 , y20902 , y20903 , y20904 , y20905 , y20906 , y20907 , y20908 , y20909 , y20910 , y20911 , y20912 , y20913 , y20914 , y20915 , y20916 , y20917 , y20918 , y20919 , y20920 , y20921 , y20922 , y20923 , y20924 , y20925 , y20926 , y20927 , y20928 , y20929 , y20930 , y20931 , y20932 , y20933 , y20934 , y20935 , y20936 , y20937 , y20938 , y20939 , y20940 , y20941 , y20942 , y20943 , y20944 , y20945 , y20946 , y20947 , y20948 , y20949 , y20950 , y20951 , y20952 , y20953 , y20954 , y20955 , y20956 , y20957 , y20958 , y20959 , y20960 , y20961 , y20962 , y20963 , y20964 , y20965 , y20966 , y20967 , y20968 , y20969 , y20970 , y20971 , y20972 , y20973 , y20974 , y20975 , y20976 , y20977 , y20978 , y20979 , y20980 , y20981 , y20982 , y20983 , y20984 , y20985 , y20986 , y20987 , y20988 , y20989 , y20990 , y20991 , y20992 , y20993 , y20994 , y20995 , y20996 , y20997 , y20998 , y20999 , y21000 , y21001 , y21002 , y21003 , y21004 , y21005 , y21006 , y21007 , y21008 , y21009 , y21010 , y21011 , y21012 , y21013 , y21014 , y21015 , y21016 , y21017 , y21018 , y21019 , y21020 , y21021 , y21022 , y21023 , y21024 , y21025 , y21026 , y21027 , y21028 , y21029 , y21030 , y21031 , y21032 , y21033 , y21034 , y21035 , y21036 , y21037 , y21038 , y21039 , y21040 , y21041 , y21042 , y21043 , y21044 , y21045 , y21046 , y21047 , y21048 , y21049 , y21050 , y21051 , y21052 , y21053 , y21054 , y21055 , y21056 , y21057 , y21058 , y21059 , y21060 , y21061 , y21062 , y21063 , y21064 , y21065 , y21066 , y21067 , y21068 , y21069 , y21070 , y21071 , y21072 , y21073 , y21074 , y21075 , y21076 , y21077 , y21078 , y21079 , y21080 , y21081 , y21082 , y21083 , y21084 , y21085 , y21086 , y21087 , y21088 , y21089 , y21090 , y21091 , y21092 , y21093 , y21094 , y21095 , y21096 , y21097 , y21098 , y21099 , y21100 , y21101 , y21102 , y21103 , y21104 , y21105 , y21106 , y21107 , y21108 , y21109 , y21110 , y21111 , y21112 , y21113 , y21114 , y21115 , y21116 , y21117 , y21118 , y21119 , y21120 , y21121 , y21122 , y21123 , y21124 , y21125 , y21126 , y21127 , y21128 , y21129 , y21130 , y21131 , y21132 , y21133 , y21134 , y21135 , y21136 , y21137 , y21138 , y21139 , y21140 , y21141 , y21142 , y21143 , y21144 , y21145 , y21146 , y21147 , y21148 , y21149 , y21150 , y21151 , y21152 , y21153 , y21154 , y21155 , y21156 , y21157 , y21158 , y21159 , y21160 , y21161 , y21162 , y21163 , y21164 , y21165 , y21166 , y21167 , y21168 , y21169 , y21170 , y21171 , y21172 , y21173 , y21174 , y21175 , y21176 , y21177 , y21178 , y21179 , y21180 , y21181 , y21182 , y21183 , y21184 , y21185 , y21186 , y21187 , y21188 , y21189 , y21190 , y21191 , y21192 , y21193 , y21194 , y21195 , y21196 , y21197 , y21198 , y21199 , y21200 , y21201 , y21202 , y21203 , y21204 , y21205 , y21206 , y21207 , y21208 , y21209 , y21210 , y21211 , y21212 , y21213 , y21214 , y21215 , y21216 , y21217 , y21218 , y21219 , y21220 , y21221 , y21222 , y21223 , y21224 , y21225 , y21226 , y21227 , y21228 , y21229 , y21230 , y21231 , y21232 , y21233 , y21234 , y21235 , y21236 , y21237 , y21238 , y21239 , y21240 , y21241 , y21242 , y21243 , y21244 , y21245 , y21246 , y21247 , y21248 , y21249 , y21250 , y21251 , y21252 , y21253 , y21254 , y21255 , y21256 , y21257 , y21258 , y21259 , y21260 , y21261 , y21262 , y21263 , y21264 , y21265 , y21266 , y21267 , y21268 , y21269 , y21270 , y21271 , y21272 , y21273 , y21274 , y21275 , y21276 , y21277 , y21278 , y21279 , y21280 , y21281 , y21282 , y21283 , y21284 , y21285 , y21286 , y21287 , y21288 , y21289 , y21290 , y21291 , y21292 , y21293 , y21294 , y21295 , y21296 , y21297 , y21298 , y21299 , y21300 , y21301 , y21302 , y21303 , y21304 , y21305 , y21306 , y21307 , y21308 , y21309 , y21310 , y21311 , y21312 , y21313 , y21314 , y21315 , y21316 , y21317 , y21318 , y21319 , y21320 , y21321 , y21322 , y21323 , y21324 , y21325 , y21326 , y21327 , y21328 , y21329 , y21330 , y21331 , y21332 , y21333 , y21334 , y21335 , y21336 , y21337 , y21338 , y21339 , y21340 , y21341 , y21342 , y21343 , y21344 , y21345 , y21346 , y21347 , y21348 , y21349 , y21350 , y21351 , y21352 , y21353 , y21354 , y21355 , y21356 , y21357 , y21358 , y21359 , y21360 , y21361 , y21362 , y21363 , y21364 , y21365 , y21366 , y21367 , y21368 , y21369 , y21370 , y21371 , y21372 , y21373 , y21374 , y21375 , y21376 , y21377 , y21378 , y21379 , y21380 , y21381 , y21382 , y21383 , y21384 , y21385 , y21386 , y21387 , y21388 , y21389 , y21390 , y21391 , y21392 , y21393 , y21394 , y21395 , y21396 , y21397 , y21398 , y21399 , y21400 , y21401 , y21402 , y21403 , y21404 , y21405 , y21406 , y21407 , y21408 , y21409 , y21410 , y21411 , y21412 , y21413 , y21414 , y21415 , y21416 , y21417 , y21418 , y21419 , y21420 , y21421 , y21422 , y21423 , y21424 , y21425 , y21426 , y21427 , y21428 , y21429 , y21430 , y21431 , y21432 , y21433 , y21434 , y21435 , y21436 , y21437 , y21438 , y21439 , y21440 , y21441 , y21442 , y21443 , y21444 , y21445 , y21446 , y21447 , y21448 , y21449 , y21450 , y21451 , y21452 , y21453 , y21454 , y21455 , y21456 , y21457 , y21458 , y21459 , y21460 , y21461 , y21462 , y21463 , y21464 , y21465 , y21466 , y21467 , y21468 , y21469 , y21470 , y21471 , y21472 , y21473 , y21474 , y21475 , y21476 , y21477 , y21478 , y21479 , y21480 , y21481 , y21482 , y21483 , y21484 , y21485 , y21486 , y21487 , y21488 , y21489 , y21490 , y21491 , y21492 , y21493 , y21494 , y21495 , y21496 , y21497 , y21498 , y21499 , y21500 , y21501 , y21502 , y21503 , y21504 , y21505 , y21506 , y21507 , y21508 , y21509 , y21510 , y21511 , y21512 , y21513 , y21514 , y21515 , y21516 , y21517 , y21518 , y21519 , y21520 , y21521 , y21522 , y21523 , y21524 , y21525 , y21526 , y21527 , y21528 , y21529 , y21530 , y21531 , y21532 , y21533 , y21534 , y21535 , y21536 , y21537 , y21538 , y21539 , y21540 , y21541 , y21542 , y21543 , y21544 , y21545 , y21546 , y21547 , y21548 , y21549 , y21550 , y21551 , y21552 , y21553 , y21554 , y21555 , y21556 , y21557 , y21558 , y21559 , y21560 , y21561 , y21562 , y21563 , y21564 , y21565 , y21566 , y21567 , y21568 , y21569 , y21570 , y21571 , y21572 , y21573 , y21574 , y21575 , y21576 , y21577 , y21578 , y21579 , y21580 , y21581 , y21582 , y21583 , y21584 , y21585 , y21586 , y21587 , y21588 , y21589 , y21590 , y21591 , y21592 , y21593 , y21594 , y21595 , y21596 , y21597 , y21598 , y21599 , y21600 , y21601 , y21602 , y21603 , y21604 , y21605 , y21606 , y21607 , y21608 , y21609 , y21610 , y21611 , y21612 , y21613 , y21614 , y21615 , y21616 , y21617 , y21618 , y21619 , y21620 , y21621 , y21622 , y21623 , y21624 , y21625 , y21626 , y21627 , y21628 , y21629 , y21630 , y21631 , y21632 , y21633 , y21634 , y21635 , y21636 , y21637 , y21638 , y21639 , y21640 , y21641 , y21642 , y21643 , y21644 , y21645 , y21646 , y21647 , y21648 , y21649 , y21650 , y21651 , y21652 , y21653 , y21654 , y21655 , y21656 , y21657 , y21658 , y21659 , y21660 , y21661 , y21662 , y21663 , y21664 , y21665 , y21666 , y21667 , y21668 , y21669 , y21670 , y21671 , y21672 , y21673 , y21674 , y21675 , y21676 , y21677 , y21678 , y21679 , y21680 , y21681 , y21682 , y21683 , y21684 , y21685 , y21686 , y21687 , y21688 , y21689 , y21690 , y21691 , y21692 , y21693 , y21694 , y21695 , y21696 , y21697 , y21698 , y21699 , y21700 , y21701 , y21702 , y21703 , y21704 , y21705 , y21706 , y21707 , y21708 , y21709 , y21710 , y21711 , y21712 , y21713 , y21714 , y21715 , y21716 , y21717 , y21718 , y21719 , y21720 , y21721 , y21722 , y21723 , y21724 , y21725 , y21726 , y21727 , y21728 , y21729 , y21730 , y21731 , y21732 , y21733 , y21734 , y21735 , y21736 , y21737 , y21738 , y21739 , y21740 , y21741 , y21742 , y21743 , y21744 , y21745 , y21746 , y21747 , y21748 , y21749 , y21750 , y21751 , y21752 , y21753 , y21754 , y21755 , y21756 , y21757 , y21758 , y21759 , y21760 , y21761 , y21762 , y21763 , y21764 , y21765 , y21766 , y21767 , y21768 , y21769 , y21770 , y21771 , y21772 , y21773 , y21774 , y21775 , y21776 , y21777 , y21778 , y21779 , y21780 , y21781 , y21782 , y21783 , y21784 , y21785 , y21786 , y21787 , y21788 , y21789 , y21790 , y21791 , y21792 , y21793 , y21794 , y21795 , y21796 , y21797 , y21798 , y21799 , y21800 , y21801 , y21802 , y21803 , y21804 , y21805 , y21806 , y21807 , y21808 , y21809 , y21810 , y21811 , y21812 , y21813 , y21814 , y21815 , y21816 , y21817 , y21818 , y21819 , y21820 , y21821 , y21822 , y21823 , y21824 , y21825 , y21826 , y21827 , y21828 , y21829 , y21830 , y21831 , y21832 , y21833 , y21834 , y21835 , y21836 , y21837 , y21838 , y21839 , y21840 , y21841 , y21842 , y21843 , y21844 , y21845 , y21846 , y21847 , y21848 , y21849 , y21850 , y21851 , y21852 , y21853 , y21854 , y21855 , y21856 , y21857 , y21858 , y21859 , y21860 , y21861 , y21862 , y21863 , y21864 , y21865 , y21866 , y21867 , y21868 , y21869 , y21870 , y21871 , y21872 , y21873 , y21874 , y21875 , y21876 , y21877 , y21878 , y21879 , y21880 , y21881 , y21882 , y21883 , y21884 , y21885 , y21886 , y21887 , y21888 , y21889 , y21890 , y21891 , y21892 , y21893 , y21894 , y21895 , y21896 , y21897 , y21898 , y21899 , y21900 , y21901 , y21902 , y21903 , y21904 , y21905 , y21906 , y21907 , y21908 , y21909 , y21910 , y21911 , y21912 , y21913 , y21914 , y21915 , y21916 , y21917 , y21918 , y21919 , y21920 , y21921 , y21922 , y21923 , y21924 , y21925 , y21926 , y21927 , y21928 , y21929 , y21930 , y21931 , y21932 , y21933 , y21934 , y21935 , y21936 , y21937 , y21938 , y21939 , y21940 , y21941 , y21942 , y21943 , y21944 , y21945 , y21946 , y21947 , y21948 , y21949 , y21950 , y21951 , y21952 , y21953 , y21954 , y21955 , y21956 , y21957 , y21958 , y21959 , y21960 , y21961 , y21962 , y21963 , y21964 , y21965 , y21966 , y21967 , y21968 , y21969 , y21970 , y21971 , y21972 , y21973 , y21974 , y21975 , y21976 , y21977 , y21978 , y21979 , y21980 , y21981 , y21982 , y21983 , y21984 , y21985 , y21986 , y21987 , y21988 , y21989 , y21990 , y21991 , y21992 , y21993 , y21994 , y21995 , y21996 , y21997 , y21998 , y21999 , y22000 , y22001 , y22002 , y22003 , y22004 , y22005 , y22006 , y22007 , y22008 , y22009 , y22010 , y22011 , y22012 , y22013 , y22014 , y22015 , y22016 , y22017 , y22018 , y22019 , y22020 , y22021 , y22022 , y22023 , y22024 , y22025 , y22026 , y22027 , y22028 , y22029 , y22030 , y22031 , y22032 , y22033 , y22034 , y22035 , y22036 , y22037 , y22038 , y22039 , y22040 , y22041 , y22042 , y22043 , y22044 , y22045 , y22046 , y22047 , y22048 , y22049 , y22050 , y22051 , y22052 , y22053 , y22054 , y22055 , y22056 , y22057 , y22058 , y22059 , y22060 , y22061 , y22062 , y22063 , y22064 , y22065 , y22066 , y22067 , y22068 , y22069 , y22070 , y22071 , y22072 , y22073 , y22074 , y22075 , y22076 , y22077 , y22078 , y22079 , y22080 , y22081 , y22082 , y22083 , y22084 , y22085 , y22086 , y22087 , y22088 , y22089 , y22090 , y22091 , y22092 , y22093 , y22094 , y22095 , y22096 , y22097 , y22098 , y22099 , y22100 , y22101 , y22102 , y22103 , y22104 , y22105 , y22106 , y22107 , y22108 , y22109 , y22110 , y22111 , y22112 , y22113 , y22114 , y22115 , y22116 , y22117 , y22118 , y22119 , y22120 , y22121 , y22122 , y22123 , y22124 , y22125 , y22126 , y22127 , y22128 , y22129 , y22130 , y22131 , y22132 , y22133 , y22134 , y22135 , y22136 , y22137 , y22138 , y22139 , y22140 , y22141 , y22142 , y22143 , y22144 , y22145 , y22146 , y22147 , y22148 , y22149 , y22150 , y22151 , y22152 , y22153 , y22154 , y22155 , y22156 , y22157 , y22158 , y22159 , y22160 , y22161 , y22162 , y22163 , y22164 , y22165 , y22166 , y22167 , y22168 , y22169 , y22170 , y22171 , y22172 , y22173 , y22174 , y22175 , y22176 , y22177 , y22178 , y22179 , y22180 , y22181 , y22182 , y22183 , y22184 , y22185 , y22186 , y22187 , y22188 , y22189 , y22190 , y22191 , y22192 , y22193 , y22194 , y22195 , y22196 , y22197 , y22198 , y22199 , y22200 , y22201 , y22202 , y22203 , y22204 , y22205 , y22206 , y22207 , y22208 , y22209 , y22210 , y22211 , y22212 , y22213 , y22214 , y22215 , y22216 , y22217 , y22218 , y22219 , y22220 , y22221 , y22222 , y22223 , y22224 , y22225 , y22226 , y22227 , y22228 , y22229 , y22230 , y22231 , y22232 , y22233 , y22234 , y22235 , y22236 , y22237 , y22238 , y22239 , y22240 , y22241 , y22242 , y22243 , y22244 , y22245 , y22246 , y22247 , y22248 , y22249 , y22250 , y22251 , y22252 , y22253 , y22254 , y22255 , y22256 , y22257 , y22258 , y22259 , y22260 , y22261 , y22262 , y22263 , y22264 , y22265 , y22266 , y22267 , y22268 , y22269 , y22270 , y22271 , y22272 , y22273 , y22274 , y22275 , y22276 , y22277 , y22278 , y22279 , y22280 , y22281 , y22282 , y22283 , y22284 , y22285 , y22286 , y22287 , y22288 , y22289 , y22290 , y22291 , y22292 , y22293 , y22294 , y22295 , y22296 , y22297 , y22298 , y22299 , y22300 , y22301 , y22302 , y22303 , y22304 , y22305 , y22306 , y22307 , y22308 , y22309 , y22310 , y22311 , y22312 , y22313 , y22314 , y22315 , y22316 , y22317 , y22318 , y22319 , y22320 , y22321 , y22322 , y22323 , y22324 , y22325 , y22326 , y22327 , y22328 , y22329 , y22330 , y22331 , y22332 , y22333 , y22334 , y22335 , y22336 , y22337 , y22338 , y22339 , y22340 , y22341 , y22342 , y22343 , y22344 , y22345 , y22346 , y22347 , y22348 , y22349 , y22350 , y22351 , y22352 , y22353 , y22354 , y22355 , y22356 , y22357 , y22358 , y22359 , y22360 , y22361 , y22362 , y22363 , y22364 , y22365 , y22366 , y22367 , y22368 , y22369 , y22370 , y22371 , y22372 , y22373 , y22374 , y22375 , y22376 , y22377 , y22378 , y22379 , y22380 , y22381 , y22382 , y22383 , y22384 , y22385 , y22386 , y22387 , y22388 , y22389 , y22390 , y22391 , y22392 , y22393 , y22394 , y22395 , y22396 , y22397 , y22398 , y22399 , y22400 , y22401 , y22402 , y22403 , y22404 , y22405 , y22406 , y22407 , y22408 , y22409 , y22410 , y22411 , y22412 , y22413 , y22414 , y22415 , y22416 , y22417 , y22418 , y22419 , y22420 , y22421 , y22422 , y22423 , y22424 , y22425 , y22426 , y22427 , y22428 , y22429 , y22430 , y22431 , y22432 , y22433 , y22434 , y22435 , y22436 , y22437 , y22438 , y22439 , y22440 , y22441 , y22442 , y22443 , y22444 , y22445 , y22446 , y22447 , y22448 , y22449 , y22450 , y22451 , y22452 , y22453 , y22454 , y22455 , y22456 , y22457 , y22458 , y22459 , y22460 , y22461 , y22462 , y22463 , y22464 , y22465 , y22466 , y22467 , y22468 , y22469 , y22470 , y22471 , y22472 , y22473 , y22474 , y22475 , y22476 , y22477 , y22478 , y22479 , y22480 , y22481 , y22482 , y22483 , y22484 , y22485 , y22486 , y22487 , y22488 , y22489 , y22490 , y22491 , y22492 , y22493 , y22494 , y22495 , y22496 , y22497 , y22498 , y22499 , y22500 , y22501 , y22502 , y22503 , y22504 , y22505 , y22506 , y22507 , y22508 , y22509 , y22510 , y22511 , y22512 , y22513 , y22514 , y22515 , y22516 , y22517 , y22518 , y22519 , y22520 , y22521 , y22522 , y22523 , y22524 , y22525 , y22526 , y22527 , y22528 , y22529 , y22530 , y22531 , y22532 , y22533 , y22534 , y22535 , y22536 , y22537 , y22538 , y22539 , y22540 , y22541 , y22542 , y22543 , y22544 , y22545 , y22546 , y22547 , y22548 , y22549 , y22550 , y22551 , y22552 , y22553 , y22554 , y22555 , y22556 , y22557 , y22558 , y22559 , y22560 , y22561 , y22562 , y22563 , y22564 , y22565 , y22566 , y22567 , y22568 , y22569 , y22570 , y22571 , y22572 , y22573 , y22574 , y22575 , y22576 , y22577 , y22578 , y22579 , y22580 , y22581 , y22582 , y22583 , y22584 , y22585 , y22586 , y22587 , y22588 , y22589 , y22590 , y22591 , y22592 , y22593 , y22594 , y22595 , y22596 , y22597 , y22598 , y22599 , y22600 , y22601 , y22602 , y22603 , y22604 , y22605 , y22606 , y22607 , y22608 , y22609 , y22610 , y22611 , y22612 , y22613 , y22614 , y22615 , y22616 , y22617 , y22618 , y22619 , y22620 , y22621 , y22622 , y22623 , y22624 , y22625 , y22626 , y22627 , y22628 , y22629 , y22630 , y22631 , y22632 , y22633 , y22634 , y22635 , y22636 , y22637 , y22638 , y22639 , y22640 , y22641 , y22642 , y22643 , y22644 , y22645 , y22646 , y22647 , y22648 , y22649 , y22650 , y22651 , y22652 , y22653 , y22654 , y22655 , y22656 , y22657 , y22658 , y22659 , y22660 , y22661 , y22662 , y22663 , y22664 , y22665 , y22666 , y22667 , y22668 , y22669 , y22670 , y22671 , y22672 , y22673 , y22674 , y22675 , y22676 , y22677 , y22678 , y22679 , y22680 , y22681 , y22682 , y22683 , y22684 , y22685 , y22686 , y22687 , y22688 , y22689 , y22690 , y22691 , y22692 , y22693 , y22694 , y22695 , y22696 , y22697 , y22698 , y22699 , y22700 , y22701 , y22702 , y22703 , y22704 , y22705 , y22706 , y22707 , y22708 , y22709 , y22710 , y22711 , y22712 , y22713 , y22714 , y22715 , y22716 , y22717 , y22718 , y22719 , y22720 , y22721 , y22722 , y22723 , y22724 , y22725 , y22726 , y22727 , y22728 , y22729 , y22730 , y22731 , y22732 , y22733 , y22734 , y22735 , y22736 , y22737 , y22738 , y22739 , y22740 , y22741 , y22742 , y22743 , y22744 , y22745 , y22746 , y22747 , y22748 , y22749 , y22750 , y22751 , y22752 , y22753 , y22754 , y22755 , y22756 , y22757 , y22758 , y22759 , y22760 , y22761 , y22762 , y22763 , y22764 , y22765 , y22766 , y22767 , y22768 , y22769 , y22770 , y22771 , y22772 , y22773 , y22774 , y22775 , y22776 , y22777 , y22778 , y22779 , y22780 , y22781 , y22782 , y22783 , y22784 , y22785 , y22786 , y22787 , y22788 , y22789 , y22790 , y22791 , y22792 , y22793 , y22794 , y22795 , y22796 , y22797 , y22798 , y22799 , y22800 , y22801 , y22802 , y22803 , y22804 , y22805 , y22806 , y22807 , y22808 , y22809 , y22810 , y22811 , y22812 , y22813 , y22814 , y22815 , y22816 , y22817 , y22818 , y22819 , y22820 , y22821 , y22822 , y22823 , y22824 , y22825 , y22826 , y22827 , y22828 , y22829 , y22830 , y22831 , y22832 , y22833 , y22834 , y22835 , y22836 , y22837 , y22838 , y22839 , y22840 , y22841 , y22842 , y22843 , y22844 , y22845 , y22846 , y22847 , y22848 , y22849 , y22850 , y22851 , y22852 , y22853 , y22854 , y22855 , y22856 , y22857 , y22858 , y22859 , y22860 , y22861 , y22862 , y22863 , y22864 , y22865 , y22866 , y22867 , y22868 , y22869 , y22870 , y22871 , y22872 , y22873 , y22874 , y22875 , y22876 , y22877 , y22878 , y22879 , y22880 , y22881 , y22882 , y22883 , y22884 , y22885 , y22886 , y22887 , y22888 , y22889 , y22890 , y22891 , y22892 , y22893 , y22894 , y22895 , y22896 , y22897 , y22898 , y22899 , y22900 , y22901 , y22902 , y22903 , y22904 , y22905 , y22906 , y22907 , y22908 , y22909 , y22910 , y22911 , y22912 , y22913 , y22914 , y22915 , y22916 , y22917 , y22918 , y22919 , y22920 , y22921 , y22922 , y22923 , y22924 , y22925 , y22926 , y22927 , y22928 , y22929 , y22930 , y22931 , y22932 , y22933 , y22934 , y22935 , y22936 , y22937 , y22938 , y22939 , y22940 , y22941 , y22942 , y22943 , y22944 , y22945 , y22946 , y22947 , y22948 , y22949 , y22950 , y22951 , y22952 , y22953 , y22954 , y22955 , y22956 , y22957 , y22958 , y22959 , y22960 , y22961 , y22962 , y22963 , y22964 , y22965 , y22966 , y22967 , y22968 , y22969 , y22970 , y22971 , y22972 , y22973 , y22974 , y22975 , y22976 , y22977 , y22978 , y22979 , y22980 , y22981 , y22982 , y22983 , y22984 , y22985 , y22986 , y22987 , y22988 , y22989 , y22990 , y22991 , y22992 , y22993 , y22994 , y22995 , y22996 , y22997 , y22998 , y22999 , y23000 , y23001 , y23002 , y23003 , y23004 , y23005 , y23006 , y23007 , y23008 , y23009 , y23010 , y23011 , y23012 , y23013 , y23014 , y23015 , y23016 , y23017 , y23018 , y23019 , y23020 , y23021 , y23022 , y23023 , y23024 , y23025 , y23026 , y23027 , y23028 , y23029 , y23030 , y23031 , y23032 , y23033 , y23034 , y23035 , y23036 , y23037 , y23038 , y23039 , y23040 , y23041 , y23042 , y23043 , y23044 , y23045 , y23046 , y23047 , y23048 , y23049 , y23050 , y23051 , y23052 , y23053 , y23054 , y23055 , y23056 , y23057 , y23058 , y23059 , y23060 , y23061 , y23062 , y23063 , y23064 , y23065 , y23066 , y23067 , y23068 , y23069 , y23070 , y23071 , y23072 , y23073 , y23074 , y23075 , y23076 , y23077 , y23078 , y23079 , y23080 , y23081 , y23082 , y23083 , y23084 , y23085 , y23086 , y23087 , y23088 , y23089 , y23090 , y23091 , y23092 , y23093 , y23094 , y23095 , y23096 , y23097 , y23098 , y23099 , y23100 , y23101 , y23102 , y23103 , y23104 , y23105 , y23106 , y23107 , y23108 , y23109 , y23110 , y23111 , y23112 , y23113 , y23114 , y23115 , y23116 , y23117 , y23118 , y23119 , y23120 , y23121 , y23122 , y23123 , y23124 , y23125 , y23126 , y23127 , y23128 , y23129 , y23130 , y23131 , y23132 , y23133 , y23134 , y23135 , y23136 , y23137 , y23138 , y23139 , y23140 , y23141 , y23142 , y23143 , y23144 , y23145 , y23146 , y23147 , y23148 , y23149 , y23150 , y23151 , y23152 , y23153 , y23154 , y23155 , y23156 , y23157 , y23158 , y23159 , y23160 , y23161 , y23162 , y23163 , y23164 , y23165 , y23166 , y23167 , y23168 , y23169 , y23170 , y23171 , y23172 , y23173 , y23174 , y23175 , y23176 , y23177 , y23178 , y23179 , y23180 , y23181 , y23182 , y23183 , y23184 , y23185 , y23186 , y23187 , y23188 , y23189 , y23190 , y23191 , y23192 , y23193 , y23194 , y23195 , y23196 , y23197 , y23198 , y23199 , y23200 , y23201 , y23202 , y23203 , y23204 , y23205 , y23206 , y23207 , y23208 , y23209 , y23210 , y23211 , y23212 , y23213 , y23214 , y23215 , y23216 , y23217 , y23218 , y23219 , y23220 , y23221 , y23222 , y23223 , y23224 , y23225 , y23226 , y23227 , y23228 , y23229 , y23230 , y23231 , y23232 , y23233 , y23234 , y23235 , y23236 , y23237 , y23238 , y23239 , y23240 , y23241 , y23242 , y23243 , y23244 , y23245 , y23246 , y23247 , y23248 , y23249 , y23250 , y23251 , y23252 , y23253 , y23254 , y23255 , y23256 , y23257 , y23258 , y23259 , y23260 , y23261 , y23262 , y23263 , y23264 , y23265 , y23266 , y23267 , y23268 , y23269 , y23270 , y23271 , y23272 , y23273 , y23274 , y23275 , y23276 , y23277 , y23278 , y23279 , y23280 , y23281 , y23282 , y23283 , y23284 , y23285 , y23286 , y23287 , y23288 , y23289 , y23290 , y23291 , y23292 , y23293 , y23294 , y23295 , y23296 , y23297 , y23298 , y23299 , y23300 , y23301 , y23302 , y23303 , y23304 , y23305 , y23306 , y23307 , y23308 , y23309 , y23310 , y23311 , y23312 , y23313 , y23314 , y23315 , y23316 , y23317 , y23318 , y23319 , y23320 , y23321 , y23322 , y23323 , y23324 , y23325 , y23326 , y23327 , y23328 , y23329 , y23330 , y23331 , y23332 , y23333 , y23334 , y23335 , y23336 , y23337 , y23338 , y23339 , y23340 , y23341 , y23342 , y23343 , y23344 , y23345 , y23346 , y23347 , y23348 , y23349 , y23350 , y23351 , y23352 , y23353 , y23354 , y23355 , y23356 , y23357 , y23358 , y23359 , y23360 , y23361 , y23362 , y23363 , y23364 , y23365 , y23366 , y23367 , y23368 , y23369 , y23370 , y23371 , y23372 , y23373 , y23374 , y23375 , y23376 , y23377 , y23378 , y23379 , y23380 , y23381 , y23382 , y23383 , y23384 , y23385 , y23386 , y23387 , y23388 , y23389 , y23390 , y23391 , y23392 , y23393 , y23394 , y23395 , y23396 , y23397 , y23398 , y23399 , y23400 , y23401 , y23402 , y23403 , y23404 , y23405 , y23406 , y23407 , y23408 , y23409 , y23410 , y23411 , y23412 , y23413 , y23414 , y23415 , y23416 , y23417 , y23418 , y23419 , y23420 , y23421 , y23422 , y23423 , y23424 , y23425 , y23426 , y23427 , y23428 , y23429 , y23430 , y23431 , y23432 , y23433 , y23434 , y23435 , y23436 , y23437 , y23438 , y23439 , y23440 , y23441 , y23442 , y23443 , y23444 , y23445 , y23446 , y23447 , y23448 , y23449 , y23450 , y23451 , y23452 , y23453 , y23454 , y23455 , y23456 , y23457 , y23458 , y23459 , y23460 , y23461 , y23462 , y23463 , y23464 , y23465 , y23466 , y23467 , y23468 , y23469 , y23470 , y23471 , y23472 , y23473 , y23474 , y23475 , y23476 , y23477 , y23478 , y23479 , y23480 , y23481 , y23482 , y23483 , y23484 , y23485 , y23486 , y23487 , y23488 , y23489 , y23490 , y23491 , y23492 , y23493 , y23494 , y23495 , y23496 , y23497 , y23498 , y23499 , y23500 , y23501 , y23502 , y23503 , y23504 , y23505 , y23506 , y23507 , y23508 , y23509 , y23510 , y23511 , y23512 , y23513 , y23514 , y23515 , y23516 , y23517 , y23518 , y23519 , y23520 , y23521 , y23522 , y23523 , y23524 , y23525 , y23526 , y23527 , y23528 , y23529 , y23530 , y23531 , y23532 , y23533 , y23534 , y23535 , y23536 , y23537 , y23538 , y23539 , y23540 , y23541 , y23542 , y23543 , y23544 , y23545 , y23546 , y23547 , y23548 , y23549 , y23550 , y23551 , y23552 , y23553 , y23554 , y23555 , y23556 , y23557 , y23558 , y23559 , y23560 , y23561 , y23562 , y23563 , y23564 , y23565 , y23566 , y23567 , y23568 , y23569 , y23570 , y23571 , y23572 , y23573 , y23574 , y23575 , y23576 , y23577 , y23578 , y23579 , y23580 , y23581 , y23582 , y23583 , y23584 , y23585 , y23586 , y23587 , y23588 , y23589 , y23590 , y23591 , y23592 , y23593 , y23594 , y23595 , y23596 , y23597 , y23598 , y23599 , y23600 , y23601 , y23602 , y23603 , y23604 , y23605 , y23606 , y23607 , y23608 , y23609 , y23610 , y23611 , y23612 , y23613 , y23614 , y23615 , y23616 , y23617 , y23618 , y23619 , y23620 , y23621 , y23622 , y23623 , y23624 , y23625 , y23626 , y23627 , y23628 , y23629 , y23630 , y23631 , y23632 , y23633 , y23634 , y23635 , y23636 , y23637 , y23638 , y23639 , y23640 , y23641 , y23642 , y23643 , y23644 , y23645 , y23646 , y23647 , y23648 , y23649 , y23650 , y23651 , y23652 , y23653 , y23654 , y23655 , y23656 , y23657 , y23658 , y23659 , y23660 , y23661 , y23662 , y23663 , y23664 , y23665 , y23666 , y23667 , y23668 , y23669 , y23670 , y23671 , y23672 , y23673 , y23674 , y23675 , y23676 , y23677 , y23678 , y23679 , y23680 , y23681 , y23682 , y23683 , y23684 , y23685 , y23686 , y23687 , y23688 , y23689 , y23690 , y23691 , y23692 , y23693 , y23694 , y23695 , y23696 , y23697 , y23698 , y23699 , y23700 , y23701 , y23702 , y23703 , y23704 , y23705 , y23706 , y23707 , y23708 , y23709 , y23710 , y23711 , y23712 , y23713 , y23714 , y23715 , y23716 , y23717 , y23718 , y23719 , y23720 , y23721 , y23722 , y23723 , y23724 , y23725 , y23726 , y23727 , y23728 , y23729 , y23730 , y23731 , y23732 , y23733 , y23734 , y23735 , y23736 , y23737 , y23738 , y23739 , y23740 , y23741 , y23742 , y23743 , y23744 , y23745 , y23746 , y23747 , y23748 , y23749 , y23750 , y23751 , y23752 , y23753 , y23754 , y23755 , y23756 , y23757 , y23758 , y23759 , y23760 , y23761 , y23762 , y23763 , y23764 , y23765 , y23766 , y23767 , y23768 , y23769 , y23770 , y23771 , y23772 , y23773 , y23774 , y23775 , y23776 , y23777 , y23778 , y23779 , y23780 , y23781 , y23782 , y23783 , y23784 , y23785 , y23786 , y23787 , y23788 , y23789 , y23790 , y23791 , y23792 , y23793 , y23794 , y23795 , y23796 , y23797 , y23798 , y23799 , y23800 , y23801 , y23802 , y23803 , y23804 , y23805 , y23806 , y23807 , y23808 , y23809 , y23810 , y23811 , y23812 , y23813 , y23814 , y23815 , y23816 , y23817 , y23818 , y23819 , y23820 , y23821 , y23822 , y23823 , y23824 , y23825 , y23826 , y23827 , y23828 , y23829 , y23830 , y23831 , y23832 , y23833 , y23834 , y23835 , y23836 , y23837 , y23838 , y23839 , y23840 , y23841 , y23842 , y23843 , y23844 , y23845 , y23846 , y23847 , y23848 , y23849 , y23850 , y23851 , y23852 , y23853 , y23854 , y23855 , y23856 , y23857 , y23858 , y23859 , y23860 , y23861 , y23862 , y23863 , y23864 , y23865 , y23866 , y23867 , y23868 , y23869 , y23870 , y23871 , y23872 , y23873 , y23874 , y23875 , y23876 , y23877 , y23878 , y23879 , y23880 , y23881 , y23882 , y23883 , y23884 , y23885 , y23886 , y23887 , y23888 , y23889 , y23890 , y23891 , y23892 , y23893 , y23894 , y23895 , y23896 , y23897 , y23898 , y23899 , y23900 , y23901 , y23902 , y23903 , y23904 , y23905 , y23906 , y23907 , y23908 , y23909 , y23910 , y23911 , y23912 , y23913 , y23914 , y23915 , y23916 , y23917 , y23918 , y23919 , y23920 , y23921 , y23922 , y23923 , y23924 , y23925 , y23926 , y23927 , y23928 , y23929 , y23930 , y23931 , y23932 , y23933 , y23934 , y23935 , y23936 , y23937 , y23938 , y23939 , y23940 , y23941 , y23942 , y23943 , y23944 , y23945 , y23946 , y23947 , y23948 , y23949 , y23950 , y23951 , y23952 , y23953 , y23954 , y23955 , y23956 , y23957 , y23958 , y23959 , y23960 , y23961 , y23962 , y23963 , y23964 , y23965 , y23966 , y23967 , y23968 , y23969 , y23970 , y23971 , y23972 , y23973 , y23974 , y23975 , y23976 , y23977 , y23978 , y23979 , y23980 , y23981 , y23982 , y23983 , y23984 , y23985 , y23986 , y23987 , y23988 , y23989 , y23990 , y23991 , y23992 , y23993 , y23994 , y23995 , y23996 , y23997 , y23998 , y23999 , y24000 , y24001 , y24002 , y24003 , y24004 , y24005 , y24006 , y24007 , y24008 , y24009 , y24010 , y24011 , y24012 , y24013 , y24014 , y24015 , y24016 , y24017 , y24018 , y24019 , y24020 , y24021 , y24022 , y24023 , y24024 , y24025 , y24026 , y24027 , y24028 , y24029 , y24030 , y24031 , y24032 , y24033 , y24034 , y24035 , y24036 , y24037 , y24038 , y24039 , y24040 , y24041 , y24042 , y24043 , y24044 , y24045 , y24046 , y24047 , y24048 , y24049 , y24050 , y24051 , y24052 , y24053 , y24054 , y24055 , y24056 , y24057 , y24058 , y24059 , y24060 , y24061 , y24062 , y24063 , y24064 , y24065 , y24066 , y24067 , y24068 , y24069 , y24070 , y24071 , y24072 , y24073 , y24074 , y24075 , y24076 , y24077 , y24078 , y24079 , y24080 , y24081 , y24082 , y24083 , y24084 , y24085 , y24086 , y24087 , y24088 , y24089 , y24090 , y24091 , y24092 , y24093 , y24094 , y24095 , y24096 , y24097 , y24098 , y24099 , y24100 , y24101 , y24102 , y24103 , y24104 , y24105 , y24106 , y24107 , y24108 , y24109 , y24110 , y24111 , y24112 , y24113 , y24114 , y24115 , y24116 , y24117 , y24118 , y24119 , y24120 , y24121 , y24122 , y24123 , y24124 , y24125 , y24126 , y24127 , y24128 , y24129 , y24130 , y24131 , y24132 , y24133 , y24134 , y24135 , y24136 , y24137 , y24138 , y24139 , y24140 , y24141 , y24142 , y24143 , y24144 , y24145 , y24146 , y24147 , y24148 , y24149 , y24150 , y24151 , y24152 , y24153 , y24154 , y24155 , y24156 , y24157 , y24158 , y24159 , y24160 , y24161 , y24162 , y24163 , y24164 , y24165 , y24166 , y24167 , y24168 , y24169 , y24170 , y24171 , y24172 , y24173 , y24174 , y24175 , y24176 , y24177 , y24178 , y24179 , y24180 , y24181 , y24182 , y24183 , y24184 , y24185 , y24186 , y24187 , y24188 , y24189 , y24190 , y24191 , y24192 , y24193 , y24194 , y24195 , y24196 , y24197 , y24198 , y24199 , y24200 , y24201 , y24202 , y24203 , y24204 , y24205 , y24206 , y24207 , y24208 , y24209 , y24210 , y24211 , y24212 , y24213 , y24214 , y24215 , y24216 , y24217 , y24218 , y24219 , y24220 , y24221 , y24222 , y24223 , y24224 , y24225 , y24226 , y24227 , y24228 , y24229 , y24230 , y24231 , y24232 , y24233 , y24234 , y24235 , y24236 , y24237 , y24238 , y24239 , y24240 , y24241 , y24242 , y24243 , y24244 , y24245 , y24246 , y24247 , y24248 , y24249 , y24250 , y24251 , y24252 , y24253 , y24254 , y24255 , y24256 , y24257 , y24258 , y24259 , y24260 , y24261 , y24262 , y24263 , y24264 , y24265 , y24266 , y24267 , y24268 , y24269 , y24270 , y24271 , y24272 , y24273 , y24274 , y24275 , y24276 , y24277 , y24278 , y24279 , y24280 , y24281 , y24282 , y24283 , y24284 , y24285 , y24286 , y24287 , y24288 , y24289 , y24290 , y24291 , y24292 , y24293 , y24294 , y24295 , y24296 , y24297 , y24298 , y24299 , y24300 , y24301 , y24302 , y24303 , y24304 , y24305 , y24306 , y24307 , y24308 , y24309 , y24310 , y24311 , y24312 , y24313 , y24314 , y24315 , y24316 , y24317 , y24318 , y24319 , y24320 , y24321 , y24322 , y24323 , y24324 , y24325 , y24326 , y24327 , y24328 , y24329 , y24330 , y24331 , y24332 , y24333 , y24334 , y24335 , y24336 , y24337 , y24338 , y24339 , y24340 , y24341 , y24342 , y24343 , y24344 , y24345 , y24346 , y24347 , y24348 , y24349 , y24350 , y24351 , y24352 , y24353 , y24354 , y24355 , y24356 , y24357 , y24358 , y24359 , y24360 , y24361 , y24362 , y24363 , y24364 , y24365 , y24366 , y24367 , y24368 , y24369 , y24370 , y24371 , y24372 , y24373 , y24374 , y24375 , y24376 , y24377 , y24378 , y24379 , y24380 , y24381 , y24382 , y24383 , y24384 , y24385 , y24386 , y24387 , y24388 , y24389 , y24390 , y24391 , y24392 , y24393 , y24394 , y24395 , y24396 , y24397 , y24398 , y24399 , y24400 , y24401 , y24402 , y24403 , y24404 , y24405 , y24406 , y24407 , y24408 , y24409 , y24410 , y24411 , y24412 , y24413 , y24414 , y24415 , y24416 , y24417 , y24418 , y24419 , y24420 , y24421 , y24422 , y24423 , y24424 , y24425 , y24426 , y24427 , y24428 , y24429 , y24430 , y24431 , y24432 , y24433 , y24434 , y24435 , y24436 , y24437 , y24438 , y24439 , y24440 , y24441 , y24442 , y24443 , y24444 , y24445 , y24446 , y24447 , y24448 , y24449 , y24450 , y24451 , y24452 , y24453 , y24454 , y24455 , y24456 , y24457 , y24458 , y24459 , y24460 , y24461 , y24462 , y24463 , y24464 , y24465 , y24466 , y24467 , y24468 , y24469 , y24470 , y24471 , y24472 , y24473 , y24474 , y24475 , y24476 , y24477 , y24478 , y24479 , y24480 , y24481 , y24482 , y24483 , y24484 , y24485 , y24486 , y24487 , y24488 , y24489 , y24490 , y24491 , y24492 , y24493 , y24494 , y24495 , y24496 , y24497 , y24498 , y24499 , y24500 , y24501 , y24502 , y24503 , y24504 , y24505 , y24506 , y24507 , y24508 , y24509 , y24510 , y24511 , y24512 , y24513 , y24514 , y24515 , y24516 , y24517 , y24518 , y24519 , y24520 , y24521 , y24522 , y24523 , y24524 , y24525 , y24526 , y24527 , y24528 , y24529 , y24530 , y24531 , y24532 , y24533 , y24534 , y24535 , y24536 , y24537 , y24538 , y24539 , y24540 , y24541 , y24542 , y24543 , y24544 , y24545 , y24546 , y24547 , y24548 , y24549 , y24550 , y24551 , y24552 , y24553 , y24554 , y24555 , y24556 , y24557 , y24558 , y24559 , y24560 , y24561 , y24562 , y24563 , y24564 , y24565 , y24566 , y24567 , y24568 , y24569 , y24570 , y24571 , y24572 , y24573 , y24574 , y24575 , y24576 , y24577 , y24578 , y24579 , y24580 , y24581 , y24582 , y24583 , y24584 , y24585 , y24586 , y24587 , y24588 , y24589 , y24590 , y24591 , y24592 , y24593 , y24594 , y24595 , y24596 , y24597 , y24598 , y24599 , y24600 , y24601 , y24602 , y24603 , y24604 , y24605 , y24606 , y24607 , y24608 , y24609 , y24610 , y24611 , y24612 , y24613 , y24614 , y24615 , y24616 , y24617 , y24618 , y24619 , y24620 , y24621 , y24622 , y24623 , y24624 , y24625 , y24626 , y24627 , y24628 , y24629 , y24630 , y24631 , y24632 , y24633 , y24634 , y24635 , y24636 , y24637 , y24638 , y24639 , y24640 , y24641 , y24642 , y24643 , y24644 , y24645 , y24646 , y24647 , y24648 , y24649 , y24650 , y24651 , y24652 , y24653 , y24654 , y24655 , y24656 , y24657 , y24658 , y24659 , y24660 , y24661 , y24662 , y24663 , y24664 , y24665 , y24666 , y24667 , y24668 , y24669 , y24670 , y24671 , y24672 , y24673 , y24674 , y24675 , y24676 , y24677 , y24678 , y24679 , y24680 , y24681 , y24682 , y24683 , y24684 , y24685 , y24686 , y24687 , y24688 , y24689 , y24690 , y24691 , y24692 , y24693 , y24694 , y24695 , y24696 , y24697 , y24698 , y24699 , y24700 , y24701 , y24702 , y24703 , y24704 , y24705 , y24706 , y24707 , y24708 , y24709 , y24710 , y24711 , y24712 , y24713 , y24714 , y24715 , y24716 , y24717 , y24718 , y24719 , y24720 , y24721 , y24722 , y24723 , y24724 , y24725 , y24726 , y24727 , y24728 , y24729 , y24730 , y24731 , y24732 , y24733 , y24734 , y24735 , y24736 , y24737 , y24738 , y24739 , y24740 , y24741 , y24742 , y24743 , y24744 , y24745 , y24746 , y24747 , y24748 , y24749 , y24750 , y24751 , y24752 , y24753 , y24754 , y24755 , y24756 , y24757 , y24758 , y24759 , y24760 , y24761 , y24762 , y24763 , y24764 , y24765 , y24766 , y24767 , y24768 , y24769 , y24770 , y24771 , y24772 , y24773 , y24774 , y24775 , y24776 , y24777 , y24778 , y24779 , y24780 , y24781 , y24782 , y24783 , y24784 , y24785 , y24786 , y24787 , y24788 , y24789 , y24790 , y24791 , y24792 , y24793 , y24794 , y24795 , y24796 , y24797 , y24798 , y24799 , y24800 , y24801 , y24802 , y24803 , y24804 , y24805 , y24806 , y24807 , y24808 , y24809 , y24810 , y24811 , y24812 , y24813 , y24814 , y24815 , y24816 , y24817 , y24818 , y24819 , y24820 , y24821 , y24822 , y24823 , y24824 , y24825 , y24826 , y24827 , y24828 , y24829 , y24830 , y24831 , y24832 , y24833 , y24834 , y24835 , y24836 , y24837 , y24838 , y24839 , y24840 , y24841 , y24842 , y24843 , y24844 , y24845 , y24846 , y24847 , y24848 , y24849 , y24850 , y24851 , y24852 , y24853 , y24854 , y24855 , y24856 , y24857 , y24858 , y24859 , y24860 , y24861 , y24862 , y24863 , y24864 , y24865 , y24866 , y24867 , y24868 , y24869 , y24870 , y24871 , y24872 , y24873 , y24874 , y24875 , y24876 , y24877 , y24878 , y24879 , y24880 , y24881 , y24882 , y24883 , y24884 , y24885 , y24886 , y24887 , y24888 , y24889 , y24890 , y24891 , y24892 , y24893 , y24894 , y24895 , y24896 , y24897 , y24898 , y24899 , y24900 , y24901 , y24902 , y24903 , y24904 , y24905 , y24906 , y24907 , y24908 , y24909 , y24910 , y24911 , y24912 , y24913 , y24914 , y24915 , y24916 , y24917 , y24918 , y24919 , y24920 , y24921 , y24922 ;
  wire n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 ;
  assign n256 = x127 ^ x119 ^ 1'b0 ;
  assign n257 = x175 & n256 ;
  assign n258 = x74 & x199 ;
  assign n259 = n258 ^ x156 ^ 1'b0 ;
  assign n260 = x98 & x147 ;
  assign n261 = n260 ^ x146 ^ 1'b0 ;
  assign n262 = x23 ^ x3 ^ 1'b0 ;
  assign n263 = x75 & n262 ;
  assign n264 = x218 ^ x202 ^ 1'b0 ;
  assign n265 = x220 & n264 ;
  assign n266 = x224 ^ x81 ^ 1'b0 ;
  assign n267 = ~n259 & n266 ;
  assign n268 = x246 ^ x19 ^ 1'b0 ;
  assign n269 = x46 & n268 ;
  assign n270 = x246 & x254 ;
  assign n271 = n270 ^ x146 ^ 1'b0 ;
  assign n272 = x141 & ~n271 ;
  assign n273 = n272 ^ x238 ^ 1'b0 ;
  assign n274 = x32 & x33 ;
  assign n275 = ~x95 & n274 ;
  assign n276 = n261 ^ x203 ^ 1'b0 ;
  assign n277 = x8 & ~n276 ;
  assign n278 = n277 ^ x5 ^ 1'b0 ;
  assign n279 = x150 ^ x125 ^ x70 ;
  assign n280 = x231 ^ x125 ^ 1'b0 ;
  assign n281 = ~n279 & n280 ;
  assign n282 = x80 & x227 ;
  assign n283 = n282 ^ x193 ^ 1'b0 ;
  assign n284 = x0 & x223 ;
  assign n285 = ~x8 & n284 ;
  assign n286 = ~x25 & x144 ;
  assign n287 = x110 ^ x105 ^ 1'b0 ;
  assign n288 = x37 & n287 ;
  assign n289 = x155 & x254 ;
  assign n290 = ~n288 & n289 ;
  assign n291 = x175 ^ x157 ^ 1'b0 ;
  assign n292 = x48 & n291 ;
  assign n293 = x47 & x231 ;
  assign n294 = n293 ^ x102 ^ 1'b0 ;
  assign n295 = x36 ^ x0 ^ 1'b0 ;
  assign n296 = x226 & n295 ;
  assign n297 = x241 ^ x237 ^ 1'b0 ;
  assign n298 = x1 & n297 ;
  assign n299 = x58 & x163 ;
  assign n300 = n299 ^ x178 ^ 1'b0 ;
  assign n301 = n300 ^ x246 ^ 1'b0 ;
  assign n302 = n298 & ~n301 ;
  assign n303 = x231 ^ x127 ^ 1'b0 ;
  assign n304 = x154 & n303 ;
  assign n305 = ( x80 & x138 ) | ( x80 & ~n304 ) | ( x138 & ~n304 ) ;
  assign n306 = x191 ^ x34 ^ 1'b0 ;
  assign n307 = x77 & n306 ;
  assign n308 = x106 & x175 ;
  assign n309 = ~x191 & n308 ;
  assign n310 = x78 & x236 ;
  assign n311 = ~x199 & n310 ;
  assign n312 = x169 & ~n300 ;
  assign n313 = n312 ^ n257 ^ 1'b0 ;
  assign n314 = x238 & ~n259 ;
  assign n315 = n314 ^ x207 ^ 1'b0 ;
  assign n316 = x2 & x135 ;
  assign n317 = ~x186 & n316 ;
  assign n318 = n294 ^ n263 ^ x42 ;
  assign n319 = x93 & ~n275 ;
  assign n320 = n319 ^ x115 ^ 1'b0 ;
  assign n321 = x113 & x249 ;
  assign n322 = n321 ^ x15 ^ 1'b0 ;
  assign n323 = x243 ^ x190 ^ 1'b0 ;
  assign n324 = x78 & ~n300 ;
  assign n325 = n324 ^ x11 ^ 1'b0 ;
  assign n326 = x105 & x196 ;
  assign n327 = ~x165 & n326 ;
  assign n328 = x18 & x158 ;
  assign n329 = n328 ^ x15 ^ 1'b0 ;
  assign n330 = x132 & x177 ;
  assign n331 = ~x125 & n330 ;
  assign n332 = n290 ^ x219 ^ 1'b0 ;
  assign n333 = x14 & ~n332 ;
  assign n334 = x118 & x203 ;
  assign n335 = ~x164 & n334 ;
  assign n336 = x181 ^ x97 ^ 1'b0 ;
  assign n337 = ~n294 & n336 ;
  assign n338 = x75 & x212 ;
  assign n339 = ~x164 & n338 ;
  assign n340 = x3 & ~n339 ;
  assign n341 = ~n267 & n340 ;
  assign n342 = x150 ^ x125 ^ 1'b0 ;
  assign n343 = ~n341 & n342 ;
  assign n344 = x35 & ~n271 ;
  assign n345 = ~x73 & n344 ;
  assign n346 = x132 & x244 ;
  assign n347 = ~x16 & n346 ;
  assign n348 = x74 & x214 ;
  assign n349 = n348 ^ x194 ^ 1'b0 ;
  assign n350 = x234 & ~n349 ;
  assign n351 = n350 ^ x13 ^ 1'b0 ;
  assign n352 = x210 ^ x79 ^ x27 ;
  assign n353 = x73 ^ x61 ^ 1'b0 ;
  assign n354 = ~n352 & n353 ;
  assign n355 = x205 ^ x158 ^ 1'b0 ;
  assign n356 = x199 & ~n355 ;
  assign n357 = ~n354 & n356 ;
  assign n358 = x203 ^ x188 ^ x53 ;
  assign n359 = x71 & x157 ;
  assign n360 = ~x163 & n359 ;
  assign n361 = ( ~x48 & x108 ) | ( ~x48 & x240 ) | ( x108 & x240 ) ;
  assign n362 = x113 & x141 ;
  assign n363 = ~x50 & n362 ;
  assign n364 = n363 ^ x115 ^ 1'b0 ;
  assign n365 = x253 & ~n364 ;
  assign n366 = ( x132 & n361 ) | ( x132 & ~n365 ) | ( n361 & ~n365 ) ;
  assign n367 = ~n360 & n366 ;
  assign n368 = n367 ^ x22 ^ 1'b0 ;
  assign n369 = n259 | n290 ;
  assign n370 = x97 | n369 ;
  assign n371 = x250 ^ x28 ^ 1'b0 ;
  assign n372 = ~n335 & n371 ;
  assign n373 = ( ~x110 & x117 ) | ( ~x110 & n265 ) | ( x117 & n265 ) ;
  assign n374 = ~n275 & n327 ;
  assign n375 = x67 & x100 ;
  assign n376 = n375 ^ x43 ^ 1'b0 ;
  assign n377 = n341 ^ x198 ^ 1'b0 ;
  assign n378 = x161 & ~n377 ;
  assign n379 = x118 & ~n325 ;
  assign n380 = ~x184 & n379 ;
  assign n381 = ( x54 & ~x239 ) | ( x54 & n380 ) | ( ~x239 & n380 ) ;
  assign n383 = x60 & x76 ;
  assign n384 = ~x45 & n383 ;
  assign n382 = x29 & x115 ;
  assign n385 = n384 ^ n382 ^ 1'b0 ;
  assign n386 = n385 ^ x33 ^ 1'b0 ;
  assign n387 = x167 & n386 ;
  assign n388 = x155 ^ x153 ^ 1'b0 ;
  assign n389 = n283 ^ x180 ^ 1'b0 ;
  assign n390 = n311 | n389 ;
  assign n391 = n388 | n390 ;
  assign n392 = n391 ^ x161 ^ 1'b0 ;
  assign n394 = x139 & ~n354 ;
  assign n393 = x51 & x187 ;
  assign n395 = n394 ^ n393 ^ 1'b0 ;
  assign n396 = x99 & ~n395 ;
  assign n397 = n396 ^ x73 ^ 1'b0 ;
  assign n402 = n267 ^ x229 ^ 1'b0 ;
  assign n403 = x108 & n402 ;
  assign n404 = x127 & n403 ;
  assign n405 = ~n305 & n404 ;
  assign n398 = n370 ^ x178 ^ 1'b0 ;
  assign n399 = x29 & n398 ;
  assign n400 = x215 & n399 ;
  assign n401 = ~x180 & n400 ;
  assign n406 = n405 ^ n401 ^ 1'b0 ;
  assign n407 = x243 & n406 ;
  assign n408 = x48 ^ x44 ^ 1'b0 ;
  assign n409 = x195 & n408 ;
  assign n410 = x17 & x227 ;
  assign n411 = n410 ^ x153 ^ 1'b0 ;
  assign n412 = x58 ^ x0 ^ 1'b0 ;
  assign n413 = ~n411 & n412 ;
  assign n414 = ~n304 & n413 ;
  assign n415 = ( x177 & n411 ) | ( x177 & ~n414 ) | ( n411 & ~n414 ) ;
  assign n416 = x207 ^ x115 ^ 1'b0 ;
  assign n417 = x41 & n416 ;
  assign n418 = n417 ^ n288 ^ x194 ;
  assign n419 = n418 ^ x31 ^ 1'b0 ;
  assign n420 = n415 & ~n419 ;
  assign n421 = n420 ^ x27 ^ 1'b0 ;
  assign n422 = x139 ^ x123 ^ 1'b0 ;
  assign n423 = x164 & n422 ;
  assign n424 = x95 & n423 ;
  assign n425 = n424 ^ x26 ^ 1'b0 ;
  assign n426 = x164 | n425 ;
  assign n427 = x159 & n372 ;
  assign n428 = n427 ^ x145 ^ 1'b0 ;
  assign n429 = x148 & x197 ;
  assign n430 = n429 ^ x105 ^ 1'b0 ;
  assign n431 = x159 & ~n430 ;
  assign n432 = n431 ^ x250 ^ 1'b0 ;
  assign n433 = x3 & x195 ;
  assign n434 = ~x183 & n433 ;
  assign n435 = x160 & x173 ;
  assign n436 = ~x142 & n435 ;
  assign n437 = x3 & x132 ;
  assign n438 = n436 & n437 ;
  assign n439 = x245 & n265 ;
  assign n440 = ~x246 & n439 ;
  assign n441 = n440 ^ x88 ^ 1'b0 ;
  assign n442 = n438 | n441 ;
  assign n443 = n366 ^ n257 ^ 1'b0 ;
  assign n444 = x6 & n443 ;
  assign n445 = ( x190 & ~x205 ) | ( x190 & x233 ) | ( ~x205 & x233 ) ;
  assign n446 = ( x44 & n354 ) | ( x44 & ~n445 ) | ( n354 & ~n445 ) ;
  assign n447 = x13 & x176 ;
  assign n448 = n447 ^ x229 ^ 1'b0 ;
  assign n449 = x179 & x198 ;
  assign n450 = n449 ^ n335 ^ 1'b0 ;
  assign n451 = x67 ^ x21 ^ 1'b0 ;
  assign n452 = ~n279 & n451 ;
  assign n453 = n261 ^ x21 ^ 1'b0 ;
  assign n454 = n281 & ~n453 ;
  assign n455 = n452 & n454 ;
  assign n456 = ~n450 & n455 ;
  assign n457 = x29 ^ x2 ^ 1'b0 ;
  assign n458 = x130 & n457 ;
  assign n459 = n387 & n458 ;
  assign n460 = ~x192 & n459 ;
  assign n461 = n305 & n460 ;
  assign n462 = x198 ^ x47 ^ 1'b0 ;
  assign n463 = x95 & n462 ;
  assign n464 = n446 ^ x17 ^ 1'b0 ;
  assign n465 = n463 & n464 ;
  assign n466 = x145 & ~n273 ;
  assign n467 = n466 ^ n349 ^ 1'b0 ;
  assign n468 = x110 ^ x44 ^ 1'b0 ;
  assign n469 = x37 & x153 ;
  assign n470 = ~n302 & n469 ;
  assign n471 = x195 & ~n470 ;
  assign n472 = ~x129 & n471 ;
  assign n473 = x78 & x122 ;
  assign n474 = ~n257 & n473 ;
  assign n475 = x30 & ~n474 ;
  assign n476 = n275 & n475 ;
  assign n477 = x44 & x185 ;
  assign n478 = n311 & n477 ;
  assign n479 = x203 & ~n368 ;
  assign n480 = n479 ^ n454 ^ 1'b0 ;
  assign n481 = x162 & ~n480 ;
  assign n482 = x245 | n478 ;
  assign n484 = x238 ^ x32 ^ 1'b0 ;
  assign n485 = x243 & n484 ;
  assign n483 = x6 & x237 ;
  assign n486 = n485 ^ n483 ^ 1'b0 ;
  assign n487 = x247 & ~n486 ;
  assign n488 = n487 ^ x174 ^ 1'b0 ;
  assign n489 = n298 ^ x96 ^ 1'b0 ;
  assign n490 = n385 & n489 ;
  assign n491 = n414 ^ x221 ^ 1'b0 ;
  assign n492 = n490 & ~n491 ;
  assign n493 = ( ~x119 & n488 ) | ( ~x119 & n492 ) | ( n488 & n492 ) ;
  assign n494 = n320 | n341 ;
  assign n495 = n494 ^ x157 ^ 1'b0 ;
  assign n496 = x246 & n288 ;
  assign n497 = n496 ^ x141 ^ 1'b0 ;
  assign n498 = x235 ^ x87 ^ 1'b0 ;
  assign n499 = x111 ^ x38 ^ 1'b0 ;
  assign n500 = ~n414 & n499 ;
  assign n501 = n500 ^ n480 ^ 1'b0 ;
  assign n502 = x225 & ~n501 ;
  assign n503 = n351 & n502 ;
  assign n504 = x195 & ~x197 ;
  assign n505 = n436 ^ n385 ^ n360 ;
  assign n507 = x138 ^ x101 ^ 1'b0 ;
  assign n508 = x70 & n507 ;
  assign n509 = ( x180 & ~x216 ) | ( x180 & n508 ) | ( ~x216 & n508 ) ;
  assign n510 = ( x89 & ~x197 ) | ( x89 & n509 ) | ( ~x197 & n509 ) ;
  assign n511 = x215 ^ x197 ^ 1'b0 ;
  assign n512 = n510 & n511 ;
  assign n513 = x180 & x210 ;
  assign n514 = ~x240 & n513 ;
  assign n515 = x79 & ~n514 ;
  assign n516 = ~x70 & n515 ;
  assign n517 = n265 & ~n516 ;
  assign n518 = ~n512 & n517 ;
  assign n506 = x36 & x251 ;
  assign n519 = n518 ^ n506 ^ 1'b0 ;
  assign n520 = x122 & x171 ;
  assign n521 = n520 ^ x45 ^ 1'b0 ;
  assign n522 = n519 | n521 ;
  assign n523 = x254 ^ x127 ^ 1'b0 ;
  assign n524 = x109 & n523 ;
  assign n525 = n378 & ~n505 ;
  assign n526 = ~n524 & n525 ;
  assign n527 = x179 & ~n259 ;
  assign n528 = n354 | n436 ;
  assign n529 = x21 & ~x98 ;
  assign n531 = x212 ^ x74 ^ 1'b0 ;
  assign n532 = ~n436 & n531 ;
  assign n530 = n307 & ~n516 ;
  assign n533 = n532 ^ n530 ^ 1'b0 ;
  assign n534 = x76 ^ x0 ^ 1'b0 ;
  assign n535 = n392 ^ n296 ^ x21 ;
  assign n536 = n535 ^ x206 ^ 1'b0 ;
  assign n537 = x38 & x78 ;
  assign n538 = n537 ^ x76 ^ 1'b0 ;
  assign n539 = ( ~x67 & n292 ) | ( ~x67 & n358 ) | ( n292 & n358 ) ;
  assign n540 = n423 & ~n486 ;
  assign n541 = n540 ^ x221 ^ 1'b0 ;
  assign n542 = ~n434 & n541 ;
  assign n543 = n257 ^ x219 ^ 1'b0 ;
  assign n544 = x11 & ~n543 ;
  assign n545 = n544 ^ x16 ^ 1'b0 ;
  assign n546 = n542 & n545 ;
  assign n547 = x58 & ~n309 ;
  assign n548 = ~x2 & n547 ;
  assign n549 = x157 & n548 ;
  assign n550 = x7 & ~x210 ;
  assign n551 = n456 & n550 ;
  assign n552 = n551 ^ x176 ^ 1'b0 ;
  assign n555 = x54 & ~n436 ;
  assign n556 = ~x0 & n555 ;
  assign n554 = x234 & n482 ;
  assign n557 = n556 ^ n554 ^ 1'b0 ;
  assign n553 = x118 & ~x242 ;
  assign n558 = n557 ^ n553 ^ 1'b0 ;
  assign n559 = x106 & ~n558 ;
  assign n560 = n341 ^ x89 ^ 1'b0 ;
  assign n561 = x74 & ~n560 ;
  assign n562 = n309 | n561 ;
  assign n563 = n458 ^ n425 ^ 1'b0 ;
  assign n564 = x12 & ~n563 ;
  assign n565 = n564 ^ n327 ^ 1'b0 ;
  assign n566 = x241 & ~n565 ;
  assign n567 = n566 ^ x108 ^ 1'b0 ;
  assign n568 = ~n329 & n567 ;
  assign n569 = n568 ^ x80 ^ 1'b0 ;
  assign n570 = n378 & n569 ;
  assign n571 = n390 & n433 ;
  assign n572 = x25 & x229 ;
  assign n573 = ~n463 & n572 ;
  assign n574 = x73 & ~x157 ;
  assign n575 = ~n573 & n574 ;
  assign n576 = x197 & ~n574 ;
  assign n577 = n576 ^ n510 ^ 1'b0 ;
  assign n578 = n577 ^ x194 ^ 1'b0 ;
  assign n579 = x10 & ~n578 ;
  assign n580 = n317 ^ x137 ^ 1'b0 ;
  assign n581 = n564 & ~n580 ;
  assign n582 = x128 ^ x4 ^ 1'b0 ;
  assign n583 = n581 & n582 ;
  assign n588 = x211 & n452 ;
  assign n589 = ~x196 & n588 ;
  assign n584 = x61 & n365 ;
  assign n585 = n345 & n584 ;
  assign n586 = n521 | n585 ;
  assign n587 = n586 ^ n265 ^ 1'b0 ;
  assign n590 = n589 ^ n587 ^ 1'b0 ;
  assign n592 = x188 & x231 ;
  assign n593 = n592 ^ n514 ^ 1'b0 ;
  assign n591 = n257 & n538 ;
  assign n594 = n593 ^ n591 ^ 1'b0 ;
  assign n595 = n577 ^ n311 ^ 1'b0 ;
  assign n596 = x44 & x181 ;
  assign n597 = n538 & n596 ;
  assign n598 = n597 ^ n320 ^ x146 ;
  assign n599 = x22 & x69 ;
  assign n600 = n430 & n599 ;
  assign n601 = n600 ^ x118 ^ 1'b0 ;
  assign n602 = x100 & ~n601 ;
  assign n606 = x230 ^ x159 ^ 1'b0 ;
  assign n607 = x123 & n606 ;
  assign n604 = x7 & n304 ;
  assign n605 = n521 & n604 ;
  assign n603 = ~x49 & x115 ;
  assign n608 = n607 ^ n605 ^ n603 ;
  assign n609 = x189 ^ x133 ^ 1'b0 ;
  assign n610 = x56 & n609 ;
  assign n611 = ( ~x74 & x197 ) | ( ~x74 & n610 ) | ( x197 & n610 ) ;
  assign n612 = x81 & n611 ;
  assign n613 = n533 & n612 ;
  assign n614 = n583 ^ x71 ^ 1'b0 ;
  assign n615 = n387 & ~n614 ;
  assign n616 = n615 ^ n373 ^ 1'b0 ;
  assign n617 = x163 & x230 ;
  assign n618 = n617 ^ n343 ^ 1'b0 ;
  assign n619 = x92 ^ x89 ^ 1'b0 ;
  assign n620 = ~n294 & n619 ;
  assign n621 = n273 ^ x204 ^ x144 ;
  assign n622 = ~n355 & n621 ;
  assign n623 = ~n620 & n622 ;
  assign n624 = x233 & n337 ;
  assign n625 = n624 ^ n265 ^ 1'b0 ;
  assign n626 = ( ~x1 & x70 ) | ( ~x1 & n625 ) | ( x70 & n625 ) ;
  assign n627 = x186 & x224 ;
  assign n628 = n627 ^ x174 ^ 1'b0 ;
  assign n629 = n366 | n628 ;
  assign n630 = x217 ^ x71 ^ 1'b0 ;
  assign n631 = n630 ^ n277 ^ x56 ;
  assign n632 = n456 ^ n440 ^ 1'b0 ;
  assign n633 = x154 & n632 ;
  assign n634 = n288 & n561 ;
  assign n635 = n634 ^ x14 ^ 1'b0 ;
  assign n636 = x34 & x191 ;
  assign n637 = n636 ^ x154 ^ 1'b0 ;
  assign n638 = n637 ^ x244 ^ x174 ;
  assign n639 = n638 ^ x241 ^ 1'b0 ;
  assign n640 = n510 & ~n608 ;
  assign n641 = ~x127 & n640 ;
  assign n642 = ~x93 & x236 ;
  assign n643 = n504 ^ n417 ^ 1'b0 ;
  assign n644 = n620 ^ x189 ^ 1'b0 ;
  assign n645 = n532 ^ n279 ^ 1'b0 ;
  assign n646 = n535 ^ x66 ^ 1'b0 ;
  assign n647 = x18 & ~n646 ;
  assign n648 = n647 ^ n521 ^ n412 ;
  assign n649 = ( x17 & ~x195 ) | ( x17 & n361 ) | ( ~x195 & n361 ) ;
  assign n650 = x28 & x171 ;
  assign n651 = n368 & n650 ;
  assign n652 = x79 & ~n651 ;
  assign n653 = n652 ^ n549 ^ 1'b0 ;
  assign n654 = n653 ^ n510 ^ 1'b0 ;
  assign n655 = n649 & ~n654 ;
  assign n658 = x78 & x102 ;
  assign n659 = n658 ^ x82 ^ 1'b0 ;
  assign n660 = x90 & x212 ;
  assign n661 = n659 & n660 ;
  assign n656 = x16 & x190 ;
  assign n657 = n656 ^ x42 ^ 1'b0 ;
  assign n662 = n661 ^ n657 ^ 1'b0 ;
  assign n663 = x150 | n339 ;
  assign n665 = x92 ^ x86 ^ 1'b0 ;
  assign n666 = x137 & n665 ;
  assign n664 = x8 & ~n261 ;
  assign n667 = n666 ^ n664 ^ 1'b0 ;
  assign n668 = n450 & ~n667 ;
  assign n669 = n663 & n668 ;
  assign n670 = x27 & ~n456 ;
  assign n671 = ~x11 & n670 ;
  assign n672 = n502 ^ x53 ^ 1'b0 ;
  assign n673 = x74 ^ x68 ^ x13 ;
  assign n674 = x187 & ~n505 ;
  assign n675 = n674 ^ n357 ^ 1'b0 ;
  assign n676 = ~n673 & n675 ;
  assign n677 = n676 ^ x75 ^ 1'b0 ;
  assign n678 = x69 & x213 ;
  assign n679 = n678 ^ n257 ^ 1'b0 ;
  assign n680 = x147 & ~n679 ;
  assign n681 = ~x132 & n680 ;
  assign n682 = n288 & ~n681 ;
  assign n683 = n677 & n682 ;
  assign n684 = n683 ^ x2 ^ 1'b0 ;
  assign n685 = n672 | n684 ;
  assign n686 = ( x133 & x227 ) | ( x133 & n261 ) | ( x227 & n261 ) ;
  assign n687 = x198 & n305 ;
  assign n688 = n687 ^ n679 ^ 1'b0 ;
  assign n689 = x154 & n688 ;
  assign n690 = ~n686 & n689 ;
  assign n691 = x14 & n690 ;
  assign n692 = n360 ^ n307 ^ 1'b0 ;
  assign n693 = x83 & ~n374 ;
  assign n694 = n692 & n693 ;
  assign n695 = x58 & x84 ;
  assign n696 = n695 ^ n361 ^ 1'b0 ;
  assign n697 = n618 ^ n583 ^ 1'b0 ;
  assign n698 = n390 | n697 ;
  assign n699 = x32 ^ x9 ^ 1'b0 ;
  assign n700 = x40 & n699 ;
  assign n701 = ~x68 & n700 ;
  assign n703 = n514 ^ x142 ^ 1'b0 ;
  assign n704 = x44 & x46 ;
  assign n705 = ~n703 & n704 ;
  assign n706 = n390 | n705 ;
  assign n707 = n706 ^ x83 ^ 1'b0 ;
  assign n702 = x187 & x206 ;
  assign n708 = n707 ^ n702 ^ 1'b0 ;
  assign n709 = n290 & ~n613 ;
  assign n710 = n616 ^ x59 ^ 1'b0 ;
  assign n712 = x68 & n524 ;
  assign n713 = n712 ^ x138 ^ 1'b0 ;
  assign n714 = x43 & ~n713 ;
  assign n715 = ~n607 & n714 ;
  assign n716 = n302 & ~n715 ;
  assign n717 = n716 ^ n411 ^ 1'b0 ;
  assign n711 = x72 & x125 ;
  assign n718 = n717 ^ n711 ^ 1'b0 ;
  assign n719 = n718 ^ n691 ^ 1'b0 ;
  assign n720 = x170 & n719 ;
  assign n721 = n390 | n589 ;
  assign n722 = x222 | n721 ;
  assign n723 = x244 ^ x186 ^ 1'b0 ;
  assign n724 = n723 ^ x50 ^ 1'b0 ;
  assign n725 = x90 & ~n352 ;
  assign n726 = x2 & ~x37 ;
  assign n727 = n397 | n616 ;
  assign n728 = x95 | n727 ;
  assign n729 = n589 ^ n302 ^ 1'b0 ;
  assign n730 = x39 & x187 ;
  assign n745 = ~x59 & n333 ;
  assign n746 = n745 ^ x8 ^ 1'b0 ;
  assign n741 = n313 ^ n278 ^ 1'b0 ;
  assign n742 = n302 & n741 ;
  assign n743 = n481 & n742 ;
  assign n744 = x175 & n743 ;
  assign n738 = x46 & x57 ;
  assign n739 = x187 & n738 ;
  assign n740 = n536 & n739 ;
  assign n747 = n746 ^ n744 ^ n740 ;
  assign n731 = x100 & x249 ;
  assign n732 = ~x153 & n731 ;
  assign n733 = ~n514 & n732 ;
  assign n734 = n593 ^ x23 ^ 1'b0 ;
  assign n735 = x56 & ~n734 ;
  assign n736 = ~x169 & n735 ;
  assign n737 = n733 | n736 ;
  assign n748 = n747 ^ n737 ^ 1'b0 ;
  assign n749 = x75 | n747 ;
  assign n750 = x72 & x233 ;
  assign n751 = x15 & ~n526 ;
  assign n752 = ~n638 & n751 ;
  assign n753 = n503 ^ x44 ^ 1'b0 ;
  assign n754 = x123 & n307 ;
  assign n755 = n754 ^ x101 ^ 1'b0 ;
  assign n756 = x219 & n755 ;
  assign n757 = n548 ^ n385 ^ 1'b0 ;
  assign n758 = n361 | n757 ;
  assign n759 = n304 ^ n278 ^ 1'b0 ;
  assign n760 = x83 & ~n759 ;
  assign n761 = n296 | n685 ;
  assign n762 = n387 ^ x46 ^ 1'b0 ;
  assign n763 = x95 & x177 ;
  assign n764 = ~x0 & n763 ;
  assign n765 = x224 & n519 ;
  assign n766 = ~x51 & n765 ;
  assign n767 = x233 & n522 ;
  assign n768 = n767 ^ x72 ^ 1'b0 ;
  assign n769 = n768 ^ n754 ^ 1'b0 ;
  assign n770 = n766 | n769 ;
  assign n771 = ~x129 & x144 ;
  assign n772 = ( x169 & n351 ) | ( x169 & n771 ) | ( n351 & n771 ) ;
  assign n773 = n750 & n772 ;
  assign n774 = ~n446 & n773 ;
  assign n775 = n500 ^ n446 ^ 1'b0 ;
  assign n776 = ~n641 & n775 ;
  assign n777 = x221 ^ x60 ^ 1'b0 ;
  assign n778 = n776 & n777 ;
  assign n779 = n597 ^ x152 ^ 1'b0 ;
  assign n780 = n478 & n779 ;
  assign n781 = x136 ^ x1 ^ 1'b0 ;
  assign n782 = n585 ^ x57 ^ 1'b0 ;
  assign n783 = x135 & n420 ;
  assign n784 = ~n782 & n783 ;
  assign n785 = x86 & ~x107 ;
  assign n786 = x57 & ~x73 ;
  assign n787 = n614 & ~n690 ;
  assign n788 = ( ~x6 & x101 ) | ( ~x6 & n313 ) | ( x101 & n313 ) ;
  assign n789 = n486 & ~n788 ;
  assign n790 = x58 & n789 ;
  assign n791 = x87 & ~n488 ;
  assign n792 = ~n331 & n510 ;
  assign n793 = n792 ^ n300 ^ 1'b0 ;
  assign n794 = n686 & n793 ;
  assign n795 = ~n791 & n794 ;
  assign n796 = n552 & ~n795 ;
  assign n797 = x91 & x185 ;
  assign n798 = n797 ^ x236 ^ 1'b0 ;
  assign n799 = x236 ^ x149 ^ 1'b0 ;
  assign n800 = ~n380 & n799 ;
  assign n801 = n736 ^ x83 ^ 1'b0 ;
  assign n802 = ~x41 & x161 ;
  assign n803 = ~n307 & n802 ;
  assign n804 = ~n313 & n561 ;
  assign n805 = ~x137 & n804 ;
  assign n806 = n495 | n805 ;
  assign n807 = x38 & n806 ;
  assign n808 = n807 ^ x203 ^ 1'b0 ;
  assign n809 = ~x111 & x252 ;
  assign n810 = ~x42 & x101 ;
  assign n811 = n810 ^ x125 ^ 1'b0 ;
  assign n812 = x32 & ~n811 ;
  assign n813 = x154 & n335 ;
  assign n814 = ~x104 & x109 ;
  assign n815 = n813 & ~n814 ;
  assign n816 = n812 & n815 ;
  assign n817 = n561 & ~n816 ;
  assign n819 = x186 & ~n474 ;
  assign n820 = ~x140 & n819 ;
  assign n818 = n445 ^ n278 ^ 1'b0 ;
  assign n821 = n820 ^ n818 ^ 1'b0 ;
  assign n822 = ( x9 & x40 ) | ( x9 & ~x202 ) | ( x40 & ~x202 ) ;
  assign n823 = n277 & n822 ;
  assign n824 = ~n519 & n823 ;
  assign n825 = n824 ^ n672 ^ 1'b0 ;
  assign n826 = x247 & ~n352 ;
  assign n827 = n826 ^ n271 ^ 1'b0 ;
  assign n828 = n789 ^ x59 ^ 1'b0 ;
  assign n829 = ( x115 & n631 ) | ( x115 & n828 ) | ( n631 & n828 ) ;
  assign n830 = n300 | n663 ;
  assign n831 = x18 & x174 ;
  assign n832 = n831 ^ n566 ^ 1'b0 ;
  assign n833 = x194 & n832 ;
  assign n834 = n587 ^ x92 ^ 1'b0 ;
  assign n835 = x150 & n834 ;
  assign n840 = x189 ^ x96 ^ x38 ;
  assign n841 = x110 & ~n840 ;
  assign n836 = ~x82 & x193 ;
  assign n837 = n395 ^ x12 ^ 1'b0 ;
  assign n838 = n836 & ~n837 ;
  assign n839 = ~n279 & n838 ;
  assign n842 = n841 ^ n839 ^ 1'b0 ;
  assign n843 = n442 ^ x156 ^ 1'b0 ;
  assign n844 = x217 & ~n843 ;
  assign n845 = x167 & n648 ;
  assign n846 = ~n844 & n845 ;
  assign n847 = n722 & ~n846 ;
  assign n848 = ~n812 & n847 ;
  assign n849 = n700 ^ n522 ^ 1'b0 ;
  assign n850 = x90 & ~n828 ;
  assign n851 = n533 & n850 ;
  assign n852 = n851 ^ n399 ^ 1'b0 ;
  assign n853 = x46 & ~n852 ;
  assign n854 = ~x33 & x108 ;
  assign n855 = n854 ^ n628 ^ x222 ;
  assign n857 = x227 & n512 ;
  assign n858 = ~n793 & n857 ;
  assign n856 = n552 & n752 ;
  assign n859 = n858 ^ n856 ^ 1'b0 ;
  assign n860 = n405 ^ x104 ^ 1'b0 ;
  assign n861 = x213 ^ x115 ^ 1'b0 ;
  assign n862 = n329 | n861 ;
  assign n863 = n648 | n673 ;
  assign n864 = x217 | n862 ;
  assign n865 = x127 & ~n279 ;
  assign n866 = n865 ^ n538 ^ 1'b0 ;
  assign n867 = ~x43 & n866 ;
  assign n868 = x210 & n265 ;
  assign n869 = n868 ^ n564 ^ 1'b0 ;
  assign n870 = n816 ^ n671 ^ 1'b0 ;
  assign n871 = n869 | n870 ;
  assign n872 = x34 & ~x219 ;
  assign n873 = x244 & n872 ;
  assign n874 = n768 & n873 ;
  assign n875 = n444 ^ x202 ^ 1'b0 ;
  assign n876 = ~n381 & n875 ;
  assign n877 = n495 ^ n277 ^ x159 ;
  assign n878 = n812 ^ x126 ^ 1'b0 ;
  assign n879 = ~n877 & n878 ;
  assign n880 = x62 & ~n879 ;
  assign n881 = n840 ^ n273 ^ 1'b0 ;
  assign n882 = x228 ^ x70 ^ 1'b0 ;
  assign n883 = x18 & n882 ;
  assign n884 = n373 ^ x246 ^ 1'b0 ;
  assign n885 = n884 ^ n651 ^ 1'b0 ;
  assign n886 = n267 & ~n885 ;
  assign n887 = x175 & ~x213 ;
  assign n888 = n860 | n887 ;
  assign n890 = n620 ^ x221 ^ 1'b0 ;
  assign n891 = ~n573 & n890 ;
  assign n889 = n296 & n593 ;
  assign n892 = n891 ^ n889 ^ 1'b0 ;
  assign n893 = n551 | n892 ;
  assign n894 = n893 ^ x57 ^ 1'b0 ;
  assign n895 = x13 & ~n894 ;
  assign n896 = x148 & n895 ;
  assign n897 = x249 ^ x163 ^ 1'b0 ;
  assign n898 = n897 ^ x156 ^ 1'b0 ;
  assign n899 = n779 & ~n898 ;
  assign n900 = n899 ^ x22 ^ 1'b0 ;
  assign n901 = x84 | n900 ;
  assign n902 = x13 & x34 ;
  assign n903 = n902 ^ x41 ^ 1'b0 ;
  assign n904 = ( ~x18 & n856 ) | ( ~x18 & n903 ) | ( n856 & n903 ) ;
  assign n905 = ~x176 & n509 ;
  assign n906 = n436 ^ x183 ^ 1'b0 ;
  assign n907 = n905 | n906 ;
  assign n910 = n267 ^ x244 ^ 1'b0 ;
  assign n911 = n385 & n910 ;
  assign n908 = n385 & ~n414 ;
  assign n909 = ~n465 & n908 ;
  assign n912 = n911 ^ n909 ^ 1'b0 ;
  assign n913 = n907 | n912 ;
  assign n914 = n300 | n358 ;
  assign n915 = n914 ^ n370 ^ 1'b0 ;
  assign n916 = ~n875 & n915 ;
  assign n917 = ~x168 & n916 ;
  assign n918 = n490 | n917 ;
  assign n919 = n417 ^ x144 ^ 1'b0 ;
  assign n920 = x115 & n919 ;
  assign n921 = x168 & n920 ;
  assign n922 = n440 ^ x108 ^ 1'b0 ;
  assign n923 = x37 & ~n922 ;
  assign n924 = ~x19 & n277 ;
  assign n925 = x5 & x23 ;
  assign n926 = n925 ^ n521 ^ 1'b0 ;
  assign n927 = x70 & ~n926 ;
  assign n928 = ~n381 & n647 ;
  assign n929 = n512 | n851 ;
  assign n930 = ( x68 & n341 ) | ( x68 & ~n438 ) | ( n341 & ~n438 ) ;
  assign n931 = x222 & ~n930 ;
  assign n932 = ~n269 & n281 ;
  assign n933 = ~n931 & n932 ;
  assign n934 = ~n394 & n933 ;
  assign n935 = n318 ^ x88 ^ 1'b0 ;
  assign n936 = x165 & n935 ;
  assign n937 = n936 ^ n360 ^ 1'b0 ;
  assign n938 = x251 & n318 ;
  assign n939 = n937 & n938 ;
  assign n940 = n581 ^ x58 ^ 1'b0 ;
  assign n941 = x88 & n940 ;
  assign n942 = ~n939 & n941 ;
  assign n943 = n942 ^ x217 ^ 1'b0 ;
  assign n944 = n587 & n943 ;
  assign n945 = n585 ^ n512 ^ 1'b0 ;
  assign n946 = n445 & ~n945 ;
  assign n947 = x236 & ~n535 ;
  assign n948 = n659 & n947 ;
  assign n949 = x19 & ~n948 ;
  assign n950 = n949 ^ n259 ^ 1'b0 ;
  assign n951 = n950 ^ n486 ^ 1'b0 ;
  assign n953 = x102 & ~n600 ;
  assign n954 = n259 & n953 ;
  assign n952 = n343 & ~n543 ;
  assign n955 = n954 ^ n952 ^ 1'b0 ;
  assign n956 = ( ~x210 & n603 ) | ( ~x210 & n955 ) | ( n603 & n955 ) ;
  assign n957 = ~x139 & x165 ;
  assign n958 = ~x42 & x167 ;
  assign n962 = n476 ^ x150 ^ 1'b0 ;
  assign n963 = n448 | n962 ;
  assign n961 = x131 & n620 ;
  assign n964 = n963 ^ n961 ^ 1'b0 ;
  assign n959 = n651 & ~n752 ;
  assign n960 = n397 & ~n959 ;
  assign n965 = n964 ^ n960 ^ 1'b0 ;
  assign n966 = n373 | n965 ;
  assign n967 = x39 | n360 ;
  assign n968 = x143 | n846 ;
  assign n969 = n968 ^ n374 ^ 1'b0 ;
  assign n970 = n686 ^ n653 ^ 1'b0 ;
  assign n971 = n552 | n970 ;
  assign n972 = ~x47 & x50 ;
  assign n973 = x167 & ~n972 ;
  assign n974 = n973 ^ n524 ^ 1'b0 ;
  assign n975 = x220 & ~n974 ;
  assign n976 = x136 & ~n600 ;
  assign n977 = ~x182 & n976 ;
  assign n978 = n977 ^ n566 ^ 1'b0 ;
  assign n979 = n975 & n978 ;
  assign n980 = x179 & ~n323 ;
  assign n981 = ~x130 & n980 ;
  assign n982 = x34 & ~n551 ;
  assign n983 = n758 & n982 ;
  assign n986 = x158 & n686 ;
  assign n987 = n986 ^ n805 ^ 1'b0 ;
  assign n984 = n384 ^ x158 ^ 1'b0 ;
  assign n985 = n411 | n984 ;
  assign n988 = n987 ^ n985 ^ 1'b0 ;
  assign n989 = x230 & n701 ;
  assign n990 = x239 ^ x205 ^ x163 ;
  assign n991 = x190 & n269 ;
  assign n992 = n990 & n991 ;
  assign n993 = x28 & x47 ;
  assign n994 = n993 ^ x147 ^ 1'b0 ;
  assign n995 = x149 & n994 ;
  assign n996 = n995 ^ n535 ^ 1'b0 ;
  assign n997 = n996 ^ n527 ^ 1'b0 ;
  assign n998 = ~n992 & n997 ;
  assign n999 = x234 & n581 ;
  assign n1000 = n990 & n999 ;
  assign n1001 = x65 & x76 ;
  assign n1002 = n514 & n1001 ;
  assign n1003 = n581 & ~n1002 ;
  assign n1004 = n1000 & n1003 ;
  assign n1005 = n771 & ~n1004 ;
  assign n1006 = n1005 ^ n663 ^ 1'b0 ;
  assign n1007 = x7 & ~n1006 ;
  assign n1008 = n844 & n899 ;
  assign n1009 = n1008 ^ n915 ^ 1'b0 ;
  assign n1010 = x231 & ~n620 ;
  assign n1011 = x191 & n1010 ;
  assign n1012 = n1011 ^ n535 ^ 1'b0 ;
  assign n1013 = n968 ^ x46 ^ 1'b0 ;
  assign n1014 = n1012 & ~n1013 ;
  assign n1015 = x205 & ~n539 ;
  assign n1016 = ~n1014 & n1015 ;
  assign n1017 = n543 ^ x150 ^ 1'b0 ;
  assign n1018 = n1017 ^ n620 ^ 1'b0 ;
  assign n1019 = n643 ^ n440 ^ 1'b0 ;
  assign n1020 = n1018 & ~n1019 ;
  assign n1021 = n1020 ^ n313 ^ 1'b0 ;
  assign n1022 = n1021 ^ n545 ^ 1'b0 ;
  assign n1023 = ~n934 & n1022 ;
  assign n1024 = n992 ^ x48 ^ 1'b0 ;
  assign n1025 = n1023 & ~n1024 ;
  assign n1026 = n292 ^ n290 ^ 1'b0 ;
  assign n1027 = n349 | n1026 ;
  assign n1028 = n616 & ~n1027 ;
  assign n1029 = n385 & n505 ;
  assign n1030 = n1028 & n1029 ;
  assign n1031 = ~x125 & n1030 ;
  assign n1032 = ~n290 & n298 ;
  assign n1033 = n1032 ^ n798 ^ 1'b0 ;
  assign n1034 = n641 ^ n450 ^ 1'b0 ;
  assign n1035 = n500 & ~n1034 ;
  assign n1036 = n598 | n603 ;
  assign n1037 = n1036 ^ x248 ^ 1'b0 ;
  assign n1038 = n426 & n994 ;
  assign n1039 = x198 ^ x151 ^ 1'b0 ;
  assign n1041 = n341 ^ x50 ^ 1'b0 ;
  assign n1042 = x169 & ~n1041 ;
  assign n1043 = n688 ^ x32 ^ 1'b0 ;
  assign n1044 = n1042 & n1043 ;
  assign n1040 = n771 ^ n673 ^ x127 ;
  assign n1045 = n1044 ^ n1040 ^ 1'b0 ;
  assign n1046 = ~n1039 & n1045 ;
  assign n1047 = n1046 ^ x113 ^ 1'b0 ;
  assign n1048 = n788 ^ n351 ^ 1'b0 ;
  assign n1049 = ~x151 & n392 ;
  assign n1050 = n1048 & n1049 ;
  assign n1051 = x214 ^ x45 ^ 1'b0 ;
  assign n1052 = x205 & n1051 ;
  assign n1053 = n1052 ^ x158 ^ 1'b0 ;
  assign n1054 = ~n533 & n1053 ;
  assign n1055 = x153 & ~n877 ;
  assign n1056 = ~n417 & n1055 ;
  assign n1057 = n994 | n1056 ;
  assign n1058 = x226 | n1057 ;
  assign n1059 = x208 ^ x63 ^ 1'b0 ;
  assign n1060 = x247 & ~n1059 ;
  assign n1061 = n311 & n1060 ;
  assign n1062 = n415 ^ x147 ^ 1'b0 ;
  assign n1063 = x21 & n1062 ;
  assign n1064 = n663 & n1063 ;
  assign n1065 = n1064 ^ n673 ^ 1'b0 ;
  assign n1066 = n623 ^ n278 ^ 1'b0 ;
  assign n1067 = n415 & ~n516 ;
  assign n1068 = ~n446 & n1067 ;
  assign n1069 = n771 ^ n380 ^ 1'b0 ;
  assign n1070 = n931 | n1069 ;
  assign n1071 = n1068 & ~n1070 ;
  assign n1072 = n1039 | n1071 ;
  assign n1073 = n1072 ^ n738 ^ 1'b0 ;
  assign n1075 = ~x66 & x114 ;
  assign n1074 = x99 & n570 ;
  assign n1076 = n1075 ^ n1074 ^ 1'b0 ;
  assign n1077 = n397 & n741 ;
  assign n1078 = n796 | n1077 ;
  assign n1079 = n1076 & ~n1078 ;
  assign n1080 = n323 & ~n440 ;
  assign n1081 = ~x158 & x181 ;
  assign n1082 = n1081 ^ n1059 ^ n456 ;
  assign n1083 = n307 ^ x233 ^ 1'b0 ;
  assign n1084 = n669 ^ x218 ^ 1'b0 ;
  assign n1085 = n1047 & ~n1084 ;
  assign n1086 = n1085 ^ x225 ^ 1'b0 ;
  assign n1087 = ~n1083 & n1086 ;
  assign n1088 = n577 ^ n397 ^ 1'b0 ;
  assign n1089 = n867 & n1088 ;
  assign n1090 = n305 & ~n497 ;
  assign n1091 = n1090 ^ n322 ^ 1'b0 ;
  assign n1092 = x1 & x120 ;
  assign n1093 = n421 & n1092 ;
  assign n1094 = ( ~n539 & n1091 ) | ( ~n539 & n1093 ) | ( n1091 & n1093 ) ;
  assign n1095 = n858 ^ n643 ^ 1'b0 ;
  assign n1096 = n1094 & ~n1095 ;
  assign n1097 = n585 | n659 ;
  assign n1098 = n1097 ^ n307 ^ 1'b0 ;
  assign n1099 = x149 & n286 ;
  assign n1100 = ~n390 & n1099 ;
  assign n1101 = x22 & ~n322 ;
  assign n1102 = n1101 ^ n744 ^ 1'b0 ;
  assign n1103 = n1100 & n1102 ;
  assign n1104 = n1103 ^ x79 ^ 1'b0 ;
  assign n1105 = ~n397 & n495 ;
  assign n1106 = n611 ^ x98 ^ 1'b0 ;
  assign n1110 = x200 ^ x153 ^ 1'b0 ;
  assign n1111 = n666 & n1110 ;
  assign n1107 = x158 & ~n381 ;
  assign n1108 = ~n373 & n1107 ;
  assign n1109 = n635 | n1108 ;
  assign n1112 = n1111 ^ n1109 ^ 1'b0 ;
  assign n1113 = n796 ^ n790 ^ 1'b0 ;
  assign n1114 = n1029 & n1113 ;
  assign n1115 = ~n671 & n1044 ;
  assign n1116 = n1115 ^ x195 ^ 1'b0 ;
  assign n1117 = ( x82 & ~n502 ) | ( x82 & n1116 ) | ( ~n502 & n1116 ) ;
  assign n1118 = x152 & n1117 ;
  assign n1119 = n829 | n1004 ;
  assign n1120 = x107 | n1119 ;
  assign n1123 = n343 & n549 ;
  assign n1124 = x254 & n1123 ;
  assign n1122 = x70 & n593 ;
  assign n1125 = n1124 ^ n1122 ^ 1'b0 ;
  assign n1121 = x177 & ~n1056 ;
  assign n1126 = n1125 ^ n1121 ^ 1'b0 ;
  assign n1127 = x103 & x151 ;
  assign n1128 = ~x83 & n1127 ;
  assign n1129 = n694 ^ n372 ^ 1'b0 ;
  assign n1130 = n1128 | n1129 ;
  assign n1131 = n1116 ^ n620 ^ 1'b0 ;
  assign n1132 = ~n539 & n607 ;
  assign n1133 = n1132 ^ n450 ^ 1'b0 ;
  assign n1134 = x107 | n1133 ;
  assign n1135 = n1134 ^ x112 ^ 1'b0 ;
  assign n1136 = n1096 ^ n842 ^ 1'b0 ;
  assign n1137 = x92 & ~n1136 ;
  assign n1138 = x72 & x227 ;
  assign n1139 = n1138 ^ n271 ^ 1'b0 ;
  assign n1140 = ~n376 & n1139 ;
  assign n1141 = ~x164 & n1140 ;
  assign n1142 = x245 & n649 ;
  assign n1143 = ~x96 & n1142 ;
  assign n1144 = x205 & n372 ;
  assign n1145 = n1144 ^ n1139 ^ 1'b0 ;
  assign n1146 = ( n813 & ~n1143 ) | ( n813 & n1145 ) | ( ~n1143 & n1145 ) ;
  assign n1147 = n1146 ^ n438 ^ 1'b0 ;
  assign n1148 = x53 & n1147 ;
  assign n1149 = x134 & ~n349 ;
  assign n1150 = n1149 ^ n748 ^ 1'b0 ;
  assign n1151 = x192 & n593 ;
  assign n1152 = ~n354 & n1151 ;
  assign n1153 = n594 | n1152 ;
  assign n1154 = n1153 ^ n841 ^ 1'b0 ;
  assign n1160 = n378 ^ x90 ^ 1'b0 ;
  assign n1155 = x2 & x241 ;
  assign n1156 = n1155 ^ x19 ^ 1'b0 ;
  assign n1157 = n1156 ^ x150 ^ 1'b0 ;
  assign n1158 = x233 & ~n1157 ;
  assign n1159 = n281 & n1158 ;
  assign n1161 = n1160 ^ n1159 ^ 1'b0 ;
  assign n1162 = n1154 & ~n1161 ;
  assign n1163 = n1162 ^ n1112 ^ 1'b0 ;
  assign n1164 = ~n1064 & n1163 ;
  assign n1165 = n551 & n1012 ;
  assign n1166 = n833 & n855 ;
  assign n1167 = n1166 ^ n734 ^ 1'b0 ;
  assign n1168 = n1035 ^ n296 ^ 1'b0 ;
  assign n1169 = n869 | n1168 ;
  assign n1170 = n395 & n866 ;
  assign n1171 = x170 & ~n768 ;
  assign n1172 = n1170 & n1171 ;
  assign n1173 = ~x156 & n876 ;
  assign n1179 = n1158 ^ x59 ^ 1'b0 ;
  assign n1180 = x96 & n1179 ;
  assign n1181 = n1180 ^ n1152 ^ 1'b0 ;
  assign n1177 = x167 & ~n508 ;
  assign n1178 = n1059 & n1177 ;
  assign n1174 = x239 & n488 ;
  assign n1175 = n709 | n1174 ;
  assign n1176 = n1035 & ~n1175 ;
  assign n1182 = n1181 ^ n1178 ^ n1176 ;
  assign n1188 = ~n671 & n708 ;
  assign n1189 = x254 ^ x113 ^ 1'b0 ;
  assign n1190 = n1188 | n1189 ;
  assign n1183 = x129 & ~x253 ;
  assign n1184 = x155 & n1183 ;
  assign n1185 = n1085 ^ x227 ^ 1'b0 ;
  assign n1186 = ~n815 & n1185 ;
  assign n1187 = ~n1184 & n1186 ;
  assign n1191 = n1190 ^ n1187 ^ 1'b0 ;
  assign n1192 = n500 ^ x59 ^ 1'b0 ;
  assign n1193 = n1192 ^ n415 ^ 1'b0 ;
  assign n1194 = n463 & ~n1193 ;
  assign n1195 = n595 ^ x251 ^ 1'b0 ;
  assign n1196 = n818 ^ x45 ^ 1'b0 ;
  assign n1197 = x152 & ~n1196 ;
  assign n1198 = x207 & n1197 ;
  assign n1199 = n618 & ~n989 ;
  assign n1200 = ~n805 & n1018 ;
  assign n1201 = n1200 ^ n625 ^ 1'b0 ;
  assign n1202 = n754 & ~n1201 ;
  assign n1203 = ~n283 & n566 ;
  assign n1204 = n1203 ^ n474 ^ 1'b0 ;
  assign n1205 = x15 & ~n300 ;
  assign n1206 = n645 & ~n1205 ;
  assign n1207 = ~x99 & n1206 ;
  assign n1208 = n1204 | n1207 ;
  assign n1209 = n936 & n1208 ;
  assign n1210 = n1209 ^ x206 ^ 1'b0 ;
  assign n1211 = x4 & n337 ;
  assign n1212 = n1211 ^ x116 ^ 1'b0 ;
  assign n1213 = n616 | n1212 ;
  assign n1214 = n1213 ^ x241 ^ 1'b0 ;
  assign n1215 = ~n1210 & n1214 ;
  assign n1216 = n1215 ^ n1159 ^ 1'b0 ;
  assign n1217 = n347 & ~n1216 ;
  assign n1223 = ~x50 & n872 ;
  assign n1218 = x110 & n412 ;
  assign n1219 = ~x41 & n1218 ;
  assign n1220 = ~n1056 & n1159 ;
  assign n1221 = n1220 ^ x203 ^ 1'b0 ;
  assign n1222 = n1219 | n1221 ;
  assign n1224 = n1223 ^ n1222 ^ 1'b0 ;
  assign n1225 = n842 | n1224 ;
  assign n1226 = x61 | n1225 ;
  assign n1227 = n879 & ~n1226 ;
  assign n1228 = n937 ^ x55 ^ 1'b0 ;
  assign n1229 = n1228 ^ n1128 ^ 1'b0 ;
  assign n1230 = n669 | n1229 ;
  assign n1231 = x75 & x157 ;
  assign n1232 = ~n540 & n1231 ;
  assign n1233 = n446 & ~n1232 ;
  assign n1234 = n1233 ^ x168 ^ 1'b0 ;
  assign n1235 = n880 & ~n1198 ;
  assign n1236 = ~x243 & n1235 ;
  assign n1237 = n610 ^ n288 ^ 1'b0 ;
  assign n1238 = ~x23 & n1237 ;
  assign n1239 = n440 & n1238 ;
  assign n1240 = n349 ^ x158 ^ 1'b0 ;
  assign n1241 = n1077 ^ n302 ^ 1'b0 ;
  assign n1242 = n1241 ^ n860 ^ x113 ;
  assign n1243 = x196 ^ x170 ^ 1'b0 ;
  assign n1244 = x138 & n292 ;
  assign n1245 = n1243 & n1244 ;
  assign n1246 = n1245 ^ n1170 ^ 1'b0 ;
  assign n1247 = n1242 & n1246 ;
  assign n1248 = ( x210 & n355 ) | ( x210 & n972 ) | ( n355 & n972 ) ;
  assign n1249 = n1044 ^ n789 ^ 1'b0 ;
  assign n1254 = n355 ^ x40 ^ 1'b0 ;
  assign n1255 = n331 | n1254 ;
  assign n1250 = n977 ^ x14 ^ 1'b0 ;
  assign n1251 = n946 & ~n1250 ;
  assign n1252 = n498 & ~n923 ;
  assign n1253 = n1251 & n1252 ;
  assign n1256 = n1255 ^ n1253 ^ 1'b0 ;
  assign n1259 = x14 & ~n1039 ;
  assign n1260 = ~x175 & n1259 ;
  assign n1257 = n577 | n871 ;
  assign n1258 = n1257 ^ n1094 ^ 1'b0 ;
  assign n1261 = n1260 ^ n1258 ^ 1'b0 ;
  assign n1262 = n618 ^ x73 ^ 1'b0 ;
  assign n1263 = x15 & x44 ;
  assign n1264 = n723 ^ x234 ^ 1'b0 ;
  assign n1265 = n454 & n540 ;
  assign n1266 = ~n844 & n1265 ;
  assign n1267 = n1264 & n1266 ;
  assign n1268 = n288 ^ x33 ^ 1'b0 ;
  assign n1269 = x115 | n1268 ;
  assign n1270 = x142 & x191 ;
  assign n1271 = n518 & n1270 ;
  assign n1272 = n1271 ^ n789 ^ 1'b0 ;
  assign n1273 = n1027 ^ x61 ^ 1'b0 ;
  assign n1274 = n782 ^ x139 ^ 1'b0 ;
  assign n1275 = n1273 & n1274 ;
  assign n1276 = ~n1272 & n1275 ;
  assign n1277 = n1276 ^ n1174 ^ 1'b0 ;
  assign n1278 = n474 | n542 ;
  assign n1279 = ~n810 & n879 ;
  assign n1280 = ~x233 & n1279 ;
  assign n1281 = x77 & ~n474 ;
  assign n1282 = ~n568 & n1281 ;
  assign n1283 = n397 | n585 ;
  assign n1284 = n1173 & ~n1283 ;
  assign n1285 = n1282 & n1284 ;
  assign n1286 = n989 ^ x225 ^ 1'b0 ;
  assign n1287 = x171 & ~n705 ;
  assign n1288 = ~n772 & n1287 ;
  assign n1289 = n907 | n1288 ;
  assign n1290 = n605 & ~n1289 ;
  assign n1291 = n675 ^ n666 ^ 1'b0 ;
  assign n1292 = x189 & n420 ;
  assign n1293 = n921 & n1292 ;
  assign n1294 = n1191 & ~n1293 ;
  assign n1295 = n1294 ^ x210 ^ 1'b0 ;
  assign n1296 = n948 ^ n677 ^ 1'b0 ;
  assign n1297 = ~n1295 & n1296 ;
  assign n1298 = n1195 ^ x76 ^ 1'b0 ;
  assign n1299 = ~x116 & n1233 ;
  assign n1300 = n1299 ^ n358 ^ 1'b0 ;
  assign n1301 = n924 & n1300 ;
  assign n1302 = n1278 ^ x96 ^ 1'b0 ;
  assign n1303 = n669 | n956 ;
  assign n1304 = n1128 & ~n1303 ;
  assign n1305 = ~n514 & n1156 ;
  assign n1309 = n504 ^ n341 ^ 1'b0 ;
  assign n1310 = n666 & n1309 ;
  assign n1306 = x2 & ~n296 ;
  assign n1307 = n1205 & n1306 ;
  assign n1308 = n1307 ^ n504 ^ x84 ;
  assign n1311 = n1310 ^ n1308 ^ 1'b0 ;
  assign n1312 = x50 & n512 ;
  assign n1313 = x113 & ~n729 ;
  assign n1314 = ~n343 & n703 ;
  assign n1315 = n641 ^ x188 ^ 1'b0 ;
  assign n1316 = n1314 | n1315 ;
  assign n1317 = n1313 & ~n1316 ;
  assign n1318 = n1317 ^ n1156 ^ 1'b0 ;
  assign n1323 = n1233 ^ n376 ^ 1'b0 ;
  assign n1324 = n539 | n1323 ;
  assign n1319 = x94 & n365 ;
  assign n1320 = ~x103 & n1319 ;
  assign n1321 = n1320 ^ n621 ^ n399 ;
  assign n1322 = ~n669 & n1321 ;
  assign n1325 = n1324 ^ n1322 ^ 1'b0 ;
  assign n1326 = n1325 ^ x149 ^ x102 ;
  assign n1327 = n1326 ^ n351 ^ 1'b0 ;
  assign n1328 = n568 ^ x25 ^ 1'b0 ;
  assign n1329 = n778 ^ n290 ^ 1'b0 ;
  assign n1330 = n1031 | n1329 ;
  assign n1331 = x94 & x107 ;
  assign n1332 = n1331 ^ x15 ^ 1'b0 ;
  assign n1333 = ( ~x105 & x175 ) | ( ~x105 & n1332 ) | ( x175 & n1332 ) ;
  assign n1334 = ~n994 & n1333 ;
  assign n1335 = n807 & n1065 ;
  assign n1336 = n1263 ^ x61 ^ 1'b0 ;
  assign n1337 = n928 ^ n559 ^ 1'b0 ;
  assign n1340 = x32 & ~n907 ;
  assign n1341 = ~n866 & n1340 ;
  assign n1342 = x73 & ~n1341 ;
  assign n1343 = n1342 ^ n688 ^ 1'b0 ;
  assign n1338 = x175 & ~n895 ;
  assign n1339 = ~x252 & n1338 ;
  assign n1344 = n1343 ^ n1339 ^ 1'b0 ;
  assign n1345 = ~n1039 & n1280 ;
  assign n1346 = x208 ^ x139 ^ 1'b0 ;
  assign n1347 = n785 ^ n672 ^ n329 ;
  assign n1348 = ~x71 & n1347 ;
  assign n1349 = n1346 & ~n1348 ;
  assign n1350 = n1349 ^ x233 ^ 1'b0 ;
  assign n1351 = x77 & ~n351 ;
  assign n1352 = n809 | n1028 ;
  assign n1353 = n320 ^ x244 ^ 1'b0 ;
  assign n1354 = n452 | n1255 ;
  assign n1355 = n958 ^ n871 ^ 1'b0 ;
  assign n1356 = n766 | n1355 ;
  assign n1357 = n1356 ^ x103 ^ 1'b0 ;
  assign n1358 = x131 & ~n1357 ;
  assign n1359 = x202 & ~n1143 ;
  assign n1360 = n1359 ^ n1271 ^ 1'b0 ;
  assign n1361 = n546 & n1360 ;
  assign n1362 = ~n698 & n806 ;
  assign n1363 = n1362 ^ x246 ^ 1'b0 ;
  assign n1364 = n387 & n581 ;
  assign n1365 = n977 & n1364 ;
  assign n1369 = x32 & ~x66 ;
  assign n1366 = ~n257 & n643 ;
  assign n1367 = n732 | n1366 ;
  assign n1368 = n915 | n1367 ;
  assign n1370 = n1369 ^ n1368 ^ x72 ;
  assign n1371 = ~n1365 & n1370 ;
  assign n1372 = ~x66 & n1371 ;
  assign n1373 = x3 & n1223 ;
  assign n1374 = n1373 ^ n1217 ^ 1'b0 ;
  assign n1375 = n259 ^ x24 ^ 1'b0 ;
  assign n1376 = n791 & ~n1375 ;
  assign n1377 = ~n460 & n1376 ;
  assign n1378 = n1377 ^ n1268 ^ 1'b0 ;
  assign n1379 = x245 & ~n331 ;
  assign n1380 = x182 | n1356 ;
  assign n1381 = x234 & n967 ;
  assign n1382 = n1176 | n1381 ;
  assign n1386 = x28 & x191 ;
  assign n1387 = ~n508 & n1386 ;
  assign n1383 = n1031 ^ n641 ^ 1'b0 ;
  assign n1384 = n887 | n1383 ;
  assign n1385 = n1384 ^ n738 ^ 1'b0 ;
  assign n1388 = n1387 ^ n1385 ^ 1'b0 ;
  assign n1389 = x165 & ~n1388 ;
  assign n1390 = ~x61 & x171 ;
  assign n1391 = n605 ^ n259 ^ x28 ;
  assign n1392 = x107 & ~n1391 ;
  assign n1393 = n1392 ^ x101 ^ 1'b0 ;
  assign n1394 = n877 ^ n581 ^ 1'b0 ;
  assign n1395 = n1393 | n1394 ;
  assign n1396 = n436 ^ x178 ^ 1'b0 ;
  assign n1397 = n378 & ~n1396 ;
  assign n1398 = n415 & ~n551 ;
  assign n1399 = n1398 ^ x90 ^ 1'b0 ;
  assign n1400 = n292 | n1399 ;
  assign n1401 = n587 ^ x112 ^ 1'b0 ;
  assign n1402 = x71 & n1401 ;
  assign n1403 = x30 & ~n472 ;
  assign n1404 = ~x146 & n1403 ;
  assign n1405 = n1044 & n1404 ;
  assign n1406 = x241 & ~n1405 ;
  assign n1407 = ~n1402 & n1406 ;
  assign n1408 = n1365 ^ n779 ^ 1'b0 ;
  assign n1409 = x138 & ~n1408 ;
  assign n1410 = ( n666 & n1280 ) | ( n666 & ~n1409 ) | ( n1280 & ~n1409 ) ;
  assign n1411 = ~n566 & n1233 ;
  assign n1412 = n1256 ^ x185 ^ 1'b0 ;
  assign n1413 = ~n1116 & n1412 ;
  assign n1414 = ~n1411 & n1413 ;
  assign n1415 = n955 & n1143 ;
  assign n1416 = x7 & x234 ;
  assign n1417 = n1416 ^ x230 ^ 1'b0 ;
  assign n1418 = n748 | n1417 ;
  assign n1419 = n1418 ^ n594 ^ 1'b0 ;
  assign n1420 = n510 & ~n1419 ;
  assign n1421 = n1405 & n1420 ;
  assign n1425 = n1326 ^ n1156 ^ 1'b0 ;
  assign n1426 = x158 & n1425 ;
  assign n1422 = n552 ^ n442 ^ 1'b0 ;
  assign n1423 = x230 & ~n1422 ;
  assign n1424 = n1325 & ~n1423 ;
  assign n1427 = n1426 ^ n1424 ^ n1385 ;
  assign n1428 = n450 ^ x111 ^ 1'b0 ;
  assign n1429 = x239 & n1428 ;
  assign n1430 = n1429 ^ x46 ^ 1'b0 ;
  assign n1431 = n1080 & n1430 ;
  assign n1432 = n456 | n1332 ;
  assign n1433 = x66 | n1432 ;
  assign n1434 = x61 & n1433 ;
  assign n1435 = n1434 ^ x167 ^ 1'b0 ;
  assign n1436 = n778 & ~n1435 ;
  assign n1437 = n638 ^ x8 ^ 1'b0 ;
  assign n1438 = x226 & n1437 ;
  assign n1439 = ~n358 & n1438 ;
  assign n1440 = n1439 ^ x222 ^ 1'b0 ;
  assign n1441 = n1440 ^ n269 ^ 1'b0 ;
  assign n1442 = n1158 & n1441 ;
  assign n1443 = ( x9 & ~n926 ) | ( x9 & n1093 ) | ( ~n926 & n1093 ) ;
  assign n1444 = n1442 & n1443 ;
  assign n1445 = n1177 & n1444 ;
  assign n1446 = n1445 ^ n1093 ^ 1'b0 ;
  assign n1447 = n598 ^ x86 ^ 1'b0 ;
  assign n1448 = n574 | n1236 ;
  assign n1449 = n1447 & ~n1448 ;
  assign n1450 = n958 ^ n701 ^ 1'b0 ;
  assign n1451 = ~n329 & n1241 ;
  assign n1452 = x191 & n724 ;
  assign n1453 = ~x9 & n1452 ;
  assign n1454 = n1191 & ~n1356 ;
  assign n1455 = ~n899 & n1454 ;
  assign n1456 = n401 | n934 ;
  assign n1457 = n841 | n1456 ;
  assign n1458 = n936 ^ n635 ^ 1'b0 ;
  assign n1459 = n1457 & ~n1458 ;
  assign n1460 = ~n1405 & n1459 ;
  assign n1461 = n1460 ^ n1288 ^ 1'b0 ;
  assign n1462 = n556 | n1028 ;
  assign n1463 = x254 | n1462 ;
  assign n1464 = n1463 ^ n1027 ^ 1'b0 ;
  assign n1466 = n858 | n1174 ;
  assign n1467 = n1305 & ~n1466 ;
  assign n1465 = n771 & n1114 ;
  assign n1468 = n1467 ^ n1465 ^ 1'b0 ;
  assign n1469 = n603 | n901 ;
  assign n1470 = n1469 ^ n351 ^ 1'b0 ;
  assign n1471 = n454 & ~n1470 ;
  assign n1472 = n983 & n1471 ;
  assign n1473 = n298 | n384 ;
  assign n1474 = n836 ^ x232 ^ x226 ;
  assign n1475 = n1474 ^ n1249 ^ x134 ;
  assign n1476 = n1016 | n1472 ;
  assign n1477 = n1476 ^ n409 ^ 1'b0 ;
  assign n1478 = n538 | n1269 ;
  assign n1479 = n1478 ^ x30 ^ 1'b0 ;
  assign n1480 = ~n728 & n1318 ;
  assign n1482 = x151 ^ x77 ^ 1'b0 ;
  assign n1483 = x180 & n1482 ;
  assign n1484 = n1483 ^ n545 ^ 1'b0 ;
  assign n1485 = n841 & ~n1484 ;
  assign n1481 = n904 ^ x196 ^ 1'b0 ;
  assign n1486 = n1485 ^ n1481 ^ 1'b0 ;
  assign n1487 = n361 & ~n1486 ;
  assign n1488 = n331 | n1324 ;
  assign n1489 = n1361 ^ n625 ^ 1'b0 ;
  assign n1490 = n1374 ^ n1025 ^ 1'b0 ;
  assign n1491 = x46 & n385 ;
  assign n1492 = n1491 ^ n478 ^ 1'b0 ;
  assign n1493 = n789 | n1391 ;
  assign n1494 = n1493 ^ x147 ^ 1'b0 ;
  assign n1495 = ~x20 & n1494 ;
  assign n1496 = n728 & ~n1339 ;
  assign n1497 = n1339 ^ n608 ^ 1'b0 ;
  assign n1498 = n420 & ~n768 ;
  assign n1499 = n1498 ^ n620 ^ 1'b0 ;
  assign n1500 = n1499 ^ n488 ^ 1'b0 ;
  assign n1501 = ~n1497 & n1500 ;
  assign n1502 = ~n709 & n1501 ;
  assign n1503 = n1387 & n1502 ;
  assign n1504 = x172 & x237 ;
  assign n1505 = ~n540 & n1504 ;
  assign n1506 = n269 | n361 ;
  assign n1507 = ( ~n983 & n1505 ) | ( ~n983 & n1506 ) | ( n1505 & n1506 ) ;
  assign n1508 = n1195 & n1507 ;
  assign n1509 = x240 & n1409 ;
  assign n1510 = ~x73 & n1509 ;
  assign n1511 = n825 | n1510 ;
  assign n1513 = n478 & ~n659 ;
  assign n1512 = n880 ^ n848 ^ n490 ;
  assign n1514 = n1513 ^ n1512 ^ x222 ;
  assign n1515 = ~n366 & n964 ;
  assign n1516 = x166 & ~n384 ;
  assign n1517 = ~n445 & n1516 ;
  assign n1518 = n939 & ~n1517 ;
  assign n1520 = n1447 ^ n1064 ^ 1'b0 ;
  assign n1521 = x249 & n1520 ;
  assign n1519 = x98 & n1195 ;
  assign n1522 = n1521 ^ n1519 ^ 1'b0 ;
  assign n1523 = x33 & ~n485 ;
  assign n1524 = n1523 ^ x203 ^ 1'b0 ;
  assign n1525 = ( x97 & n1007 ) | ( x97 & ~n1239 ) | ( n1007 & ~n1239 ) ;
  assign n1526 = x231 & ~n669 ;
  assign n1527 = ~n915 & n1526 ;
  assign n1528 = x105 ^ x86 ^ 1'b0 ;
  assign n1529 = n1528 ^ n594 ^ n476 ;
  assign n1530 = x58 & ~n840 ;
  assign n1531 = n766 & n1530 ;
  assign n1532 = x34 & ~n1531 ;
  assign n1533 = n1227 & n1532 ;
  assign n1534 = n607 & ~n805 ;
  assign n1535 = ~n540 & n1534 ;
  assign n1536 = n278 ^ x207 ^ 1'b0 ;
  assign n1537 = n1100 | n1536 ;
  assign n1538 = x188 & ~n1537 ;
  assign n1539 = ( ~x58 & x151 ) | ( ~x58 & n502 ) | ( x151 & n502 ) ;
  assign n1540 = x121 & n1539 ;
  assign n1543 = n789 ^ x151 ^ 1'b0 ;
  assign n1544 = x163 & ~n1543 ;
  assign n1545 = n791 & n1544 ;
  assign n1546 = n1545 ^ n621 ^ 1'b0 ;
  assign n1547 = n337 & ~n1546 ;
  assign n1548 = n1182 & n1547 ;
  assign n1541 = x180 | n1031 ;
  assign n1542 = ~n1172 & n1541 ;
  assign n1549 = n1548 ^ n1542 ^ 1'b0 ;
  assign n1550 = n778 ^ x34 ^ 1'b0 ;
  assign n1551 = ~n363 & n1550 ;
  assign n1552 = ~n1522 & n1551 ;
  assign n1553 = ~x159 & n1552 ;
  assign n1554 = x144 & x178 ;
  assign n1555 = n825 & n1554 ;
  assign n1556 = n1555 ^ n1224 ^ 1'b0 ;
  assign n1557 = n698 | n1348 ;
  assign n1558 = ~n556 & n568 ;
  assign n1559 = n1558 ^ x213 ^ 1'b0 ;
  assign n1560 = n718 ^ x57 ^ 1'b0 ;
  assign n1561 = n1139 & ~n1440 ;
  assign n1562 = ~x24 & n1561 ;
  assign n1563 = n1356 | n1562 ;
  assign n1564 = n1563 ^ n1135 ^ 1'b0 ;
  assign n1565 = x164 ^ x128 ^ 1'b0 ;
  assign n1566 = ~n981 & n1565 ;
  assign n1567 = ~n736 & n1566 ;
  assign n1568 = ~x106 & n1567 ;
  assign n1569 = n728 | n1568 ;
  assign n1570 = n349 ^ x177 ^ 1'b0 ;
  assign n1571 = n1570 ^ n836 ^ 1'b0 ;
  assign n1572 = n681 & ~n1571 ;
  assign n1573 = n1052 ^ n815 ^ 1'b0 ;
  assign n1574 = n1573 ^ n286 ^ 1'b0 ;
  assign n1575 = n734 | n1574 ;
  assign n1576 = ~n1572 & n1575 ;
  assign n1577 = n924 ^ n302 ^ 1'b0 ;
  assign n1578 = ~n1399 & n1577 ;
  assign n1579 = ( ~n577 & n1472 ) | ( ~n577 & n1578 ) | ( n1472 & n1578 ) ;
  assign n1580 = n1450 ^ n411 ^ 1'b0 ;
  assign n1585 = n323 | n341 ;
  assign n1586 = n341 & ~n1585 ;
  assign n1581 = x143 & x164 ;
  assign n1582 = ~x143 & n1581 ;
  assign n1583 = n337 & ~n1582 ;
  assign n1584 = n1582 & n1583 ;
  assign n1587 = n1586 ^ n1584 ^ 1'b0 ;
  assign n1588 = n448 ^ n360 ^ 1'b0 ;
  assign n1589 = n461 & ~n1000 ;
  assign n1590 = x114 & ~n1116 ;
  assign n1591 = ~n463 & n1590 ;
  assign n1592 = n844 ^ n761 ^ 1'b0 ;
  assign n1593 = n1139 & ~n1592 ;
  assign n1594 = n434 ^ x75 ^ 1'b0 ;
  assign n1600 = n795 ^ x28 ^ 1'b0 ;
  assign n1598 = x185 & n891 ;
  assign n1599 = n830 & n1598 ;
  assign n1595 = x248 ^ x48 ^ 1'b0 ;
  assign n1596 = n607 & n1595 ;
  assign n1597 = n1596 ^ n323 ^ 1'b0 ;
  assign n1601 = n1600 ^ n1599 ^ n1597 ;
  assign n1602 = n1601 ^ x191 ^ 1'b0 ;
  assign n1603 = n1249 ^ n918 ^ 1'b0 ;
  assign n1604 = n1602 & n1603 ;
  assign n1605 = ~x239 & n1604 ;
  assign n1606 = n854 ^ n556 ^ 1'b0 ;
  assign n1607 = n1029 & n1325 ;
  assign n1608 = ~n776 & n1607 ;
  assign n1609 = n1608 ^ n859 ^ 1'b0 ;
  assign n1610 = n1606 | n1609 ;
  assign n1611 = n860 ^ n637 ^ 1'b0 ;
  assign n1612 = x101 & n365 ;
  assign n1613 = ~n1226 & n1612 ;
  assign n1614 = n700 | n789 ;
  assign n1615 = n1010 ^ n629 ^ 1'b0 ;
  assign n1616 = ~n683 & n1615 ;
  assign n1617 = n1616 ^ n957 ^ 1'b0 ;
  assign n1618 = ~n1423 & n1617 ;
  assign n1619 = n1223 ^ n259 ^ 1'b0 ;
  assign n1620 = n1594 ^ n621 ^ 1'b0 ;
  assign n1621 = n772 & n1214 ;
  assign n1622 = n1002 ^ n858 ^ 1'b0 ;
  assign n1623 = n705 ^ x254 ^ 1'b0 ;
  assign n1624 = n1223 ^ n638 ^ 1'b0 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = n1622 | n1625 ;
  assign n1627 = x246 & ~n521 ;
  assign n1628 = n1627 ^ n594 ^ 1'b0 ;
  assign n1629 = ~n574 & n1628 ;
  assign n1630 = n1182 | n1629 ;
  assign n1631 = ~n323 & n926 ;
  assign n1632 = n931 & n1631 ;
  assign n1633 = x18 | n1632 ;
  assign n1634 = ( x12 & x144 ) | ( x12 & n1633 ) | ( x144 & n1633 ) ;
  assign n1635 = ~n1310 & n1634 ;
  assign n1636 = n949 ^ n930 ^ 1'b0 ;
  assign n1637 = n1438 & ~n1636 ;
  assign n1638 = n294 ^ x149 ^ 1'b0 ;
  assign n1639 = x75 & n1638 ;
  assign n1640 = n432 ^ x132 ^ 1'b0 ;
  assign n1641 = n1541 & ~n1640 ;
  assign n1642 = ( x140 & n1201 ) | ( x140 & ~n1641 ) | ( n1201 & ~n1641 ) ;
  assign n1643 = x143 & ~n637 ;
  assign n1644 = ~n1228 & n1643 ;
  assign n1645 = n1638 ^ n542 ^ 1'b0 ;
  assign n1646 = n1644 | n1645 ;
  assign n1647 = n1646 ^ n1128 ^ 1'b0 ;
  assign n1648 = n1642 & n1647 ;
  assign n1649 = ~n526 & n1360 ;
  assign n1650 = n1649 ^ n1018 ^ 1'b0 ;
  assign n1651 = n1299 ^ n1236 ^ 1'b0 ;
  assign n1652 = x205 & n707 ;
  assign n1653 = n1652 ^ x154 ^ 1'b0 ;
  assign n1654 = ~n341 & n1653 ;
  assign n1656 = n1082 | n1269 ;
  assign n1655 = x160 & n1378 ;
  assign n1657 = n1656 ^ n1655 ^ 1'b0 ;
  assign n1658 = n950 ^ n807 ^ 1'b0 ;
  assign n1659 = n1158 & n1237 ;
  assign n1660 = ~n787 & n1659 ;
  assign n1661 = n561 & n1660 ;
  assign n1662 = ~n1623 & n1661 ;
  assign n1663 = n1662 ^ n476 ^ 1'b0 ;
  assign n1665 = n1629 ^ x43 ^ 1'b0 ;
  assign n1666 = ~n1152 & n1665 ;
  assign n1667 = n1666 ^ n987 ^ 1'b0 ;
  assign n1664 = ~n722 & n1389 ;
  assign n1668 = n1667 ^ n1664 ^ 1'b0 ;
  assign n1669 = n493 | n637 ;
  assign n1670 = n288 | n1669 ;
  assign n1671 = ~n951 & n1670 ;
  assign n1672 = n1633 ^ n543 ^ 1'b0 ;
  assign n1673 = n1004 & n1159 ;
  assign n1674 = n1175 ^ n1130 ^ 1'b0 ;
  assign n1675 = ~n352 & n1674 ;
  assign n1676 = n821 | n1339 ;
  assign n1677 = n1676 ^ n432 ^ 1'b0 ;
  assign n1678 = n927 & ~n1677 ;
  assign n1679 = ~n388 & n1205 ;
  assign n1680 = n1679 ^ x198 ^ 1'b0 ;
  assign n1681 = x141 & ~x209 ;
  assign n1682 = n760 & ~n1681 ;
  assign n1683 = n1682 ^ n1271 ^ 1'b0 ;
  assign n1684 = x170 & n1683 ;
  assign n1685 = x63 & ~n1684 ;
  assign n1686 = ( n614 & n1100 ) | ( n614 & ~n1347 ) | ( n1100 & ~n1347 ) ;
  assign n1687 = x180 & ~n1314 ;
  assign n1688 = n1687 ^ n671 ^ 1'b0 ;
  assign n1689 = n595 | n977 ;
  assign n1690 = n1611 ^ n518 ^ 1'b0 ;
  assign n1691 = n743 ^ n733 ^ 1'b0 ;
  assign n1692 = ~n669 & n1691 ;
  assign n1693 = n692 & n1692 ;
  assign n1694 = n452 ^ n446 ^ n405 ;
  assign n1695 = ~n1172 & n1694 ;
  assign n1696 = n846 & n1695 ;
  assign n1697 = n911 & ~n1029 ;
  assign n1698 = n1694 & n1697 ;
  assign n1699 = n279 | n573 ;
  assign n1700 = n409 | n1699 ;
  assign n1701 = x66 & ~n859 ;
  assign n1702 = n1700 & n1701 ;
  assign n1703 = ~n1525 & n1702 ;
  assign n1704 = x20 | n432 ;
  assign n1705 = n1190 | n1704 ;
  assign n1706 = n671 & ~n1705 ;
  assign n1707 = n1706 ^ n1487 ^ 1'b0 ;
  assign n1712 = x29 & n277 ;
  assign n1713 = n1712 ^ n907 ^ 1'b0 ;
  assign n1708 = x252 & ~n1243 ;
  assign n1709 = n1708 ^ n305 ^ 1'b0 ;
  assign n1710 = x37 & n1709 ;
  assign n1711 = n1611 | n1710 ;
  assign n1714 = n1713 ^ n1711 ^ 1'b0 ;
  assign n1715 = x223 & n1549 ;
  assign n1716 = x31 & n1256 ;
  assign n1717 = ~x87 & n1716 ;
  assign n1718 = n620 | n1717 ;
  assign n1719 = n1174 ^ n1016 ^ 1'b0 ;
  assign n1720 = ~n1503 & n1719 ;
  assign n1722 = x169 & ~n715 ;
  assign n1723 = n651 & n1722 ;
  assign n1721 = x61 & ~n374 ;
  assign n1724 = n1723 ^ n1721 ^ 1'b0 ;
  assign n1725 = n1724 ^ n1313 ^ 1'b0 ;
  assign n1726 = n899 & ~n1272 ;
  assign n1727 = ~n1054 & n1726 ;
  assign n1728 = ( ~x244 & n907 ) | ( ~x244 & n1539 ) | ( n907 & n1539 ) ;
  assign n1729 = n1718 & ~n1728 ;
  assign n1730 = x212 & ~n381 ;
  assign n1731 = n1730 ^ n548 ^ 1'b0 ;
  assign n1732 = ~n607 & n791 ;
  assign n1733 = n403 & ~n1243 ;
  assign n1734 = n1269 | n1733 ;
  assign n1735 = n1734 ^ n776 ^ 1'b0 ;
  assign n1736 = n1358 ^ n1192 ^ 1'b0 ;
  assign n1737 = n430 | n635 ;
  assign n1738 = n941 | n1737 ;
  assign n1739 = n987 ^ n354 ^ 1'b0 ;
  assign n1740 = n1739 ^ n543 ^ 1'b0 ;
  assign n1741 = ~n835 & n1740 ;
  assign n1742 = x173 | n774 ;
  assign n1743 = n503 & n1742 ;
  assign n1744 = ~x128 & n502 ;
  assign n1745 = n1258 ^ n926 ^ x140 ;
  assign n1746 = n1378 ^ x137 ^ x55 ;
  assign n1747 = n420 & ~n1461 ;
  assign n1748 = n1065 ^ x22 ^ 1'b0 ;
  assign n1749 = ~n828 & n1748 ;
  assign n1756 = n277 & n841 ;
  assign n1757 = n1756 ^ n968 ^ 1'b0 ;
  assign n1750 = n510 & ~n963 ;
  assign n1751 = n637 & n1750 ;
  assign n1752 = n1212 | n1751 ;
  assign n1753 = n1752 ^ n1660 ^ 1'b0 ;
  assign n1754 = ~n296 & n1753 ;
  assign n1755 = n1644 | n1754 ;
  assign n1758 = n1757 ^ n1755 ^ 1'b0 ;
  assign n1759 = n638 ^ x151 ^ 1'b0 ;
  assign n1760 = ~n994 & n1759 ;
  assign n1761 = n1760 ^ x5 ^ 1'b0 ;
  assign n1762 = n1761 ^ n1182 ^ 1'b0 ;
  assign n1763 = x158 & n867 ;
  assign n1764 = n1763 ^ n1651 ^ 1'b0 ;
  assign n1765 = n747 ^ x26 ^ 1'b0 ;
  assign n1766 = n1765 ^ n1376 ^ 1'b0 ;
  assign n1767 = x194 | n551 ;
  assign n1768 = n1767 ^ n1369 ^ 1'b0 ;
  assign n1769 = n956 | n1768 ;
  assign n1770 = x189 & n1769 ;
  assign n1771 = n548 | n1405 ;
  assign n1772 = n1771 ^ n381 ^ 1'b0 ;
  assign n1773 = n1237 ^ n871 ^ 1'b0 ;
  assign n1776 = n562 & ~n607 ;
  assign n1777 = n1776 ^ n913 ^ 1'b0 ;
  assign n1774 = n718 | n1017 ;
  assign n1775 = n1139 | n1774 ;
  assign n1778 = n1777 ^ n1775 ^ 1'b0 ;
  assign n1779 = n1773 & ~n1778 ;
  assign n1780 = n1000 ^ n302 ^ 1'b0 ;
  assign n1781 = n1368 & n1780 ;
  assign n1782 = ~n1411 & n1781 ;
  assign n1783 = n780 & n942 ;
  assign n1786 = ~x135 & x248 ;
  assign n1787 = n1173 & n1786 ;
  assign n1784 = n688 & ~n954 ;
  assign n1785 = ~x108 & n1784 ;
  assign n1788 = n1787 ^ n1785 ^ 1'b0 ;
  assign n1789 = n598 | n740 ;
  assign n1790 = n1789 ^ n815 ^ 1'b0 ;
  assign n1791 = n345 & ~n1790 ;
  assign n1792 = ~n597 & n886 ;
  assign n1793 = n420 & ~n1501 ;
  assign n1794 = n605 ^ n486 ^ 1'b0 ;
  assign n1795 = x232 & n1794 ;
  assign n1796 = x32 & n1795 ;
  assign n1797 = n1796 ^ n1205 ^ 1'b0 ;
  assign n1798 = x51 & n927 ;
  assign n1799 = n1798 ^ x17 ^ 1'b0 ;
  assign n1800 = n698 | n1027 ;
  assign n1801 = n1799 & ~n1800 ;
  assign n1802 = n388 ^ x248 ^ 1'b0 ;
  assign n1803 = n1802 ^ n1788 ^ 1'b0 ;
  assign n1804 = n1134 & ~n1393 ;
  assign n1805 = ~n415 & n1804 ;
  assign n1806 = ~n1332 & n1562 ;
  assign n1807 = n1302 & n1806 ;
  assign n1808 = n1807 ^ n1568 ^ 1'b0 ;
  assign n1809 = ~n307 & n1637 ;
  assign n1810 = n365 & ~n1103 ;
  assign n1811 = ~n673 & n1442 ;
  assign n1812 = n1811 ^ x31 ^ 1'b0 ;
  assign n1813 = n946 ^ x140 ^ 1'b0 ;
  assign n1814 = n911 & n1813 ;
  assign n1815 = n1619 | n1814 ;
  assign n1816 = x98 & ~n963 ;
  assign n1817 = n1816 ^ n1470 ^ 1'b0 ;
  assign n1818 = n1093 & n1817 ;
  assign n1819 = ~x64 & n809 ;
  assign n1820 = n894 | n1819 ;
  assign n1821 = n917 ^ n672 ^ 1'b0 ;
  assign n1822 = n1679 & n1821 ;
  assign n1823 = ~n864 & n1822 ;
  assign n1824 = n1823 ^ n859 ^ 1'b0 ;
  assign n1825 = ( n345 & n1117 ) | ( n345 & ~n1824 ) | ( n1117 & ~n1824 ) ;
  assign n1826 = n1025 & n1441 ;
  assign n1827 = ~n481 & n1826 ;
  assign n1828 = n683 & n1827 ;
  assign n1829 = n915 ^ x242 ^ 1'b0 ;
  assign n1830 = n1829 ^ x181 ^ 1'b0 ;
  assign n1831 = x213 & n1830 ;
  assign n1832 = ~n692 & n1831 ;
  assign n1833 = x157 & ~n621 ;
  assign n1834 = ~n1196 & n1833 ;
  assign n1835 = n1807 ^ n985 ^ 1'b0 ;
  assign n1836 = n797 | n1541 ;
  assign n1837 = n1438 ^ n1100 ^ 1'b0 ;
  assign n1838 = x30 & n500 ;
  assign n1839 = n1838 ^ n454 ^ 1'b0 ;
  assign n1840 = n641 & ~n1839 ;
  assign n1841 = n1282 & n1286 ;
  assign n1845 = n992 ^ x238 ^ 1'b0 ;
  assign n1842 = n608 | n628 ;
  assign n1843 = n1842 ^ n964 ^ 1'b0 ;
  assign n1844 = x246 & n1843 ;
  assign n1846 = n1845 ^ n1844 ^ 1'b0 ;
  assign n1847 = x205 ^ x84 ^ 1'b0 ;
  assign n1848 = n1847 ^ n1803 ^ 1'b0 ;
  assign n1849 = n1397 & n1848 ;
  assign n1850 = ~x59 & n1826 ;
  assign n1851 = x49 & ~n1438 ;
  assign n1852 = x184 ^ x149 ^ 1'b0 ;
  assign n1853 = ~n1851 & n1852 ;
  assign n1854 = n1047 & ~n1853 ;
  assign n1855 = n934 ^ n931 ^ n669 ;
  assign n1856 = n1855 ^ n1239 ^ n374 ;
  assign n1857 = n860 ^ x96 ^ 1'b0 ;
  assign n1858 = x93 | n1857 ;
  assign n1859 = n1858 ^ n1016 ^ 1'b0 ;
  assign n1860 = n1376 ^ x8 ^ 1'b0 ;
  assign n1861 = n924 & n1860 ;
  assign n1862 = n709 | n1828 ;
  assign n1863 = n1862 ^ n1272 ^ 1'b0 ;
  assign n1864 = ( x132 & x177 ) | ( x132 & ~n1671 ) | ( x177 & ~n1671 ) ;
  assign n1865 = n607 ^ n325 ^ 1'b0 ;
  assign n1866 = n1864 & n1865 ;
  assign n1867 = n446 & n1638 ;
  assign n1868 = n378 ^ x217 ^ 1'b0 ;
  assign n1869 = ~n748 & n1868 ;
  assign n1870 = n409 & n1869 ;
  assign n1871 = n1870 ^ x165 ^ 1'b0 ;
  assign n1872 = n1871 ^ n275 ^ x80 ;
  assign n1873 = x232 & ~n681 ;
  assign n1874 = x73 & x97 ;
  assign n1875 = ~n1029 & n1874 ;
  assign n1876 = n1875 ^ n707 ^ 1'b0 ;
  assign n1877 = n1313 & ~n1876 ;
  assign n1878 = x131 & n1877 ;
  assign n1879 = n430 & n1878 ;
  assign n1880 = x81 & ~n1324 ;
  assign n1881 = n1444 & n1880 ;
  assign n1882 = n357 & n1881 ;
  assign n1883 = n994 ^ n318 ^ 1'b0 ;
  assign n1884 = n1883 ^ x76 ^ 1'b0 ;
  assign n1885 = ~n1882 & n1884 ;
  assign n1886 = x239 & n608 ;
  assign n1887 = n428 ^ x100 ^ 1'b0 ;
  assign n1888 = n854 & ~n1887 ;
  assign n1889 = ~n971 & n1888 ;
  assign n1890 = n1889 ^ n1626 ^ 1'b0 ;
  assign n1891 = n1890 ^ n261 ^ 1'b0 ;
  assign n1892 = n1438 & ~n1891 ;
  assign n1893 = n361 ^ x227 ^ 1'b0 ;
  assign n1894 = n1208 & n1251 ;
  assign n1895 = x245 & n318 ;
  assign n1896 = ~n730 & n1895 ;
  assign n1897 = n1896 ^ n1269 ^ 1'b0 ;
  assign n1898 = n1091 | n1632 ;
  assign n1899 = n1288 ^ n540 ^ 1'b0 ;
  assign n1900 = ( ~x147 & n975 ) | ( ~x147 & n1899 ) | ( n975 & n1899 ) ;
  assign n1901 = n707 & ~n1725 ;
  assign n1902 = n454 & ~n1288 ;
  assign n1903 = n1902 ^ x254 ^ 1'b0 ;
  assign n1904 = x124 | n1903 ;
  assign n1905 = n1224 & ~n1904 ;
  assign n1906 = x205 & ~n1905 ;
  assign n1907 = n1906 ^ n313 ^ 1'b0 ;
  assign n1908 = n1709 ^ n1016 ^ 1'b0 ;
  assign n1909 = ~n1907 & n1908 ;
  assign n1911 = x164 & n1523 ;
  assign n1912 = n1911 ^ n1288 ^ 1'b0 ;
  assign n1910 = n259 | n1056 ;
  assign n1913 = n1912 ^ n1910 ^ 1'b0 ;
  assign n1914 = n1523 & ~n1913 ;
  assign n1915 = n1442 ^ n724 ^ 1'b0 ;
  assign n1916 = ~n281 & n1915 ;
  assign n1918 = n1260 ^ n490 ^ 1'b0 ;
  assign n1919 = n1903 | n1918 ;
  assign n1920 = n1919 ^ n497 ^ 1'b0 ;
  assign n1917 = n814 ^ n493 ^ 1'b0 ;
  assign n1921 = n1920 ^ n1917 ^ 1'b0 ;
  assign n1922 = ~n1133 & n1921 ;
  assign n1923 = n307 | n380 ;
  assign n1924 = ~n290 & n1263 ;
  assign n1925 = n1924 ^ n1195 ^ 1'b0 ;
  assign n1926 = n1923 | n1925 ;
  assign n1927 = n1524 | n1926 ;
  assign n1928 = n1156 & ~n1927 ;
  assign n1929 = n528 & ~n1928 ;
  assign n1930 = n1608 ^ n761 ^ 1'b0 ;
  assign n1931 = n388 & n1666 ;
  assign n1932 = x16 | n842 ;
  assign n1934 = n874 ^ n838 ^ 1'b0 ;
  assign n1935 = x172 & ~n1934 ;
  assign n1933 = n918 & n1029 ;
  assign n1936 = n1935 ^ n1933 ^ 1'b0 ;
  assign n1937 = x75 & x235 ;
  assign n1938 = ~n503 & n1775 ;
  assign n1939 = n1551 ^ n814 ^ 1'b0 ;
  assign n1940 = n1939 ^ n445 ^ 1'b0 ;
  assign n1941 = ~n1527 & n1940 ;
  assign n1942 = x102 & ~n1006 ;
  assign n1943 = n1942 ^ n1760 ^ 1'b0 ;
  assign n1944 = n896 & n1943 ;
  assign n1945 = n512 & n924 ;
  assign n1946 = n822 & ~n1939 ;
  assign n1947 = n1946 ^ n691 ^ 1'b0 ;
  assign n1948 = ( ~n858 & n965 ) | ( ~n858 & n1333 ) | ( n965 & n1333 ) ;
  assign n1949 = n1948 ^ n1318 ^ 1'b0 ;
  assign n1950 = n1724 ^ x48 ^ 1'b0 ;
  assign n1951 = x144 | n534 ;
  assign n1952 = n1226 | n1522 ;
  assign n1953 = ( x102 & x142 ) | ( x102 & ~x191 ) | ( x142 & ~x191 ) ;
  assign n1954 = ~n840 & n1953 ;
  assign n1955 = n1954 ^ n365 ^ 1'b0 ;
  assign n1956 = n1091 & ~n1955 ;
  assign n1957 = ~n426 & n1956 ;
  assign n1958 = n1957 ^ n1075 ^ 1'b0 ;
  assign n1959 = n524 & ~n1958 ;
  assign n1963 = ~n805 & n923 ;
  assign n1964 = n1963 ^ n465 ^ 1'b0 ;
  assign n1960 = n1114 & n1869 ;
  assign n1961 = ~n1264 & n1960 ;
  assign n1962 = n1372 | n1961 ;
  assign n1965 = n1964 ^ n1962 ^ 1'b0 ;
  assign n1966 = n378 ^ n333 ^ 1'b0 ;
  assign n1967 = n318 & n1966 ;
  assign n1968 = n911 ^ x186 ^ x43 ;
  assign n1969 = n1968 ^ n715 ^ 1'b0 ;
  assign n1972 = ~x64 & x196 ;
  assign n1970 = ~n352 & n363 ;
  assign n1971 = x170 & n1970 ;
  assign n1973 = n1972 ^ n1971 ^ 1'b0 ;
  assign n1974 = x22 & n325 ;
  assign n1975 = x59 & x129 ;
  assign n1976 = n1975 ^ x152 ^ 1'b0 ;
  assign n1977 = n891 & n1976 ;
  assign n1978 = n1977 ^ n438 ^ 1'b0 ;
  assign n1979 = n1974 | n1978 ;
  assign n1980 = n467 & n909 ;
  assign n1981 = n1980 ^ x228 ^ 1'b0 ;
  assign n1982 = x18 & n1429 ;
  assign n1983 = n275 & n1982 ;
  assign n1984 = n988 ^ n798 ^ 1'b0 ;
  assign n1985 = x115 & n1984 ;
  assign n1986 = n1985 ^ n1684 ^ 1'b0 ;
  assign n1987 = n707 & ~n1986 ;
  assign n1988 = n1987 ^ n1883 ^ 1'b0 ;
  assign n1989 = x73 & ~n1928 ;
  assign n1990 = n1989 ^ n1133 ^ 1'b0 ;
  assign n1991 = n1819 ^ n1326 ^ 1'b0 ;
  assign n1992 = n1991 ^ n1399 ^ 1'b0 ;
  assign n1993 = n1760 & n1767 ;
  assign n1994 = ~n1953 & n1993 ;
  assign n1995 = n553 | n1994 ;
  assign n1996 = x75 | n1995 ;
  assign n1997 = ~n796 & n1996 ;
  assign n1998 = n1992 & n1997 ;
  assign n1999 = n1626 & n1998 ;
  assign n2000 = n1769 | n1845 ;
  assign n2001 = n2000 ^ n1099 ^ 1'b0 ;
  assign n2002 = ~n472 & n1594 ;
  assign n2003 = n2002 ^ n985 ^ 1'b0 ;
  assign n2004 = n1849 ^ x81 ^ 1'b0 ;
  assign n2005 = n932 & ~n951 ;
  assign n2006 = n2005 ^ n1854 ^ 1'b0 ;
  assign n2007 = n1243 ^ x226 ^ 1'b0 ;
  assign n2008 = n1629 & ~n2007 ;
  assign n2009 = n1002 ^ n385 ^ 1'b0 ;
  assign n2010 = n581 & ~n2009 ;
  assign n2011 = n2010 ^ n327 ^ 1'b0 ;
  assign n2012 = n2011 ^ n543 ^ 1'b0 ;
  assign n2013 = x98 ^ x90 ^ x68 ;
  assign n2014 = n1096 & n2013 ;
  assign n2015 = x251 ^ x158 ^ x15 ;
  assign n2016 = n2014 | n2015 ;
  assign n2017 = n2016 ^ n813 ^ 1'b0 ;
  assign n2018 = n2017 ^ x157 ^ x70 ;
  assign n2019 = n2018 ^ x10 ^ 1'b0 ;
  assign n2020 = n1143 ^ x84 ^ 1'b0 ;
  assign n2021 = n1068 | n2020 ;
  assign n2033 = x194 ^ x44 ^ 1'b0 ;
  assign n2034 = n1120 & n2033 ;
  assign n2022 = n1230 | n1474 ;
  assign n2023 = x190 & ~n535 ;
  assign n2024 = n2023 ^ x52 ^ 1'b0 ;
  assign n2025 = n1023 & ~n2024 ;
  assign n2026 = n2025 ^ n257 ^ 1'b0 ;
  assign n2027 = n2026 ^ x170 ^ 1'b0 ;
  assign n2028 = ~n285 & n2027 ;
  assign n2029 = n2028 ^ n911 ^ 1'b0 ;
  assign n2030 = n2022 | n2029 ;
  assign n2031 = n2030 ^ n784 ^ 1'b0 ;
  assign n2032 = n1169 | n2031 ;
  assign n2035 = n2034 ^ n2032 ^ 1'b0 ;
  assign n2036 = ~n341 & n836 ;
  assign n2037 = n2036 ^ n793 ^ 1'b0 ;
  assign n2038 = n1018 & n2037 ;
  assign n2039 = x202 ^ x64 ^ 1'b0 ;
  assign n2040 = n2039 ^ n1896 ^ 1'b0 ;
  assign n2041 = n2040 ^ n1328 ^ 1'b0 ;
  assign n2042 = n347 | n2041 ;
  assign n2043 = n2042 ^ x67 ^ 1'b0 ;
  assign n2044 = x3 & ~n2043 ;
  assign n2045 = n1459 ^ x51 ^ 1'b0 ;
  assign n2046 = ~n1320 & n2045 ;
  assign n2047 = n1599 | n1654 ;
  assign n2048 = n1194 ^ n901 ^ 1'b0 ;
  assign n2049 = ~n322 & n987 ;
  assign n2050 = n2049 ^ n994 ^ 1'b0 ;
  assign n2051 = n2050 ^ n1904 ^ 1'b0 ;
  assign n2052 = n2048 & ~n2051 ;
  assign n2053 = n2052 ^ n480 ^ 1'b0 ;
  assign n2054 = x4 & n1330 ;
  assign n2055 = ~x204 & n787 ;
  assign n2056 = n1496 ^ n1316 ^ 1'b0 ;
  assign n2057 = x233 & ~n2056 ;
  assign n2058 = ~x67 & n644 ;
  assign n2059 = n1833 ^ x187 ^ 1'b0 ;
  assign n2060 = n1810 & ~n2059 ;
  assign n2061 = n855 ^ x2 ^ 1'b0 ;
  assign n2062 = n1400 & n1770 ;
  assign n2063 = n1635 | n2062 ;
  assign n2064 = n394 & ~n1227 ;
  assign n2065 = n2064 ^ n1251 ^ 1'b0 ;
  assign n2066 = n2065 ^ n1566 ^ 1'b0 ;
  assign n2067 = n1126 | n1553 ;
  assign n2068 = n2067 ^ x173 ^ 1'b0 ;
  assign n2069 = x186 & ~n1116 ;
  assign n2070 = n863 & n2069 ;
  assign n2071 = ~n533 & n1075 ;
  assign n2072 = n930 ^ n838 ^ x138 ;
  assign n2073 = n2072 ^ n559 ^ 1'b0 ;
  assign n2074 = n1506 ^ n593 ^ n357 ;
  assign n2075 = n1146 & n2074 ;
  assign n2076 = n2075 ^ x252 ^ 1'b0 ;
  assign n2077 = n1788 ^ n1318 ^ 1'b0 ;
  assign n2078 = n1252 & n2077 ;
  assign n2079 = n1164 ^ n849 ^ 1'b0 ;
  assign n2080 = n749 | n2079 ;
  assign n2081 = x234 & ~n318 ;
  assign n2082 = n2081 ^ n1378 ^ 1'b0 ;
  assign n2083 = n1457 & n1541 ;
  assign n2084 = x159 & n595 ;
  assign n2085 = ~x4 & n2084 ;
  assign n2086 = n2085 ^ x251 ^ 1'b0 ;
  assign n2087 = n1453 | n2086 ;
  assign n2088 = ~n795 & n836 ;
  assign n2089 = n2088 ^ n733 ^ 1'b0 ;
  assign n2090 = n2089 ^ n1326 ^ 1'b0 ;
  assign n2091 = x235 & ~n2090 ;
  assign n2092 = x105 & n2091 ;
  assign n2093 = n2092 ^ n948 ^ 1'b0 ;
  assign n2094 = n2014 ^ x244 ^ 1'b0 ;
  assign n2095 = n836 & ~n2094 ;
  assign n2096 = n556 | n1183 ;
  assign n2097 = n2095 | n2096 ;
  assign n2098 = ~n546 & n2097 ;
  assign n2099 = n661 ^ x64 ^ 1'b0 ;
  assign n2100 = ( ~x160 & n292 ) | ( ~x160 & n2099 ) | ( n292 & n2099 ) ;
  assign n2101 = ~n1108 & n1654 ;
  assign n2102 = n2100 & n2101 ;
  assign n2103 = x39 & n2102 ;
  assign n2104 = n568 & n2103 ;
  assign n2105 = n2104 ^ n2097 ^ 1'b0 ;
  assign n2106 = x128 & ~n825 ;
  assign n2107 = n2106 ^ n1829 ^ 1'b0 ;
  assign n2108 = n2107 ^ n2080 ^ 1'b0 ;
  assign n2109 = ~n2105 & n2108 ;
  assign n2110 = n450 & n1071 ;
  assign n2111 = n874 | n2110 ;
  assign n2112 = n1564 | n2111 ;
  assign n2113 = ( n445 & n909 ) | ( n445 & n2112 ) | ( n909 & n2112 ) ;
  assign n2114 = n1906 ^ x232 ^ 1'b0 ;
  assign n2115 = n828 | n1819 ;
  assign n2116 = n842 ^ n585 ^ 1'b0 ;
  assign n2117 = n2079 ^ x125 ^ 1'b0 ;
  assign n2122 = n399 ^ x223 ^ 1'b0 ;
  assign n2123 = n1757 ^ x201 ^ 1'b0 ;
  assign n2124 = ~n2122 & n2123 ;
  assign n2118 = n931 ^ n671 ^ 1'b0 ;
  assign n2119 = x226 & n2118 ;
  assign n2120 = ~n1762 & n2119 ;
  assign n2121 = n1047 & ~n2120 ;
  assign n2125 = n2124 ^ n2121 ^ 1'b0 ;
  assign n2126 = x23 | n635 ;
  assign n2127 = n1997 | n2126 ;
  assign n2128 = x164 & ~n1268 ;
  assign n2129 = n2128 ^ n317 ^ 1'b0 ;
  assign n2130 = n730 ^ n500 ^ 1'b0 ;
  assign n2131 = ~n677 & n2130 ;
  assign n2132 = ~n896 & n2131 ;
  assign n2133 = n2129 & ~n2132 ;
  assign n2134 = n801 ^ n528 ^ 1'b0 ;
  assign n2135 = ~n444 & n2134 ;
  assign n2136 = n2133 & n2135 ;
  assign n2137 = x178 & ~n1449 ;
  assign n2138 = n2137 ^ n1098 ^ 1'b0 ;
  assign n2139 = x101 & ~n1232 ;
  assign n2140 = n2138 & n2139 ;
  assign n2141 = n992 | n1606 ;
  assign n2142 = n2141 ^ n633 ^ 1'b0 ;
  assign n2143 = n1634 | n2142 ;
  assign n2144 = x23 & x185 ;
  assign n2145 = n2144 ^ x116 ^ 1'b0 ;
  assign n2146 = n2145 ^ x58 ^ 1'b0 ;
  assign n2147 = n1847 & ~n2146 ;
  assign n2148 = n2147 ^ n1851 ^ 1'b0 ;
  assign n2149 = n2119 & ~n2148 ;
  assign n2150 = n1979 ^ n1832 ^ 1'b0 ;
  assign n2151 = n1285 | n1651 ;
  assign n2152 = n2151 ^ n901 ^ 1'b0 ;
  assign n2153 = x105 | n1324 ;
  assign n2154 = n766 ^ n388 ^ 1'b0 ;
  assign n2155 = n791 & n2154 ;
  assign n2156 = x138 & ~n1751 ;
  assign n2157 = ~n1029 & n2156 ;
  assign n2158 = n2157 ^ n415 ^ 1'b0 ;
  assign n2159 = n793 ^ n286 ^ x229 ;
  assign n2160 = n1262 & n2159 ;
  assign n2161 = n2160 ^ n333 ^ 1'b0 ;
  assign n2162 = n1179 ^ n683 ^ 1'b0 ;
  assign n2163 = n1566 ^ x251 ^ 1'b0 ;
  assign n2164 = x31 & n2163 ;
  assign n2165 = n681 | n2164 ;
  assign n2166 = x235 ^ x144 ^ 1'b0 ;
  assign n2167 = ~n2165 & n2166 ;
  assign n2168 = n1481 & n2167 ;
  assign n2169 = n1818 ^ n1411 ^ n390 ;
  assign n2171 = x92 & n1411 ;
  assign n2172 = n2171 ^ x219 ^ 1'b0 ;
  assign n2170 = n472 | n829 ;
  assign n2173 = n2172 ^ n2170 ^ 1'b0 ;
  assign n2174 = n812 ^ x0 ^ 1'b0 ;
  assign n2175 = ~x115 & n2174 ;
  assign n2176 = n1863 ^ n734 ^ 1'b0 ;
  assign n2177 = n2175 & n2176 ;
  assign n2178 = n1247 ^ x203 ^ 1'b0 ;
  assign n2179 = n1757 & n2178 ;
  assign n2180 = n1249 & n2179 ;
  assign n2181 = n557 | n1391 ;
  assign n2182 = n1108 ^ n432 ^ 1'b0 ;
  assign n2183 = ~n1212 & n2182 ;
  assign n2184 = x186 & n2183 ;
  assign n2185 = x208 & ~n2184 ;
  assign n2186 = n729 & ~n1568 ;
  assign n2187 = n1438 ^ x77 ^ 1'b0 ;
  assign n2188 = ~n2042 & n2138 ;
  assign n2189 = n1767 ^ x68 ^ 1'b0 ;
  assign n2190 = ~n535 & n2189 ;
  assign n2191 = n1941 & ~n2190 ;
  assign n2192 = x94 & x177 ;
  assign n2193 = n2192 ^ x139 ^ 1'b0 ;
  assign n2194 = n2193 ^ n779 ^ 1'b0 ;
  assign n2195 = n1236 ^ n522 ^ 1'b0 ;
  assign n2196 = n2195 ^ n1990 ^ 1'b0 ;
  assign n2197 = n2194 & n2196 ;
  assign n2198 = x92 & ~n279 ;
  assign n2199 = n2198 ^ n613 ^ 1'b0 ;
  assign n2200 = n2199 ^ x154 ^ 1'b0 ;
  assign n2201 = x253 & n2200 ;
  assign n2202 = n2201 ^ n524 ^ 1'b0 ;
  assign n2203 = n1784 & n2202 ;
  assign n2204 = n1058 & n1134 ;
  assign n2205 = n2204 ^ n1953 ^ 1'b0 ;
  assign n2206 = n317 | n691 ;
  assign n2207 = n2205 & ~n2206 ;
  assign n2208 = ( ~x132 & n942 ) | ( ~x132 & n2207 ) | ( n942 & n2207 ) ;
  assign n2209 = n1890 & ~n2117 ;
  assign n2210 = n2209 ^ n1501 ^ 1'b0 ;
  assign n2211 = n733 ^ x81 ^ 1'b0 ;
  assign n2212 = n1098 & ~n2211 ;
  assign n2213 = n1765 ^ x247 ^ 1'b0 ;
  assign n2214 = n756 & n2213 ;
  assign n2215 = ~n710 & n2214 ;
  assign n2216 = n2212 | n2215 ;
  assign n2217 = x218 & ~n859 ;
  assign n2218 = n776 & ~n1068 ;
  assign n2219 = x4 & ~n2218 ;
  assign n2220 = n1402 ^ x173 ^ 1'b0 ;
  assign n2221 = ~n2219 & n2220 ;
  assign n2222 = n2221 ^ x242 ^ 1'b0 ;
  assign n2223 = x228 & n2222 ;
  assign n2224 = ~n1939 & n2223 ;
  assign n2225 = n425 & n2224 ;
  assign n2226 = x47 & ~n456 ;
  assign n2227 = n2226 ^ n903 ^ 1'b0 ;
  assign n2228 = n2227 ^ n1952 ^ 1'b0 ;
  assign n2229 = n1025 ^ n909 ^ 1'b0 ;
  assign n2230 = n1245 | n2229 ;
  assign n2231 = n458 & ~n2230 ;
  assign n2232 = n2228 & n2231 ;
  assign n2234 = x162 & ~n551 ;
  assign n2235 = ~n779 & n2234 ;
  assign n2236 = n378 & ~n2235 ;
  assign n2237 = n2236 ^ n2148 ^ 1'b0 ;
  assign n2238 = n278 | n2237 ;
  assign n2239 = x139 | n2238 ;
  assign n2240 = n2239 ^ n500 ^ 1'b0 ;
  assign n2241 = ~x1 & n2240 ;
  assign n2233 = x239 & ~n1039 ;
  assign n2242 = n2241 ^ n2233 ^ 1'b0 ;
  assign n2243 = n2008 | n2242 ;
  assign n2244 = ~n361 & n1221 ;
  assign n2245 = ~n954 & n2244 ;
  assign n2246 = n2245 ^ n1996 ^ 1'b0 ;
  assign n2248 = n871 & n1226 ;
  assign n2249 = x184 | n2248 ;
  assign n2247 = ~x242 & n461 ;
  assign n2250 = n2249 ^ n2247 ^ 1'b0 ;
  assign n2251 = x76 & x204 ;
  assign n2252 = n478 & n2251 ;
  assign n2253 = n376 | n2252 ;
  assign n2254 = n1160 & ~n2253 ;
  assign n2255 = n2138 ^ n642 ^ 1'b0 ;
  assign n2256 = n2254 | n2255 ;
  assign n2257 = ( x63 & ~n2250 ) | ( x63 & n2256 ) | ( ~n2250 & n2256 ) ;
  assign n2258 = n730 & ~n2120 ;
  assign n2259 = ~n1916 & n2258 ;
  assign n2260 = n981 ^ n909 ^ 1'b0 ;
  assign n2262 = n1850 ^ n720 ^ 1'b0 ;
  assign n2263 = ~n1776 & n2262 ;
  assign n2261 = ( n1131 & n2022 ) | ( n1131 & n2148 ) | ( n2022 & n2148 ) ;
  assign n2264 = n2263 ^ n2261 ^ 1'b0 ;
  assign n2265 = x150 & n655 ;
  assign n2266 = n2265 ^ n610 ^ 1'b0 ;
  assign n2267 = n1094 | n2266 ;
  assign n2268 = n833 & n2267 ;
  assign n2269 = n2268 ^ n325 ^ 1'b0 ;
  assign n2270 = x191 ^ x13 ^ 1'b0 ;
  assign n2271 = n637 ^ x61 ^ 1'b0 ;
  assign n2272 = n888 | n2271 ;
  assign n2273 = n854 & n1202 ;
  assign n2274 = x181 & ~n1277 ;
  assign n2275 = ( n621 & n1479 ) | ( n621 & n1875 ) | ( n1479 & n1875 ) ;
  assign n2276 = n503 ^ x152 ^ x129 ;
  assign n2277 = n2276 ^ n917 ^ 1'b0 ;
  assign n2278 = x112 & n2277 ;
  assign n2279 = n2278 ^ x33 ^ 1'b0 ;
  assign n2280 = x66 & n2279 ;
  assign n2281 = n1656 & n2280 ;
  assign n2282 = x199 & n666 ;
  assign n2283 = ~n936 & n2282 ;
  assign n2284 = n1847 & ~n1863 ;
  assign n2285 = n2283 & n2284 ;
  assign n2286 = n497 ^ x87 ^ 1'b0 ;
  assign n2287 = x125 | n1957 ;
  assign n2288 = n793 & ~n1239 ;
  assign n2289 = ~n2287 & n2288 ;
  assign n2290 = n2289 ^ x39 ^ 1'b0 ;
  assign n2291 = n1668 & ~n2290 ;
  assign n2292 = n1195 & ~n2291 ;
  assign n2293 = n432 ^ n337 ^ 1'b0 ;
  assign n2294 = ~n788 & n1809 ;
  assign n2295 = n2293 & n2294 ;
  assign n2296 = n1551 | n2181 ;
  assign n2297 = n827 & ~n1563 ;
  assign n2298 = n2297 ^ n1890 ^ 1'b0 ;
  assign n2299 = n478 & ~n2298 ;
  assign n2300 = n2299 ^ n1740 ^ 1'b0 ;
  assign n2301 = n1245 | n2300 ;
  assign n2302 = n2037 ^ n921 ^ x226 ;
  assign n2303 = n1224 & ~n1414 ;
  assign n2304 = x193 & ~n710 ;
  assign n2305 = n456 | n1467 ;
  assign n2306 = x174 & n2305 ;
  assign n2307 = n1077 ^ n320 ^ 1'b0 ;
  assign n2308 = n1291 ^ n278 ^ 1'b0 ;
  assign n2309 = n542 & n2308 ;
  assign n2310 = n2309 ^ n2237 ^ 1'b0 ;
  assign n2311 = ~n1477 & n2159 ;
  assign n2314 = n1272 ^ x155 ^ 1'b0 ;
  assign n2312 = n1159 | n1261 ;
  assign n2313 = n895 & n2312 ;
  assign n2315 = n2314 ^ n2313 ^ 1'b0 ;
  assign n2318 = n1483 ^ n842 ^ 1'b0 ;
  assign n2319 = ~x245 & n1847 ;
  assign n2320 = n2319 ^ n2145 ^ n1139 ;
  assign n2321 = ~n2318 & n2320 ;
  assign n2322 = n1886 & n2321 ;
  assign n2323 = n360 | n2322 ;
  assign n2324 = n2323 ^ n1158 ^ 1'b0 ;
  assign n2316 = n307 ^ x154 ^ 1'b0 ;
  assign n2317 = n1762 & ~n2316 ;
  assign n2325 = n2324 ^ n2317 ^ 1'b0 ;
  assign n2326 = ~n623 & n2072 ;
  assign n2327 = n436 | n1343 ;
  assign n2328 = n392 | n2327 ;
  assign n2330 = n600 & ~n1009 ;
  assign n2329 = n1062 & n2148 ;
  assign n2331 = n2330 ^ n2329 ^ 1'b0 ;
  assign n2332 = x83 & ~n436 ;
  assign n2333 = ~n1972 & n2332 ;
  assign n2334 = x182 ^ x64 ^ 1'b0 ;
  assign n2335 = x222 & n1409 ;
  assign n2336 = ( n2333 & n2334 ) | ( n2333 & n2335 ) | ( n2334 & n2335 ) ;
  assign n2337 = n1112 & n2336 ;
  assign n2338 = ~n333 & n2337 ;
  assign n2339 = n2331 & ~n2338 ;
  assign n2340 = ~n2328 & n2339 ;
  assign n2341 = n296 | n430 ;
  assign n2342 = n2341 ^ n1679 ^ 1'b0 ;
  assign n2343 = n387 ^ x205 ^ 1'b0 ;
  assign n2344 = n2343 ^ n2068 ^ 1'b0 ;
  assign n2345 = n2342 & ~n2344 ;
  assign n2347 = n527 & n1262 ;
  assign n2348 = n1243 & n2347 ;
  assign n2349 = n725 ^ n510 ^ 1'b0 ;
  assign n2350 = x140 & n2349 ;
  assign n2351 = ~n2348 & n2350 ;
  assign n2346 = x237 & n1978 ;
  assign n2352 = n2351 ^ n2346 ^ 1'b0 ;
  assign n2353 = n460 | n2230 ;
  assign n2354 = n782 | n2353 ;
  assign n2355 = ~n2237 & n2354 ;
  assign n2356 = n2355 ^ n286 ^ 1'b0 ;
  assign n2357 = x102 & n1271 ;
  assign n2358 = ( x76 & n1139 ) | ( x76 & ~n2357 ) | ( n1139 & ~n2357 ) ;
  assign n2359 = n2157 ^ n436 ^ 1'b0 ;
  assign n2360 = n2145 ^ n741 ^ 1'b0 ;
  assign n2361 = n2359 & ~n2360 ;
  assign n2362 = n1976 & n2361 ;
  assign n2363 = n2358 & ~n2362 ;
  assign n2364 = n2363 ^ n1941 ^ 1'b0 ;
  assign n2365 = n691 ^ n395 ^ 1'b0 ;
  assign n2366 = n1091 & n2365 ;
  assign n2367 = x74 & ~n2318 ;
  assign n2369 = n1961 ^ x76 ^ 1'b0 ;
  assign n2370 = n1525 & n2369 ;
  assign n2368 = ( n300 & n822 ) | ( n300 & n1205 ) | ( n822 & n1205 ) ;
  assign n2371 = n2370 ^ n2368 ^ 1'b0 ;
  assign n2372 = n1942 ^ n648 ^ 1'b0 ;
  assign n2373 = x55 & n2372 ;
  assign n2374 = n1820 ^ n1228 ^ 1'b0 ;
  assign n2375 = n611 & ~n651 ;
  assign n2376 = n2375 ^ n671 ^ 1'b0 ;
  assign n2377 = n2376 ^ x156 ^ 1'b0 ;
  assign n2378 = n2048 & n2377 ;
  assign n2379 = n649 & n2103 ;
  assign n2380 = n2336 ^ n2034 ^ 1'b0 ;
  assign n2381 = ~n1606 & n2143 ;
  assign n2382 = ~x73 & n2381 ;
  assign n2383 = ~n387 & n1540 ;
  assign n2384 = n1753 & n2383 ;
  assign n2385 = ( n259 & n311 ) | ( n259 & n1237 ) | ( n311 & n1237 ) ;
  assign n2386 = n875 ^ n320 ^ 1'b0 ;
  assign n2387 = x156 ^ x92 ^ 1'b0 ;
  assign n2388 = ~n808 & n1521 ;
  assign n2389 = n2387 & n2388 ;
  assign n2390 = n2386 | n2389 ;
  assign n2391 = n2385 & ~n2390 ;
  assign n2392 = x51 | n1212 ;
  assign n2393 = n2074 ^ n559 ^ 1'b0 ;
  assign n2394 = n2393 ^ n1560 ^ x68 ;
  assign n2395 = n2392 & ~n2394 ;
  assign n2396 = n368 ^ x1 ^ 1'b0 ;
  assign n2397 = n2395 & n2396 ;
  assign n2398 = n570 & n2358 ;
  assign n2399 = ~n2336 & n2398 ;
  assign n2400 = x68 | n2399 ;
  assign n2401 = n420 & ~n548 ;
  assign n2402 = n2401 ^ n1760 ^ 1'b0 ;
  assign n2403 = n888 | n2402 ;
  assign n2404 = ( x72 & ~n948 ) | ( x72 & n2403 ) | ( ~n948 & n2403 ) ;
  assign n2405 = n556 ^ x66 ^ 1'b0 ;
  assign n2406 = n1818 & ~n2405 ;
  assign n2407 = ~n909 & n1374 ;
  assign n2408 = n2407 ^ n2047 ^ 1'b0 ;
  assign n2409 = ~n300 & n1241 ;
  assign n2414 = n655 ^ n625 ^ 1'b0 ;
  assign n2415 = n2414 ^ n698 ^ x40 ;
  assign n2416 = ~n744 & n2415 ;
  assign n2417 = n2416 ^ n1610 ^ 1'b0 ;
  assign n2410 = n1413 ^ n395 ^ 1'b0 ;
  assign n2411 = x55 & ~n2410 ;
  assign n2412 = n1228 & ~n2411 ;
  assign n2413 = n2124 & n2412 ;
  assign n2418 = n2417 ^ n2413 ^ 1'b0 ;
  assign n2419 = n2291 ^ n1510 ^ 1'b0 ;
  assign n2420 = n454 & ~n2419 ;
  assign n2421 = ( x148 & n351 ) | ( x148 & ~n521 ) | ( n351 & ~n521 ) ;
  assign n2422 = x170 & ~n1369 ;
  assign n2423 = n2422 ^ n1039 ^ 1'b0 ;
  assign n2424 = n2421 & n2423 ;
  assign n2425 = n1451 & n2424 ;
  assign n2426 = n1335 ^ n415 ^ 1'b0 ;
  assign n2427 = n700 ^ n661 ^ 1'b0 ;
  assign n2428 = n2427 ^ n1977 ^ 1'b0 ;
  assign n2429 = x62 & x95 ;
  assign n2430 = n2429 ^ x213 ^ 1'b0 ;
  assign n2431 = n370 & n2430 ;
  assign n2432 = ~n872 & n2431 ;
  assign n2433 = n2432 ^ n772 ^ 1'b0 ;
  assign n2434 = ~n1704 & n2433 ;
  assign n2435 = n2318 & n2434 ;
  assign n2436 = n685 ^ x182 ^ 1'b0 ;
  assign n2437 = n750 & n2385 ;
  assign n2438 = n814 & n2437 ;
  assign n2439 = n1126 & ~n2085 ;
  assign n2440 = ~x178 & n730 ;
  assign n2441 = n2319 ^ n729 ^ 1'b0 ;
  assign n2442 = n2441 ^ n879 ^ 1'b0 ;
  assign n2443 = n597 | n2442 ;
  assign n2444 = n2266 ^ x186 ^ 1'b0 ;
  assign n2445 = n1864 & ~n2444 ;
  assign n2446 = ~n2443 & n2445 ;
  assign n2447 = n2446 ^ n657 ^ 1'b0 ;
  assign n2450 = ~x129 & n807 ;
  assign n2448 = n1511 ^ n840 ^ 1'b0 ;
  assign n2449 = n815 | n2448 ;
  assign n2451 = n2450 ^ n2449 ^ 1'b0 ;
  assign n2452 = n2394 ^ n1820 ^ 1'b0 ;
  assign n2453 = x65 & n2452 ;
  assign n2454 = n472 & n2453 ;
  assign n2455 = ~n335 & n897 ;
  assign n2456 = n1777 | n1920 ;
  assign n2457 = n2455 & ~n2456 ;
  assign n2458 = n2057 ^ n528 ^ 1'b0 ;
  assign n2459 = n2044 & n2458 ;
  assign n2460 = x254 & n1733 ;
  assign n2461 = n401 | n2460 ;
  assign n2462 = n2461 ^ n2387 ^ 1'b0 ;
  assign n2463 = n2462 ^ x220 ^ 1'b0 ;
  assign n2464 = n1112 & n1277 ;
  assign n2465 = ( n1596 & n1677 ) | ( n1596 & n2464 ) | ( n1677 & n2464 ) ;
  assign n2466 = n452 & n867 ;
  assign n2467 = n846 ^ x31 ^ 1'b0 ;
  assign n2468 = n869 | n2467 ;
  assign n2469 = n2447 | n2468 ;
  assign n2470 = n734 ^ n425 ^ x178 ;
  assign n2471 = n728 & ~n2470 ;
  assign n2472 = n2471 ^ n1441 ^ 1'b0 ;
  assign n2473 = ~n1285 & n2472 ;
  assign n2474 = n1271 & n2473 ;
  assign n2476 = ~n557 & n1179 ;
  assign n2477 = n1237 | n2476 ;
  assign n2475 = x230 | n965 ;
  assign n2478 = n2477 ^ n2475 ^ 1'b0 ;
  assign n2479 = x146 & n2478 ;
  assign n2480 = n2479 ^ n1243 ^ 1'b0 ;
  assign n2481 = n768 ^ x126 ^ 1'b0 ;
  assign n2482 = n1258 & ~n2481 ;
  assign n2483 = n305 & n969 ;
  assign n2484 = n2483 ^ n2018 ^ 1'b0 ;
  assign n2485 = ~n1282 & n1324 ;
  assign n2486 = n2184 & ~n2485 ;
  assign n2487 = n821 ^ n713 ^ 1'b0 ;
  assign n2488 = n263 & n1831 ;
  assign n2489 = n2488 ^ n1970 ^ 1'b0 ;
  assign n2490 = n1733 | n2489 ;
  assign n2491 = n2490 ^ n1517 ^ 1'b0 ;
  assign n2492 = n1926 ^ n1360 ^ 1'b0 ;
  assign n2493 = n597 ^ n510 ^ 1'b0 ;
  assign n2494 = n828 | n2493 ;
  assign n2495 = n2494 ^ n534 ^ 1'b0 ;
  assign n2496 = n2495 ^ n1570 ^ 1'b0 ;
  assign n2497 = x244 & n1514 ;
  assign n2498 = n2497 ^ x244 ^ 1'b0 ;
  assign n2499 = x74 & ~n683 ;
  assign n2500 = n2499 ^ n2412 ^ 1'b0 ;
  assign n2501 = n2359 ^ n302 ^ 1'b0 ;
  assign n2502 = n1720 & n2501 ;
  assign n2503 = x6 & ~x100 ;
  assign n2504 = n450 ^ n395 ^ 1'b0 ;
  assign n2505 = x60 & ~n2504 ;
  assign n2506 = n2505 ^ n2024 ^ 1'b0 ;
  assign n2507 = n1020 & ~n2506 ;
  assign n2508 = n2507 ^ n815 ^ 1'b0 ;
  assign n2509 = ~n1620 & n1973 ;
  assign n2510 = n798 & n2509 ;
  assign n2511 = ~n325 & n2510 ;
  assign n2512 = n642 & n844 ;
  assign n2513 = n1145 & n2512 ;
  assign n2514 = n807 & ~n2513 ;
  assign n2515 = n2514 ^ n936 ^ 1'b0 ;
  assign n2516 = ~n1358 & n1379 ;
  assign n2517 = ~n679 & n909 ;
  assign n2518 = n1828 ^ n686 ^ 1'b0 ;
  assign n2519 = n924 & ~n2492 ;
  assign n2520 = n323 | n503 ;
  assign n2521 = x53 | n2520 ;
  assign n2522 = n1992 & n2521 ;
  assign n2523 = n637 & n2522 ;
  assign n2524 = n833 | n1694 ;
  assign n2525 = x123 & ~n2524 ;
  assign n2526 = n2525 ^ n456 ^ 1'b0 ;
  assign n2527 = x90 & ~x182 ;
  assign n2533 = n1217 & n1487 ;
  assign n2534 = n1751 & n2533 ;
  assign n2535 = x170 & n859 ;
  assign n2536 = n2535 ^ n966 ^ 1'b0 ;
  assign n2537 = ( x48 & x60 ) | ( x48 & n972 ) | ( x60 & n972 ) ;
  assign n2538 = n2537 ^ n1531 ^ 1'b0 ;
  assign n2539 = n2536 | n2538 ;
  assign n2540 = n2162 | n2539 ;
  assign n2541 = n2534 & ~n2540 ;
  assign n2528 = n872 ^ n281 ^ 1'b0 ;
  assign n2529 = n2528 ^ n415 ^ 1'b0 ;
  assign n2530 = n352 | n2529 ;
  assign n2531 = n1252 | n2530 ;
  assign n2532 = x50 & n2531 ;
  assign n2542 = n2541 ^ n2532 ^ 1'b0 ;
  assign n2543 = n1754 ^ n509 ^ 1'b0 ;
  assign n2544 = n1718 & ~n2543 ;
  assign n2545 = x151 & ~n296 ;
  assign n2546 = ~x22 & n2545 ;
  assign n2547 = n2546 ^ n1204 ^ 1'b0 ;
  assign n2548 = n688 ^ n385 ^ 1'b0 ;
  assign n2549 = n2548 ^ n1596 ^ 1'b0 ;
  assign n2550 = n1559 ^ n1490 ^ n304 ;
  assign n2552 = ~n535 & n782 ;
  assign n2553 = ~n1020 & n2552 ;
  assign n2551 = n1328 & ~n1980 ;
  assign n2554 = n2553 ^ n2551 ^ 1'b0 ;
  assign n2555 = x8 & ~n2227 ;
  assign n2556 = n1272 ^ n529 ^ 1'b0 ;
  assign n2557 = ~n2555 & n2556 ;
  assign n2558 = n2132 ^ x195 ^ 1'b0 ;
  assign n2559 = n1361 ^ x149 ^ 1'b0 ;
  assign n2560 = n2558 & ~n2559 ;
  assign n2561 = ~n2557 & n2560 ;
  assign n2562 = n1829 ^ n1297 ^ 1'b0 ;
  assign n2563 = n818 & n1358 ;
  assign n2564 = n2563 ^ n1667 ^ 1'b0 ;
  assign n2565 = n625 ^ n418 ^ 1'b0 ;
  assign n2566 = n2565 ^ n426 ^ x64 ;
  assign n2567 = n669 | n2566 ;
  assign n2568 = n685 & ~n2567 ;
  assign n2574 = n738 ^ x226 ^ 1'b0 ;
  assign n2575 = n1970 & n2574 ;
  assign n2576 = n2575 ^ n1472 ^ 1'b0 ;
  assign n2569 = n828 ^ x97 ^ 1'b0 ;
  assign n2570 = ~n529 & n2569 ;
  assign n2571 = n637 & n2570 ;
  assign n2572 = n425 & ~n2571 ;
  assign n2573 = ~n672 & n2572 ;
  assign n2577 = n2576 ^ n2573 ^ 1'b0 ;
  assign n2578 = n2493 | n2577 ;
  assign n2579 = x240 & n884 ;
  assign n2580 = ~n1133 & n1492 ;
  assign n2581 = ~n2579 & n2580 ;
  assign n2582 = n1304 & ~n2581 ;
  assign n2583 = n2342 & n2582 ;
  assign n2584 = n2578 & n2583 ;
  assign n2585 = n2584 ^ n1492 ^ 1'b0 ;
  assign n2586 = x176 & ~n1286 ;
  assign n2587 = ( x154 & n444 ) | ( x154 & n806 ) | ( n444 & n806 ) ;
  assign n2591 = n401 & n550 ;
  assign n2589 = n669 ^ n273 ^ 1'b0 ;
  assign n2588 = n1167 & ~n2239 ;
  assign n2590 = n2589 ^ n2588 ^ 1'b0 ;
  assign n2592 = n2591 ^ n2590 ^ 1'b0 ;
  assign n2593 = x240 & ~n2592 ;
  assign n2595 = x59 & n644 ;
  assign n2596 = ~n298 & n2595 ;
  assign n2597 = n2596 ^ n1824 ^ n747 ;
  assign n2598 = ~n1588 & n1920 ;
  assign n2599 = ~n2597 & n2598 ;
  assign n2594 = x208 & n1446 ;
  assign n2600 = n2599 ^ n2594 ^ 1'b0 ;
  assign n2601 = n1710 ^ x199 ^ 1'b0 ;
  assign n2602 = n2600 & ~n2601 ;
  assign n2603 = ~n518 & n1268 ;
  assign n2604 = n2603 ^ n1633 ^ 1'b0 ;
  assign n2605 = n2604 ^ x222 ^ 1'b0 ;
  assign n2606 = n343 & n2605 ;
  assign n2607 = n2606 ^ n1096 ^ 1'b0 ;
  assign n2608 = x181 & ~n1266 ;
  assign n2609 = n764 & n2608 ;
  assign n2610 = n1697 ^ n1616 ^ 1'b0 ;
  assign n2611 = n2474 ^ n1068 ^ 1'b0 ;
  assign n2612 = n1102 ^ n490 ^ 1'b0 ;
  assign n2613 = x48 & ~n2612 ;
  assign n2614 = n2613 ^ x104 ^ 1'b0 ;
  assign n2615 = x33 & n2614 ;
  assign n2616 = n1299 & ~n2615 ;
  assign n2617 = n1383 & ~n1703 ;
  assign n2618 = n2617 ^ n2015 ^ 1'b0 ;
  assign n2619 = n354 & n1541 ;
  assign n2620 = n2619 ^ n2116 ^ 1'b0 ;
  assign n2621 = x178 & n302 ;
  assign n2622 = n2621 ^ x84 ^ 1'b0 ;
  assign n2623 = ~n1124 & n2622 ;
  assign n2624 = ~n2457 & n2623 ;
  assign n2625 = n1578 ^ n368 ^ 1'b0 ;
  assign n2626 = n1304 | n2625 ;
  assign n2627 = n643 & n2626 ;
  assign n2628 = n1882 ^ n1769 ^ 1'b0 ;
  assign n2629 = x111 & n2628 ;
  assign n2630 = n526 & n1944 ;
  assign n2632 = n345 ^ x80 ^ 1'b0 ;
  assign n2633 = n2632 ^ n2569 ^ 1'b0 ;
  assign n2631 = n844 & ~n2003 ;
  assign n2634 = n2633 ^ n2631 ^ 1'b0 ;
  assign n2635 = x231 & n2397 ;
  assign n2636 = n2485 & n2635 ;
  assign n2637 = n720 & ~n1614 ;
  assign n2638 = n1062 ^ x184 ^ 1'b0 ;
  assign n2639 = ~n623 & n2638 ;
  assign n2640 = n749 ^ x30 ^ 1'b0 ;
  assign n2641 = n519 & ~n1729 ;
  assign n2642 = n2641 ^ n800 ^ 1'b0 ;
  assign n2643 = n307 | n2098 ;
  assign n2644 = n1957 | n2643 ;
  assign n2645 = ~n772 & n797 ;
  assign n2646 = ~n959 & n2645 ;
  assign n2647 = n2646 ^ x218 ^ 1'b0 ;
  assign n2648 = n729 & n1544 ;
  assign n2649 = x220 & n818 ;
  assign n2650 = ~n2648 & n2649 ;
  assign n2651 = n539 ^ x20 ^ 1'b0 ;
  assign n2652 = x109 & n2651 ;
  assign n2653 = ~x191 & n2652 ;
  assign n2654 = x167 & n1784 ;
  assign n2655 = n729 & n2654 ;
  assign n2656 = x141 & ~n2655 ;
  assign n2657 = ~n1570 & n2656 ;
  assign n2658 = n1667 ^ n1183 ^ 1'b0 ;
  assign n2659 = n1833 ^ n1481 ^ 1'b0 ;
  assign n2660 = n1035 & n2659 ;
  assign n2661 = ~n2658 & n2660 ;
  assign n2662 = x40 & n1920 ;
  assign n2663 = n2661 & n2662 ;
  assign n2664 = x179 | n2663 ;
  assign n2665 = ~n2657 & n2664 ;
  assign n2666 = n2637 ^ n1724 ^ 1'b0 ;
  assign n2667 = x131 & ~n2666 ;
  assign n2668 = n754 & n1835 ;
  assign n2669 = n1854 & n2668 ;
  assign n2670 = n2131 ^ n1866 ^ x124 ;
  assign n2671 = n583 & ~n2670 ;
  assign n2672 = ~n723 & n1352 ;
  assign n2673 = n1797 & ~n2672 ;
  assign n2674 = ~n278 & n2673 ;
  assign n2675 = n2674 ^ n320 ^ 1'b0 ;
  assign n2676 = ~n832 & n1407 ;
  assign n2677 = n1732 ^ n1621 ^ 1'b0 ;
  assign n2680 = n1387 ^ x28 ^ 1'b0 ;
  assign n2681 = n820 & n2680 ;
  assign n2678 = n1148 & ~n2517 ;
  assign n2679 = ~n401 & n2678 ;
  assign n2682 = n2681 ^ n2679 ^ 1'b0 ;
  assign n2683 = n288 ^ x224 ^ 1'b0 ;
  assign n2684 = x134 & n2683 ;
  assign n2685 = n2684 ^ n875 ^ 1'b0 ;
  assign n2686 = n2685 ^ n2497 ^ n323 ;
  assign n2687 = n579 ^ x233 ^ 1'b0 ;
  assign n2688 = n2440 & n2687 ;
  assign n2689 = ~n1264 & n2688 ;
  assign n2690 = n345 | n1772 ;
  assign n2691 = x242 | n2690 ;
  assign n2695 = n590 & n2112 ;
  assign n2696 = n2098 & n2695 ;
  assign n2692 = n557 | n2298 ;
  assign n2693 = n994 | n2692 ;
  assign n2694 = n895 & n2693 ;
  assign n2697 = n2696 ^ n2694 ^ 1'b0 ;
  assign n2698 = n454 ^ x8 ^ 1'b0 ;
  assign n2699 = ~x70 & n833 ;
  assign n2700 = n956 & n2699 ;
  assign n2701 = ( x24 & ~n1837 ) | ( x24 & n1957 ) | ( ~n1837 & n1957 ) ;
  assign n2702 = x62 | n1485 ;
  assign n2703 = n1188 | n1747 ;
  assign n2704 = n2703 ^ n642 ^ 1'b0 ;
  assign n2705 = ~n1840 & n2704 ;
  assign n2706 = ~n1431 & n2705 ;
  assign n2707 = n1108 ^ n956 ^ 1'b0 ;
  assign n2708 = n2482 ^ x178 ^ 1'b0 ;
  assign n2709 = n2065 | n2708 ;
  assign n2710 = n343 & ~n1393 ;
  assign n2711 = n705 & n2710 ;
  assign n2712 = n2711 ^ n2376 ^ 1'b0 ;
  assign n2713 = n1926 | n2712 ;
  assign n2714 = n1158 | n2713 ;
  assign n2715 = x223 & ~n1091 ;
  assign n2716 = n666 & n963 ;
  assign n2717 = n2715 | n2716 ;
  assign n2718 = n2717 ^ n1786 ^ 1'b0 ;
  assign n2719 = x125 & n2718 ;
  assign n2720 = ~n2714 & n2719 ;
  assign n2722 = ~x231 & n1415 ;
  assign n2721 = x183 & n1979 ;
  assign n2723 = n2722 ^ n2721 ^ 1'b0 ;
  assign n2724 = ~n1143 & n2723 ;
  assign n2725 = n2724 ^ n1330 ^ 1'b0 ;
  assign n2728 = n1070 | n2081 ;
  assign n2729 = n2558 ^ n1515 ^ 1'b0 ;
  assign n2730 = n2728 & n2729 ;
  assign n2726 = n269 & n1914 ;
  assign n2727 = n2726 ^ n1252 ^ 1'b0 ;
  assign n2731 = n2730 ^ n2727 ^ x62 ;
  assign n2732 = x228 & ~n358 ;
  assign n2733 = ~x194 & n2732 ;
  assign n2734 = n2733 ^ n937 ^ 1'b0 ;
  assign n2735 = ~n1004 & n2734 ;
  assign n2736 = n1997 ^ n679 ^ 1'b0 ;
  assign n2737 = n2735 & n2736 ;
  assign n2738 = x251 & n2597 ;
  assign n2739 = n2738 ^ n1091 ^ 1'b0 ;
  assign n2740 = ( x114 & n1173 ) | ( x114 & ~n1819 ) | ( n1173 & ~n1819 ) ;
  assign n2741 = n2739 & n2740 ;
  assign n2742 = n399 & ~n2264 ;
  assign n2743 = ~n891 & n2742 ;
  assign n2744 = n1839 ^ n1468 ^ n1311 ;
  assign n2745 = n985 ^ n351 ^ 1'b0 ;
  assign n2746 = n1937 & ~n2745 ;
  assign n2748 = x24 & x80 ;
  assign n2749 = n2748 ^ x247 ^ 1'b0 ;
  assign n2747 = n2420 ^ n420 ^ 1'b0 ;
  assign n2750 = n2749 ^ n2747 ^ 1'b0 ;
  assign n2751 = n662 & ~n1126 ;
  assign n2752 = n503 & n2751 ;
  assign n2753 = n2336 & ~n2752 ;
  assign n2754 = n2753 ^ n1172 ^ 1'b0 ;
  assign n2755 = n2531 & ~n2754 ;
  assign n2759 = n374 ^ x175 ^ 1'b0 ;
  assign n2760 = n1728 | n2759 ;
  assign n2757 = n461 ^ x212 ^ 1'b0 ;
  assign n2758 = n1029 & ~n2757 ;
  assign n2761 = n2760 ^ n2758 ^ 1'b0 ;
  assign n2756 = n552 & ~n1230 ;
  assign n2762 = n2761 ^ n2756 ^ 1'b0 ;
  assign n2763 = n2762 ^ x192 ^ 1'b0 ;
  assign n2764 = ~n1221 & n2763 ;
  assign n2765 = x8 & x144 ;
  assign n2766 = n840 | n2765 ;
  assign n2767 = n613 ^ x90 ^ 1'b0 ;
  assign n2768 = n2050 & ~n2767 ;
  assign n2769 = n320 & n1714 ;
  assign n2770 = ( ~n2616 & n2768 ) | ( ~n2616 & n2769 ) | ( n2768 & n2769 ) ;
  assign n2771 = n685 | n813 ;
  assign n2772 = n1346 | n2771 ;
  assign n2773 = x29 & ~n2305 ;
  assign n2774 = ~n2772 & n2773 ;
  assign n2775 = n2328 & ~n2333 ;
  assign n2776 = n1531 & n2775 ;
  assign n2777 = n2776 ^ n2310 ^ 1'b0 ;
  assign n2778 = n2507 & ~n2777 ;
  assign n2779 = n948 & n1715 ;
  assign n2782 = n2241 ^ n1283 ^ 1'b0 ;
  assign n2783 = n2782 ^ n1529 ^ 1'b0 ;
  assign n2784 = n1506 & ~n2783 ;
  assign n2781 = ~n1068 & n1178 ;
  assign n2785 = n2784 ^ n2781 ^ 1'b0 ;
  assign n2780 = x60 & ~n1988 ;
  assign n2786 = n2785 ^ n2780 ^ 1'b0 ;
  assign n2787 = n1468 | n1572 ;
  assign n2788 = x136 & ~n1314 ;
  assign n2789 = n2788 ^ x234 ^ 1'b0 ;
  assign n2790 = ~n532 & n1062 ;
  assign n2791 = n2789 & n2790 ;
  assign n2792 = ~n1117 & n1814 ;
  assign n2793 = ~n946 & n2792 ;
  assign n2794 = n1757 ^ n1192 ^ 1'b0 ;
  assign n2795 = n2794 ^ n1494 ^ 1'b0 ;
  assign n2796 = n1654 & ~n2795 ;
  assign n2797 = n1846 & n2796 ;
  assign n2798 = n2797 ^ n2596 ^ 1'b0 ;
  assign n2799 = n1190 & ~n2590 ;
  assign n2800 = n345 & n1564 ;
  assign n2801 = ~n1442 & n2800 ;
  assign n2802 = n2159 ^ n1414 ^ 1'b0 ;
  assign n2803 = n929 | n2802 ;
  assign n2804 = ~x95 & n738 ;
  assign n2808 = n864 | n1562 ;
  assign n2809 = n2808 ^ n1102 ^ 1'b0 ;
  assign n2805 = n337 & ~n1269 ;
  assign n2806 = n2805 ^ n1663 ^ 1'b0 ;
  assign n2807 = n2806 ^ n2314 ^ 1'b0 ;
  assign n2810 = n2809 ^ n2807 ^ 1'b0 ;
  assign n2811 = n2804 | n2810 ;
  assign n2812 = x160 & ~n2811 ;
  assign n2815 = n454 ^ x44 ^ 1'b0 ;
  assign n2816 = x235 & n2815 ;
  assign n2817 = x132 & n2816 ;
  assign n2818 = n2817 ^ n421 ^ 1'b0 ;
  assign n2819 = n2575 | n2818 ;
  assign n2813 = n969 & n1195 ;
  assign n2814 = ~n2684 & n2813 ;
  assign n2820 = n2819 ^ n2814 ^ n1258 ;
  assign n2821 = n772 & n1646 ;
  assign n2822 = n2821 ^ n2352 ^ 1'b0 ;
  assign n2823 = n358 | n813 ;
  assign n2824 = x199 | n2823 ;
  assign n2825 = x52 & ~n2824 ;
  assign n2826 = ( ~n872 & n2426 ) | ( ~n872 & n2825 ) | ( n2426 & n2825 ) ;
  assign n2827 = n2814 ^ n2728 ^ n2498 ;
  assign n2828 = ~n1531 & n2437 ;
  assign n2829 = n1343 | n1499 ;
  assign n2830 = n2829 ^ n1080 ^ 1'b0 ;
  assign n2832 = n728 & n1249 ;
  assign n2833 = ~n1539 & n2832 ;
  assign n2834 = n1923 | n2833 ;
  assign n2835 = n2834 ^ n1066 ^ 1'b0 ;
  assign n2831 = x195 | n1188 ;
  assign n2836 = n2835 ^ n2831 ^ 1'b0 ;
  assign n2837 = x132 | n2731 ;
  assign n2838 = n647 & ~n1196 ;
  assign n2839 = n1977 ^ x181 ^ 1'b0 ;
  assign n2840 = x163 & ~n1348 ;
  assign n2841 = n2840 ^ n1822 ^ 1'b0 ;
  assign n2842 = n2239 ^ x29 ^ 1'b0 ;
  assign n2843 = n1120 & ~n2842 ;
  assign n2844 = ~n2008 & n2843 ;
  assign n2845 = n1977 & ~n2615 ;
  assign n2846 = x65 | n355 ;
  assign n2847 = n1974 ^ n1160 ^ 1'b0 ;
  assign n2848 = n1713 & n2847 ;
  assign n2849 = n1546 & n2848 ;
  assign n2850 = ~x160 & n2185 ;
  assign n2851 = n2850 ^ n2185 ^ n296 ;
  assign n2852 = x29 & ~x182 ;
  assign n2854 = n766 ^ n709 ^ 1'b0 ;
  assign n2853 = ~n955 & n1444 ;
  assign n2855 = n2854 ^ n2853 ^ 1'b0 ;
  assign n2856 = n2852 & n2855 ;
  assign n2857 = ~n2208 & n2856 ;
  assign n2858 = n444 | n600 ;
  assign n2859 = n1160 | n1417 ;
  assign n2860 = n2858 & ~n2859 ;
  assign n2861 = x84 & n1928 ;
  assign n2862 = n1096 & ~n2861 ;
  assign n2863 = n2860 & n2862 ;
  assign n2864 = n1272 ^ n387 ^ 1'b0 ;
  assign n2865 = x99 & ~n2864 ;
  assign n2866 = n2863 & n2865 ;
  assign n2867 = n2866 ^ n2285 ^ 1'b0 ;
  assign n2868 = n927 & ~n1333 ;
  assign n2869 = n2819 ^ n2164 ^ 1'b0 ;
  assign n2870 = n2869 ^ n594 ^ 1'b0 ;
  assign n2871 = n1271 & n1700 ;
  assign n2872 = ~x160 & n1736 ;
  assign n2873 = ~n259 & n472 ;
  assign n2874 = x169 & ~n2873 ;
  assign n2875 = n2874 ^ n796 ^ 1'b0 ;
  assign n2876 = n2117 ^ x235 ^ 1'b0 ;
  assign n2877 = n1178 & ~n2876 ;
  assign n2878 = n2877 ^ n1158 ^ 1'b0 ;
  assign n2885 = ( ~n597 & n760 ) | ( ~n597 & n1341 ) | ( n760 & n1341 ) ;
  assign n2882 = ~n347 & n420 ;
  assign n2883 = n309 & n2882 ;
  assign n2884 = n949 | n2883 ;
  assign n2886 = n2885 ^ n2884 ^ 1'b0 ;
  assign n2879 = n2842 ^ n1782 ^ 1'b0 ;
  assign n2880 = n577 | n2879 ;
  assign n2881 = n2429 | n2880 ;
  assign n2887 = n2886 ^ n2881 ^ 1'b0 ;
  assign n2888 = n470 ^ n444 ^ 1'b0 ;
  assign n2889 = n2205 | n2888 ;
  assign n2890 = n347 | n2889 ;
  assign n2891 = n1103 & ~n2400 ;
  assign n2892 = n2890 & n2891 ;
  assign n2896 = x224 ^ x10 ^ 1'b0 ;
  assign n2893 = n2110 ^ n1633 ^ n608 ;
  assign n2894 = x175 & n2893 ;
  assign n2895 = ~x237 & n2894 ;
  assign n2897 = n2896 ^ n2895 ^ 1'b0 ;
  assign n2898 = n630 & ~n1438 ;
  assign n2899 = ~n296 & n2898 ;
  assign n2900 = n2899 ^ n1339 ^ 1'b0 ;
  assign n2901 = ( x160 & n607 ) | ( x160 & n2547 ) | ( n607 & n2547 ) ;
  assign n2902 = n474 & n867 ;
  assign n2903 = x157 | n351 ;
  assign n2904 = x136 | n2903 ;
  assign n2905 = ~n307 & n2904 ;
  assign n2906 = n2905 ^ n2765 ^ 1'b0 ;
  assign n2907 = n1955 ^ n1463 ^ 1'b0 ;
  assign n2908 = n2492 & ~n2907 ;
  assign n2909 = n1251 | n1288 ;
  assign n2910 = n1085 & ~n2909 ;
  assign n2911 = n2441 ^ n1608 ^ 1'b0 ;
  assign n2912 = ~n1654 & n2273 ;
  assign n2913 = n320 & ~n585 ;
  assign n2914 = n2913 ^ x205 ^ 1'b0 ;
  assign n2915 = n1137 & ~n2914 ;
  assign n2916 = n2912 & n2915 ;
  assign n2917 = x130 & n1262 ;
  assign n2918 = n2917 ^ n1016 ^ 1'b0 ;
  assign n2919 = n1234 ^ n701 ^ 1'b0 ;
  assign n2920 = ~n1441 & n2919 ;
  assign n2921 = ~n2918 & n2920 ;
  assign n2922 = n2921 ^ n263 ^ 1'b0 ;
  assign n2928 = n1152 ^ x149 ^ 1'b0 ;
  assign n2929 = n614 & n2928 ;
  assign n2930 = n420 & ~n2929 ;
  assign n2931 = n2930 ^ n2129 ^ 1'b0 ;
  assign n2924 = n1210 ^ n985 ^ 1'b0 ;
  assign n2925 = n1765 & ~n2924 ;
  assign n2923 = n1173 & n1523 ;
  assign n2926 = n2925 ^ n2923 ^ 1'b0 ;
  assign n2927 = n1825 & ~n2926 ;
  assign n2932 = n2931 ^ n2927 ^ 1'b0 ;
  assign n2933 = n1326 ^ n595 ^ 1'b0 ;
  assign n2934 = n2057 & ~n2933 ;
  assign n2935 = n320 & n2934 ;
  assign n2936 = n2175 & n2935 ;
  assign n2937 = n1836 | n2727 ;
  assign n2938 = n2508 & ~n2937 ;
  assign n2941 = n1116 ^ x204 ^ 1'b0 ;
  assign n2939 = n2218 ^ n442 ^ 1'b0 ;
  assign n2940 = ~n2566 & n2939 ;
  assign n2942 = n2941 ^ n2940 ^ 1'b0 ;
  assign n2943 = ~n329 & n1325 ;
  assign n2944 = ~n1670 & n2943 ;
  assign n2945 = n1307 | n2205 ;
  assign n2946 = n1165 & ~n2945 ;
  assign n2947 = n869 | n1400 ;
  assign n2948 = n2947 ^ n1096 ^ 1'b0 ;
  assign n2949 = n2948 ^ n2740 ^ 1'b0 ;
  assign n2950 = n2946 | n2949 ;
  assign n2951 = n2944 & ~n2950 ;
  assign n2952 = n1232 | n1295 ;
  assign n2953 = n1111 | n2952 ;
  assign n2954 = n327 & n2953 ;
  assign n2955 = n2954 ^ n1602 ^ 1'b0 ;
  assign n2956 = ~n651 & n1050 ;
  assign n2957 = n1470 & n2956 ;
  assign n2958 = n1749 ^ x73 ^ 1'b0 ;
  assign n2959 = ~n2228 & n2958 ;
  assign n2960 = n1116 ^ x26 ^ 1'b0 ;
  assign n2961 = n1901 & ~n2960 ;
  assign n2962 = n753 & n2947 ;
  assign n2963 = n1773 & n2962 ;
  assign n2964 = ~n1846 & n2963 ;
  assign n2965 = n286 ^ x112 ^ 1'b0 ;
  assign n2966 = n281 & n2965 ;
  assign n2967 = n2966 ^ n1242 ^ 1'b0 ;
  assign n2968 = ~n832 & n2967 ;
  assign n2969 = n2106 & ~n2811 ;
  assign n2970 = n2969 ^ x89 ^ 1'b0 ;
  assign n2971 = n797 & ~n2970 ;
  assign n2972 = n2971 ^ n875 ^ 1'b0 ;
  assign n2974 = x133 & n269 ;
  assign n2975 = ~x27 & n2974 ;
  assign n2973 = ~x26 & x124 ;
  assign n2976 = n2975 ^ n2973 ^ 1'b0 ;
  assign n2977 = n732 ^ x155 ^ x0 ;
  assign n2978 = ~n859 & n2977 ;
  assign n2981 = ~n726 & n2169 ;
  assign n2982 = ~x235 & n2981 ;
  assign n2979 = n343 & n1360 ;
  assign n2980 = n2322 & n2979 ;
  assign n2983 = n2982 ^ n2980 ^ n2711 ;
  assign n2985 = n974 ^ x24 ^ 1'b0 ;
  assign n2984 = n1751 | n2769 ;
  assign n2986 = n2985 ^ n2984 ^ 1'b0 ;
  assign n2987 = ~x14 & n1888 ;
  assign n2988 = n2987 ^ n1776 ^ 1'b0 ;
  assign n2989 = ~n1680 & n2988 ;
  assign n2990 = ~n2352 & n2989 ;
  assign n2991 = n1974 & ~n2990 ;
  assign n2992 = n915 & n1424 ;
  assign n2993 = ~n2604 & n2992 ;
  assign n2994 = x226 & n710 ;
  assign n2995 = n2993 & n2994 ;
  assign n2996 = x151 & ~n663 ;
  assign n2997 = n2996 ^ x39 ^ 1'b0 ;
  assign n2998 = ( n420 & n1616 ) | ( n420 & n2997 ) | ( n1616 & n2997 ) ;
  assign n2999 = ~n2995 & n2998 ;
  assign n3000 = n2999 ^ n620 ^ 1'b0 ;
  assign n3001 = n2017 ^ n1117 ^ n325 ;
  assign n3002 = ~n1272 & n3001 ;
  assign n3003 = n3002 ^ x112 ^ 1'b0 ;
  assign n3004 = n688 & n1757 ;
  assign n3005 = ~n1313 & n3004 ;
  assign n3006 = n3005 ^ n2752 ^ n998 ;
  assign n3007 = n401 | n1298 ;
  assign n3008 = n3007 ^ x43 ^ 1'b0 ;
  assign n3009 = n3008 ^ n1399 ^ 1'b0 ;
  assign n3010 = n3009 ^ n700 ^ 1'b0 ;
  assign n3011 = ~n539 & n3010 ;
  assign n3012 = n3011 ^ n2668 ^ 1'b0 ;
  assign n3013 = n3006 | n3012 ;
  assign n3014 = n725 & n2019 ;
  assign n3015 = n2366 ^ n1802 ^ 1'b0 ;
  assign n3016 = n2491 ^ n1451 ^ 1'b0 ;
  assign n3017 = n959 ^ n456 ^ 1'b0 ;
  assign n3018 = n766 ^ x179 ^ 1'b0 ;
  assign n3019 = n1566 ^ n801 ^ 1'b0 ;
  assign n3020 = n3018 & n3019 ;
  assign n3021 = n2596 & n2687 ;
  assign n3022 = ( ~n500 & n3020 ) | ( ~n500 & n3021 ) | ( n3020 & n3021 ) ;
  assign n3023 = x226 & ~n1143 ;
  assign n3024 = n785 & n3023 ;
  assign n3025 = n3024 ^ n666 ^ 1'b0 ;
  assign n3026 = x174 & ~n3025 ;
  assign n3027 = n666 & ~n3008 ;
  assign n3028 = ~n724 & n2011 ;
  assign n3030 = n1419 ^ n292 ^ 1'b0 ;
  assign n3031 = ( n838 & n1658 ) | ( n838 & n3030 ) | ( n1658 & n3030 ) ;
  assign n3032 = n3031 ^ n2008 ^ 1'b0 ;
  assign n3029 = n1059 | n2842 ;
  assign n3033 = n3032 ^ n3029 ^ 1'b0 ;
  assign n3034 = ~n1898 & n1953 ;
  assign n3035 = n3034 ^ n2606 ^ 1'b0 ;
  assign n3036 = n1617 & n3035 ;
  assign n3037 = x81 | n1000 ;
  assign n3038 = n3037 ^ n1252 ^ 1'b0 ;
  assign n3039 = n2523 | n3038 ;
  assign n3040 = n781 & n1713 ;
  assign n3041 = n292 & n1433 ;
  assign n3042 = ~n1996 & n3041 ;
  assign n3043 = ~n374 & n1198 ;
  assign n3044 = n2106 & ~n3043 ;
  assign n3045 = n3042 & n3044 ;
  assign n3046 = ~n474 & n2639 ;
  assign n3047 = n1780 ^ x151 ^ 1'b0 ;
  assign n3048 = n1473 | n2696 ;
  assign n3049 = n3048 ^ n2228 ^ 1'b0 ;
  assign n3050 = ~n450 & n1047 ;
  assign n3051 = n323 ^ x101 ^ 1'b0 ;
  assign n3052 = n3050 | n3051 ;
  assign n3053 = n2079 ^ n1905 ^ 1'b0 ;
  assign n3054 = n3053 ^ n2668 ^ 1'b0 ;
  assign n3055 = n397 & n1696 ;
  assign n3057 = n397 & ~n1539 ;
  assign n3058 = x139 & ~n3057 ;
  assign n3059 = ~n1173 & n3058 ;
  assign n3056 = ~n1517 & n2312 ;
  assign n3060 = n3059 ^ n3056 ^ 1'b0 ;
  assign n3061 = n2581 ^ n907 ^ 1'b0 ;
  assign n3062 = ~n414 & n3061 ;
  assign n3063 = x35 & ~n521 ;
  assign n3064 = ~n3062 & n3063 ;
  assign n3065 = x182 & n1133 ;
  assign n3066 = x137 & n3065 ;
  assign n3067 = ~n595 & n3066 ;
  assign n3068 = n723 & ~n3067 ;
  assign n3069 = n1754 ^ n1426 ^ n770 ;
  assign n3070 = n358 | n557 ;
  assign n3071 = n3070 ^ n801 ^ 1'b0 ;
  assign n3072 = n3071 ^ n1050 ^ 1'b0 ;
  assign n3073 = n2314 & n3072 ;
  assign n3074 = ( x48 & n1082 ) | ( x48 & ~n1154 ) | ( n1082 & ~n1154 ) ;
  assign n3075 = n2585 ^ n320 ^ 1'b0 ;
  assign n3076 = n3074 | n3075 ;
  assign n3077 = n840 | n1170 ;
  assign n3078 = n3077 ^ n448 ^ 1'b0 ;
  assign n3079 = x17 & ~n3078 ;
  assign n3080 = n589 & n3079 ;
  assign n3081 = n508 & ~n2582 ;
  assign n3082 = n1517 ^ n1131 ^ 1'b0 ;
  assign n3085 = x28 & x231 ;
  assign n3086 = n3085 ^ n1775 ^ 1'b0 ;
  assign n3087 = n2807 ^ x199 ^ 1'b0 ;
  assign n3088 = ~n3086 & n3087 ;
  assign n3089 = n2578 | n3088 ;
  assign n3083 = n2712 ^ n923 ^ 1'b0 ;
  assign n3084 = ~n983 & n3083 ;
  assign n3090 = n3089 ^ n3084 ^ 1'b0 ;
  assign n3091 = ( n992 & ~n1407 ) | ( n992 & n1693 ) | ( ~n1407 & n1693 ) ;
  assign n3092 = n3091 ^ n2871 ^ 1'b0 ;
  assign n3093 = n1890 & ~n3092 ;
  assign n3094 = ~n1785 & n3093 ;
  assign n3095 = ~n1682 & n3094 ;
  assign n3096 = n1639 ^ n532 ^ 1'b0 ;
  assign n3097 = x31 & n3096 ;
  assign n3098 = x48 & n3097 ;
  assign n3099 = n3098 ^ n1540 ^ 1'b0 ;
  assign n3100 = ~n1988 & n3099 ;
  assign n3101 = n2179 & n2865 ;
  assign n3102 = n3101 ^ n2087 ^ 1'b0 ;
  assign n3103 = x73 & n2145 ;
  assign n3104 = n3103 ^ x14 ^ 1'b0 ;
  assign n3105 = n3102 & n3104 ;
  assign n3112 = x220 & ~n1694 ;
  assign n3106 = n611 & n666 ;
  assign n3107 = ~n257 & n3106 ;
  assign n3108 = n1684 & n1802 ;
  assign n3109 = n3108 ^ x24 ^ 1'b0 ;
  assign n3110 = n2015 | n3109 ;
  assign n3111 = n3107 & ~n3110 ;
  assign n3113 = n3112 ^ n3111 ^ 1'b0 ;
  assign n3114 = n320 | n3113 ;
  assign n3115 = n1378 & ~n1749 ;
  assign n3116 = n605 ^ n331 ^ 1'b0 ;
  assign n3117 = n616 & ~n2343 ;
  assign n3118 = n623 & n2669 ;
  assign n3119 = n2334 ^ n2093 ^ n1459 ;
  assign n3120 = ~n271 & n3119 ;
  assign n3121 = ~x22 & x89 ;
  assign n3122 = n3120 & n3121 ;
  assign n3123 = n1653 ^ n869 ^ 1'b0 ;
  assign n3124 = n3123 ^ n360 ^ 1'b0 ;
  assign n3125 = n360 | n2228 ;
  assign n3126 = n3125 ^ n1751 ^ 1'b0 ;
  assign n3127 = n2352 ^ n1419 ^ 1'b0 ;
  assign n3128 = n1506 & n3127 ;
  assign n3129 = n1143 ^ x73 ^ 1'b0 ;
  assign n3130 = n1152 | n3129 ;
  assign n3131 = n399 & ~n3130 ;
  assign n3132 = n3131 ^ x232 ^ 1'b0 ;
  assign n3133 = n1832 & n2893 ;
  assign n3134 = n556 & n3133 ;
  assign n3135 = n3132 & ~n3134 ;
  assign n3136 = n1738 & n2739 ;
  assign n3137 = x199 & n616 ;
  assign n3138 = n630 & ~n3137 ;
  assign n3139 = n781 & n3138 ;
  assign n3140 = n3139 ^ n1079 ^ 1'b0 ;
  assign n3141 = n1671 & n3140 ;
  assign n3142 = n3141 ^ n2103 ^ 1'b0 ;
  assign n3143 = n1411 ^ n460 ^ 1'b0 ;
  assign n3144 = ( n1108 & n1979 ) | ( n1108 & n3143 ) | ( n1979 & n3143 ) ;
  assign n3147 = ~n585 & n2133 ;
  assign n3148 = n3147 ^ n1996 ^ 1'b0 ;
  assign n3149 = n1028 & ~n3148 ;
  assign n3150 = n2140 & n3149 ;
  assign n3145 = n613 | n749 ;
  assign n3146 = n3145 ^ n345 ^ 1'b0 ;
  assign n3151 = n3150 ^ n3146 ^ 1'b0 ;
  assign n3152 = ~n1453 & n3151 ;
  assign n3153 = n1427 ^ x156 ^ 1'b0 ;
  assign n3154 = n1701 | n2842 ;
  assign n3157 = n1736 & n2201 ;
  assign n3158 = n1727 & n3157 ;
  assign n3155 = n2916 ^ n1173 ^ 1'b0 ;
  assign n3156 = n1758 & ~n3155 ;
  assign n3159 = n3158 ^ n3156 ^ 1'b0 ;
  assign n3160 = ~n862 & n1212 ;
  assign n3161 = n841 & ~n3160 ;
  assign n3162 = n3161 ^ n2747 ^ 1'b0 ;
  assign n3163 = n1839 ^ n1684 ^ 1'b0 ;
  assign n3164 = n566 & n3163 ;
  assign n3165 = n3164 ^ n2772 ^ 1'b0 ;
  assign n3166 = x15 & ~n1646 ;
  assign n3167 = n2953 & n3001 ;
  assign n3168 = ~n1746 & n2342 ;
  assign n3169 = n3168 ^ n1573 ^ 1'b0 ;
  assign n3170 = n380 ^ n261 ^ 1'b0 ;
  assign n3171 = ~n363 & n3170 ;
  assign n3172 = n641 | n1658 ;
  assign n3173 = n3172 ^ n2997 ^ 1'b0 ;
  assign n3174 = x68 & ~n3173 ;
  assign n3175 = n3174 ^ n2491 ^ 1'b0 ;
  assign n3176 = ~x111 & x221 ;
  assign n3177 = n1494 & n3176 ;
  assign n3178 = n710 & n3177 ;
  assign n3179 = n3178 ^ n1588 ^ 1'b0 ;
  assign n3180 = ~x92 & n3179 ;
  assign n3181 = n1877 ^ n370 ^ 1'b0 ;
  assign n3182 = n1298 ^ n1093 ^ 1'b0 ;
  assign n3183 = n644 & n2071 ;
  assign n3184 = ~n1539 & n3183 ;
  assign n3185 = n1350 ^ n614 ^ 1'b0 ;
  assign n3186 = ~n1449 & n3185 ;
  assign n3187 = n2324 ^ n1365 ^ 1'b0 ;
  assign n3188 = n3187 ^ n1613 ^ 1'b0 ;
  assign n3189 = n3186 & n3188 ;
  assign n3190 = n1383 ^ n1125 ^ 1'b0 ;
  assign n3191 = x27 & n3190 ;
  assign n3192 = n1974 & n3191 ;
  assign n3193 = n3192 ^ n1739 ^ 1'b0 ;
  assign n3194 = n1181 & ~n1683 ;
  assign n3195 = n3194 ^ n836 ^ 1'b0 ;
  assign n3196 = n1172 ^ n1093 ^ 1'b0 ;
  assign n3197 = n3195 | n3196 ;
  assign n3198 = ( ~x216 & n1803 ) | ( ~x216 & n3197 ) | ( n1803 & n3197 ) ;
  assign n3199 = n1833 | n2531 ;
  assign n3200 = n2961 ^ n705 ^ n553 ;
  assign n3202 = x135 & ~n456 ;
  assign n3203 = n3202 ^ n1845 ^ 1'b0 ;
  assign n3201 = x226 & n570 ;
  assign n3204 = n3203 ^ n3201 ^ 1'b0 ;
  assign n3205 = n1593 & ~n3204 ;
  assign n3206 = n3205 ^ n921 ^ 1'b0 ;
  assign n3207 = n1242 & n3206 ;
  assign n3208 = n2505 ^ x133 ^ 1'b0 ;
  assign n3209 = n2613 & n3208 ;
  assign n3210 = n946 & ~n3209 ;
  assign n3211 = ~n1335 & n3210 ;
  assign n3212 = n3211 ^ n1028 ^ 1'b0 ;
  assign n3213 = ~n2571 & n3212 ;
  assign n3214 = n456 & ~n758 ;
  assign n3215 = ~n2015 & n3214 ;
  assign n3216 = ~x213 & n3215 ;
  assign n3217 = ( ~n1324 & n3142 ) | ( ~n1324 & n3216 ) | ( n3142 & n3216 ) ;
  assign n3220 = n987 ^ n575 ^ 1'b0 ;
  assign n3221 = n1682 & n3220 ;
  assign n3218 = x163 & ~n1510 ;
  assign n3219 = n3218 ^ n1757 ^ 1'b0 ;
  assign n3222 = n3221 ^ n3219 ^ 1'b0 ;
  assign n3223 = n904 | n3222 ;
  assign n3224 = n2172 ^ n1985 ^ x22 ;
  assign n3225 = n805 | n3107 ;
  assign n3226 = x183 | n3225 ;
  assign n3227 = n3132 & n3226 ;
  assign n3228 = n994 & n2079 ;
  assign n3229 = n3228 ^ n725 ^ 1'b0 ;
  assign n3230 = n883 | n3229 ;
  assign n3231 = n532 & n3230 ;
  assign n3232 = ~n607 & n3231 ;
  assign n3233 = n2185 & ~n3232 ;
  assign n3234 = n983 & n3233 ;
  assign n3235 = x42 & ~n1983 ;
  assign n3236 = n2908 & ~n3235 ;
  assign n3237 = n2264 & n3236 ;
  assign n3238 = n514 ^ n434 ^ 1'b0 ;
  assign n3239 = x246 & n3238 ;
  assign n3240 = ~n337 & n3239 ;
  assign n3241 = n2723 ^ n2114 ^ 1'b0 ;
  assign n3242 = n3240 & ~n3241 ;
  assign n3243 = n283 | n3162 ;
  assign n3244 = n305 ^ x141 ^ 1'b0 ;
  assign n3245 = ~n1172 & n3244 ;
  assign n3246 = n2024 ^ n1788 ^ 1'b0 ;
  assign n3247 = x49 & ~n3246 ;
  assign n3248 = n3100 | n3247 ;
  assign n3249 = n1073 & n1618 ;
  assign n3250 = n2414 & ~n3249 ;
  assign n3255 = n649 ^ n546 ^ 1'b0 ;
  assign n3253 = n1183 ^ x201 ^ 1'b0 ;
  assign n3254 = n647 & ~n3253 ;
  assign n3256 = n3255 ^ n3254 ^ x214 ;
  assign n3251 = n2247 ^ n1600 ^ n1188 ;
  assign n3252 = ( ~n990 & n1198 ) | ( ~n990 & n3251 ) | ( n1198 & n3251 ) ;
  assign n3257 = n3256 ^ n3252 ^ 1'b0 ;
  assign n3258 = n2782 ^ n1971 ^ 1'b0 ;
  assign n3259 = ~n2257 & n2431 ;
  assign n3260 = n3259 ^ n1713 ^ 1'b0 ;
  assign n3261 = n1512 & ~n1893 ;
  assign n3262 = n3261 ^ n2089 ^ 1'b0 ;
  assign n3263 = n349 ^ x82 ^ 1'b0 ;
  assign n3264 = n333 & ~n3263 ;
  assign n3265 = ~n2715 & n3264 ;
  assign n3266 = n557 | n1704 ;
  assign n3267 = n3266 ^ n2630 ^ n2438 ;
  assign n3268 = x192 | n948 ;
  assign n3269 = n3043 ^ n300 ^ 1'b0 ;
  assign n3270 = ~x112 & n1282 ;
  assign n3271 = n700 & n3270 ;
  assign n3272 = n3269 & n3271 ;
  assign n3273 = n1012 & ~n3272 ;
  assign n3274 = n3268 & n3273 ;
  assign n3275 = n1065 | n1488 ;
  assign n3277 = n2610 ^ n1646 ^ 1'b0 ;
  assign n3276 = n2266 | n3223 ;
  assign n3278 = n3277 ^ n3276 ^ 1'b0 ;
  assign n3279 = n2040 ^ n610 ^ 1'b0 ;
  assign n3280 = x245 & ~n3279 ;
  assign n3281 = n1700 & ~n2340 ;
  assign n3282 = n3280 & n3281 ;
  assign n3283 = n3282 ^ n836 ^ 1'b0 ;
  assign n3284 = n589 ^ n559 ^ 1'b0 ;
  assign n3285 = n3284 ^ n2480 ^ 1'b0 ;
  assign n3286 = n2054 | n3285 ;
  assign n3287 = n3286 ^ n2361 ^ 1'b0 ;
  assign n3288 = n917 & n1114 ;
  assign n3291 = x195 & ~n1680 ;
  assign n3292 = n3291 ^ x6 ^ 1'b0 ;
  assign n3289 = ~n1062 & n2423 ;
  assign n3290 = ~x6 & n3289 ;
  assign n3293 = n3292 ^ n3290 ^ 1'b0 ;
  assign n3294 = n3288 & ~n3293 ;
  assign n3295 = ~x45 & n1154 ;
  assign n3296 = ~n1606 & n3295 ;
  assign n3297 = n3296 ^ n954 ^ 1'b0 ;
  assign n3298 = n855 ^ x186 ^ 1'b0 ;
  assign n3299 = n1228 ^ n956 ^ 1'b0 ;
  assign n3300 = x63 & ~n3299 ;
  assign n3301 = x60 & n3300 ;
  assign n3302 = n1563 & n3301 ;
  assign n3303 = n1694 & n3302 ;
  assign n3304 = n304 & ~n1932 ;
  assign n3305 = n3304 ^ n1449 ^ 1'b0 ;
  assign n3306 = n2668 ^ n1611 ^ 1'b0 ;
  assign n3307 = ~n1709 & n3306 ;
  assign n3308 = ~n1064 & n1474 ;
  assign n3309 = n1056 | n3308 ;
  assign n3310 = n1195 & ~n3309 ;
  assign n3311 = n1974 ^ n637 ^ 1'b0 ;
  assign n3312 = ~n758 & n3311 ;
  assign n3313 = n3312 ^ n2466 ^ n490 ;
  assign n3314 = n1164 & n2505 ;
  assign n3315 = x158 & n3314 ;
  assign n3316 = n3315 ^ n2845 ^ 1'b0 ;
  assign n3317 = n535 | n2254 ;
  assign n3318 = n3195 & ~n3317 ;
  assign n3319 = n486 & n1164 ;
  assign n3320 = n1125 & n2824 ;
  assign n3321 = n3319 & n3320 ;
  assign n3322 = n370 & ~n3314 ;
  assign n3323 = n1333 ^ n766 ^ x158 ;
  assign n3324 = n573 & ~n3323 ;
  assign n3325 = n3324 ^ n3050 ^ 1'b0 ;
  assign n3326 = n2342 & n3325 ;
  assign n3327 = n498 & n1899 ;
  assign n3328 = n3327 ^ n1537 ^ 1'b0 ;
  assign n3329 = n1160 & ~n3328 ;
  assign n3330 = n1544 | n1673 ;
  assign n3331 = n3330 ^ n329 ^ 1'b0 ;
  assign n3332 = n3331 ^ n1255 ^ 1'b0 ;
  assign n3333 = n315 ^ n296 ^ 1'b0 ;
  assign n3334 = n468 | n1749 ;
  assign n3335 = ~n438 & n3334 ;
  assign n3336 = n3335 ^ n510 ^ 1'b0 ;
  assign n3337 = x31 & n1517 ;
  assign n3338 = n2249 & ~n2566 ;
  assign n3339 = n3338 ^ x77 ^ 1'b0 ;
  assign n3340 = n1463 & n3109 ;
  assign n3341 = n3031 ^ n556 ^ 1'b0 ;
  assign n3342 = n1869 & ~n3341 ;
  assign n3343 = x28 & n3342 ;
  assign n3344 = n607 & ~n1017 ;
  assign n3345 = ~n772 & n3344 ;
  assign n3346 = n1914 | n3345 ;
  assign n3347 = n1378 & ~n2757 ;
  assign n3348 = ~x231 & n3347 ;
  assign n3349 = n3348 ^ n1637 ^ 1'b0 ;
  assign n3350 = n3349 ^ n2423 ^ 1'b0 ;
  assign n3351 = ~n733 & n3350 ;
  assign n3352 = ~n956 & n1795 ;
  assign n3353 = n3352 ^ n3082 ^ 1'b0 ;
  assign n3355 = n1399 ^ n257 ^ 1'b0 ;
  assign n3354 = n1819 & n2819 ;
  assign n3356 = n3355 ^ n3354 ^ 1'b0 ;
  assign n3357 = n1738 & ~n3137 ;
  assign n3358 = n1131 & ~n3357 ;
  assign n3359 = n2314 & n3358 ;
  assign n3360 = n2774 & n3359 ;
  assign n3361 = n779 ^ x129 ^ 1'b0 ;
  assign n3362 = n3361 ^ n2846 ^ 1'b0 ;
  assign n3364 = n570 & ~n871 ;
  assign n3363 = n562 & n2429 ;
  assign n3365 = n3364 ^ n3363 ^ 1'b0 ;
  assign n3366 = n3365 ^ n538 ^ 1'b0 ;
  assign n3367 = ~n1263 & n3366 ;
  assign n3368 = n895 ^ x149 ^ 1'b0 ;
  assign n3375 = n1037 & n1707 ;
  assign n3376 = ~n1247 & n3375 ;
  assign n3369 = n2441 ^ n1318 ^ 1'b0 ;
  assign n3370 = n1981 & ~n3369 ;
  assign n3371 = n969 & n1196 ;
  assign n3372 = n3371 ^ n917 ^ 1'b0 ;
  assign n3373 = n3370 & n3372 ;
  assign n3374 = ~x103 & n3373 ;
  assign n3377 = n3376 ^ n3374 ^ 1'b0 ;
  assign n3378 = n3368 & ~n3377 ;
  assign n3379 = n1540 & n2201 ;
  assign n3380 = ~n1560 & n2358 ;
  assign n3381 = n1093 & n3380 ;
  assign n3382 = ~x42 & n2475 ;
  assign n3383 = n3381 & n3382 ;
  assign n3384 = n2181 | n2833 ;
  assign n3385 = n1693 & ~n3384 ;
  assign n3386 = n762 | n3385 ;
  assign n3387 = x238 | n797 ;
  assign n3388 = n1038 & n3308 ;
  assign n3389 = ~n2013 & n2725 ;
  assign n3390 = n3171 & ~n3389 ;
  assign n3391 = n1793 & n3297 ;
  assign n3392 = n3391 ^ x67 ^ 1'b0 ;
  assign n3393 = ~n430 & n577 ;
  assign n3394 = n546 & n942 ;
  assign n3395 = ~n801 & n3394 ;
  assign n3396 = n1787 & ~n3224 ;
  assign n3397 = n3396 ^ n1539 ^ 1'b0 ;
  assign n3398 = n3397 ^ n1656 ^ 1'b0 ;
  assign n3399 = ~n3395 & n3398 ;
  assign n3401 = n1170 | n1447 ;
  assign n3402 = n3401 ^ n1646 ^ 1'b0 ;
  assign n3400 = n1463 & ~n2455 ;
  assign n3403 = n3402 ^ n3400 ^ 1'b0 ;
  assign n3404 = n2500 ^ n2254 ^ x89 ;
  assign n3405 = ~n641 & n3404 ;
  assign n3406 = n3405 ^ n915 ^ 1'b0 ;
  assign n3407 = n1736 & n3406 ;
  assign n3408 = ( ~n553 & n844 ) | ( ~n553 & n1224 ) | ( n844 & n1224 ) ;
  assign n3409 = n2073 ^ x15 ^ 1'b0 ;
  assign n3410 = n2990 ^ n583 ^ 1'b0 ;
  assign n3411 = n1137 ^ n948 ^ 1'b0 ;
  assign n3412 = n701 | n3411 ;
  assign n3413 = n1985 & n3412 ;
  assign n3414 = n3165 & ~n3413 ;
  assign n3415 = n1077 | n3402 ;
  assign n3416 = n1822 | n3204 ;
  assign n3417 = x129 & n2083 ;
  assign n3419 = ~n1633 & n3050 ;
  assign n3418 = ~n1638 & n2012 ;
  assign n3420 = n3419 ^ n3418 ^ 1'b0 ;
  assign n3421 = n2271 ^ n753 ^ 1'b0 ;
  assign n3422 = n602 & n3421 ;
  assign n3423 = ~n1829 & n3422 ;
  assign n3424 = n3043 ^ x52 ^ 1'b0 ;
  assign n3425 = x154 | n937 ;
  assign n3426 = n3425 ^ x37 ^ 1'b0 ;
  assign n3427 = n3426 ^ n1779 ^ 1'b0 ;
  assign n3428 = n564 & n3427 ;
  assign n3429 = n2989 ^ n1148 ^ 1'b0 ;
  assign n3430 = ~n3428 & n3429 ;
  assign n3431 = n2474 ^ n1481 ^ 1'b0 ;
  assign n3432 = x101 & ~n2089 ;
  assign n3433 = x238 | n1031 ;
  assign n3434 = n1736 & ~n3433 ;
  assign n3436 = n798 & n1050 ;
  assign n3437 = n3436 ^ n1733 ^ 1'b0 ;
  assign n3435 = ~n2301 & n2328 ;
  assign n3438 = n3437 ^ n3435 ^ 1'b0 ;
  assign n3439 = n1120 ^ x207 ^ 1'b0 ;
  assign n3440 = ~n3035 & n3439 ;
  assign n3441 = n1093 ^ n381 ^ 1'b0 ;
  assign n3442 = n2414 & ~n3441 ;
  assign n3443 = n3417 ^ n877 ^ 1'b0 ;
  assign n3444 = n2916 ^ n392 ^ 1'b0 ;
  assign n3445 = ~x12 & n3444 ;
  assign n3446 = n3445 ^ n300 ^ 1'b0 ;
  assign n3447 = n288 ^ x76 ^ 1'b0 ;
  assign n3448 = n3447 ^ n2681 ^ x18 ;
  assign n3449 = x91 & ~n1313 ;
  assign n3450 = n666 & ~n3449 ;
  assign n3451 = n3450 ^ n987 ^ 1'b0 ;
  assign n3452 = n3451 ^ n1832 ^ 1'b0 ;
  assign n3453 = n3452 ^ n1622 ^ n1441 ;
  assign n3454 = n3453 ^ n1269 ^ 1'b0 ;
  assign n3455 = n341 | n641 ;
  assign n3456 = n1125 | n3455 ;
  assign n3457 = ~n1304 & n3456 ;
  assign n3458 = n3457 ^ n2562 ^ 1'b0 ;
  assign n3459 = n2040 & ~n2083 ;
  assign n3460 = n1282 | n3095 ;
  assign n3461 = n3459 & ~n3460 ;
  assign n3462 = n805 | n2440 ;
  assign n3463 = n593 & n3462 ;
  assign n3464 = n679 | n1280 ;
  assign n3465 = n3464 ^ n397 ^ 1'b0 ;
  assign n3466 = ~x65 & x242 ;
  assign n3467 = n3465 & n3466 ;
  assign n3468 = n1689 | n2027 ;
  assign n3469 = n3468 ^ n709 ^ x176 ;
  assign n3471 = n1635 & n1814 ;
  assign n3472 = ~n1694 & n3471 ;
  assign n3470 = x207 | n1925 ;
  assign n3473 = n3472 ^ n3470 ^ 1'b0 ;
  assign n3474 = n3473 ^ x245 ^ 1'b0 ;
  assign n3475 = n2749 | n3474 ;
  assign n3476 = n1423 | n3475 ;
  assign n3477 = n710 ^ x43 ^ 1'b0 ;
  assign n3478 = x219 & ~n2872 ;
  assign n3479 = n3176 & n3478 ;
  assign n3480 = n1621 | n2247 ;
  assign n3481 = ~n1859 & n3480 ;
  assign n3482 = n1174 | n2757 ;
  assign n3483 = n3482 ^ n966 ^ 1'b0 ;
  assign n3484 = n296 & n3483 ;
  assign n3485 = x124 & n345 ;
  assign n3488 = n325 & n333 ;
  assign n3486 = n1217 & ~n2402 ;
  assign n3487 = n3486 ^ n1372 ^ 1'b0 ;
  assign n3489 = n3488 ^ n3487 ^ 1'b0 ;
  assign n3490 = n3489 ^ x54 ^ 1'b0 ;
  assign n3491 = n3485 & ~n3490 ;
  assign n3492 = n3112 | n3308 ;
  assign n3493 = n1822 ^ n1058 ^ 1'b0 ;
  assign n3494 = x159 & ~n1611 ;
  assign n3495 = n3494 ^ n1776 ^ 1'b0 ;
  assign n3496 = n3493 & ~n3495 ;
  assign n3497 = x99 & x177 ;
  assign n3498 = n3497 ^ x54 ^ 1'b0 ;
  assign n3499 = x67 & n3498 ;
  assign n3500 = n1126 ^ x5 ^ 1'b0 ;
  assign n3501 = n1135 | n3500 ;
  assign n3502 = n3308 | n3501 ;
  assign n3503 = n3502 ^ n1903 ^ 1'b0 ;
  assign n3504 = ~n700 & n3414 ;
  assign n3505 = n1805 & n3504 ;
  assign n3506 = x87 & ~n476 ;
  assign n3507 = n3506 ^ n1638 ^ 1'b0 ;
  assign n3508 = n3507 ^ n2555 ^ 1'b0 ;
  assign n3509 = n2165 | n3508 ;
  assign n3510 = ~n748 & n1286 ;
  assign n3511 = n1241 & n3510 ;
  assign n3512 = n981 ^ n581 ^ 1'b0 ;
  assign n3513 = ~n3353 & n3512 ;
  assign n3514 = n3511 & n3513 ;
  assign n3515 = n2465 ^ n1068 ^ 1'b0 ;
  assign n3516 = n1490 | n3515 ;
  assign n3517 = n3047 & ~n3176 ;
  assign n3518 = n3517 ^ n1653 ^ 1'b0 ;
  assign n3519 = n1955 | n2849 ;
  assign n3520 = n2455 & ~n3519 ;
  assign n3521 = x160 | n3520 ;
  assign n3522 = n1961 ^ n770 ^ 1'b0 ;
  assign n3523 = n277 ^ x83 ^ 1'b0 ;
  assign n3524 = n490 & n3523 ;
  assign n3525 = n3524 ^ n307 ^ 1'b0 ;
  assign n3526 = n3522 & ~n3525 ;
  assign n3527 = n3288 ^ x62 ^ 1'b0 ;
  assign n3528 = n3527 ^ n3154 ^ 1'b0 ;
  assign n3529 = ~n810 & n2120 ;
  assign n3530 = ~n309 & n887 ;
  assign n3531 = n956 | n3530 ;
  assign n3532 = n1335 & ~n3055 ;
  assign n3533 = n965 ^ n607 ^ 1'b0 ;
  assign n3534 = ~n707 & n2291 ;
  assign n3535 = n2908 & n3534 ;
  assign n3536 = ~n2665 & n3535 ;
  assign n3537 = x207 & ~n397 ;
  assign n3538 = ~n1143 & n2825 ;
  assign n3539 = ~n3537 & n3538 ;
  assign n3540 = n325 & n3441 ;
  assign n3541 = n2804 & ~n3540 ;
  assign n3542 = ( ~n724 & n1182 ) | ( ~n724 & n1233 ) | ( n1182 & n1233 ) ;
  assign n3543 = n3112 | n3542 ;
  assign n3544 = n2219 ^ n1521 ^ 1'b0 ;
  assign n3545 = n1326 | n3544 ;
  assign n3546 = n1134 & n2165 ;
  assign n3547 = n1237 & ~n3546 ;
  assign n3548 = n3545 & n3547 ;
  assign n3549 = x83 & ~n2223 ;
  assign n3550 = ~n1061 & n1909 ;
  assign n3551 = n3550 ^ n516 ^ 1'b0 ;
  assign n3552 = ~n446 & n1037 ;
  assign n3553 = ~n669 & n3552 ;
  assign n3554 = ~x56 & n3553 ;
  assign n3555 = n3551 & ~n3554 ;
  assign n3556 = n772 & ~n3074 ;
  assign n3557 = n2370 ^ n892 ^ 1'b0 ;
  assign n3558 = x148 & ~n3557 ;
  assign n3559 = n1263 ^ n675 ^ 1'b0 ;
  assign n3560 = n1438 & ~n1926 ;
  assign n3561 = ~n452 & n3560 ;
  assign n3562 = n2972 ^ n2026 ^ n1850 ;
  assign n3563 = n2292 & n3562 ;
  assign n3564 = n1025 & n1038 ;
  assign n3565 = ~n720 & n3564 ;
  assign n3566 = n3565 ^ n2276 ^ 1'b0 ;
  assign n3567 = x95 | n3566 ;
  assign n3568 = n919 & n2611 ;
  assign n3569 = n3568 ^ n983 ^ 1'b0 ;
  assign n3571 = n1481 & n1525 ;
  assign n3572 = n784 | n3571 ;
  assign n3573 = n3203 | n3572 ;
  assign n3570 = x89 & ~n1957 ;
  assign n3574 = n3573 ^ n3570 ^ 1'b0 ;
  assign n3575 = n3574 ^ n3062 ^ n1920 ;
  assign n3576 = n271 | n2584 ;
  assign n3577 = n3177 ^ n2017 ^ n844 ;
  assign n3578 = n3577 ^ n2571 ^ 1'b0 ;
  assign n3579 = n482 & ~n1080 ;
  assign n3580 = ~n1654 & n3579 ;
  assign n3581 = ~n1904 & n2993 ;
  assign n3582 = ~n1731 & n3581 ;
  assign n3587 = n318 & n1814 ;
  assign n3588 = ~n559 & n3587 ;
  assign n3589 = n1969 & ~n3588 ;
  assign n3583 = ~n1387 & n2858 ;
  assign n3584 = ~n2252 & n3583 ;
  assign n3585 = n3134 & n3584 ;
  assign n3586 = n3143 & ~n3585 ;
  assign n3590 = n3589 ^ n3586 ^ 1'b0 ;
  assign n3591 = x112 | n833 ;
  assign n3592 = n460 | n3591 ;
  assign n3593 = n1262 & ~n3592 ;
  assign n3605 = n787 & n2768 ;
  assign n3606 = ~x253 & n3605 ;
  assign n3594 = x89 & x162 ;
  assign n3595 = n3594 ^ x182 ^ 1'b0 ;
  assign n3596 = n647 ^ x122 ^ 1'b0 ;
  assign n3597 = ~n3595 & n3596 ;
  assign n3598 = n1833 | n2528 ;
  assign n3599 = n734 & ~n3598 ;
  assign n3600 = n3599 ^ n2510 ^ 1'b0 ;
  assign n3601 = ~n2009 & n3600 ;
  assign n3602 = n1461 & n3601 ;
  assign n3603 = ~n3597 & n3602 ;
  assign n3604 = n3603 ^ n2765 ^ 1'b0 ;
  assign n3607 = n3606 ^ n3604 ^ 1'b0 ;
  assign n3608 = n2199 & ~n3607 ;
  assign n3609 = n3219 | n3488 ;
  assign n3610 = n3609 ^ n378 ^ 1'b0 ;
  assign n3611 = n1639 ^ x217 ^ 1'b0 ;
  assign n3612 = n3610 & n3611 ;
  assign n3613 = ~x27 & n3612 ;
  assign n3614 = n3195 ^ n669 ^ 1'b0 ;
  assign n3615 = x181 & n926 ;
  assign n3616 = n3615 ^ n1626 ^ 1'b0 ;
  assign n3617 = ~n1227 & n3616 ;
  assign n3618 = n1919 & n3617 ;
  assign n3619 = n3255 ^ n529 ^ 1'b0 ;
  assign n3620 = n3618 | n3619 ;
  assign n3621 = ( ~n1160 & n3614 ) | ( ~n1160 & n3620 ) | ( n3614 & n3620 ) ;
  assign n3622 = n1312 ^ n927 ^ n841 ;
  assign n3623 = x86 & ~n1673 ;
  assign n3624 = ~n3622 & n3623 ;
  assign n3625 = n3624 ^ n2671 ^ 1'b0 ;
  assign n3626 = n3625 ^ n688 ^ 1'b0 ;
  assign n3627 = x54 & ~n1703 ;
  assign n3628 = ~n552 & n3627 ;
  assign n3629 = n1390 | n3628 ;
  assign n3630 = n1529 ^ n1159 ^ n840 ;
  assign n3631 = n2107 & n2153 ;
  assign n3632 = ~n2082 & n3631 ;
  assign n3633 = x81 & ~n1016 ;
  assign n3634 = n3633 ^ n1096 ^ 1'b0 ;
  assign n3635 = n3634 ^ n1047 ^ 1'b0 ;
  assign n3636 = n361 & ~n1904 ;
  assign n3637 = n1021 | n2645 ;
  assign n3638 = n3637 ^ n283 ^ 1'b0 ;
  assign n3639 = n3636 & ~n3638 ;
  assign n3640 = x62 & n807 ;
  assign n3641 = ~n3639 & n3640 ;
  assign n3644 = ~n366 & n836 ;
  assign n3645 = n3644 ^ n278 ^ 1'b0 ;
  assign n3642 = n1444 & ~n3069 ;
  assign n3643 = n3642 ^ n3214 ^ 1'b0 ;
  assign n3646 = n3645 ^ n3643 ^ 1'b0 ;
  assign n3647 = n972 | n3646 ;
  assign n3648 = ~n1845 & n3187 ;
  assign n3649 = n1411 ^ n809 ^ 1'b0 ;
  assign n3650 = n3649 ^ n2472 ^ 1'b0 ;
  assign n3651 = n1639 & ~n3650 ;
  assign n3654 = n1521 ^ x127 ^ 1'b0 ;
  assign n3655 = ~n732 & n3654 ;
  assign n3652 = n1477 & n1898 ;
  assign n3653 = ~n3567 & n3652 ;
  assign n3656 = n3655 ^ n3653 ^ 1'b0 ;
  assign n3657 = n518 | n3536 ;
  assign n3658 = n1014 & ~n1777 ;
  assign n3659 = n3658 ^ x93 ^ 1'b0 ;
  assign n3660 = n1855 ^ n394 ^ 1'b0 ;
  assign n3661 = n3659 | n3660 ;
  assign n3662 = n1378 & n3661 ;
  assign n3663 = n2267 & ~n3662 ;
  assign n3664 = n3663 ^ n2273 ^ 1'b0 ;
  assign n3665 = n2650 ^ n1396 ^ 1'b0 ;
  assign n3666 = n2076 | n3665 ;
  assign n3667 = n856 & ~n3666 ;
  assign n3668 = n1939 ^ n1295 ^ 1'b0 ;
  assign n3669 = n3031 & n3668 ;
  assign n3670 = x241 & ~n3669 ;
  assign n3671 = ( ~n2158 & n2319 ) | ( ~n2158 & n2866 ) | ( n2319 & n2866 ) ;
  assign n3672 = ( n1242 & n3512 ) | ( n1242 & n3671 ) | ( n3512 & n3671 ) ;
  assign n3673 = n2203 ^ x160 ^ 1'b0 ;
  assign n3674 = n583 & n1020 ;
  assign n3675 = n3673 & n3674 ;
  assign n3676 = n3675 ^ n639 ^ 1'b0 ;
  assign n3677 = n605 | n1027 ;
  assign n3678 = n3677 ^ x18 ^ 1'b0 ;
  assign n3679 = ( ~n1192 & n1463 ) | ( ~n1192 & n3678 ) | ( n1463 & n3678 ) ;
  assign n3680 = n482 & n3679 ;
  assign n3681 = n3680 ^ x31 ^ 1'b0 ;
  assign n3682 = n1139 & n1670 ;
  assign n3683 = n3682 ^ n1167 ^ 1'b0 ;
  assign n3684 = n3105 & ~n3683 ;
  assign n3685 = ~n1766 & n3684 ;
  assign n3686 = n1343 | n2099 ;
  assign n3687 = n3686 ^ n1738 ^ 1'b0 ;
  assign n3688 = n3687 ^ x112 ^ 1'b0 ;
  assign n3689 = ~n1236 & n2529 ;
  assign n3690 = ~n1383 & n2119 ;
  assign n3691 = n1463 & n3690 ;
  assign n3692 = n3691 ^ n1859 ^ 1'b0 ;
  assign n3694 = x42 ^ x23 ^ 1'b0 ;
  assign n3693 = n1413 & n2367 ;
  assign n3695 = n3694 ^ n3693 ^ 1'b0 ;
  assign n3696 = n1126 ^ n930 ^ 1'b0 ;
  assign n3697 = n2411 & ~n3696 ;
  assign n3698 = ~n3613 & n3697 ;
  assign n3699 = n2527 ^ n2517 ^ 1'b0 ;
  assign n3700 = n2195 & n3699 ;
  assign n3701 = n1025 & n3700 ;
  assign n3702 = n3701 ^ n1828 ^ 1'b0 ;
  assign n3703 = n2964 ^ n2926 ^ 1'b0 ;
  assign n3704 = n1929 ^ n833 ^ 1'b0 ;
  assign n3705 = n2822 & ~n3704 ;
  assign n3706 = n2739 ^ x232 ^ 1'b0 ;
  assign n3707 = n718 | n3706 ;
  assign n3708 = n2435 | n3707 ;
  assign n3709 = n271 & ~n3708 ;
  assign n3710 = ~n887 & n2110 ;
  assign n3711 = n3038 ^ n666 ^ 1'b0 ;
  assign n3712 = n1094 ^ x141 ^ 1'b0 ;
  assign n3713 = ~n1546 & n3712 ;
  assign n3714 = n3713 ^ n1591 ^ 1'b0 ;
  assign n3715 = n1368 ^ n760 ^ 1'b0 ;
  assign n3716 = n325 | n3250 ;
  assign n3717 = n3645 & ~n3716 ;
  assign n3718 = ~n579 & n3717 ;
  assign n3719 = n707 & ~n954 ;
  assign n3720 = n3719 ^ n2916 ^ 1'b0 ;
  assign n3721 = ~n1549 & n1566 ;
  assign n3722 = n1953 ^ n840 ^ 1'b0 ;
  assign n3723 = n1337 | n3722 ;
  assign n3724 = n3430 ^ n343 ^ 1'b0 ;
  assign n3725 = n1846 & ~n3724 ;
  assign n3726 = ( n426 & n1441 ) | ( n426 & ~n3604 ) | ( n1441 & ~n3604 ) ;
  assign n3727 = n1791 | n1875 ;
  assign n3728 = n987 & n2277 ;
  assign n3729 = n3728 ^ n1747 ^ 1'b0 ;
  assign n3730 = n2761 & n2848 ;
  assign n3731 = ~n3729 & n3730 ;
  assign n3732 = n2715 ^ x76 ^ 1'b0 ;
  assign n3733 = ~n3731 & n3732 ;
  assign n3734 = n294 | n476 ;
  assign n3735 = n3734 ^ n1715 ^ 1'b0 ;
  assign n3736 = ~x93 & x128 ;
  assign n3737 = n3395 ^ n2750 ^ 1'b0 ;
  assign n3738 = ~n3736 & n3737 ;
  assign n3739 = ~n3735 & n3738 ;
  assign n3740 = x250 & n1969 ;
  assign n3741 = n3171 ^ n2122 ^ 1'b0 ;
  assign n3742 = n3740 & n3741 ;
  assign n3743 = n1457 & n1638 ;
  assign n3744 = n3743 ^ n2728 ^ 1'b0 ;
  assign n3745 = n3744 ^ n1311 ^ 1'b0 ;
  assign n3747 = n964 ^ n450 ^ n286 ;
  assign n3746 = n620 | n2553 ;
  assign n3748 = n3747 ^ n3746 ^ 1'b0 ;
  assign n3749 = n3630 ^ n2218 ^ x208 ;
  assign n3750 = ~x186 & n2975 ;
  assign n3751 = n3499 ^ n1546 ^ 1'b0 ;
  assign n3753 = n1162 ^ x68 ^ x3 ;
  assign n3752 = x175 & ~n1694 ;
  assign n3754 = n3753 ^ n3752 ^ 1'b0 ;
  assign n3755 = n2558 ^ x39 ^ 1'b0 ;
  assign n3756 = ~n3434 & n3750 ;
  assign n3757 = n337 & n2602 ;
  assign n3758 = n2135 & n3757 ;
  assign n3759 = n3250 | n3758 ;
  assign n3760 = n2765 & n3321 ;
  assign n3761 = n822 | n1093 ;
  assign n3762 = n3761 ^ n3694 ^ n1473 ;
  assign n3763 = n2435 ^ n571 ^ 1'b0 ;
  assign n3764 = n3116 ^ n2129 ^ 1'b0 ;
  assign n3765 = ~n526 & n1162 ;
  assign n3766 = ~n2872 & n3765 ;
  assign n3767 = n1679 | n2038 ;
  assign n3768 = x38 & ~n3767 ;
  assign n3769 = ~n1148 & n2786 ;
  assign n3770 = n1223 & n3769 ;
  assign n3771 = n1723 | n3348 ;
  assign n3772 = n2155 | n3771 ;
  assign n3773 = n1075 | n2739 ;
  assign n3777 = n800 & n1094 ;
  assign n3778 = ~x234 & n3777 ;
  assign n3774 = n867 ^ n430 ^ 1'b0 ;
  assign n3775 = n3774 ^ n1740 ^ 1'b0 ;
  assign n3776 = ~n313 & n3775 ;
  assign n3779 = n3778 ^ n3776 ^ 1'b0 ;
  assign n3780 = ~n815 & n1909 ;
  assign n3781 = ~n1217 & n1564 ;
  assign n3782 = n2119 & n3227 ;
  assign n3783 = n3483 & n3782 ;
  assign n3784 = ~n2747 & n3783 ;
  assign n3785 = n1769 ^ n642 ^ 1'b0 ;
  assign n3786 = n3499 & ~n3785 ;
  assign n3788 = n950 ^ n805 ^ 1'b0 ;
  assign n3789 = n1929 & n3788 ;
  assign n3787 = n1137 & ~n1285 ;
  assign n3790 = n3789 ^ n3787 ^ 1'b0 ;
  assign n3791 = n373 | n3790 ;
  assign n3792 = n2175 ^ x60 ^ 1'b0 ;
  assign n3793 = x39 | n273 ;
  assign n3794 = ~n3736 & n3793 ;
  assign n3795 = n2179 & ~n3165 ;
  assign n3796 = n468 | n2259 ;
  assign n3797 = ~n1812 & n2857 ;
  assign n3798 = ~n1014 & n3797 ;
  assign n3799 = ~n2186 & n3798 ;
  assign n3800 = n626 ^ n333 ^ 1'b0 ;
  assign n3801 = n3116 & ~n3800 ;
  assign n3802 = ~n3799 & n3801 ;
  assign n3803 = n1413 ^ n1314 ^ 1'b0 ;
  assign n3804 = n3388 & n3803 ;
  assign n3805 = ~n1374 & n3804 ;
  assign n3806 = n548 | n907 ;
  assign n3807 = n3806 ^ n2063 ^ 1'b0 ;
  assign n3808 = n2546 ^ n1202 ^ x51 ;
  assign n3809 = n3808 ^ n1405 ^ n1111 ;
  assign n3810 = n2962 ^ n2936 ^ 1'b0 ;
  assign n3811 = ( x50 & ~n975 ) | ( x50 & n2261 ) | ( ~n975 & n2261 ) ;
  assign n3812 = n996 & n1731 ;
  assign n3813 = n3812 ^ n1969 ^ 1'b0 ;
  assign n3814 = n1214 & n2696 ;
  assign n3815 = n3814 ^ n430 ^ 1'b0 ;
  assign n3816 = n3813 & n3815 ;
  assign n3817 = n3158 | n3816 ;
  assign n3818 = ~n456 & n1186 ;
  assign n3819 = n1632 & n3818 ;
  assign n3820 = n3819 ^ n2480 ^ 1'b0 ;
  assign n3832 = n1646 ^ n909 ^ 1'b0 ;
  assign n3827 = n951 ^ x231 ^ 1'b0 ;
  assign n3826 = ~n2576 & n3143 ;
  assign n3828 = n3827 ^ n3826 ^ 1'b0 ;
  assign n3821 = x217 & ~n1569 ;
  assign n3822 = ~n1325 & n3821 ;
  assign n3823 = n1365 & ~n3822 ;
  assign n3824 = n3823 ^ n3465 ^ 1'b0 ;
  assign n3825 = n3824 ^ n2168 ^ n1343 ;
  assign n3829 = n3828 ^ n3825 ^ 1'b0 ;
  assign n3830 = n3015 & n3829 ;
  assign n3831 = ~n605 & n3830 ;
  assign n3833 = n3832 ^ n3831 ^ 1'b0 ;
  assign n3834 = n2309 ^ n1709 ^ 1'b0 ;
  assign n3835 = ~n830 & n1330 ;
  assign n3836 = n3835 ^ n2447 ^ 1'b0 ;
  assign n3837 = n1112 ^ n894 ^ 1'b0 ;
  assign n3838 = x175 & n3837 ;
  assign n3839 = n2686 & n3838 ;
  assign n3840 = n2364 | n3839 ;
  assign n3841 = n3840 ^ n1472 ^ 1'b0 ;
  assign n3842 = ~x143 & n1549 ;
  assign n3843 = n1264 & n2904 ;
  assign n3844 = n3843 ^ n1840 ^ 1'b0 ;
  assign n3845 = n3844 ^ n1379 ^ 1'b0 ;
  assign n3848 = ~n296 & n543 ;
  assign n3846 = n1510 ^ n1007 ^ 1'b0 ;
  assign n3847 = ~n653 & n3846 ;
  assign n3849 = n3848 ^ n3847 ^ 1'b0 ;
  assign n3850 = n294 | n3849 ;
  assign n3851 = n2916 ^ n1693 ^ 1'b0 ;
  assign n3852 = n2112 & n3851 ;
  assign n3853 = n354 & ~n1746 ;
  assign n3854 = n577 & n3853 ;
  assign n3855 = n2142 ^ n2099 ^ 1'b0 ;
  assign n3856 = n3855 ^ n2338 ^ n1077 ;
  assign n3857 = n3289 ^ n2819 ^ 1'b0 ;
  assign n3858 = ~n3076 & n3857 ;
  assign n3859 = n2652 & ~n3858 ;
  assign n3860 = n3128 & ~n3551 ;
  assign n3861 = n1038 & n2129 ;
  assign n3862 = n3861 ^ n917 ^ 1'b0 ;
  assign n3863 = n3862 ^ n620 ^ 1'b0 ;
  assign n3864 = n880 & ~n2035 ;
  assign n3865 = n3864 ^ n2358 ^ 1'b0 ;
  assign n3866 = n3863 | n3865 ;
  assign n3867 = x155 & ~n1077 ;
  assign n3868 = n3867 ^ n1025 ^ 1'b0 ;
  assign n3869 = n3868 ^ n3533 ^ 1'b0 ;
  assign n3870 = ~n2314 & n3869 ;
  assign n3871 = n2855 ^ n1002 ^ 1'b0 ;
  assign n3872 = x28 | n3871 ;
  assign n3873 = n1139 ^ n683 ^ 1'b0 ;
  assign n3874 = n3057 | n3873 ;
  assign n3875 = ~n2021 & n3874 ;
  assign n3877 = ~n1423 & n2947 ;
  assign n3876 = n1106 & n2593 ;
  assign n3878 = n3877 ^ n3876 ^ 1'b0 ;
  assign n3879 = n1299 & n1864 ;
  assign n3880 = n1332 & n1890 ;
  assign n3881 = n3880 ^ n1440 ^ 1'b0 ;
  assign n3882 = x25 & n1028 ;
  assign n3883 = n3881 | n3882 ;
  assign n3884 = n832 | n1385 ;
  assign n3885 = n662 ^ n417 ^ 1'b0 ;
  assign n3886 = ~n1733 & n3885 ;
  assign n3887 = ~n2427 & n3886 ;
  assign n3888 = n3884 & n3887 ;
  assign n3889 = n866 & n1444 ;
  assign n3890 = n1207 & n3889 ;
  assign n3891 = n3890 ^ n2302 ^ 1'b0 ;
  assign n3892 = ~n2371 & n3563 ;
  assign n3893 = n3892 ^ n838 ^ 1'b0 ;
  assign n3894 = n3071 ^ n2819 ^ 1'b0 ;
  assign n3895 = ~n1499 & n3894 ;
  assign n3898 = n1461 & ~n2794 ;
  assign n3899 = ~n3361 & n3898 ;
  assign n3900 = n1847 ^ n1134 ^ 1'b0 ;
  assign n3901 = ~n3899 & n3900 ;
  assign n3896 = n1093 | n1383 ;
  assign n3897 = n3219 | n3896 ;
  assign n3902 = n3901 ^ n3897 ^ 1'b0 ;
  assign n3903 = n663 & n2621 ;
  assign n3904 = n3902 & n3903 ;
  assign n3905 = n3904 ^ n1727 ^ 1'b0 ;
  assign n3906 = ( n1312 & ~n3895 ) | ( n1312 & n3905 ) | ( ~n3895 & n3905 ) ;
  assign n3907 = n1769 | n1936 ;
  assign n3908 = n3907 ^ n2350 ^ 1'b0 ;
  assign n3909 = n2618 & n3908 ;
  assign n3910 = n1366 & n3909 ;
  assign n3911 = n2314 & ~n3910 ;
  assign n3912 = x101 & ~n1064 ;
  assign n3913 = n3912 ^ n2110 ^ 1'b0 ;
  assign n3914 = n3451 ^ n3216 ^ 1'b0 ;
  assign n3915 = n1178 | n2338 ;
  assign n3916 = n2672 & n3915 ;
  assign n3917 = n2841 & n3916 ;
  assign n3918 = n2586 ^ n1501 ^ 1'b0 ;
  assign n3919 = ~n1083 & n3918 ;
  assign n3920 = n3284 & n3919 ;
  assign n3921 = ~n651 & n1521 ;
  assign n3922 = ~n3872 & n3921 ;
  assign n3923 = n3436 ^ n2423 ^ 1'b0 ;
  assign n3924 = n2075 & ~n3923 ;
  assign n3925 = n3616 & n3924 ;
  assign n3927 = n1785 ^ x73 ^ 1'b0 ;
  assign n3928 = x230 & ~n3927 ;
  assign n3926 = n1521 ^ n1191 ^ 1'b0 ;
  assign n3929 = n3928 ^ n3926 ^ 1'b0 ;
  assign n3930 = x8 & n343 ;
  assign n3931 = n278 & n3930 ;
  assign n3932 = n2853 ^ n2561 ^ 1'b0 ;
  assign n3933 = ~n3931 & n3932 ;
  assign n3934 = ~n1988 & n3933 ;
  assign n3935 = ~n3929 & n3934 ;
  assign n3936 = x2 & n3935 ;
  assign n3937 = n1931 & ~n3459 ;
  assign n3938 = n3937 ^ n3856 ^ 1'b0 ;
  assign n3939 = ~x29 & n2119 ;
  assign n3940 = ( ~n741 & n1793 ) | ( ~n741 & n3939 ) | ( n1793 & n3939 ) ;
  assign n3941 = n1152 & ~n3727 ;
  assign n3942 = ~n968 & n3941 ;
  assign n3943 = n3942 ^ n1985 ^ 1'b0 ;
  assign n3944 = n286 | n2266 ;
  assign n3945 = x205 | n3944 ;
  assign n3946 = ~n2223 & n3945 ;
  assign n3947 = n2789 ^ n1111 ^ 1'b0 ;
  assign n3948 = n3947 ^ n2716 ^ 1'b0 ;
  assign n3949 = ~n949 & n3637 ;
  assign n3950 = n514 & n3949 ;
  assign n3951 = n923 & ~n3740 ;
  assign n3952 = n2975 ^ n374 ^ 1'b0 ;
  assign n3953 = n611 & ~n3952 ;
  assign n3954 = n3953 ^ n3761 ^ 1'b0 ;
  assign n3955 = x109 & ~n3954 ;
  assign n3956 = ~n3189 & n3955 ;
  assign n3959 = n2166 & n2539 ;
  assign n3957 = ( x189 & n269 ) | ( x189 & n552 ) | ( n269 & n552 ) ;
  assign n3958 = x41 & n3957 ;
  assign n3960 = n3959 ^ n3958 ^ 1'b0 ;
  assign n3961 = ~n498 & n1692 ;
  assign n3962 = n3961 ^ n3333 ^ 1'b0 ;
  assign n3963 = n470 | n3962 ;
  assign n3964 = n3791 & ~n3963 ;
  assign n3965 = ~n1641 & n3855 ;
  assign n3966 = n3589 ^ n3090 ^ 1'b0 ;
  assign n3967 = n1780 ^ n581 ^ 1'b0 ;
  assign n3968 = n1808 & n3967 ;
  assign n3969 = n884 & n3968 ;
  assign n3970 = ~n1360 & n3969 ;
  assign n3971 = n3295 ^ n1866 ^ 1'b0 ;
  assign n3972 = n761 ^ x160 ^ 1'b0 ;
  assign n3973 = n1104 | n3972 ;
  assign n3974 = n1262 & ~n3973 ;
  assign n3975 = ~n2037 & n3830 ;
  assign n3976 = n3975 ^ n1658 ^ 1'b0 ;
  assign n3977 = ~n1236 & n1336 ;
  assign n3978 = n937 & n3977 ;
  assign n3979 = ( x61 & ~n448 ) | ( x61 & n789 ) | ( ~n448 & n789 ) ;
  assign n3980 = n1904 ^ n1049 ^ 1'b0 ;
  assign n3981 = ~n3979 & n3980 ;
  assign n3982 = ~n3978 & n3981 ;
  assign n3983 = n1843 & n2714 ;
  assign n3984 = n3983 ^ n611 ^ 1'b0 ;
  assign n3985 = n415 & n1268 ;
  assign n3986 = n1601 & ~n3985 ;
  assign n3987 = n1350 | n3986 ;
  assign n3988 = n3987 ^ n1023 ^ 1'b0 ;
  assign n3989 = ( n774 & ~n1740 ) | ( n774 & n2665 ) | ( ~n1740 & n2665 ) ;
  assign n3990 = x65 & n1969 ;
  assign n3991 = n3989 & n3990 ;
  assign n3992 = x160 & n1604 ;
  assign n3993 = x157 & n3992 ;
  assign n3994 = n666 | n2890 ;
  assign n3995 = n3014 | n3158 ;
  assign n3996 = n3670 ^ n2324 ^ 1'b0 ;
  assign n3997 = x222 & ~n3302 ;
  assign n3998 = ~n1214 & n3997 ;
  assign n3999 = n550 & n3511 ;
  assign n4000 = x237 & ~n1693 ;
  assign n4001 = ~n3999 & n4000 ;
  assign n4002 = ~n2655 & n3528 ;
  assign n4003 = n1573 & n3865 ;
  assign n4004 = n2207 ^ n2161 ^ 1'b0 ;
  assign n4005 = ~n3910 & n4004 ;
  assign n4006 = n1436 ^ x124 ^ 1'b0 ;
  assign n4007 = n4006 ^ x147 ^ 1'b0 ;
  assign n4008 = x36 & ~n4007 ;
  assign n4009 = ( n278 & n637 ) | ( n278 & n1709 ) | ( n637 & n1709 ) ;
  assign n4010 = n3071 ^ n1856 ^ 1'b0 ;
  assign n4011 = n3209 & ~n4010 ;
  assign n4012 = ~n1707 & n4011 ;
  assign n4013 = n3773 ^ n347 ^ 1'b0 ;
  assign n4014 = n2715 & n2962 ;
  assign n4015 = n2925 ^ n2718 ^ 1'b0 ;
  assign n4016 = n3859 | n4015 ;
  assign n4017 = n2765 ^ n548 ^ 1'b0 ;
  assign n4018 = n3488 | n4017 ;
  assign n4019 = n1021 | n4018 ;
  assign n4020 = n4019 ^ n2689 ^ 1'b0 ;
  assign n4021 = n3723 & ~n3855 ;
  assign n4022 = n1252 | n3641 ;
  assign n4023 = n631 | n2254 ;
  assign n4024 = n1540 | n4023 ;
  assign n4025 = ~n985 & n1150 ;
  assign n4026 = n4025 ^ n2099 ^ 1'b0 ;
  assign n4027 = ( n2358 & n2955 ) | ( n2358 & ~n4026 ) | ( n2955 & ~n4026 ) ;
  assign n4028 = n444 ^ n397 ^ 1'b0 ;
  assign n4029 = n1914 | n4028 ;
  assign n4030 = n779 & ~n1059 ;
  assign n4031 = n4030 ^ n2099 ^ 1'b0 ;
  assign n4032 = n4031 ^ n1158 ^ 1'b0 ;
  assign n4033 = n1135 | n4032 ;
  assign n4034 = n2648 | n4033 ;
  assign n4035 = n2333 ^ n1159 ^ x4 ;
  assign n4036 = x218 | n2670 ;
  assign n4037 = n4036 ^ n468 ^ 1'b0 ;
  assign n4038 = n553 ^ n349 ^ 1'b0 ;
  assign n4039 = n649 & n4038 ;
  assign n4040 = x209 & n4039 ;
  assign n4041 = n4040 ^ n2098 ^ n1328 ;
  assign n4042 = n1485 & ~n4006 ;
  assign n4043 = ~n4041 & n4042 ;
  assign n4044 = n875 | n1690 ;
  assign n4045 = n4044 ^ n1968 ^ 1'b0 ;
  assign n4046 = n3863 ^ x150 ^ 1'b0 ;
  assign n4047 = ~n1606 & n4046 ;
  assign n4048 = x14 | n505 ;
  assign n4049 = n4048 ^ n1159 ^ 1'b0 ;
  assign n4050 = n4047 & n4049 ;
  assign n4051 = ~n2947 & n4050 ;
  assign n4052 = ~x81 & n2577 ;
  assign n4053 = n4052 ^ n2386 ^ 1'b0 ;
  assign n4054 = ~x155 & n4053 ;
  assign n4055 = n4054 ^ n1517 ^ 1'b0 ;
  assign n4057 = n1251 & ~n2281 ;
  assign n4058 = n4057 ^ n2132 ^ 1'b0 ;
  assign n4056 = n442 | n4001 ;
  assign n4059 = n4058 ^ n4056 ^ 1'b0 ;
  assign n4060 = n286 ^ x150 ^ 1'b0 ;
  assign n4061 = x67 & ~n4060 ;
  assign n4062 = ~n3099 & n4061 ;
  assign n4063 = ~n639 & n4062 ;
  assign n4064 = n1178 & ~n1879 ;
  assign n4065 = n2599 & n4064 ;
  assign n4066 = n4065 ^ n3516 ^ 1'b0 ;
  assign n4067 = n988 ^ x108 ^ 1'b0 ;
  assign n4068 = n3102 ^ x44 ^ 1'b0 ;
  assign n4069 = n1732 & ~n4068 ;
  assign n4070 = n1549 & n2040 ;
  assign n4071 = n4070 ^ n1784 ^ 1'b0 ;
  assign n4072 = n4071 ^ n3432 ^ 1'b0 ;
  assign n4073 = n296 & ~n4072 ;
  assign n4074 = n4073 ^ x3 ^ 1'b0 ;
  assign n4075 = n1754 | n3727 ;
  assign n4076 = n4075 ^ n1521 ^ 1'b0 ;
  assign n4077 = n1409 | n3759 ;
  assign n4078 = n575 & n3495 ;
  assign n4079 = n4078 ^ n3575 ^ 1'b0 ;
  assign n4080 = n1485 | n2037 ;
  assign n4081 = n951 | n2870 ;
  assign n4082 = x226 & ~n3292 ;
  assign n4083 = ~n1429 & n4082 ;
  assign n4084 = n3546 ^ x53 ^ 1'b0 ;
  assign n4085 = n772 & ~n2105 ;
  assign n4086 = n4085 ^ n1784 ^ 1'b0 ;
  assign n4087 = ~n2854 & n4086 ;
  assign n4088 = x76 & ~n2426 ;
  assign n4089 = n4087 & n4088 ;
  assign n4090 = x232 & ~n1650 ;
  assign n4091 = n4090 ^ n3822 ^ 1'b0 ;
  assign n4092 = ~n1002 & n1125 ;
  assign n4093 = x77 & n4092 ;
  assign n4094 = n4093 ^ n3024 ^ 1'b0 ;
  assign n4095 = n521 | n1632 ;
  assign n4096 = n4095 ^ n963 ^ 1'b0 ;
  assign n4097 = n1056 ^ n1006 ^ 1'b0 ;
  assign n4098 = ~n551 & n4097 ;
  assign n4099 = n4098 ^ n2012 ^ 1'b0 ;
  assign n4100 = ( n2257 & n2689 ) | ( n2257 & ~n4099 ) | ( n2689 & ~n4099 ) ;
  assign n4101 = n3590 | n4100 ;
  assign n4102 = n3692 ^ n2591 ^ 1'b0 ;
  assign n4103 = n1337 & ~n4102 ;
  assign n4104 = n574 | n577 ;
  assign n4105 = n2404 ^ n1738 ^ 1'b0 ;
  assign n4106 = ~n4104 & n4105 ;
  assign n4107 = ~x135 & n4106 ;
  assign n4108 = n1344 & n2778 ;
  assign n4110 = x130 & ~n1568 ;
  assign n4111 = n4110 ^ n2261 ^ 1'b0 ;
  assign n4109 = n323 | n1378 ;
  assign n4112 = n4111 ^ n4109 ^ n590 ;
  assign n4113 = n2978 ^ n1560 ^ 1'b0 ;
  assign n4114 = x81 & n1653 ;
  assign n4115 = n311 & n4114 ;
  assign n4116 = n4115 ^ n1314 ^ 1'b0 ;
  assign n4117 = n915 & n1411 ;
  assign n4118 = n315 ^ x85 ^ 1'b0 ;
  assign n4119 = ~n4117 & n4118 ;
  assign n4120 = ( x230 & ~n444 ) | ( x230 & n2898 ) | ( ~n444 & n2898 ) ;
  assign n4121 = n1527 ^ n497 ^ 1'b0 ;
  assign n4122 = x18 & n4121 ;
  assign n4123 = n1216 ^ n1170 ^ 1'b0 ;
  assign n4124 = x102 & n4123 ;
  assign n4125 = ~n2889 & n4124 ;
  assign n4126 = ~x246 & n4125 ;
  assign n4127 = n4122 & ~n4126 ;
  assign n4128 = n4127 ^ n3606 ^ 1'b0 ;
  assign n4129 = ( n4054 & n4120 ) | ( n4054 & n4128 ) | ( n4120 & n4128 ) ;
  assign n4130 = n399 | n3981 ;
  assign n4131 = n1667 | n4130 ;
  assign n4132 = n1686 & ~n4131 ;
  assign n4133 = n1400 ^ n285 ^ 1'b0 ;
  assign n4134 = n390 & ~n4133 ;
  assign n4135 = n1009 | n4134 ;
  assign n4136 = n2001 | n4135 ;
  assign n4137 = n3076 ^ n423 ^ 1'b0 ;
  assign n4138 = n1599 | n4137 ;
  assign n4139 = ~n983 & n2893 ;
  assign n4140 = n4139 ^ n2589 ^ 1'b0 ;
  assign n4141 = ~n1232 & n3031 ;
  assign n4142 = n4141 ^ n281 ^ 1'b0 ;
  assign n4143 = ( n3479 & n4140 ) | ( n3479 & n4142 ) | ( n4140 & n4142 ) ;
  assign n4144 = n1266 ^ x34 ^ 1'b0 ;
  assign n4145 = n1646 | n1907 ;
  assign n4146 = n766 | n4145 ;
  assign n4147 = n4146 ^ n1882 ^ 1'b0 ;
  assign n4148 = n2241 & n2431 ;
  assign n4149 = n4148 ^ n2175 ^ 1'b0 ;
  assign n4150 = n2879 ^ x70 ^ 1'b0 ;
  assign n4151 = ~n2869 & n4150 ;
  assign n4152 = n2042 ^ n341 ^ 1'b0 ;
  assign n4153 = ~n1527 & n2212 ;
  assign n4154 = ~n4152 & n4153 ;
  assign n4155 = n4151 & ~n4154 ;
  assign n4156 = n4155 ^ n1485 ^ 1'b0 ;
  assign n4157 = n1912 | n2715 ;
  assign n4158 = n2658 ^ x7 ^ 1'b0 ;
  assign n4159 = ~n1042 & n4158 ;
  assign n4160 = n4157 & ~n4159 ;
  assign n4161 = n399 & n4160 ;
  assign n4162 = n352 ^ n325 ^ 1'b0 ;
  assign n4163 = n4162 ^ n2886 ^ 1'b0 ;
  assign n4164 = n1952 & ~n4163 ;
  assign n4165 = n1239 | n2318 ;
  assign n4166 = x112 & ~n4165 ;
  assign n4167 = n1062 & ~n2252 ;
  assign n4168 = n4166 & n4167 ;
  assign n4169 = ~n1075 & n1888 ;
  assign n4170 = n1190 | n1628 ;
  assign n4171 = n2277 ^ n1328 ^ 1'b0 ;
  assign n4172 = ~n4170 & n4171 ;
  assign n4173 = ~n1757 & n4172 ;
  assign n4174 = n456 ^ x95 ^ 1'b0 ;
  assign n4175 = n585 | n4174 ;
  assign n4176 = x186 | n4175 ;
  assign n4177 = n3583 ^ n3100 ^ x115 ;
  assign n4178 = n1111 | n4177 ;
  assign n4179 = n1903 ^ n347 ^ 1'b0 ;
  assign n4180 = n3886 & ~n4179 ;
  assign n4181 = n1795 ^ n653 ^ 1'b0 ;
  assign n4182 = n2878 & n4181 ;
  assign n4183 = n4182 ^ n581 ^ 1'b0 ;
  assign n4185 = x24 & ~n1709 ;
  assign n4184 = n2648 & ~n3505 ;
  assign n4186 = n4185 ^ n4184 ^ 1'b0 ;
  assign n4187 = n4186 ^ n4067 ^ 1'b0 ;
  assign n4188 = n3986 | n4187 ;
  assign n4189 = n460 | n1376 ;
  assign n4190 = ~n327 & n2278 ;
  assign n4191 = ~n2071 & n4190 ;
  assign n4192 = n409 & n4191 ;
  assign n4193 = n1824 & n4192 ;
  assign n4194 = n2804 | n4193 ;
  assign n4195 = x53 | n4194 ;
  assign n4196 = ~n790 & n4195 ;
  assign n4197 = n4196 ^ n1409 ^ 1'b0 ;
  assign n4198 = x199 & ~n3033 ;
  assign n4199 = n4198 ^ n2081 ^ n1983 ;
  assign n4200 = ~n307 & n969 ;
  assign n4201 = n4200 ^ n899 ^ 1'b0 ;
  assign n4202 = n2350 ^ n1569 ^ 1'b0 ;
  assign n4203 = n1777 | n4202 ;
  assign n4204 = n3287 & ~n4203 ;
  assign n4205 = x199 | n4204 ;
  assign n4206 = n787 & n896 ;
  assign n4207 = n614 & n4206 ;
  assign n4208 = n1404 & ~n3632 ;
  assign n4209 = n1183 ^ x125 ^ 1'b0 ;
  assign n4210 = n4209 ^ n2825 ^ 1'b0 ;
  assign n4211 = n589 | n4210 ;
  assign n4212 = x95 & ~n3284 ;
  assign n4213 = n4212 ^ n4176 ^ 1'b0 ;
  assign n4214 = n4168 ^ n1405 ^ 1'b0 ;
  assign n4215 = n1732 & ~n3451 ;
  assign n4216 = ~n574 & n4215 ;
  assign n4217 = ~n1431 & n4216 ;
  assign n4220 = n1707 | n2306 ;
  assign n4218 = ~n1202 & n2597 ;
  assign n4219 = n4218 ^ n981 ^ 1'b0 ;
  assign n4221 = n4220 ^ n4219 ^ 1'b0 ;
  assign n4222 = n2273 & ~n4221 ;
  assign n4223 = n4222 ^ n2681 ^ 1'b0 ;
  assign n4224 = ~n2148 & n2704 ;
  assign n4225 = n4224 ^ n806 ^ 1'b0 ;
  assign n4226 = n1169 | n4225 ;
  assign n4227 = n4226 ^ n2755 ^ 1'b0 ;
  assign n4235 = x167 & n3524 ;
  assign n4236 = n4235 ^ n698 ^ 1'b0 ;
  assign n4237 = n3481 & ~n4236 ;
  assign n4228 = ~n423 & n3186 ;
  assign n4229 = n1757 & n4228 ;
  assign n4230 = n1861 ^ n1784 ^ 1'b0 ;
  assign n4231 = n485 & n4230 ;
  assign n4232 = n1339 & n4231 ;
  assign n4233 = n288 | n4232 ;
  assign n4234 = n4229 & n4233 ;
  assign n4238 = n4237 ^ n4234 ^ 1'b0 ;
  assign n4239 = x60 & n2929 ;
  assign n4240 = n2395 ^ n349 ^ 1'b0 ;
  assign n4241 = x53 & ~n4240 ;
  assign n4242 = n296 | n1468 ;
  assign n4243 = ( ~n3733 & n4241 ) | ( ~n3733 & n4242 ) | ( n4241 & n4242 ) ;
  assign n4244 = ~x21 & n1541 ;
  assign n4245 = n1191 & n4244 ;
  assign n4246 = n4245 ^ n1974 ^ 1'b0 ;
  assign n4247 = n1194 & ~n4246 ;
  assign n4248 = n1117 | n4159 ;
  assign n4249 = n4248 ^ n296 ^ 1'b0 ;
  assign n4250 = n4249 ^ n3436 ^ 1'b0 ;
  assign n4251 = n1916 & ~n4250 ;
  assign n4252 = n2645 & ~n3546 ;
  assign n4253 = n4252 ^ n1658 ^ 1'b0 ;
  assign n4254 = n835 & n2517 ;
  assign n4255 = n381 & n4254 ;
  assign n4256 = n1337 | n4255 ;
  assign n4257 = ~x154 & n3065 ;
  assign n4258 = n639 | n4257 ;
  assign n4259 = n4257 ^ x186 ^ 1'b0 ;
  assign n4260 = n3524 & ~n4259 ;
  assign n4266 = n1075 ^ n1027 ^ 1'b0 ;
  assign n4267 = n1324 | n4266 ;
  assign n4268 = n4267 ^ n1152 ^ x196 ;
  assign n4261 = n3899 ^ n1173 ^ 1'b0 ;
  assign n4262 = ~n709 & n2507 ;
  assign n4263 = n1903 & n4262 ;
  assign n4264 = n4263 ^ n2169 ^ 1'b0 ;
  assign n4265 = n4261 & ~n4264 ;
  assign n4269 = n4268 ^ n4265 ^ 1'b0 ;
  assign n4270 = ~n2581 & n4269 ;
  assign n4271 = n384 | n862 ;
  assign n4272 = ( n482 & n895 ) | ( n482 & ~n4271 ) | ( n895 & ~n4271 ) ;
  assign n4273 = n4272 ^ n1252 ^ n345 ;
  assign n4274 = n3522 & ~n4273 ;
  assign n4275 = n1693 ^ n1307 ^ 1'b0 ;
  assign n4276 = n1560 & n4275 ;
  assign n4277 = n918 & n2074 ;
  assign n4278 = n4277 ^ n1141 ^ 1'b0 ;
  assign n4279 = ( x251 & n1787 ) | ( x251 & ~n3428 ) | ( n1787 & ~n3428 ) ;
  assign n4280 = x252 & n4279 ;
  assign n4281 = ~n1252 & n4280 ;
  assign n4282 = n2263 ^ n2155 ^ 1'b0 ;
  assign n4283 = n3373 & n4282 ;
  assign n4284 = n4283 ^ n3126 ^ 1'b0 ;
  assign n4285 = n1148 & ~n1575 ;
  assign n4286 = n4285 ^ n753 ^ 1'b0 ;
  assign n4287 = n4286 ^ n1007 ^ 1'b0 ;
  assign n4288 = n1217 & n1228 ;
  assign n4289 = n4288 ^ x218 ^ 1'b0 ;
  assign n4290 = n2158 & ~n4289 ;
  assign n4291 = n4290 ^ n3645 ^ n3083 ;
  assign n4293 = x9 & ~x109 ;
  assign n4294 = ( n1833 & n4061 ) | ( n1833 & ~n4293 ) | ( n4061 & ~n4293 ) ;
  assign n4292 = n2109 & n2320 ;
  assign n4295 = n4294 ^ n4292 ^ 1'b0 ;
  assign n4296 = n1255 | n4295 ;
  assign n4297 = n2990 ^ n779 ^ 1'b0 ;
  assign n4298 = n2970 ^ n1907 ^ 1'b0 ;
  assign n4299 = n1363 ^ n692 ^ 1'b0 ;
  assign n4300 = ~n1337 & n4299 ;
  assign n4301 = x214 & ~n4300 ;
  assign n4302 = n1210 & ~n4301 ;
  assign n4303 = n1610 ^ n436 ^ 1'b0 ;
  assign n4304 = ~n2872 & n4303 ;
  assign n4305 = n1920 & ~n2207 ;
  assign n4306 = ~n2855 & n4305 ;
  assign n4307 = n1407 ^ n508 ^ 1'b0 ;
  assign n4308 = n3499 | n4307 ;
  assign n4309 = n3245 ^ x226 ^ 1'b0 ;
  assign n4310 = n3387 & n4309 ;
  assign n4312 = n1328 ^ n1068 ^ 1'b0 ;
  assign n4313 = n3512 & ~n4312 ;
  assign n4311 = ~n397 & n1479 ;
  assign n4314 = n4313 ^ n4311 ^ 1'b0 ;
  assign n4315 = n2166 & n2702 ;
  assign n4316 = n1952 ^ x106 ^ 1'b0 ;
  assign n4317 = ~n2793 & n3379 ;
  assign n4318 = n2205 & n4317 ;
  assign n4319 = ~n1684 & n3667 ;
  assign n4320 = n4319 ^ n3226 ^ 1'b0 ;
  assign n4321 = n4213 & n4320 ;
  assign n4322 = n605 & ~n3204 ;
  assign n4323 = ~x43 & n4322 ;
  assign n4324 = x186 & ~n3287 ;
  assign n4325 = n4324 ^ n2593 ^ 1'b0 ;
  assign n4326 = n2985 ^ n1148 ^ 1'b0 ;
  assign n4327 = n4326 ^ n1252 ^ 1'b0 ;
  assign n4328 = ( ~x35 & x156 ) | ( ~x35 & n1888 ) | ( x156 & n1888 ) ;
  assign n4329 = ~n1190 & n4328 ;
  assign n4330 = n2576 ^ n1455 ^ 1'b0 ;
  assign n4331 = ~n2145 & n4330 ;
  assign n4332 = ~n977 & n4331 ;
  assign n4333 = n3868 & n4332 ;
  assign n4334 = n267 & ~n2270 ;
  assign n4335 = n4334 ^ n2604 ^ 1'b0 ;
  assign n4336 = n4333 | n4335 ;
  assign n4337 = n1608 ^ n657 ^ 1'b0 ;
  assign n4338 = ~n1605 & n4337 ;
  assign n4339 = x59 | n3488 ;
  assign n4340 = n1441 & ~n4339 ;
  assign n4341 = ( n335 & ~n4267 ) | ( n335 & n4340 ) | ( ~n4267 & n4340 ) ;
  assign n4342 = n4341 ^ n1872 ^ 1'b0 ;
  assign n4343 = n2314 & n4342 ;
  assign n4344 = n1226 & n2263 ;
  assign n4345 = n4344 ^ n551 ^ 1'b0 ;
  assign n4346 = n1646 & n4345 ;
  assign n4347 = n4346 ^ x165 ^ 1'b0 ;
  assign n4348 = ~n1061 & n4347 ;
  assign n4349 = n1775 & n4348 ;
  assign n4350 = ~n380 & n1564 ;
  assign n4351 = n3269 ^ n2267 ^ x130 ;
  assign n4352 = ( ~n1690 & n1732 ) | ( ~n1690 & n4351 ) | ( n1732 & n4351 ) ;
  assign n4353 = n4352 ^ x152 ^ 1'b0 ;
  assign n4354 = ~n846 & n4353 ;
  assign n4355 = ~n3767 & n4354 ;
  assign n4356 = n4355 ^ n669 ^ 1'b0 ;
  assign n4357 = n1920 ^ n372 ^ 1'b0 ;
  assign n4358 = n2571 | n4357 ;
  assign n4359 = n4356 & ~n4358 ;
  assign n4360 = ~n4352 & n4359 ;
  assign n4361 = n4350 | n4360 ;
  assign n4364 = n1697 ^ n397 ^ 1'b0 ;
  assign n4362 = x167 & n1268 ;
  assign n4363 = ~n456 & n4362 ;
  assign n4365 = n4364 ^ n4363 ^ 1'b0 ;
  assign n4366 = n2686 | n4365 ;
  assign n4367 = x218 & ~n2643 ;
  assign n4368 = n4367 ^ n1080 ^ 1'b0 ;
  assign n4369 = n1242 & ~n3412 ;
  assign n4370 = n4369 ^ n3312 ^ 1'b0 ;
  assign n4371 = n4370 ^ n2985 ^ 1'b0 ;
  assign n4372 = n2863 | n4371 ;
  assign n4373 = ~n1642 & n2624 ;
  assign n4374 = n524 & ~n2259 ;
  assign n4375 = n4374 ^ n1980 ^ 1'b0 ;
  assign n4376 = n1405 & n4375 ;
  assign n4377 = n888 & n2076 ;
  assign n4378 = x236 & n4377 ;
  assign n4379 = n4243 ^ x157 ^ 1'b0 ;
  assign n4380 = x184 & ~n4379 ;
  assign n4381 = n2368 ^ n2087 ^ 1'b0 ;
  assign n4382 = n3503 | n4381 ;
  assign n4383 = x245 & n1742 ;
  assign n4384 = n4383 ^ n1064 ^ 1'b0 ;
  assign n4385 = n663 & n4384 ;
  assign n4386 = n366 | n4385 ;
  assign n4387 = n667 | n1503 ;
  assign n4388 = x63 | n4387 ;
  assign n4389 = n1525 ^ n1178 ^ 1'b0 ;
  assign n4390 = ( n1339 & ~n4388 ) | ( n1339 & n4389 ) | ( ~n4388 & n4389 ) ;
  assign n4391 = n1784 ^ x135 ^ 1'b0 ;
  assign n4392 = n1237 & n4391 ;
  assign n4393 = n271 & n4392 ;
  assign n4394 = n4132 | n4393 ;
  assign n4395 = n2351 | n4394 ;
  assign n4396 = n2081 ^ n1857 ^ 1'b0 ;
  assign n4397 = n730 & n1344 ;
  assign n4398 = n4397 ^ n480 ^ 1'b0 ;
  assign n4399 = n3076 ^ n1657 ^ 1'b0 ;
  assign n4400 = n395 | n4151 ;
  assign n4411 = n3298 ^ n1093 ^ 1'b0 ;
  assign n4401 = n2858 ^ n358 ^ 1'b0 ;
  assign n4402 = ~n2387 & n4401 ;
  assign n4403 = n271 | n1851 ;
  assign n4404 = n392 | n4403 ;
  assign n4405 = n3713 & n4404 ;
  assign n4406 = n4405 ^ n855 ^ 1'b0 ;
  assign n4407 = n4402 & ~n4406 ;
  assign n4408 = n4407 ^ n2274 ^ 1'b0 ;
  assign n4409 = n2102 & ~n4408 ;
  assign n4410 = n1556 & n4409 ;
  assign n4412 = n4411 ^ n4410 ^ 1'b0 ;
  assign n4413 = n2519 ^ n269 ^ 1'b0 ;
  assign n4414 = n3619 & n4413 ;
  assign n4415 = n294 | n1630 ;
  assign n4416 = n4415 ^ n2336 ^ 1'b0 ;
  assign n4417 = n1167 | n2869 ;
  assign n4418 = n1330 ^ n688 ^ 1'b0 ;
  assign n4420 = n1654 ^ n463 ^ 1'b0 ;
  assign n4419 = n760 & n1075 ;
  assign n4421 = n4420 ^ n4419 ^ 1'b0 ;
  assign n4422 = n4421 ^ n1348 ^ 1'b0 ;
  assign n4423 = n1120 | n3459 ;
  assign n4424 = ~n987 & n3903 ;
  assign n4425 = n1511 ^ x171 ^ 1'b0 ;
  assign n4426 = ( n1685 & n1961 ) | ( n1685 & n2626 ) | ( n1961 & n2626 ) ;
  assign n4427 = n4426 ^ n1023 ^ 1'b0 ;
  assign n4428 = ~n4425 & n4427 ;
  assign n4429 = n934 | n2979 ;
  assign n4430 = n4429 ^ n754 ^ 1'b0 ;
  assign n4431 = n2539 | n3947 ;
  assign n4432 = n1923 ^ n432 ^ 1'b0 ;
  assign n4433 = x123 | n4197 ;
  assign n4434 = n3388 & ~n4433 ;
  assign n4435 = ~n877 & n2412 ;
  assign n4436 = n4435 ^ n824 ^ 1'b0 ;
  assign n4437 = x154 ^ x151 ^ 1'b0 ;
  assign n4438 = n1483 & n4437 ;
  assign n4439 = n1700 & n1959 ;
  assign n4440 = ~n271 & n4439 ;
  assign n4441 = n1974 & n2412 ;
  assign n4442 = ~n4260 & n4441 ;
  assign n4443 = n4442 ^ n1010 ^ 1'b0 ;
  assign n4444 = n4440 | n4443 ;
  assign n4445 = ( n267 & n2022 ) | ( n267 & ~n3412 ) | ( n2022 & ~n3412 ) ;
  assign n4446 = ~n3711 & n4445 ;
  assign n4447 = n4446 ^ x207 ^ 1'b0 ;
  assign n4448 = ~x219 & n2314 ;
  assign n4449 = n1521 ^ n733 ^ 1'b0 ;
  assign n4450 = n4249 ^ x67 ^ 1'b0 ;
  assign n4451 = ~n4054 & n4450 ;
  assign n4452 = ( n2267 & ~n3409 ) | ( n2267 & n3945 ) | ( ~n3409 & n3945 ) ;
  assign n4453 = ~n2210 & n3959 ;
  assign n4454 = n4453 ^ n4304 ^ 1'b0 ;
  assign n4455 = n1326 | n2134 ;
  assign n4458 = n1510 | n1836 ;
  assign n4459 = n4458 ^ n4058 ^ 1'b0 ;
  assign n4456 = n1571 ^ n279 ^ 1'b0 ;
  assign n4457 = ~n3117 & n4456 ;
  assign n4460 = n4459 ^ n4457 ^ 1'b0 ;
  assign n4463 = x56 & ~n3606 ;
  assign n4464 = n2836 & n4463 ;
  assign n4461 = n1824 ^ n538 ^ 1'b0 ;
  assign n4462 = n485 & n4461 ;
  assign n4465 = n4464 ^ n4462 ^ 1'b0 ;
  assign n4466 = n3746 ^ n1864 ^ 1'b0 ;
  assign n4467 = ( x226 & ~n1192 ) | ( x226 & n2819 ) | ( ~n1192 & n2819 ) ;
  assign n4468 = n1376 ^ n361 ^ 1'b0 ;
  assign n4469 = n3552 & n4468 ;
  assign n4470 = ~n583 & n4469 ;
  assign n4471 = n1010 | n3542 ;
  assign n4472 = n4471 ^ n1740 ^ 1'b0 ;
  assign n4473 = n4470 & n4472 ;
  assign n4474 = n1635 & n3929 ;
  assign n4475 = ~n3694 & n4474 ;
  assign n4476 = n1629 ^ n488 ^ n279 ;
  assign n4477 = n1400 & ~n4476 ;
  assign n4478 = n4477 ^ n2954 ^ 1'b0 ;
  assign n4479 = n4478 ^ n2898 ^ n1378 ;
  assign n4480 = n444 & n3626 ;
  assign n4483 = n3637 ^ n2003 ^ 1'b0 ;
  assign n4481 = n420 | n1382 ;
  assign n4482 = n4278 & n4481 ;
  assign n4484 = n4483 ^ n4482 ^ 1'b0 ;
  assign n4485 = n561 & n789 ;
  assign n4486 = n3420 ^ n3148 ^ 1'b0 ;
  assign n4487 = ~n4485 & n4486 ;
  assign n4488 = n975 ^ n926 ^ 1'b0 ;
  assign n4489 = n4488 ^ n3195 ^ 1'b0 ;
  assign n4490 = n1059 ^ n536 ^ 1'b0 ;
  assign n4491 = n3794 | n4490 ;
  assign n4492 = n381 | n4491 ;
  assign n4493 = n4492 ^ n1622 ^ 1'b0 ;
  assign n4494 = n963 | n2146 ;
  assign n4495 = n4494 ^ n285 ^ 1'b0 ;
  assign n4496 = n4495 ^ n337 ^ 1'b0 ;
  assign n4497 = n4496 ^ n1354 ^ 1'b0 ;
  assign n4498 = ~n3407 & n4375 ;
  assign n4499 = n1777 | n4242 ;
  assign n4500 = x182 | n729 ;
  assign n4501 = n2079 & n3721 ;
  assign n4502 = n1546 ^ x96 ^ 1'b0 ;
  assign n4503 = x111 | n4502 ;
  assign n4504 = x83 & n2684 ;
  assign n4505 = ~x24 & n4504 ;
  assign n4506 = n573 | n4505 ;
  assign n4507 = n4208 ^ x14 ^ 1'b0 ;
  assign n4508 = n701 ^ n445 ^ 1'b0 ;
  assign n4509 = n3879 & ~n4508 ;
  assign n4510 = ~n474 & n4283 ;
  assign n4512 = n2746 ^ n372 ^ 1'b0 ;
  assign n4511 = x16 & n1622 ;
  assign n4513 = n4512 ^ n4511 ^ 1'b0 ;
  assign n4514 = n2331 & ~n2500 ;
  assign n4515 = x62 & n4514 ;
  assign n4516 = ( n994 & n4513 ) | ( n994 & n4515 ) | ( n4513 & n4515 ) ;
  assign n4517 = n1762 & n3361 ;
  assign n4518 = n4517 ^ n1953 ^ 1'b0 ;
  assign n4519 = n1291 | n4518 ;
  assign n4520 = n4519 ^ n2065 ^ 1'b0 ;
  assign n4521 = n1258 & n1928 ;
  assign n4522 = n281 & ~n577 ;
  assign n4523 = n1320 & n4522 ;
  assign n4524 = n2896 ^ n1007 ^ 1'b0 ;
  assign n4525 = n4523 & n4524 ;
  assign n4526 = ~n4521 & n4525 ;
  assign n4527 = n2796 & ~n3575 ;
  assign n4528 = n4527 ^ n1263 ^ 1'b0 ;
  assign n4529 = ~n2093 & n4528 ;
  assign n4530 = n989 ^ x231 ^ 1'b0 ;
  assign n4531 = n1190 | n2853 ;
  assign n4532 = n1312 & ~n4531 ;
  assign n4533 = n4532 ^ n1298 ^ 1'b0 ;
  assign n4534 = n2273 & n4533 ;
  assign n4535 = n4530 & n4534 ;
  assign n4536 = n1828 & n4535 ;
  assign n4537 = n4536 ^ x25 ^ 1'b0 ;
  assign n4538 = n771 | n3446 ;
  assign n4539 = n2305 ^ n390 ^ 1'b0 ;
  assign n4540 = n4538 | n4539 ;
  assign n4541 = n607 & ~n633 ;
  assign n4542 = n2480 & ~n4541 ;
  assign n4543 = n4542 ^ n3890 ^ 1'b0 ;
  assign n4544 = x34 | n2403 ;
  assign n4545 = n754 ^ x12 ^ 1'b0 ;
  assign n4546 = n4545 ^ n602 ^ 1'b0 ;
  assign n4547 = n304 & ~n2513 ;
  assign n4548 = n4547 ^ n4024 ^ 1'b0 ;
  assign n4549 = x142 | n628 ;
  assign n4550 = n2106 ^ n637 ^ 1'b0 ;
  assign n4551 = n3203 & n4550 ;
  assign n4552 = n3703 & n4551 ;
  assign n4553 = x243 & ~n432 ;
  assign n4554 = n4553 ^ n3770 ^ n1314 ;
  assign n4555 = n4122 | n4554 ;
  assign n4556 = ~n363 & n1656 ;
  assign n4557 = n985 | n1497 ;
  assign n4558 = n1505 & ~n4557 ;
  assign n4559 = n4558 ^ n1370 ^ 1'b0 ;
  assign n4560 = n4556 | n4559 ;
  assign n4561 = n3355 ^ x112 ^ 1'b0 ;
  assign n4562 = x34 & ~n4561 ;
  assign n4563 = n1108 | n2760 ;
  assign n4564 = n2239 | n4563 ;
  assign n4565 = n2826 & n4564 ;
  assign n4566 = n3124 ^ n2382 ^ 1'b0 ;
  assign n4567 = n987 & n1961 ;
  assign n4568 = n3910 & n4567 ;
  assign n4569 = ~n2632 & n2899 ;
  assign n4570 = n4569 ^ n4143 ^ 1'b0 ;
  assign n4571 = n830 & n4570 ;
  assign n4572 = x128 & n3467 ;
  assign n4573 = ~n2621 & n4572 ;
  assign n4574 = n708 | n1167 ;
  assign n4575 = n859 ^ x91 ^ 1'b0 ;
  assign n4576 = ~n4111 & n4575 ;
  assign n4577 = n2099 & ~n4576 ;
  assign n4578 = n593 & ~n2304 ;
  assign n4579 = n726 ^ n474 ^ 1'b0 ;
  assign n4580 = x15 | n4579 ;
  assign n4581 = n1252 & ~n4580 ;
  assign n4582 = n4578 & n4581 ;
  assign n4583 = n3694 & ~n4582 ;
  assign n4584 = n3137 & n4583 ;
  assign n4585 = n2397 & n2687 ;
  assign n4586 = ~n2309 & n4585 ;
  assign n4587 = n1150 | n1660 ;
  assign n4588 = n3626 ^ n1689 ^ 1'b0 ;
  assign n4589 = n4587 & n4588 ;
  assign n4590 = n4589 ^ n4260 ^ n1335 ;
  assign n4591 = x97 & n833 ;
  assign n4592 = n4591 ^ n808 ^ 1'b0 ;
  assign n4593 = n830 ^ n349 ^ 1'b0 ;
  assign n4594 = n2896 & n4593 ;
  assign n4595 = ~n2354 & n4594 ;
  assign n4596 = n2482 ^ n2014 ^ 1'b0 ;
  assign n4597 = n1693 | n3986 ;
  assign n4598 = n4597 ^ n1546 ^ 1'b0 ;
  assign n4599 = n3741 & ~n4598 ;
  assign n4600 = n3332 & n4599 ;
  assign n4601 = ~n1236 & n4600 ;
  assign n4602 = n445 | n1339 ;
  assign n4603 = n3622 ^ n1207 ^ 1'b0 ;
  assign n4604 = n4602 | n4603 ;
  assign n4605 = n4604 ^ n2562 ^ 1'b0 ;
  assign n4608 = n2929 ^ n1879 ^ 1'b0 ;
  assign n4606 = ~n2893 & n2976 ;
  assign n4607 = n2814 | n4606 ;
  assign n4609 = n4608 ^ n4607 ^ 1'b0 ;
  assign n4610 = ~n1343 & n2865 ;
  assign n4611 = n4610 ^ n1507 ^ 1'b0 ;
  assign n4612 = n3498 ^ x123 ^ 1'b0 ;
  assign n4613 = n2546 | n4612 ;
  assign n4614 = n3957 & ~n4613 ;
  assign n4615 = n4611 & n4614 ;
  assign n4616 = n4615 ^ n3248 ^ n1894 ;
  assign n4617 = n931 & ~n3848 ;
  assign n4618 = ~n758 & n1970 ;
  assign n4619 = ~n1082 & n1853 ;
  assign n4620 = n4582 | n4619 ;
  assign n4621 = ~n989 & n4451 ;
  assign n4622 = n4621 ^ n3611 ^ 1'b0 ;
  assign n4623 = n1757 ^ x84 ^ 1'b0 ;
  assign n4624 = n349 | n4623 ;
  assign n4625 = n1064 & ~n4624 ;
  assign n4626 = ~n3006 & n4625 ;
  assign n4627 = n3057 | n4626 ;
  assign n4633 = x51 & n1992 ;
  assign n4634 = n2941 & n4633 ;
  assign n4635 = n1673 | n4634 ;
  assign n4636 = n4635 ^ n3187 ^ 1'b0 ;
  assign n4629 = n2134 ^ n926 ^ 1'b0 ;
  assign n4630 = ( x45 & n597 ) | ( x45 & ~n4629 ) | ( n597 & ~n4629 ) ;
  assign n4628 = n271 & n3481 ;
  assign n4631 = n4630 ^ n4628 ^ 1'b0 ;
  assign n4632 = ~n2168 & n4631 ;
  assign n4637 = n4636 ^ n4632 ^ n1499 ;
  assign n4638 = n1145 ^ x183 ^ 1'b0 ;
  assign n4639 = ~n1723 & n2935 ;
  assign n4640 = n4638 & n4639 ;
  assign n4641 = n4640 ^ n2352 ^ 1'b0 ;
  assign n4642 = n1245 ^ n1169 ^ 1'b0 ;
  assign n4643 = x21 & n4642 ;
  assign n4644 = n833 & ~n4643 ;
  assign n4645 = x177 | n1305 ;
  assign n4646 = n849 & n4645 ;
  assign n4647 = ~n3636 & n4646 ;
  assign n4648 = n1114 | n4647 ;
  assign n4649 = ~n2391 & n4648 ;
  assign n4650 = ~n4644 & n4649 ;
  assign n4651 = n2247 ^ n528 ^ 1'b0 ;
  assign n4652 = n1643 & ~n4651 ;
  assign n4653 = n4652 ^ n4190 ^ 1'b0 ;
  assign n4655 = x74 & n456 ;
  assign n4654 = n556 | n3086 ;
  assign n4656 = n4655 ^ n4654 ^ 1'b0 ;
  assign n4657 = n4656 ^ x170 ^ 1'b0 ;
  assign n4658 = n1540 & ~n2848 ;
  assign n4659 = n1273 & n1446 ;
  assign n4660 = n320 & n4659 ;
  assign n4661 = n1646 ^ n903 ^ 1'b0 ;
  assign n4662 = ~n1474 & n4122 ;
  assign n4663 = n4662 ^ n867 ^ 1'b0 ;
  assign n4664 = n4047 & n4663 ;
  assign n4665 = n1802 ^ n1332 ^ 1'b0 ;
  assign n4666 = n1040 & ~n4665 ;
  assign n4667 = n3000 | n4584 ;
  assign n4668 = n4666 | n4667 ;
  assign n4671 = n1181 ^ n998 ^ 1'b0 ;
  assign n4672 = n2575 ^ n1593 ^ 1'b0 ;
  assign n4673 = n4671 & n4672 ;
  assign n4669 = n1618 & ~n3307 ;
  assign n4670 = n1038 & ~n4669 ;
  assign n4674 = n4673 ^ n4670 ^ 1'b0 ;
  assign n4675 = n337 & ~n1955 ;
  assign n4676 = n478 & n4675 ;
  assign n4677 = ( n1715 & n2354 ) | ( n1715 & ~n2766 ) | ( n2354 & ~n2766 ) ;
  assign n4678 = n4215 ^ n559 ^ 1'b0 ;
  assign n4679 = n4145 | n4678 ;
  assign n4680 = n4679 ^ n3307 ^ 1'b0 ;
  assign n4683 = n1038 & n2640 ;
  assign n4684 = ~n561 & n4683 ;
  assign n4681 = ~n1979 & n4530 ;
  assign n4682 = n4681 ^ n3046 ^ 1'b0 ;
  assign n4685 = n4684 ^ n4682 ^ 1'b0 ;
  assign n4686 = n490 | n815 ;
  assign n4687 = n4686 ^ n3588 ^ 1'b0 ;
  assign n4688 = n2899 & n4687 ;
  assign n4689 = ~n4322 & n4688 ;
  assign n4690 = n3020 & n3223 ;
  assign n4691 = n1082 | n3485 ;
  assign n4692 = ~x115 & n4691 ;
  assign n4693 = n4692 ^ n673 ^ 1'b0 ;
  assign n4694 = n1696 ^ n1546 ^ 1'b0 ;
  assign n4695 = ~n2711 & n4694 ;
  assign n4696 = n2892 | n4236 ;
  assign n4698 = ~x102 & n446 ;
  assign n4697 = ~n1646 & n3816 ;
  assign n4699 = n4698 ^ n4697 ^ 1'b0 ;
  assign n4700 = n4696 & n4699 ;
  assign n4701 = n608 & ~n2799 ;
  assign n4702 = n924 & ~n3575 ;
  assign n4703 = ~n4144 & n4702 ;
  assign n4704 = n2315 ^ x194 ^ 1'b0 ;
  assign n4705 = n2496 & ~n4704 ;
  assign n4706 = n2146 ^ x80 ^ 1'b0 ;
  assign n4707 = n3000 | n4706 ;
  assign n4708 = n3936 ^ n1594 ^ 1'b0 ;
  assign n4709 = n294 & ~n1195 ;
  assign n4710 = n304 & ~n4709 ;
  assign n4711 = n4710 ^ n3656 ^ 1'b0 ;
  assign n4714 = n4024 ^ n1822 ^ 1'b0 ;
  assign n4712 = n3193 & n3237 ;
  assign n4713 = ~n2333 & n4712 ;
  assign n4715 = n4714 ^ n4713 ^ 1'b0 ;
  assign n4716 = ~n2235 & n4304 ;
  assign n4717 = n793 & n2693 ;
  assign n4718 = n2006 & n4717 ;
  assign n4719 = n4718 ^ n4653 ^ 1'b0 ;
  assign n4723 = n2873 ^ n1775 ^ 1'b0 ;
  assign n4720 = x222 ^ x24 ^ 1'b0 ;
  assign n4721 = ~n2037 & n4720 ;
  assign n4722 = n4308 & n4721 ;
  assign n4724 = n4723 ^ n4722 ^ 1'b0 ;
  assign n4725 = n1477 ^ n866 ^ 1'b0 ;
  assign n4726 = ~n628 & n4725 ;
  assign n4727 = n2806 | n4726 ;
  assign n4728 = ~x71 & n1554 ;
  assign n4729 = n4728 ^ n3043 ^ 1'b0 ;
  assign n4730 = ~x123 & x156 ;
  assign n4731 = n4730 ^ n2261 ^ 1'b0 ;
  assign n4732 = x150 & ~n3939 ;
  assign n4733 = n2836 & n4732 ;
  assign n4734 = n4629 ^ n1405 ^ 1'b0 ;
  assign n4735 = n825 & ~n1727 ;
  assign n4736 = ~n2932 & n4735 ;
  assign n4737 = n2746 | n4736 ;
  assign n4738 = ~n1523 & n2652 ;
  assign n4739 = ( n1337 & n2624 ) | ( n1337 & ~n2761 ) | ( n2624 & ~n2761 ) ;
  assign n4740 = n4580 ^ n3514 ^ 1'b0 ;
  assign n4741 = ~n4739 & n4740 ;
  assign n4743 = n317 | n1707 ;
  assign n4742 = n869 | n3024 ;
  assign n4744 = n4743 ^ n4742 ^ 1'b0 ;
  assign n4745 = n3984 & ~n4744 ;
  assign n4746 = x231 & ~n3774 ;
  assign n4747 = n4746 ^ n2947 ^ 1'b0 ;
  assign n4748 = n4208 ^ n283 ^ 1'b0 ;
  assign n4749 = n936 & ~n4748 ;
  assign n4750 = n1483 ^ n651 ^ 1'b0 ;
  assign n4751 = ~n803 & n4750 ;
  assign n4752 = n3811 | n4751 ;
  assign n4753 = n4752 ^ n2393 ^ 1'b0 ;
  assign n4754 = n403 & n1139 ;
  assign n4755 = n4754 ^ n1531 ^ 1'b0 ;
  assign n4756 = n4755 ^ n720 ^ 1'b0 ;
  assign n4757 = n2731 & n4756 ;
  assign n4758 = n936 & n1165 ;
  assign n4759 = n4758 ^ n1365 ^ 1'b0 ;
  assign n4760 = n2747 & n4759 ;
  assign n4762 = n1025 & n3469 ;
  assign n4763 = n4762 ^ n2910 ^ 1'b0 ;
  assign n4761 = ~n2009 & n4290 ;
  assign n4764 = n4763 ^ n4761 ^ 1'b0 ;
  assign n4765 = ~n1443 & n4652 ;
  assign n4766 = ~n1605 & n4765 ;
  assign n4767 = n2750 & n3581 ;
  assign n4768 = n1738 & ~n4767 ;
  assign n4769 = n4768 ^ n1366 ^ 1'b0 ;
  assign n4770 = ~n1449 & n4769 ;
  assign n4771 = n4491 & n4770 ;
  assign n4772 = n3219 ^ n2011 ^ 1'b0 ;
  assign n4773 = ~n2807 & n4772 ;
  assign n4774 = x238 & ~n840 ;
  assign n4775 = n4774 ^ x144 ^ 1'b0 ;
  assign n4776 = n3187 | n4775 ;
  assign n4777 = ( ~n732 & n2186 ) | ( ~n732 & n2718 ) | ( n2186 & n2718 ) ;
  assign n4778 = n4084 ^ n1909 ^ 1'b0 ;
  assign n4779 = n4777 & n4778 ;
  assign n4780 = n4378 ^ n1264 ^ n1075 ;
  assign n4781 = n3489 ^ n2426 ^ 1'b0 ;
  assign n4782 = n3428 & n4781 ;
  assign n4784 = n1397 | n2384 ;
  assign n4783 = n540 & ~n626 ;
  assign n4785 = n4784 ^ n4783 ^ 1'b0 ;
  assign n4786 = n677 | n1961 ;
  assign n4787 = n2314 | n4786 ;
  assign n4788 = n4787 ^ n2452 ^ 1'b0 ;
  assign n4789 = n3090 | n3673 ;
  assign n4790 = x202 & x218 ;
  assign n4791 = n4790 ^ n1575 ^ 1'b0 ;
  assign n4792 = n4791 ^ n598 ^ 1'b0 ;
  assign n4793 = n4734 & ~n4792 ;
  assign n4794 = n2675 ^ n2469 ^ 1'b0 ;
  assign n4795 = ~n556 & n2839 ;
  assign n4796 = n1840 & n4795 ;
  assign n4797 = n1266 & n2658 ;
  assign n4798 = ~n1837 & n4797 ;
  assign n4799 = n4798 ^ n2926 ^ 1'b0 ;
  assign n4802 = n672 ^ n540 ^ 1'b0 ;
  assign n4800 = ~n1419 & n1571 ;
  assign n4801 = n2257 & n4800 ;
  assign n4803 = n4802 ^ n4801 ^ n1414 ;
  assign n4804 = n4803 ^ n1572 ^ 1'b0 ;
  assign n4805 = n647 & n1661 ;
  assign n4806 = ~n723 & n4805 ;
  assign n4807 = n3727 | n4138 ;
  assign n4808 = n4806 & ~n4807 ;
  assign n4810 = n1345 & ~n2465 ;
  assign n4811 = n4810 ^ n1080 ^ 1'b0 ;
  assign n4809 = n897 & ~n1824 ;
  assign n4812 = n4811 ^ n4809 ^ 1'b0 ;
  assign n4814 = n928 & n1970 ;
  assign n4813 = n749 & ~n2505 ;
  assign n4815 = n4814 ^ n4813 ^ 1'b0 ;
  assign n4816 = n3871 ^ n2593 ^ 1'b0 ;
  assign n4817 = n1935 ^ n840 ^ 1'b0 ;
  assign n4818 = n1419 | n4817 ;
  assign n4819 = n4818 ^ n4166 ^ 1'b0 ;
  assign n4820 = n1076 ^ x65 ^ 1'b0 ;
  assign n4821 = n3118 & ~n4820 ;
  assign n4822 = n557 & ~n3447 ;
  assign n4823 = ~n2589 & n4822 ;
  assign n4824 = ~n4821 & n4823 ;
  assign n4825 = x42 | n1126 ;
  assign n4826 = n4825 ^ n3107 ^ 1'b0 ;
  assign n4827 = n1646 & ~n4826 ;
  assign n4828 = ~x7 & n4827 ;
  assign n4829 = ~n448 & n2543 ;
  assign n4830 = n4169 ^ x20 ^ 1'b0 ;
  assign n4831 = ~n4829 & n4830 ;
  assign n4832 = n1671 ^ n957 ^ 1'b0 ;
  assign n4833 = x159 & n4832 ;
  assign n4834 = ~n3430 & n4833 ;
  assign n4835 = ~n2303 & n2397 ;
  assign n4836 = n3143 & ~n3950 ;
  assign n4837 = n3906 ^ n2428 ^ 1'b0 ;
  assign n4838 = n1164 & n4837 ;
  assign n4839 = n2855 & n3735 ;
  assign n4840 = n4839 ^ n3116 ^ 1'b0 ;
  assign n4841 = n2132 & n4840 ;
  assign n4842 = n1932 & ~n3336 ;
  assign n4843 = n1243 & n4842 ;
  assign n4844 = n3039 ^ n877 ^ 1'b0 ;
  assign n4845 = ~n4843 & n4844 ;
  assign n4846 = n2696 ^ n1643 ^ 1'b0 ;
  assign n4847 = ~n3505 & n3800 ;
  assign n4848 = ~n2221 & n4847 ;
  assign n4849 = x226 & n3543 ;
  assign n4850 = n2061 | n2246 ;
  assign n4851 = n4092 & ~n4850 ;
  assign n4852 = x59 & n2143 ;
  assign n4853 = n2100 & n4852 ;
  assign n4854 = n1337 ^ n460 ^ 1'b0 ;
  assign n4855 = ~n2416 & n4854 ;
  assign n4856 = n4172 & ~n4855 ;
  assign n4857 = n4856 ^ n2302 ^ 1'b0 ;
  assign n4858 = x208 & ~n713 ;
  assign n4859 = n4545 & n4858 ;
  assign n4860 = n4859 ^ n3492 ^ 1'b0 ;
  assign n4861 = ~n774 & n1808 ;
  assign n4862 = n4861 ^ n3622 ^ 1'b0 ;
  assign n4863 = n4862 ^ n859 ^ 1'b0 ;
  assign n4864 = ~n963 & n3255 ;
  assign n4865 = n4864 ^ n2022 ^ 1'b0 ;
  assign n4866 = n3028 & ~n4865 ;
  assign n4867 = n3800 ^ n726 ^ 1'b0 ;
  assign n4868 = n480 & ~n1417 ;
  assign n4869 = ~n474 & n4868 ;
  assign n4870 = n4869 ^ n955 ^ 1'b0 ;
  assign n4871 = n4867 & ~n4870 ;
  assign n4872 = n2439 & ~n3331 ;
  assign n4873 = n4799 ^ n4797 ^ 1'b0 ;
  assign n4874 = ~n343 & n1593 ;
  assign n4875 = n1507 ^ n390 ^ 1'b0 ;
  assign n4876 = n2399 | n2529 ;
  assign n4877 = n4876 ^ n3779 ^ 1'b0 ;
  assign n4878 = x9 & n4031 ;
  assign n4879 = ~n4310 & n4878 ;
  assign n4880 = n4688 ^ n1400 ^ 1'b0 ;
  assign n4881 = x141 & n4880 ;
  assign n4882 = x24 | x207 ;
  assign n4883 = ~n4263 & n4509 ;
  assign n4884 = ~n4882 & n4883 ;
  assign n4885 = n4582 ^ n401 ^ 1'b0 ;
  assign n4886 = ~n4372 & n4885 ;
  assign n4887 = n2883 ^ n607 ^ 1'b0 ;
  assign n4888 = n1413 & ~n4887 ;
  assign n4889 = n3773 | n4888 ;
  assign n4890 = x63 & n2089 ;
  assign n4891 = ~n2416 & n4890 ;
  assign n4892 = n4099 ^ n754 ^ 1'b0 ;
  assign n4893 = ~n4891 & n4892 ;
  assign n4894 = n436 & n4893 ;
  assign n4895 = ~n347 & n366 ;
  assign n4896 = n4895 ^ n979 ^ 1'b0 ;
  assign n4897 = x160 | n858 ;
  assign n4898 = n4897 ^ n4126 ^ 1'b0 ;
  assign n4899 = ~n4896 & n4898 ;
  assign n4900 = n1118 | n4899 ;
  assign n4901 = n2497 | n4900 ;
  assign n4902 = n3177 & ~n3599 ;
  assign n4903 = n4902 ^ n1907 ^ 1'b0 ;
  assign n4904 = n579 & n4903 ;
  assign n4905 = n666 & n4402 ;
  assign n4906 = n4905 ^ n3313 ^ 1'b0 ;
  assign n4907 = n4904 & ~n4906 ;
  assign n4908 = n3847 ^ n2760 ^ 1'b0 ;
  assign n4909 = n4907 & ~n4908 ;
  assign n4910 = n1514 & ~n2395 ;
  assign n4912 = n797 & ~n1706 ;
  assign n4913 = n4912 ^ n1658 ^ 1'b0 ;
  assign n4914 = n1739 & n4913 ;
  assign n4911 = n3698 ^ n3459 ^ 1'b0 ;
  assign n4915 = n4914 ^ n4911 ^ 1'b0 ;
  assign n4916 = n552 | n4915 ;
  assign n4917 = n4630 ^ n3449 ^ 1'b0 ;
  assign n4918 = x44 & n1025 ;
  assign n4919 = n339 & n4918 ;
  assign n4920 = n2604 | n4919 ;
  assign n4921 = n1158 & n4326 ;
  assign n4922 = n3139 & n4921 ;
  assign n4923 = ( n3132 & n4920 ) | ( n3132 & n4922 ) | ( n4920 & n4922 ) ;
  assign n4925 = n1248 & n2345 ;
  assign n4926 = n4925 ^ n587 ^ 1'b0 ;
  assign n4924 = n1496 & ~n1835 ;
  assign n4927 = n4926 ^ n4924 ^ 1'b0 ;
  assign n4930 = ~n1666 & n3221 ;
  assign n4931 = n2766 & ~n4930 ;
  assign n4932 = ~n2333 & n4931 ;
  assign n4928 = n502 | n694 ;
  assign n4929 = ~n4515 & n4928 ;
  assign n4933 = n4932 ^ n4929 ^ 1'b0 ;
  assign n4941 = n4215 ^ n915 ^ x203 ;
  assign n4942 = x6 & n4172 ;
  assign n4943 = n4941 & n4942 ;
  assign n4934 = n647 & n3123 ;
  assign n4935 = ( x16 & ~n493 ) | ( x16 & n4934 ) | ( ~n493 & n4934 ) ;
  assign n4936 = n4935 ^ n2487 ^ 1'b0 ;
  assign n4937 = n4936 ^ n3789 ^ 1'b0 ;
  assign n4938 = n1602 & ~n4937 ;
  assign n4939 = n4938 ^ n1298 ^ 1'b0 ;
  assign n4940 = n4939 ^ n3518 ^ 1'b0 ;
  assign n4944 = n4943 ^ n4940 ^ n1241 ;
  assign n4945 = x85 & n1981 ;
  assign n4946 = n4945 ^ n4430 ^ n2568 ;
  assign n4947 = n1644 | n3943 ;
  assign n4948 = n2078 | n4947 ;
  assign n4949 = n1221 | n1415 ;
  assign n4950 = ~n2852 & n4949 ;
  assign n4951 = n4950 ^ n2804 ^ 1'b0 ;
  assign n4952 = n1865 ^ n460 ^ 1'b0 ;
  assign n4953 = x5 & ~n4952 ;
  assign n4954 = n4953 ^ n3521 ^ 1'b0 ;
  assign n4955 = x103 & ~n4954 ;
  assign n4956 = n2055 ^ n1261 ^ 1'b0 ;
  assign n4957 = n736 | n4956 ;
  assign n4958 = n3935 | n4957 ;
  assign n4959 = n4958 ^ n4618 ^ 1'b0 ;
  assign n4960 = ( ~n1130 & n3186 ) | ( ~n1130 & n3855 ) | ( n3186 & n3855 ) ;
  assign n4961 = n3648 ^ n288 ^ 1'b0 ;
  assign n4962 = n1021 & ~n4281 ;
  assign n4963 = x127 & ~n3514 ;
  assign n4964 = n4963 ^ n3551 ^ 1'b0 ;
  assign n4965 = ~n3781 & n4964 ;
  assign n4966 = n2112 ^ n1330 ^ 1'b0 ;
  assign n4967 = n4965 | n4966 ;
  assign n4968 = n415 & n4967 ;
  assign n4969 = x120 & x166 ;
  assign n4970 = n4969 ^ n1675 ^ 1'b0 ;
  assign n4971 = n1540 | n3355 ;
  assign n4972 = ~n486 & n2534 ;
  assign n4973 = ~n895 & n4668 ;
  assign n4974 = ~n4972 & n4973 ;
  assign n4975 = n345 | n820 ;
  assign n4976 = n1688 | n4975 ;
  assign n4977 = n4976 ^ n1383 ^ 1'b0 ;
  assign n4978 = x230 & n4977 ;
  assign n4979 = ( n4797 & ~n4826 ) | ( n4797 & n4978 ) | ( ~n4826 & n4978 ) ;
  assign n4980 = n2460 & ~n3711 ;
  assign n4984 = ~n1806 & n3314 ;
  assign n4985 = n2769 & n4984 ;
  assign n4981 = ~n1435 & n1700 ;
  assign n4982 = n4981 ^ n2391 ^ 1'b0 ;
  assign n4983 = n2319 & ~n4982 ;
  assign n4986 = n4985 ^ n4983 ^ 1'b0 ;
  assign n4987 = n4032 ^ n3419 ^ 1'b0 ;
  assign n4988 = x151 & ~n4987 ;
  assign n4989 = n3507 & ~n4988 ;
  assign n4990 = n3637 ^ n1700 ^ 1'b0 ;
  assign n4991 = n602 & n4990 ;
  assign n4992 = n4063 ^ n1353 ^ 1'b0 ;
  assign n4993 = n3057 & ~n4992 ;
  assign n4995 = x73 & ~n3186 ;
  assign n4996 = n1415 & n4644 ;
  assign n4997 = n4996 ^ n1154 ^ 1'b0 ;
  assign n4998 = n4995 | n4997 ;
  assign n4999 = n4998 ^ n3366 ^ 1'b0 ;
  assign n4994 = n3356 & ~n4475 ;
  assign n5000 = n4999 ^ n4994 ^ 1'b0 ;
  assign n5001 = n3511 | n3877 ;
  assign n5002 = n5001 ^ n955 ^ 1'b0 ;
  assign n5003 = n265 & ~n573 ;
  assign n5004 = ~x223 & n5003 ;
  assign n5005 = n5004 ^ n2387 ^ 1'b0 ;
  assign n5006 = ( x21 & n493 ) | ( x21 & ~n5005 ) | ( n493 & ~n5005 ) ;
  assign n5007 = n2242 ^ x178 ^ 1'b0 ;
  assign n5008 = n2879 | n5007 ;
  assign n5009 = n647 & n1353 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = n5010 ^ n3756 ^ 1'b0 ;
  assign n5012 = n614 | n5011 ;
  assign n5013 = n1429 ^ x81 ^ 1'b0 ;
  assign n5014 = ~n1903 & n3028 ;
  assign n5015 = n3669 ^ n2241 ^ 1'b0 ;
  assign n5016 = n5015 ^ x239 ^ 1'b0 ;
  assign n5017 = n5016 ^ n2794 ^ 1'b0 ;
  assign n5018 = ~n2241 & n3945 ;
  assign n5019 = n4077 ^ n880 ^ 1'b0 ;
  assign n5020 = ~n2208 & n5019 ;
  assign n5021 = n1635 & ~n3953 ;
  assign n5022 = x229 & n1242 ;
  assign n5023 = n5022 ^ n2459 ^ 1'b0 ;
  assign n5024 = n1910 ^ n903 ^ 1'b0 ;
  assign n5025 = n3429 | n4695 ;
  assign n5026 = n1907 | n3552 ;
  assign n5027 = n1622 & ~n2201 ;
  assign n5028 = n2968 & ~n5027 ;
  assign n5029 = n5028 ^ n1347 ^ 1'b0 ;
  assign n5030 = n972 ^ n532 ^ 1'b0 ;
  assign n5031 = n5030 ^ n1976 ^ 1'b0 ;
  assign n5032 = n1399 & n1549 ;
  assign n5033 = ~n539 & n5032 ;
  assign n5034 = n5031 & n5033 ;
  assign n5035 = n637 ^ x20 ^ 1'b0 ;
  assign n5036 = ~n5034 & n5035 ;
  assign n5037 = n4671 ^ n862 ^ 1'b0 ;
  assign n5038 = x85 & ~n5037 ;
  assign n5039 = ~n3089 & n3902 ;
  assign n5040 = n5039 ^ n3059 ^ 1'b0 ;
  assign n5041 = n5038 & ~n5040 ;
  assign n5042 = n5041 ^ n3670 ^ 1'b0 ;
  assign n5043 = ~n3688 & n4157 ;
  assign n5044 = n3226 & ~n4804 ;
  assign n5045 = n5044 ^ n4263 ^ 1'b0 ;
  assign n5046 = n4794 ^ n2223 ^ 1'b0 ;
  assign n5047 = n5045 & n5046 ;
  assign n5048 = n1622 & ~n2270 ;
  assign n5049 = n409 & n1483 ;
  assign n5050 = ~n5048 & n5049 ;
  assign n5051 = n4641 & n4688 ;
  assign n5052 = n5050 & n5051 ;
  assign n5053 = x46 & ~n715 ;
  assign n5054 = n5053 ^ n2921 ^ 1'b0 ;
  assign n5055 = n3266 ^ n1512 ^ 1'b0 ;
  assign n5056 = n1405 | n5055 ;
  assign n5057 = n1572 & ~n5056 ;
  assign n5058 = n1356 ^ n746 ^ 1'b0 ;
  assign n5059 = n2287 & n5058 ;
  assign n5060 = n1112 & n5059 ;
  assign n5061 = n1828 | n5060 ;
  assign n5062 = ( n2539 & n5057 ) | ( n2539 & ~n5061 ) | ( n5057 & ~n5061 ) ;
  assign n5063 = n683 | n1369 ;
  assign n5064 = n5063 ^ n3862 ^ 1'b0 ;
  assign n5065 = ~n713 & n3255 ;
  assign n5066 = n5065 ^ n2916 ^ 1'b0 ;
  assign n5067 = n3858 ^ n320 ^ 1'b0 ;
  assign n5068 = n2768 | n3365 ;
  assign n5069 = n4350 ^ n3065 ^ n2124 ;
  assign n5070 = ~n2707 & n3054 ;
  assign n5071 = n1914 ^ n452 ^ 1'b0 ;
  assign n5072 = n4935 ^ n4384 ^ n3001 ;
  assign n5073 = n3462 ^ n2676 ^ 1'b0 ;
  assign n5074 = n4156 & n5073 ;
  assign n5075 = n4039 ^ n2824 ^ 1'b0 ;
  assign n5076 = n1643 & n5075 ;
  assign n5077 = x217 & n493 ;
  assign n5078 = n5077 ^ x118 ^ 1'b0 ;
  assign n5079 = n5076 & ~n5078 ;
  assign n5080 = n5079 ^ n552 ^ 1'b0 ;
  assign n5081 = ~n3187 & n5080 ;
  assign n5082 = n4806 ^ n2636 ^ 1'b0 ;
  assign n5083 = n3235 ^ n2819 ^ 1'b0 ;
  assign n5084 = x206 & ~n1925 ;
  assign n5085 = ~n5083 & n5084 ;
  assign n5086 = n4603 ^ n4580 ^ 1'b0 ;
  assign n5087 = ~n2676 & n5086 ;
  assign n5088 = n5087 ^ n3158 ^ 1'b0 ;
  assign n5089 = n2677 ^ n2303 ^ 1'b0 ;
  assign n5092 = x200 & x211 ;
  assign n5093 = n1108 & n5092 ;
  assign n5090 = n3694 ^ n978 ^ 1'b0 ;
  assign n5091 = n5090 ^ n1135 ^ n974 ;
  assign n5094 = n5093 ^ n5091 ^ 1'b0 ;
  assign n5095 = n3614 ^ n1112 ^ 1'b0 ;
  assign n5096 = n635 | n5095 ;
  assign n5097 = n1556 | n5096 ;
  assign n5098 = n5097 ^ n630 ^ 1'b0 ;
  assign n5099 = ~n1059 & n5098 ;
  assign n5100 = n1441 | n1447 ;
  assign n5101 = n1419 | n5100 ;
  assign n5102 = n4668 ^ n842 ^ 1'b0 ;
  assign n5103 = n5101 | n5102 ;
  assign n5104 = n1929 ^ n505 ^ 1'b0 ;
  assign n5105 = n2842 | n5104 ;
  assign n5106 = n472 ^ x103 ^ 1'b0 ;
  assign n5107 = n5105 & n5106 ;
  assign n5108 = n4035 ^ n3850 ^ 1'b0 ;
  assign n5109 = n2658 ^ n1160 ^ 1'b0 ;
  assign n5110 = n1971 & ~n5109 ;
  assign n5111 = n1054 & ~n3387 ;
  assign n5112 = n354 | n1703 ;
  assign n5113 = x187 & x217 ;
  assign n5114 = n4910 & n5113 ;
  assign n5115 = n2195 & ~n2515 ;
  assign n5116 = n4919 & n5115 ;
  assign n5117 = n2865 & ~n4276 ;
  assign n5118 = n5117 ^ n3679 ^ 1'b0 ;
  assign n5119 = n4851 ^ n2737 ^ 1'b0 ;
  assign n5120 = ~n380 & n438 ;
  assign n5121 = n1840 | n2798 ;
  assign n5122 = ~n3727 & n5121 ;
  assign n5124 = n1358 & ~n4888 ;
  assign n5123 = n2855 & ~n3091 ;
  assign n5125 = n5124 ^ n5123 ^ 1'b0 ;
  assign n5126 = n1160 & n4198 ;
  assign n5127 = n3588 ^ n1784 ^ 1'b0 ;
  assign n5128 = n1152 | n5127 ;
  assign n5129 = n3758 ^ n863 ^ 1'b0 ;
  assign n5131 = n540 & ~n1245 ;
  assign n5132 = ~n2376 & n5131 ;
  assign n5130 = n394 & n649 ;
  assign n5133 = n5132 ^ n5130 ^ 1'b0 ;
  assign n5134 = ~n3591 & n5133 ;
  assign n5135 = n1358 & n5134 ;
  assign n5136 = n2976 & ~n3144 ;
  assign n5137 = n4185 ^ n1976 ^ 1'b0 ;
  assign n5138 = n1450 ^ x196 ^ 1'b0 ;
  assign n5139 = n5138 ^ n2528 ^ 1'b0 ;
  assign n5140 = n1743 & ~n4743 ;
  assign n5141 = ~n663 & n5140 ;
  assign n5142 = ~n2098 & n5106 ;
  assign n5143 = ~n5141 & n5142 ;
  assign n5144 = n3257 ^ n594 ^ 1'b0 ;
  assign n5145 = n4334 & ~n4813 ;
  assign n5146 = n3278 ^ n2325 ^ 1'b0 ;
  assign n5147 = ~n2487 & n5146 ;
  assign n5148 = n4505 & n5147 ;
  assign n5149 = n3035 | n4540 ;
  assign n5150 = n5149 ^ n4627 ^ 1'b0 ;
  assign n5151 = n5059 ^ n1441 ^ 1'b0 ;
  assign n5152 = n1096 & n5151 ;
  assign n5154 = n1787 ^ x21 ^ 1'b0 ;
  assign n5153 = ~n840 & n1825 ;
  assign n5155 = n5154 ^ n5153 ^ 1'b0 ;
  assign n5156 = n4465 ^ n3828 ^ 1'b0 ;
  assign n5157 = n430 | n5156 ;
  assign n5158 = x218 | n3153 ;
  assign n5159 = n3294 | n5158 ;
  assign n5160 = n3986 & n5159 ;
  assign n5161 = n3349 & n5154 ;
  assign n5162 = ~x236 & n5161 ;
  assign n5163 = n5140 & ~n5162 ;
  assign n5164 = n1393 | n1514 ;
  assign n5165 = n966 & n5164 ;
  assign n5166 = ~n1614 & n5165 ;
  assign n5167 = n1866 ^ x41 ^ 1'b0 ;
  assign n5168 = n2521 & ~n5167 ;
  assign n5169 = ~n738 & n5168 ;
  assign n5170 = n4663 ^ n4319 ^ n709 ;
  assign n5171 = n4611 ^ n1723 ^ n929 ;
  assign n5172 = ~n2024 & n5171 ;
  assign n5173 = n5172 ^ n892 ^ 1'b0 ;
  assign n5174 = n2618 ^ n1267 ^ 1'b0 ;
  assign n5175 = n3855 & n5174 ;
  assign n5176 = n4290 & n4731 ;
  assign n5177 = ~n1326 & n3312 ;
  assign n5178 = n3601 & n5177 ;
  assign n5179 = ~n1252 & n5178 ;
  assign n5180 = n1850 & n2696 ;
  assign n5181 = ( n3554 & ~n5179 ) | ( n3554 & n5180 ) | ( ~n5179 & n5180 ) ;
  assign n5182 = n3005 ^ n1593 ^ 1'b0 ;
  assign n5183 = n2870 ^ x116 ^ 1'b0 ;
  assign n5184 = n5182 & ~n5183 ;
  assign n5185 = n4061 & n5184 ;
  assign n5186 = n4012 ^ n705 ^ 1'b0 ;
  assign n5187 = n1727 | n5186 ;
  assign n5188 = ~n1533 & n5187 ;
  assign n5189 = n317 & n3054 ;
  assign n5190 = n1522 & ~n4091 ;
  assign n5191 = n1964 ^ n1809 ^ 1'b0 ;
  assign n5192 = x151 & n4229 ;
  assign n5194 = n1784 | n3365 ;
  assign n5193 = n403 & ~n2447 ;
  assign n5195 = n5194 ^ n5193 ^ n4707 ;
  assign n5196 = n1672 ^ n724 ^ 1'b0 ;
  assign n5197 = n2223 & ~n3551 ;
  assign n5198 = n5197 ^ n2173 ^ 1'b0 ;
  assign n5199 = ~n3018 & n3524 ;
  assign n5200 = n892 | n5199 ;
  assign n5201 = n486 ^ x62 ^ 1'b0 ;
  assign n5202 = ~n1285 & n2263 ;
  assign n5203 = n1613 & n5202 ;
  assign n5204 = n1277 ^ n1214 ^ 1'b0 ;
  assign n5205 = ~n718 & n5204 ;
  assign n5206 = x204 & n5205 ;
  assign n5207 = n5203 & n5206 ;
  assign n5208 = n4263 ^ n1330 ^ 1'b0 ;
  assign n5209 = n5208 ^ n2640 ^ 1'b0 ;
  assign n5211 = n4244 ^ n1820 ^ n1663 ;
  assign n5210 = n3361 ^ n836 ^ 1'b0 ;
  assign n5212 = n5211 ^ n5210 ^ 1'b0 ;
  assign n5213 = n4484 | n5212 ;
  assign n5214 = x24 & x136 ;
  assign n5215 = ~n4888 & n5214 ;
  assign n5216 = n1822 & n3421 ;
  assign n5217 = n5215 & n5216 ;
  assign n5218 = ( x222 & n3678 ) | ( x222 & ~n5217 ) | ( n3678 & ~n5217 ) ;
  assign n5222 = n2920 ^ n2861 ^ n420 ;
  assign n5219 = n481 | n1690 ;
  assign n5220 = n288 | n5219 ;
  assign n5221 = x177 & n5220 ;
  assign n5223 = n5222 ^ n5221 ^ 1'b0 ;
  assign n5224 = ~n766 & n4122 ;
  assign n5225 = n5224 ^ n1698 ^ 1'b0 ;
  assign n5226 = ~n1488 & n5225 ;
  assign n5227 = ~n2591 & n5226 ;
  assign n5228 = n3869 ^ n1829 ^ 1'b0 ;
  assign n5229 = ~n1080 & n5228 ;
  assign n5230 = n1713 & n4244 ;
  assign n5231 = n5230 ^ n3746 ^ 1'b0 ;
  assign n5232 = n5231 ^ n1271 ^ 1'b0 ;
  assign n5233 = n3219 ^ n941 ^ n521 ;
  assign n5234 = n2597 ^ n771 ^ 1'b0 ;
  assign n5235 = n1463 & n5234 ;
  assign n5236 = ~n1158 & n5235 ;
  assign n5237 = ~n4502 & n5236 ;
  assign n5238 = n5233 & n5237 ;
  assign n5239 = ~x37 & n2203 ;
  assign n5240 = n5239 ^ n2741 ^ 1'b0 ;
  assign n5241 = n320 | n5240 ;
  assign n5242 = n5241 ^ n686 ^ 1'b0 ;
  assign n5243 = n3928 ^ n2812 ^ 1'b0 ;
  assign n5244 = n2135 & ~n5243 ;
  assign n5245 = ~n2024 & n3534 ;
  assign n5246 = ~n4671 & n5245 ;
  assign n5247 = n2011 & ~n2207 ;
  assign n5248 = ~x36 & n5247 ;
  assign n5249 = n2942 & ~n5248 ;
  assign n5250 = n5249 ^ n3124 ^ 1'b0 ;
  assign n5251 = n1745 | n5250 ;
  assign n5252 = n5251 ^ n3959 ^ 1'b0 ;
  assign n5253 = n488 & n2227 ;
  assign n5254 = n750 & ~n5253 ;
  assign n5255 = n5254 ^ n3669 ^ 1'b0 ;
  assign n5256 = n281 | n1623 ;
  assign n5257 = n5256 ^ n4257 ^ 1'b0 ;
  assign n5260 = n1970 & n1985 ;
  assign n5261 = n5260 ^ n651 ^ 1'b0 ;
  assign n5258 = n1684 & ~n1689 ;
  assign n5259 = n4271 & n5258 ;
  assign n5262 = n5261 ^ n5259 ^ n2013 ;
  assign n5263 = n341 & ~n2541 ;
  assign n5264 = n1358 & n3721 ;
  assign n5265 = n5264 ^ n4420 ^ 1'b0 ;
  assign n5266 = n1252 & n2715 ;
  assign n5267 = n2394 ^ x141 ^ 1'b0 ;
  assign n5268 = n649 & n5267 ;
  assign n5269 = n2606 & n5268 ;
  assign n5270 = ~n281 & n5269 ;
  assign n5271 = ~n5266 & n5270 ;
  assign n5272 = n5118 | n5271 ;
  assign n5273 = ~n430 & n1849 ;
  assign n5274 = n4930 ^ n2235 ^ 1'b0 ;
  assign n5275 = n1772 & ~n5274 ;
  assign n5276 = n996 & n5275 ;
  assign n5277 = ~n5273 & n5276 ;
  assign n5278 = n325 ^ x78 ^ 1'b0 ;
  assign n5279 = n5278 ^ n2575 ^ 1'b0 ;
  assign n5280 = ( ~n887 & n3856 ) | ( ~n887 & n5279 ) | ( n3856 & n5279 ) ;
  assign n5282 = ~n3961 & n4964 ;
  assign n5281 = ~n1305 & n2778 ;
  assign n5283 = n5282 ^ n5281 ^ 1'b0 ;
  assign n5284 = n5283 ^ n1693 ^ 1'b0 ;
  assign n5285 = n2153 & n4720 ;
  assign n5286 = ~n421 & n1541 ;
  assign n5287 = n2115 & n5286 ;
  assign n5288 = n3361 & ~n5287 ;
  assign n5289 = n1449 | n1644 ;
  assign n5290 = n1339 & ~n5289 ;
  assign n5291 = n5255 ^ n1174 ^ 1'b0 ;
  assign n5292 = n2855 & n5291 ;
  assign n5293 = n1739 | n1770 ;
  assign n5294 = x91 | n5293 ;
  assign n5295 = n3888 ^ n1809 ^ 1'b0 ;
  assign n5296 = n5294 & ~n5295 ;
  assign n5297 = ~n1415 & n5296 ;
  assign n5298 = n1864 & n5297 ;
  assign n5299 = x84 & ~n3465 ;
  assign n5300 = n4997 & n5299 ;
  assign n5301 = n3959 ^ n3160 ^ 1'b0 ;
  assign n5302 = x42 & ~n5301 ;
  assign n5303 = n5119 ^ n3908 ^ 1'b0 ;
  assign n5304 = n5275 ^ n1087 ^ 1'b0 ;
  assign n5305 = n1451 & ~n4205 ;
  assign n5306 = n3863 ^ n2322 ^ 1'b0 ;
  assign n5307 = n2675 & ~n5306 ;
  assign n5308 = n5307 ^ n3947 ^ n1654 ;
  assign n5309 = ~n4175 & n5308 ;
  assign n5310 = ~n320 & n5309 ;
  assign n5311 = n5310 ^ n967 ^ 1'b0 ;
  assign n5312 = n1738 & n4663 ;
  assign n5313 = n1961 ^ x50 ^ 1'b0 ;
  assign n5314 = n1442 & ~n5313 ;
  assign n5315 = n5314 ^ n1148 ^ 1'b0 ;
  assign n5316 = ~n2895 & n5315 ;
  assign n5317 = n5316 ^ n4880 ^ n1044 ;
  assign n5318 = x131 & x198 ;
  assign n5319 = ~x198 & n5318 ;
  assign n5320 = x230 & n5319 ;
  assign n5321 = n482 & ~n5320 ;
  assign n5322 = n5320 & n5321 ;
  assign n5323 = n1738 & ~n5322 ;
  assign n5324 = n5323 ^ n4639 ^ 1'b0 ;
  assign n5325 = n875 | n5324 ;
  assign n5326 = ~x11 & n452 ;
  assign n5327 = n1361 & ~n5326 ;
  assign n5328 = n5327 ^ x222 ^ 1'b0 ;
  assign n5329 = n3908 ^ n1777 ^ 1'b0 ;
  assign n5330 = n4882 & ~n5329 ;
  assign n5331 = n905 & n4367 ;
  assign n5332 = n5225 ^ n4570 ^ 1'b0 ;
  assign n5333 = x251 & ~n3618 ;
  assign n5334 = n5333 ^ n698 ^ 1'b0 ;
  assign n5335 = n5334 ^ n5166 ^ 1'b0 ;
  assign n5336 = n797 | n5335 ;
  assign n5337 = n2620 ^ n2062 ^ 1'b0 ;
  assign n5338 = n2011 & n2964 ;
  assign n5339 = n1160 & n3902 ;
  assign n5340 = n5339 ^ x176 ^ 1'b0 ;
  assign n5341 = n5045 & n5340 ;
  assign n5342 = n1854 ^ n445 ^ 1'b0 ;
  assign n5343 = n1058 & n5342 ;
  assign n5344 = ( n4242 & n5083 ) | ( n4242 & ~n5343 ) | ( n5083 & ~n5343 ) ;
  assign n5345 = n1442 ^ n320 ^ 1'b0 ;
  assign n5346 = x234 & ~n5345 ;
  assign n5347 = n1152 | n5346 ;
  assign n5348 = n2459 ^ n1635 ^ 1'b0 ;
  assign n5349 = n2352 ^ n2315 ^ 1'b0 ;
  assign n5350 = x221 & n5349 ;
  assign n5351 = n5343 ^ n3715 ^ 1'b0 ;
  assign n5352 = n5351 ^ n4319 ^ 1'b0 ;
  assign n5353 = n3973 | n5352 ;
  assign n5354 = n1409 ^ n965 ^ 1'b0 ;
  assign n5355 = n2093 ^ n1052 ^ 1'b0 ;
  assign n5356 = n5355 ^ n700 ^ 1'b0 ;
  assign n5357 = ~n1803 & n5356 ;
  assign n5358 = n4775 ^ n4507 ^ 1'b0 ;
  assign n5359 = n2723 ^ n1234 ^ 1'b0 ;
  assign n5360 = n3039 | n5359 ;
  assign n5361 = ~n2180 & n2518 ;
  assign n5362 = n5361 ^ n357 ^ 1'b0 ;
  assign n5363 = n5360 | n5362 ;
  assign n5364 = n4920 & n5363 ;
  assign n5365 = ~n672 & n4076 ;
  assign n5366 = n5365 ^ n2426 ^ 1'b0 ;
  assign n5367 = n2991 & ~n3822 ;
  assign n5368 = n5367 ^ n2099 ^ 1'b0 ;
  assign n5369 = ( ~n672 & n5246 ) | ( ~n672 & n5368 ) | ( n5246 & n5368 ) ;
  assign n5370 = ~x214 & n1217 ;
  assign n5371 = n675 & n5370 ;
  assign n5372 = n1028 & n5371 ;
  assign n5373 = n4684 ^ n2643 ^ 1'b0 ;
  assign n5374 = n1508 & n1903 ;
  assign n5375 = n4896 & n5374 ;
  assign n5376 = n5375 ^ n3148 ^ 1'b0 ;
  assign n5377 = n3784 | n5376 ;
  assign n5378 = n445 | n5377 ;
  assign n5379 = n5378 ^ n2624 ^ 1'b0 ;
  assign n5380 = n1037 & n2587 ;
  assign n5381 = n5380 ^ n5355 ^ 1'b0 ;
  assign n5382 = n1464 ^ n403 ^ 1'b0 ;
  assign n5383 = n5382 ^ n897 ^ 1'b0 ;
  assign n5384 = ~n285 & n5383 ;
  assign n5385 = n3472 ^ n963 ^ 1'b0 ;
  assign n5386 = n4919 & n5385 ;
  assign n5387 = n1879 ^ n698 ^ 1'b0 ;
  assign n5389 = n3740 ^ n1743 ^ 1'b0 ;
  assign n5388 = n528 & n3437 ;
  assign n5390 = n5389 ^ n5388 ^ 1'b0 ;
  assign n5391 = n5390 ^ n2517 ^ 1'b0 ;
  assign n5392 = ~x70 & n5391 ;
  assign n5393 = ( n803 & ~n905 ) | ( n803 & n2660 ) | ( ~n905 & n2660 ) ;
  assign n5394 = n320 & n2824 ;
  assign n5395 = n366 | n5394 ;
  assign n5396 = n5395 ^ n2001 ^ 1'b0 ;
  assign n5397 = n3385 | n4188 ;
  assign n5398 = n5397 ^ n4826 ^ 1'b0 ;
  assign n5399 = n5398 ^ n4677 ^ 1'b0 ;
  assign n5400 = n566 & ~n2370 ;
  assign n5401 = n1372 ^ n677 ^ 1'b0 ;
  assign n5402 = n2296 ^ n1473 ^ 1'b0 ;
  assign n5403 = n3270 & n5402 ;
  assign n5404 = ~n5401 & n5403 ;
  assign n5405 = n5404 ^ n4197 ^ 1'b0 ;
  assign n5406 = x60 ^ x26 ^ 1'b0 ;
  assign n5407 = x3 & n5406 ;
  assign n5408 = n1544 & n5407 ;
  assign n5409 = n1410 | n1896 ;
  assign n5410 = n2039 | n5409 ;
  assign n5411 = n3207 | n5410 ;
  assign n5412 = n5411 ^ n5056 ^ n2426 ;
  assign n5413 = n3874 & n4238 ;
  assign n5414 = n2190 ^ n1149 ^ 1'b0 ;
  assign n5415 = n5414 ^ x11 ^ 1'b0 ;
  assign n5416 = n2175 ^ n1455 ^ 1'b0 ;
  assign n5417 = n2629 & ~n5416 ;
  assign n5418 = n1085 & ~n5417 ;
  assign n5419 = x155 & n3433 ;
  assign n5420 = n399 & n4928 ;
  assign n5421 = n3593 ^ n1715 ^ 1'b0 ;
  assign n5422 = n4934 | n5421 ;
  assign n5423 = x2 | n2254 ;
  assign n5424 = n2420 & ~n2470 ;
  assign n5425 = ~n4333 & n5424 ;
  assign n5426 = ~n5205 & n5425 ;
  assign n5427 = n1846 & ~n3836 ;
  assign n5428 = n552 & ~n3520 ;
  assign n5429 = ~n5350 & n5428 ;
  assign n5430 = ~n2787 & n3179 ;
  assign n5431 = n5430 ^ n1822 ^ 1'b0 ;
  assign n5432 = ~n273 & n4128 ;
  assign n5433 = n5432 ^ x206 ^ 1'b0 ;
  assign n5434 = n4354 ^ n2315 ^ 1'b0 ;
  assign n5435 = n1724 & ~n5434 ;
  assign n5436 = n3530 ^ n409 ^ 1'b0 ;
  assign n5437 = n2134 & n5436 ;
  assign n5438 = n1266 & n5437 ;
  assign n5439 = ~n5435 & n5438 ;
  assign n5440 = n1426 & ~n3038 ;
  assign n5441 = n1792 ^ n1210 ^ 1'b0 ;
  assign n5442 = n5440 | n5441 ;
  assign n5443 = n5442 ^ n4758 ^ 1'b0 ;
  assign n5444 = ( n1847 & ~n1980 ) | ( n1847 & n2062 ) | ( ~n1980 & n2062 ) ;
  assign n5445 = ~n3880 & n5444 ;
  assign n5446 = n5445 ^ n1875 ^ 1'b0 ;
  assign n5447 = ~n4701 & n5446 ;
  assign n5448 = n4527 ^ n2733 ^ 1'b0 ;
  assign n5449 = x113 & n365 ;
  assign n5450 = n5449 ^ x11 ^ 1'b0 ;
  assign n5451 = n1683 ^ n1205 ^ 1'b0 ;
  assign n5452 = n2990 & n5451 ;
  assign n5453 = n3331 ^ n2630 ^ 1'b0 ;
  assign n5454 = n5452 & ~n5453 ;
  assign n5455 = n2012 & n5454 ;
  assign n5456 = n5450 & n5455 ;
  assign n5457 = n4368 ^ n924 ^ 1'b0 ;
  assign n5458 = ~n821 & n1341 ;
  assign n5459 = x30 & n4822 ;
  assign n5460 = n3780 & n5459 ;
  assign n5461 = n1361 & ~n3834 ;
  assign n5462 = n1875 & n5461 ;
  assign n5463 = n5462 ^ n3154 ^ 1'b0 ;
  assign n5464 = n5463 ^ n2124 ^ 1'b0 ;
  assign n5467 = n2569 ^ n1660 ^ x234 ;
  assign n5468 = ~n397 & n2131 ;
  assign n5469 = n5467 & n5468 ;
  assign n5470 = ~n1353 & n5469 ;
  assign n5471 = n1571 | n5470 ;
  assign n5465 = n394 ^ x190 ^ 1'b0 ;
  assign n5466 = ~x85 & n5465 ;
  assign n5472 = n5471 ^ n5466 ^ 1'b0 ;
  assign n5473 = n1914 & n2348 ;
  assign n5474 = n5039 ^ n1070 ^ 1'b0 ;
  assign n5475 = n5473 & ~n5474 ;
  assign n5476 = n445 & n1304 ;
  assign n5477 = n1464 & n1617 ;
  assign n5478 = n5477 ^ x68 ^ 1'b0 ;
  assign n5479 = n1736 & n5478 ;
  assign n5480 = n1018 & n1045 ;
  assign n5481 = ~x26 & n5480 ;
  assign n5482 = n5481 ^ n335 ^ 1'b0 ;
  assign n5483 = ~n810 & n5482 ;
  assign n5484 = ~n4497 & n5483 ;
  assign n5485 = ~n2944 & n3868 ;
  assign n5486 = n5485 ^ n263 ^ 1'b0 ;
  assign n5487 = n5486 ^ x98 ^ 1'b0 ;
  assign n5496 = n3263 ^ n1106 ^ n1066 ;
  assign n5497 = n1727 & n5496 ;
  assign n5498 = n5497 ^ n4666 ^ 1'b0 ;
  assign n5499 = n363 | n1568 ;
  assign n5500 = n5499 ^ x3 ^ 1'b0 ;
  assign n5501 = n2920 & ~n5500 ;
  assign n5502 = x237 & ~n5501 ;
  assign n5503 = n5502 ^ n1656 ^ 1'b0 ;
  assign n5504 = ( n2948 & n5498 ) | ( n2948 & ~n5503 ) | ( n5498 & ~n5503 ) ;
  assign n5493 = n1267 | n1272 ;
  assign n5490 = ( n815 & n840 ) | ( n815 & ~n1093 ) | ( n840 & ~n1093 ) ;
  assign n5491 = n2706 | n5490 ;
  assign n5492 = n1814 | n5491 ;
  assign n5494 = n5493 ^ n5492 ^ n2872 ;
  assign n5495 = n3484 & ~n5494 ;
  assign n5488 = n1877 & n5097 ;
  assign n5489 = n5488 ^ n3803 ^ 1'b0 ;
  assign n5505 = n5504 ^ n5495 ^ n5489 ;
  assign n5506 = n1841 ^ n1202 ^ 1'b0 ;
  assign n5507 = x89 | n5506 ;
  assign n5508 = n602 & ~n3828 ;
  assign n5509 = n357 | n1818 ;
  assign n5510 = n5509 ^ x33 ^ 1'b0 ;
  assign n5511 = n2910 ^ n2252 ^ 1'b0 ;
  assign n5512 = n1125 & ~n5511 ;
  assign n5513 = n4166 | n5505 ;
  assign n5514 = n5513 ^ n3509 ^ 1'b0 ;
  assign n5515 = n981 | n4440 ;
  assign n5516 = n3340 & ~n5515 ;
  assign n5517 = ~n2642 & n3481 ;
  assign n5518 = ~n3393 & n5517 ;
  assign n5519 = x38 | n954 ;
  assign n5520 = n5519 ^ n5330 ^ 1'b0 ;
  assign n5521 = n5518 | n5520 ;
  assign n5522 = ~x38 & n2158 ;
  assign n5523 = n5522 ^ n3507 ^ 1'b0 ;
  assign n5524 = x46 & ~n3707 ;
  assign n5525 = n5524 ^ n2394 ^ 1'b0 ;
  assign n5526 = n5525 ^ n3970 ^ 1'b0 ;
  assign n5527 = ~x103 & n5526 ;
  assign n5528 = n3891 | n4075 ;
  assign n5529 = n5527 | n5528 ;
  assign n5530 = n3890 ^ n3336 ^ 1'b0 ;
  assign n5531 = ~n2857 & n5530 ;
  assign n5532 = n4538 ^ n3720 ^ 1'b0 ;
  assign n5533 = n795 | n5532 ;
  assign n5534 = n5533 ^ n4855 ^ 1'b0 ;
  assign n5535 = n1451 ^ n669 ^ 1'b0 ;
  assign n5536 = ~n4390 & n5535 ;
  assign n5537 = ~n5535 & n5536 ;
  assign n5538 = n3622 & ~n4203 ;
  assign n5539 = n4203 & n5538 ;
  assign n5540 = x237 & n891 ;
  assign n5541 = n2998 & n5540 ;
  assign n5542 = ~n5540 & n5541 ;
  assign n5543 = n1417 | n5542 ;
  assign n5544 = n1417 & ~n5543 ;
  assign n5545 = n5539 | n5544 ;
  assign n5546 = n4673 & ~n5545 ;
  assign n5547 = n5537 & n5546 ;
  assign n5548 = n5510 | n5547 ;
  assign n5549 = n5548 ^ n1512 ^ 1'b0 ;
  assign n5550 = n4675 ^ n1438 ^ 1'b0 ;
  assign n5551 = n4261 & n5550 ;
  assign n5552 = n307 | n5057 ;
  assign n5553 = n3088 | n5085 ;
  assign n5554 = n4602 ^ x27 ^ 1'b0 ;
  assign n5555 = x210 & ~n5554 ;
  assign n5556 = n1680 ^ n1626 ^ 1'b0 ;
  assign n5557 = n2561 & n5556 ;
  assign n5558 = n1920 ^ n445 ^ 1'b0 ;
  assign n5559 = n2254 & n5558 ;
  assign n5560 = n2904 ^ n2037 ^ 1'b0 ;
  assign n5561 = n4686 ^ n1239 ^ 1'b0 ;
  assign n5562 = x189 & n5561 ;
  assign n5563 = n5562 ^ n3284 ^ 1'b0 ;
  assign n5564 = n3874 ^ n1877 ^ 1'b0 ;
  assign n5565 = ~n934 & n5278 ;
  assign n5566 = n5565 ^ n1512 ^ 1'b0 ;
  assign n5567 = n5566 ^ n2350 ^ 1'b0 ;
  assign n5568 = ~n1402 & n1413 ;
  assign n5569 = n5568 ^ n493 ^ 1'b0 ;
  assign n5570 = n5293 & ~n5569 ;
  assign n5571 = n3111 & n5570 ;
  assign n5576 = x65 & ~n3910 ;
  assign n5577 = n2037 & n5576 ;
  assign n5575 = n2333 | n4783 ;
  assign n5572 = n1661 ^ n1393 ^ 1'b0 ;
  assign n5573 = n583 & n5572 ;
  assign n5574 = n5573 ^ n2274 ^ 1'b0 ;
  assign n5578 = n5577 ^ n5575 ^ n5574 ;
  assign n5579 = n4763 ^ n2408 ^ 1'b0 ;
  assign n5580 = n3592 & ~n4862 ;
  assign n5581 = n4103 ^ n2232 ^ 1'b0 ;
  assign n5582 = ~n3114 & n5581 ;
  assign n5583 = n5582 ^ n4632 ^ 1'b0 ;
  assign n5584 = n1202 & ~n3729 ;
  assign n5585 = n5584 ^ x62 ^ 1'b0 ;
  assign n5586 = x177 & ~n5585 ;
  assign n5587 = n3647 ^ n2475 ^ 1'b0 ;
  assign n5588 = x69 & n625 ;
  assign n5589 = n5588 ^ n1146 ^ 1'b0 ;
  assign n5590 = ~n1255 & n5589 ;
  assign n5591 = n4731 ^ x130 ^ 1'b0 ;
  assign n5592 = ( n1351 & n3456 ) | ( n1351 & n5591 ) | ( n3456 & n5591 ) ;
  assign n5593 = n1421 | n5162 ;
  assign n5594 = ~n2165 & n5593 ;
  assign n5595 = n5594 ^ n5447 ^ 1'b0 ;
  assign n5596 = n360 ^ x190 ^ 1'b0 ;
  assign n5597 = x151 & ~n5596 ;
  assign n5598 = n1970 & ~n5597 ;
  assign n5599 = n5598 ^ n2966 ^ 1'b0 ;
  assign n5600 = n1042 & n5599 ;
  assign n5601 = n1925 ^ n1424 ^ x63 ;
  assign n5602 = ~n1188 & n5184 ;
  assign n5603 = ~x222 & n5602 ;
  assign n5604 = n4333 ^ n3616 ^ 1'b0 ;
  assign n5605 = n4097 ^ n3256 ^ 1'b0 ;
  assign n5606 = n1553 | n5605 ;
  assign n5607 = n1961 & n4773 ;
  assign n5608 = n3081 ^ n2085 ^ 1'b0 ;
  assign n5609 = n2508 ^ n1252 ^ 1'b0 ;
  assign n5610 = n1080 & ~n5609 ;
  assign n5611 = ~n894 & n5610 ;
  assign n5612 = ~n450 & n5611 ;
  assign n5613 = n2848 ^ n631 ^ n288 ;
  assign n5614 = x6 & n259 ;
  assign n5615 = ~n1736 & n5614 ;
  assign n5616 = n5615 ^ n3181 ^ 1'b0 ;
  assign n5617 = n3882 | n5616 ;
  assign n5618 = n5613 | n5617 ;
  assign n5619 = n4481 ^ n3628 ^ 1'b0 ;
  assign n5625 = ~x181 & n3634 ;
  assign n5621 = n510 & ~n1343 ;
  assign n5622 = n5621 ^ n4118 ^ 1'b0 ;
  assign n5623 = ~n4459 & n5622 ;
  assign n5624 = n5623 ^ n651 ^ 1'b0 ;
  assign n5620 = n3169 ^ n2762 ^ 1'b0 ;
  assign n5626 = n5625 ^ n5624 ^ n5620 ;
  assign n5627 = n4198 & n4336 ;
  assign n5628 = n644 ^ x219 ^ 1'b0 ;
  assign n5629 = n2415 & n5628 ;
  assign n5630 = ~n1728 & n5629 ;
  assign n5631 = n4804 & n5630 ;
  assign n5632 = n4705 ^ n2138 ^ 1'b0 ;
  assign n5633 = n3924 & ~n5632 ;
  assign n5634 = n2210 | n3221 ;
  assign n5635 = ~n1369 & n3074 ;
  assign n5636 = n1249 | n5635 ;
  assign n5637 = n3537 & n5636 ;
  assign n5638 = n5637 ^ n2524 ^ 1'b0 ;
  assign n5639 = n372 & ~n5638 ;
  assign n5640 = n2447 & ~n3681 ;
  assign n5641 = ~n2411 & n5640 ;
  assign n5642 = n5641 ^ n4109 ^ 1'b0 ;
  assign n5643 = n3207 & ~n5642 ;
  assign n5644 = n2575 ^ n663 ^ 1'b0 ;
  assign n5645 = n1240 & n5644 ;
  assign n5646 = ~n966 & n3979 ;
  assign n5647 = n1247 & n5646 ;
  assign n5648 = n963 & n5647 ;
  assign n5649 = n5645 & ~n5648 ;
  assign n5650 = ~n2279 & n5649 ;
  assign n5651 = n5458 ^ n1249 ^ n1223 ;
  assign n5652 = n5093 ^ n1393 ^ 1'b0 ;
  assign n5653 = n2336 & n5652 ;
  assign n5654 = n1192 | n5653 ;
  assign n5655 = ~n2278 & n3156 ;
  assign n5656 = n5655 ^ n3581 ^ 1'b0 ;
  assign n5657 = n1738 & n3833 ;
  assign n5658 = n2487 & n5657 ;
  assign n5659 = n1684 & ~n4484 ;
  assign n5660 = n2562 ^ n1983 ^ 1'b0 ;
  assign n5661 = n4720 ^ n1549 ^ 1'b0 ;
  assign n5662 = n5125 & n5661 ;
  assign n5663 = n2736 & n4177 ;
  assign n5664 = ~n2379 & n5663 ;
  assign n5665 = n653 | n1941 ;
  assign n5666 = x62 & n5665 ;
  assign n5667 = n5664 & n5666 ;
  assign n5668 = n3242 & n3573 ;
  assign n5669 = n5668 ^ n1546 ^ 1'b0 ;
  assign n5670 = n3925 ^ n2681 ^ x223 ;
  assign n5671 = n3729 & ~n5670 ;
  assign n5672 = n465 & n836 ;
  assign n5673 = n5294 & n5672 ;
  assign n5674 = n5673 ^ n472 ^ 1'b0 ;
  assign n5675 = n4417 & ~n5674 ;
  assign n5676 = n1818 ^ n1760 ^ 1'b0 ;
  assign n5677 = x25 & ~n1343 ;
  assign n5678 = n1339 & n5677 ;
  assign n5679 = n4613 ^ n1499 ^ 1'b0 ;
  assign n5680 = ~n614 & n4953 ;
  assign n5681 = n5679 & n5680 ;
  assign n5682 = ( ~n5351 & n5678 ) | ( ~n5351 & n5681 ) | ( n5678 & n5681 ) ;
  assign n5683 = n372 & ~n717 ;
  assign n5684 = n683 | n1212 ;
  assign n5685 = n703 | n5684 ;
  assign n5686 = ~n5683 & n5685 ;
  assign n5687 = ~n949 & n5686 ;
  assign n5688 = n5687 ^ n2191 ^ 1'b0 ;
  assign n5689 = n1112 & n2896 ;
  assign n5690 = n5689 ^ n2562 ^ 1'b0 ;
  assign n5691 = n5690 ^ n2557 ^ 1'b0 ;
  assign n5692 = n376 ^ x24 ^ 1'b0 ;
  assign n5693 = n3107 & ~n5692 ;
  assign n5694 = ~n4868 & n5693 ;
  assign n5695 = ~n3381 & n5694 ;
  assign n5696 = n4316 ^ n2228 ^ 1'b0 ;
  assign n5697 = n5696 ^ n1979 ^ 1'b0 ;
  assign n5698 = n5695 & n5697 ;
  assign n5699 = ~n1620 & n3499 ;
  assign n5700 = n5699 ^ n5372 ^ 1'b0 ;
  assign n5701 = n1125 ^ x50 ^ 1'b0 ;
  assign n5702 = n5701 ^ n1549 ^ 1'b0 ;
  assign n5703 = n743 | n1890 ;
  assign n5704 = ~x89 & n2159 ;
  assign n5705 = n5704 ^ n3342 ^ 1'b0 ;
  assign n5706 = n5703 & ~n5705 ;
  assign n5707 = n1661 & ~n4147 ;
  assign n5708 = n4236 ^ n3305 ^ 1'b0 ;
  assign n5709 = n3980 & n5708 ;
  assign n5710 = n5688 & n5709 ;
  assign n5711 = ~n5707 & n5710 ;
  assign n5712 = n1228 & ~n4172 ;
  assign n5713 = n2484 ^ n2157 ^ 1'b0 ;
  assign n5714 = n1941 & n5713 ;
  assign n5715 = n3099 | n5714 ;
  assign n5716 = n2597 & ~n3822 ;
  assign n5717 = n5716 ^ n4865 ^ 1'b0 ;
  assign n5718 = ~n3264 & n5717 ;
  assign n5719 = n4653 ^ n1354 ^ 1'b0 ;
  assign n5720 = ~n577 & n3203 ;
  assign n5721 = x254 | n4520 ;
  assign n5722 = n5721 ^ n3863 ^ 1'b0 ;
  assign n5723 = n1686 | n1701 ;
  assign n5724 = n5722 & n5723 ;
  assign n5725 = n5724 ^ n3267 ^ 1'b0 ;
  assign n5726 = n5720 & ~n5725 ;
  assign n5727 = n2920 ^ n923 ^ 1'b0 ;
  assign n5728 = x115 | n5727 ;
  assign n5729 = ( ~x183 & n1690 ) | ( ~x183 & n4483 ) | ( n1690 & n4483 ) ;
  assign n5730 = n4124 & n4177 ;
  assign n5732 = n2492 ^ n1549 ^ 1'b0 ;
  assign n5733 = n1931 & n5732 ;
  assign n5734 = n4065 ^ n2932 ^ 1'b0 ;
  assign n5735 = n5733 & n5734 ;
  assign n5736 = n5735 ^ n4177 ^ 1'b0 ;
  assign n5731 = n415 & ~n1620 ;
  assign n5737 = n5736 ^ n5731 ^ 1'b0 ;
  assign n5738 = n1667 ^ x35 ^ 1'b0 ;
  assign n5739 = n3468 | n5738 ;
  assign n5740 = n5739 ^ n4688 ^ 1'b0 ;
  assign n5741 = n1787 & ~n4475 ;
  assign n5742 = n5741 ^ n3360 ^ 1'b0 ;
  assign n5743 = ~n286 & n5540 ;
  assign n5744 = n5743 ^ x76 ^ 1'b0 ;
  assign n5745 = n884 & n5744 ;
  assign n5746 = n5745 ^ n4084 ^ 1'b0 ;
  assign n5747 = n5746 ^ x171 ^ 1'b0 ;
  assign n5748 = n5573 & ~n5747 ;
  assign n5749 = n4048 & n5748 ;
  assign n5750 = n5749 ^ x58 ^ 1'b0 ;
  assign n5751 = n1990 & n2187 ;
  assign n5752 = n3647 | n5751 ;
  assign n5753 = n4909 & ~n5752 ;
  assign n5754 = n5753 ^ n1743 ^ 1'b0 ;
  assign n5755 = x223 & n3993 ;
  assign n5756 = n3076 & n5646 ;
  assign n5757 = n5756 ^ n614 ^ 1'b0 ;
  assign n5758 = n5199 & n5757 ;
  assign n5759 = ( n992 & n2714 ) | ( n992 & n3799 ) | ( n2714 & n3799 ) ;
  assign n5760 = x132 & ~n875 ;
  assign n5761 = n5760 ^ n1297 ^ 1'b0 ;
  assign n5762 = n3216 ^ n1419 ^ 1'b0 ;
  assign n5763 = n734 & n3437 ;
  assign n5764 = ~n300 & n5763 ;
  assign n5765 = n5764 ^ n1510 ^ 1'b0 ;
  assign n5766 = n5765 ^ n3304 ^ 1'b0 ;
  assign n5767 = n3169 | n5766 ;
  assign n5768 = x69 | n651 ;
  assign n5769 = n2561 & n5414 ;
  assign n5770 = n5768 & n5769 ;
  assign n5771 = n2827 & ~n3636 ;
  assign n5773 = n1613 ^ n1354 ^ 1'b0 ;
  assign n5774 = ~n1883 & n5773 ;
  assign n5772 = n966 & ~n2704 ;
  assign n5775 = n5774 ^ n5772 ^ 1'b0 ;
  assign n5776 = n3345 ^ n1957 ^ 1'b0 ;
  assign n5777 = n5776 ^ n5568 ^ 1'b0 ;
  assign n5778 = n4787 & ~n5777 ;
  assign n5779 = n2164 & ~n5778 ;
  assign n5780 = ~n761 & n4926 ;
  assign n5781 = n5780 ^ n2709 ^ 1'b0 ;
  assign n5782 = ~n1316 & n5781 ;
  assign n5783 = n5782 ^ n4648 ^ 1'b0 ;
  assign n5784 = n522 | n691 ;
  assign n5785 = n2632 | n2700 ;
  assign n5786 = n5785 ^ n744 ^ 1'b0 ;
  assign n5787 = n4161 & n5786 ;
  assign n5788 = n5787 ^ n4251 ^ 1'b0 ;
  assign n5789 = n1907 | n5788 ;
  assign n5790 = n5789 ^ n2403 ^ 1'b0 ;
  assign n5791 = n1746 ^ x25 ^ 1'b0 ;
  assign n5792 = n5791 ^ n3082 ^ n2305 ;
  assign n5793 = n1236 & n3743 ;
  assign n5794 = ~n623 & n5793 ;
  assign n5795 = n5794 ^ n2760 ^ 1'b0 ;
  assign n5796 = n1571 ^ n1302 ^ 1'b0 ;
  assign n5797 = n1828 | n4484 ;
  assign n5798 = n5797 ^ n294 ^ 1'b0 ;
  assign n5799 = n1099 ^ x24 ^ 1'b0 ;
  assign n5800 = n4452 & n5346 ;
  assign n5801 = ~n5799 & n5800 ;
  assign n5802 = n2138 & ~n5801 ;
  assign n5803 = n744 & ~n1307 ;
  assign n5804 = n5803 ^ n1298 ^ 1'b0 ;
  assign n5805 = n5804 ^ n3759 ^ 1'b0 ;
  assign n5806 = n3240 & ~n5805 ;
  assign n5807 = ~x254 & n1038 ;
  assign n5808 = n5807 ^ n4801 ^ 1'b0 ;
  assign n5809 = n860 ^ n315 ^ 1'b0 ;
  assign n5810 = x219 & ~n1134 ;
  assign n5811 = ~n2852 & n5810 ;
  assign n5812 = n5811 ^ n1517 ^ 1'b0 ;
  assign n5816 = ~n3590 & n4701 ;
  assign n5817 = ~n4152 & n5816 ;
  assign n5813 = n701 | n1820 ;
  assign n5814 = n2879 & ~n5813 ;
  assign n5815 = n2271 | n5814 ;
  assign n5818 = n5817 ^ n5815 ^ 1'b0 ;
  assign n5819 = n1100 & ~n2358 ;
  assign n5820 = n994 & n4279 ;
  assign n5821 = ~n5819 & n5820 ;
  assign n5822 = n795 | n5217 ;
  assign n5823 = n5822 ^ n3766 ^ 1'b0 ;
  assign n5824 = ~n4168 & n4454 ;
  assign n5825 = n5823 & n5824 ;
  assign n5826 = n5825 ^ n5036 ^ 1'b0 ;
  assign n5827 = n5826 ^ n1158 ^ 1'b0 ;
  assign n5828 = ~n5821 & n5827 ;
  assign n5829 = n3353 | n4363 ;
  assign n5830 = n5829 ^ n2604 ^ 1'b0 ;
  assign n5831 = n2449 | n3750 ;
  assign n5832 = n5831 ^ n2425 ^ 1'b0 ;
  assign n5833 = n5832 ^ n1159 ^ 1'b0 ;
  assign n5834 = n2044 & n2046 ;
  assign n5835 = n600 & n5834 ;
  assign n5836 = n3957 ^ x239 ^ 1'b0 ;
  assign n5837 = ~x195 & n5836 ;
  assign n5838 = ~n2853 & n5837 ;
  assign n5839 = x204 & n5838 ;
  assign n5840 = ~n4172 & n5839 ;
  assign n5841 = n5835 | n5840 ;
  assign n5842 = n5841 ^ x101 ^ 1'b0 ;
  assign n5843 = n1875 & n5314 ;
  assign n5844 = n570 | n1339 ;
  assign n5845 = n1856 ^ n1128 ^ 1'b0 ;
  assign n5846 = ( ~n4115 & n4749 ) | ( ~n4115 & n5845 ) | ( n4749 & n5845 ) ;
  assign n5847 = x66 & ~n3189 ;
  assign n5848 = n5236 | n5847 ;
  assign n5849 = ( n1255 & n2312 ) | ( n1255 & ~n2328 ) | ( n2312 & ~n2328 ) ;
  assign n5850 = n1080 | n5849 ;
  assign n5851 = n5850 ^ n4541 ^ 1'b0 ;
  assign n5852 = n2599 & ~n4992 ;
  assign n5853 = ( ~n385 & n1942 ) | ( ~n385 & n3419 ) | ( n1942 & n3419 ) ;
  assign n5854 = n3746 & n5268 ;
  assign n5855 = n5854 ^ n1070 ^ 1'b0 ;
  assign n5856 = n366 & n5855 ;
  assign n5857 = ~n5853 & n5856 ;
  assign n5858 = n4116 ^ x229 ^ 1'b0 ;
  assign n5859 = ~n3759 & n5858 ;
  assign n5860 = n3736 | n4399 ;
  assign n5861 = n2811 ^ n1767 ^ x130 ;
  assign n5862 = n2065 & n5493 ;
  assign n5863 = ~n5690 & n5862 ;
  assign n5864 = n4370 & n5863 ;
  assign n5865 = ( n696 & n2293 ) | ( n696 & ~n2761 ) | ( n2293 & ~n2761 ) ;
  assign n5866 = x127 & ~n994 ;
  assign n5867 = n5865 & n5866 ;
  assign n5868 = n331 | n5867 ;
  assign n5869 = n3039 & ~n5868 ;
  assign n5870 = n5869 ^ n5136 ^ 1'b0 ;
  assign n5871 = n3998 | n4166 ;
  assign n5872 = n5871 ^ n3869 ^ 1'b0 ;
  assign n5873 = n2735 & ~n5129 ;
  assign n5874 = ~n4777 & n5873 ;
  assign n5875 = n4821 ^ n3060 ^ 1'b0 ;
  assign n5876 = x239 & n2431 ;
  assign n5877 = n669 | n5876 ;
  assign n5883 = n1165 | n2642 ;
  assign n5878 = n2367 & n3847 ;
  assign n5879 = ~n1085 & n5878 ;
  assign n5880 = ~n1738 & n2135 ;
  assign n5881 = n5880 ^ n3256 ^ 1'b0 ;
  assign n5882 = ~n5879 & n5881 ;
  assign n5884 = n5883 ^ n5882 ^ 1'b0 ;
  assign n5885 = n5032 & ~n5884 ;
  assign n5886 = n860 & n1014 ;
  assign n5887 = ~n269 & n5886 ;
  assign n5888 = ~n339 & n3943 ;
  assign n5889 = n1666 & n5888 ;
  assign n5890 = ~n2068 & n5889 ;
  assign n5891 = n1383 & ~n1474 ;
  assign n5892 = ~n1451 & n2207 ;
  assign n5893 = n387 & n1922 ;
  assign n5894 = n2909 & n5893 ;
  assign n5895 = ~n2991 & n5894 ;
  assign n5896 = n709 | n967 ;
  assign n5897 = n3304 & n5896 ;
  assign n5898 = n1268 ^ n1237 ^ 1'b0 ;
  assign n5899 = x208 & n1383 ;
  assign n5900 = n5899 ^ n842 ^ 1'b0 ;
  assign n5901 = n3751 ^ x158 ^ 1'b0 ;
  assign n5902 = n5900 & ~n5901 ;
  assign n5903 = n3715 | n3995 ;
  assign n5904 = n5902 & ~n5903 ;
  assign n5905 = x226 & ~n5819 ;
  assign n5906 = n2310 ^ n2079 ^ 1'b0 ;
  assign n5907 = n2820 & n5906 ;
  assign n5908 = n5907 ^ n5644 ^ 1'b0 ;
  assign n5909 = n1841 & ~n4743 ;
  assign n5910 = n766 | n1910 ;
  assign n5911 = n5909 | n5910 ;
  assign n5912 = n602 ^ n593 ^ 1'b0 ;
  assign n5913 = n2820 & n5912 ;
  assign n5914 = n5911 & ~n5913 ;
  assign n5915 = n4040 & n4562 ;
  assign n5916 = n3420 & n4777 ;
  assign n5917 = n2217 & n5916 ;
  assign n5918 = n1568 & n5917 ;
  assign n5919 = ~n3175 & n3878 ;
  assign n5920 = ~n832 & n5919 ;
  assign n5921 = x47 & x120 ;
  assign n5922 = n5920 & n5921 ;
  assign n5923 = n1896 ^ n528 ^ 1'b0 ;
  assign n5924 = n992 | n5923 ;
  assign n5925 = n4428 | n5924 ;
  assign n5926 = ~x151 & n3694 ;
  assign n5927 = n1261 ^ n669 ^ 1'b0 ;
  assign n5928 = n2841 ^ n2076 ^ 1'b0 ;
  assign n5929 = n5928 ^ x242 ^ 1'b0 ;
  assign n5930 = n3995 & ~n5929 ;
  assign n5931 = n5930 ^ n3286 ^ 1'b0 ;
  assign n5932 = n4982 ^ n1353 ^ 1'b0 ;
  assign n5933 = ~n2295 & n5932 ;
  assign n5934 = n3524 & n5933 ;
  assign n5935 = n5934 ^ n1727 ^ 1'b0 ;
  assign n5936 = n2024 ^ x65 ^ 1'b0 ;
  assign n5937 = n5692 | n5936 ;
  assign n5938 = ~x34 & n607 ;
  assign n5939 = n5938 ^ n4213 ^ 1'b0 ;
  assign n5940 = ~n5937 & n5939 ;
  assign n5941 = n1883 & n3356 ;
  assign n5942 = ~x65 & n5941 ;
  assign n5943 = n2187 & ~n4742 ;
  assign n5944 = ~n456 & n2879 ;
  assign n5945 = ~n3290 & n5944 ;
  assign n5946 = n4936 | n5945 ;
  assign n5947 = n5283 ^ x206 ^ 1'b0 ;
  assign n5948 = n5734 & n5947 ;
  assign n5949 = n2338 ^ n1859 ^ 1'b0 ;
  assign n5950 = ~n3790 & n5949 ;
  assign n5951 = n5950 ^ n4931 ^ 1'b0 ;
  assign n5952 = x169 & ~n5951 ;
  assign n5953 = n5952 ^ n1632 ^ 1'b0 ;
  assign n5954 = n1738 ^ x228 ^ 1'b0 ;
  assign n5955 = n4632 & n5954 ;
  assign n5956 = n2796 & n5955 ;
  assign n5957 = n4431 ^ n273 ^ 1'b0 ;
  assign n5958 = x179 & ~n2216 ;
  assign n5959 = n4613 ^ x203 ^ 1'b0 ;
  assign n5960 = ~n2470 & n2718 ;
  assign n5961 = n5960 ^ n3181 ^ 1'b0 ;
  assign n5962 = n3357 & n5961 ;
  assign n5963 = ~x84 & n5962 ;
  assign n5968 = n1285 ^ n1099 ^ n1081 ;
  assign n5967 = ~n1440 & n2392 ;
  assign n5969 = n5968 ^ n5967 ^ 1'b0 ;
  assign n5964 = n1320 ^ n1126 ^ 1'b0 ;
  assign n5965 = n5175 ^ n2085 ^ 1'b0 ;
  assign n5966 = ~n5964 & n5965 ;
  assign n5970 = n5969 ^ n5966 ^ 1'b0 ;
  assign n5971 = n880 ^ n821 ^ 1'b0 ;
  assign n5972 = ~n5826 & n5971 ;
  assign n5973 = n1849 ^ n1531 ^ x16 ;
  assign n5974 = n891 & ~n3200 ;
  assign n5975 = ~n545 & n3316 ;
  assign n5976 = ~n2328 & n5975 ;
  assign n5977 = n1600 & ~n4812 ;
  assign n5980 = n2590 ^ n2115 ^ 1'b0 ;
  assign n5981 = n5763 & ~n5980 ;
  assign n5982 = n5981 ^ n3798 ^ 1'b0 ;
  assign n5978 = n1614 ^ n1312 ^ 1'b0 ;
  assign n5979 = n1390 & n5978 ;
  assign n5983 = n5982 ^ n5979 ^ 1'b0 ;
  assign n5984 = n2312 & ~n2336 ;
  assign n5985 = n2395 & ~n2871 ;
  assign n5986 = n5054 ^ x191 ^ 1'b0 ;
  assign n5987 = ~n5985 & n5986 ;
  assign n5988 = n5984 & n5987 ;
  assign n5989 = n841 & ~n4889 ;
  assign n5990 = n2102 ^ n296 ^ x160 ;
  assign n5991 = n5990 ^ n2035 ^ 1'b0 ;
  assign n5992 = n4913 ^ n4203 ^ 1'b0 ;
  assign n5993 = n5991 & ~n5992 ;
  assign n5994 = n1890 | n2609 ;
  assign n5995 = n5994 ^ n2765 ^ 1'b0 ;
  assign n5996 = ~n2352 & n5995 ;
  assign n6002 = n3083 ^ n1618 ^ 1'b0 ;
  assign n5998 = x174 & n442 ;
  assign n5999 = n2177 & n2526 ;
  assign n6000 = n5998 & n5999 ;
  assign n5997 = x181 & ~n4568 ;
  assign n6001 = n6000 ^ n5997 ^ 1'b0 ;
  assign n6003 = n6002 ^ n6001 ^ 1'b0 ;
  assign n6004 = n3250 ^ x106 ^ 1'b0 ;
  assign n6005 = n4375 | n6004 ;
  assign n6006 = n1506 ^ n851 ^ 1'b0 ;
  assign n6007 = ~n472 & n6006 ;
  assign n6008 = n6007 ^ n343 ^ 1'b0 ;
  assign n6009 = ( x127 & n1522 ) | ( x127 & ~n3823 ) | ( n1522 & ~n3823 ) ;
  assign n6010 = ~n514 & n5819 ;
  assign n6013 = ~n920 & n2784 ;
  assign n6014 = n6013 ^ n2485 ^ 1'b0 ;
  assign n6015 = n5840 & n6014 ;
  assign n6011 = n4183 ^ n1648 ^ 1'b0 ;
  assign n6012 = n1832 & ~n6011 ;
  assign n6016 = n6015 ^ n6012 ^ 1'b0 ;
  assign n6017 = ~n6010 & n6016 ;
  assign n6018 = n5370 ^ n1732 ^ 1'b0 ;
  assign n6019 = n4755 ^ x227 ^ 1'b0 ;
  assign n6020 = n3577 ^ n493 ^ 1'b0 ;
  assign n6021 = n6020 ^ n3619 ^ 1'b0 ;
  assign n6022 = ~n6019 & n6021 ;
  assign n6023 = n4313 ^ n2639 ^ 1'b0 ;
  assign n6024 = n1865 | n6023 ;
  assign n6025 = n4113 | n6024 ;
  assign n6026 = n918 & n4041 ;
  assign n6027 = n281 | n1239 ;
  assign n6028 = n6027 ^ n2997 ^ 1'b0 ;
  assign n6029 = n6028 ^ n1256 ^ 1'b0 ;
  assign n6030 = n1741 | n6029 ;
  assign n6031 = n3715 & ~n6030 ;
  assign n6032 = n911 ^ x87 ^ 1'b0 ;
  assign n6033 = n1081 | n6032 ;
  assign n6034 = x216 & ~n503 ;
  assign n6035 = x17 & n6034 ;
  assign n6036 = n6035 ^ n2575 ^ 1'b0 ;
  assign n6037 = n956 | n6036 ;
  assign n6038 = n4764 | n6037 ;
  assign n6039 = n760 | n2873 ;
  assign n6040 = n392 | n6039 ;
  assign n6041 = n6040 ^ n3095 ^ 1'b0 ;
  assign n6042 = ~n3580 & n6041 ;
  assign n6043 = ~n2961 & n6042 ;
  assign n6044 = n2018 ^ x51 ^ 1'b0 ;
  assign n6045 = ~n4260 & n6044 ;
  assign n6046 = n2557 ^ n492 ^ 1'b0 ;
  assign n6047 = n4644 & n6046 ;
  assign n6048 = n6047 ^ n3495 ^ 1'b0 ;
  assign n6049 = n6045 & ~n6048 ;
  assign n6050 = n5555 ^ n3266 ^ n3175 ;
  assign n6051 = n305 & n5974 ;
  assign n6052 = ~n3621 & n4564 ;
  assign n6053 = n452 & n1831 ;
  assign n6054 = n1965 | n3407 ;
  assign n6055 = n3520 ^ n317 ^ 1'b0 ;
  assign n6056 = n2610 ^ n920 ^ 1'b0 ;
  assign n6057 = x22 & n2310 ;
  assign n6058 = n6056 & n6057 ;
  assign n6059 = n789 | n4671 ;
  assign n6060 = n6059 ^ n294 ^ 1'b0 ;
  assign n6061 = n500 & n3812 ;
  assign n6062 = n4920 ^ n4919 ^ n2968 ;
  assign n6063 = n6061 | n6062 ;
  assign n6064 = n6060 | n6063 ;
  assign n6065 = n3748 ^ n1939 ^ 1'b0 ;
  assign n6066 = n1736 & n6065 ;
  assign n6067 = ~n3562 & n6066 ;
  assign n6068 = n4437 & ~n5166 ;
  assign n6069 = n4520 | n6068 ;
  assign n6070 = n6069 ^ n4716 ^ 1'b0 ;
  assign n6071 = ( ~n726 & n1214 ) | ( ~n726 & n3321 ) | ( n1214 & n3321 ) ;
  assign n6072 = n1148 & n3562 ;
  assign n6073 = ~n6071 & n6072 ;
  assign n6074 = ~n4214 & n4999 ;
  assign n6075 = ( ~n1223 & n3940 ) | ( ~n1223 & n6074 ) | ( n3940 & n6074 ) ;
  assign n6076 = n3501 ^ n577 ^ 1'b0 ;
  assign n6077 = ~n2761 & n4354 ;
  assign n6078 = ~n6076 & n6077 ;
  assign n6079 = ~n992 & n2854 ;
  assign n6080 = n6079 ^ n5279 ^ 1'b0 ;
  assign n6081 = n2816 ^ n2249 ^ 1'b0 ;
  assign n6082 = n6081 ^ n2597 ^ 1'b0 ;
  assign n6083 = n6082 ^ n5390 ^ 1'b0 ;
  assign n6084 = n1361 ^ n963 ^ 1'b0 ;
  assign n6085 = ~n4314 & n6084 ;
  assign n6086 = x200 & n6085 ;
  assign n6087 = n6086 ^ n4865 ^ 1'b0 ;
  assign n6088 = n2185 ^ n1560 ^ 1'b0 ;
  assign n6089 = ~n2591 & n6088 ;
  assign n6090 = n2024 | n5583 ;
  assign n6091 = n6089 | n6090 ;
  assign n6092 = n4499 ^ n2474 ^ 1'b0 ;
  assign n6093 = n5990 & n6092 ;
  assign n6094 = n6093 ^ n5555 ^ 1'b0 ;
  assign n6095 = n2187 & ~n2195 ;
  assign n6096 = n5614 ^ n724 ^ 1'b0 ;
  assign n6097 = x23 | n3102 ;
  assign n6098 = n2429 & ~n5853 ;
  assign n6099 = n1347 ^ n376 ^ 1'b0 ;
  assign n6100 = x241 & ~n6099 ;
  assign n6101 = n3914 ^ n2642 ^ 1'b0 ;
  assign n6102 = n1710 | n6101 ;
  assign n6103 = n2546 | n3067 ;
  assign n6104 = n3252 & ~n6103 ;
  assign n6105 = n581 & n1765 ;
  assign n6106 = n6105 ^ n2142 ^ 1'b0 ;
  assign n6107 = n6106 ^ n1278 ^ 1'b0 ;
  assign n6108 = ~n1718 & n6107 ;
  assign n6109 = x195 & n6108 ;
  assign n6110 = ~n3675 & n6109 ;
  assign n6111 = ~n1327 & n3348 ;
  assign n6112 = n623 | n6111 ;
  assign n6113 = n5105 | n6112 ;
  assign n6114 = n3965 | n6113 ;
  assign n6115 = n2741 & ~n4952 ;
  assign n6116 = ~x130 & n6115 ;
  assign n6117 = n4384 ^ n598 ^ 1'b0 ;
  assign n6118 = n1776 | n4707 ;
  assign n6119 = n3057 & ~n5507 ;
  assign n6120 = x162 ^ x112 ^ 1'b0 ;
  assign n6121 = n944 & ~n6120 ;
  assign n6122 = n1111 & n6121 ;
  assign n6123 = n380 & n6122 ;
  assign n6124 = n2015 | n6123 ;
  assign n6125 = n6124 ^ n2093 ^ 1'b0 ;
  assign n6126 = n495 & n1380 ;
  assign n6127 = ~n587 & n6126 ;
  assign n6128 = n3438 | n6127 ;
  assign n6129 = n2140 | n5450 ;
  assign n6130 = n6128 | n6129 ;
  assign n6131 = n3480 & ~n6130 ;
  assign n6132 = n2657 | n5490 ;
  assign n6133 = n1697 & ~n6132 ;
  assign n6134 = ~n3735 & n6133 ;
  assign n6135 = x228 & ~n1324 ;
  assign n6136 = ~n2886 & n6135 ;
  assign n6137 = n5876 ^ n2076 ^ 1'b0 ;
  assign n6138 = n2314 & ~n6137 ;
  assign n6139 = n6138 ^ n2011 ^ 1'b0 ;
  assign n6140 = n1765 & n6139 ;
  assign n6141 = n5728 ^ n2384 ^ 1'b0 ;
  assign n6142 = n4398 & n6141 ;
  assign n6143 = n6142 ^ n3694 ^ 1'b0 ;
  assign n6145 = n1497 & n2438 ;
  assign n6144 = n2367 & n3720 ;
  assign n6146 = n6145 ^ n6144 ^ 1'b0 ;
  assign n6147 = ~n1124 & n2893 ;
  assign n6148 = n2235 ^ n1091 ^ 1'b0 ;
  assign n6149 = n6147 | n6148 ;
  assign n6150 = n6149 ^ n349 ^ 1'b0 ;
  assign n6151 = ~n5476 & n6150 ;
  assign n6152 = n698 | n4180 ;
  assign n6153 = x124 & n6152 ;
  assign n6154 = n6153 ^ n4720 ^ 1'b0 ;
  assign n6155 = n357 | n2949 ;
  assign n6156 = n5654 & ~n6155 ;
  assign n6157 = ~n959 & n1544 ;
  assign n6158 = n6157 ^ x86 ^ 1'b0 ;
  assign n6159 = ~n2022 & n2600 ;
  assign n6160 = ~n4313 & n6159 ;
  assign n6161 = n6160 ^ n1196 ^ 1'b0 ;
  assign n6162 = n780 & ~n3458 ;
  assign n6163 = n5622 & ~n6162 ;
  assign n6164 = ~n1358 & n6163 ;
  assign n6165 = x55 & n909 ;
  assign n6166 = n6165 ^ n1234 ^ 1'b0 ;
  assign n6167 = n1405 & ~n6166 ;
  assign n6168 = ~n481 & n6145 ;
  assign n6169 = ~n6167 & n6168 ;
  assign n6170 = ~n6164 & n6169 ;
  assign n6171 = n4310 ^ n956 ^ 1'b0 ;
  assign n6172 = n6032 & n6171 ;
  assign n6175 = n3052 ^ n1831 ^ 1'b0 ;
  assign n6176 = n1936 | n6175 ;
  assign n6177 = n2879 | n6176 ;
  assign n6178 = n6177 ^ n2812 ^ 1'b0 ;
  assign n6173 = n1959 ^ n1569 ^ 1'b0 ;
  assign n6174 = n6173 ^ n903 ^ 1'b0 ;
  assign n6179 = n6178 ^ n6174 ^ 1'b0 ;
  assign n6180 = ~n1071 & n2698 ;
  assign n6181 = n1602 & ~n1980 ;
  assign n6182 = n6181 ^ n1957 ^ 1'b0 ;
  assign n6183 = n4136 & n6182 ;
  assign n6184 = n6183 ^ n1031 ^ 1'b0 ;
  assign n6185 = n5344 ^ n5331 ^ 1'b0 ;
  assign n6186 = n6184 & ~n6185 ;
  assign n6187 = n526 & n1926 ;
  assign n6188 = n1883 | n2776 ;
  assign n6189 = n6188 ^ n5304 ^ 1'b0 ;
  assign n6190 = n1805 & ~n6189 ;
  assign n6191 = n5424 ^ n273 ^ 1'b0 ;
  assign n6192 = ( n3379 & ~n4268 ) | ( n3379 & n4338 ) | ( ~n4268 & n4338 ) ;
  assign n6193 = n6192 ^ n5167 ^ 1'b0 ;
  assign n6194 = n3736 ^ n3130 ^ 1'b0 ;
  assign n6195 = n6194 ^ n3045 ^ 1'b0 ;
  assign n6196 = n3800 & ~n5978 ;
  assign n6197 = n4516 ^ n1610 ^ 1'b0 ;
  assign n6198 = n505 | n6197 ;
  assign n6200 = n1490 | n2048 ;
  assign n6199 = n3123 ^ n801 ^ 1'b0 ;
  assign n6201 = n6200 ^ n6199 ^ 1'b0 ;
  assign n6202 = x33 & n6201 ;
  assign n6203 = n6202 ^ n1435 ^ 1'b0 ;
  assign n6207 = ~n666 & n787 ;
  assign n6208 = n6207 ^ n4115 ^ 1'b0 ;
  assign n6209 = ~n1564 & n6208 ;
  assign n6204 = n4997 ^ x228 ^ 1'b0 ;
  assign n6205 = n3571 | n6204 ;
  assign n6206 = n3939 | n6205 ;
  assign n6210 = n6209 ^ n6206 ^ 1'b0 ;
  assign n6211 = n1935 & n3419 ;
  assign n6212 = n6211 ^ x19 ^ 1'b0 ;
  assign n6213 = n966 | n6212 ;
  assign n6214 = n4087 ^ n3569 ^ 1'b0 ;
  assign n6215 = n1544 & ~n6214 ;
  assign n6216 = n6215 ^ n5152 ^ 1'b0 ;
  assign n6217 = n1866 & ~n6216 ;
  assign n6218 = n418 & n445 ;
  assign n6219 = n3001 & n6218 ;
  assign n6220 = n3773 & n6219 ;
  assign n6221 = n4276 & ~n6220 ;
  assign n6222 = n3910 & n6221 ;
  assign n6224 = n2585 & n3449 ;
  assign n6225 = n6224 ^ n1890 ^ 1'b0 ;
  assign n6226 = n1181 & n6225 ;
  assign n6227 = n3287 | n6226 ;
  assign n6228 = n5437 | n6227 ;
  assign n6223 = ~n3850 & n5392 ;
  assign n6229 = n6228 ^ n6223 ^ 1'b0 ;
  assign n6235 = ~n625 & n3467 ;
  assign n6236 = n6235 ^ n296 ^ 1'b0 ;
  assign n6237 = n4014 & ~n6236 ;
  assign n6238 = n6237 ^ n2782 ^ 1'b0 ;
  assign n6230 = x148 & ~n2637 ;
  assign n6231 = n6230 ^ n1047 ^ 1'b0 ;
  assign n6232 = x74 & ~n5776 ;
  assign n6233 = ~n2366 & n6232 ;
  assign n6234 = n6231 | n6233 ;
  assign n6239 = n6238 ^ n6234 ^ 1'b0 ;
  assign n6240 = n1888 & ~n2929 ;
  assign n6241 = n6240 ^ n1709 ^ 1'b0 ;
  assign n6242 = n2480 & n6241 ;
  assign n6243 = n6242 ^ n1594 ^ 1'b0 ;
  assign n6244 = n5756 | n6243 ;
  assign n6245 = n3614 & ~n6244 ;
  assign n6246 = x98 & ~n2870 ;
  assign n6247 = ~n2334 & n3186 ;
  assign n6248 = n2452 | n6247 ;
  assign n6249 = n6248 ^ n1014 ^ 1'b0 ;
  assign n6250 = n6246 & ~n6249 ;
  assign n6251 = n3206 & ~n4695 ;
  assign n6252 = ~n985 & n6251 ;
  assign n6253 = n979 ^ n946 ^ 1'b0 ;
  assign n6254 = n1629 & ~n4742 ;
  assign n6255 = ( n637 & ~n3204 ) | ( n637 & n4637 ) | ( ~n3204 & n4637 ) ;
  assign n6256 = ~n3593 & n6255 ;
  assign n6257 = n2613 ^ n2083 ^ n1546 ;
  assign n6258 = n4582 & ~n6257 ;
  assign n6259 = n4932 ^ n2293 ^ 1'b0 ;
  assign n6260 = n3995 & n5503 ;
  assign n6261 = ~n4857 & n6260 ;
  assign n6262 = n2587 | n3217 ;
  assign n6263 = n2331 & ~n6262 ;
  assign n6264 = n744 & ~n5937 ;
  assign n6265 = n5017 ^ n4307 ^ 1'b0 ;
  assign n6266 = n3984 & n6265 ;
  assign n6267 = n2183 & ~n3961 ;
  assign n6268 = n2164 & ~n3593 ;
  assign n6269 = n1099 | n5471 ;
  assign n6270 = n3556 | n6269 ;
  assign n6271 = n5225 ^ n4272 ^ 1'b0 ;
  assign n6272 = n6271 ^ n3902 ^ 1'b0 ;
  assign n6273 = n450 & n6272 ;
  assign n6274 = n620 & n3747 ;
  assign n6275 = n836 & ~n1450 ;
  assign n6276 = ~n2908 & n6275 ;
  assign n6277 = n1489 & ~n2715 ;
  assign n6278 = n3160 & n6277 ;
  assign n6279 = n3214 & n6278 ;
  assign n6280 = n2103 & ~n6279 ;
  assign n6281 = n5271 & n6280 ;
  assign n6282 = n595 & ~n740 ;
  assign n6283 = ~n928 & n6282 ;
  assign n6284 = n6283 ^ n2611 ^ 1'b0 ;
  assign n6285 = n791 & ~n6284 ;
  assign n6286 = n1639 & ~n6285 ;
  assign n6287 = n5076 ^ n4694 ^ x87 ;
  assign n6288 = n2175 & n2807 ;
  assign n6289 = n6288 ^ n2947 ^ 1'b0 ;
  assign n6290 = ~n770 & n6289 ;
  assign n6291 = ~n5317 & n6290 ;
  assign n6292 = ~n6287 & n6291 ;
  assign n6293 = n545 & ~n1529 ;
  assign n6294 = x169 & ~n6293 ;
  assign n6295 = ~n3361 & n6294 ;
  assign n6296 = n5781 & n6295 ;
  assign n6297 = n482 | n937 ;
  assign n6298 = n1720 ^ n1644 ^ 1'b0 ;
  assign n6299 = n3581 & ~n6298 ;
  assign n6300 = ~n5252 & n6299 ;
  assign n6301 = n2517 & ~n3134 ;
  assign n6302 = n6301 ^ n5943 ^ 1'b0 ;
  assign n6303 = n1746 & n5709 ;
  assign n6304 = n3365 ^ n1594 ^ 1'b0 ;
  assign n6305 = ~n4637 & n6304 ;
  assign n6306 = n3292 ^ n2399 ^ 1'b0 ;
  assign n6307 = n4720 & n6306 ;
  assign n6308 = n6307 ^ n621 ^ 1'b0 ;
  assign n6310 = x126 & n1905 ;
  assign n6311 = ~n1139 & n6310 ;
  assign n6309 = ~n901 & n3601 ;
  assign n6312 = n6311 ^ n6309 ^ 1'b0 ;
  assign n6313 = n1729 ^ n724 ^ 1'b0 ;
  assign n6314 = n5552 ^ x86 ^ 1'b0 ;
  assign n6315 = n6313 | n6314 ;
  assign n6316 = n1740 & n4047 ;
  assign n6317 = n6316 ^ n1729 ^ 1'b0 ;
  assign n6318 = n6317 ^ n1353 ^ 1'b0 ;
  assign n6319 = ~n1387 & n6318 ;
  assign n6320 = n1709 & ~n3043 ;
  assign n6321 = n6320 ^ x90 ^ 1'b0 ;
  assign n6322 = n6319 & ~n6321 ;
  assign n6323 = n4324 ^ n2786 ^ 1'b0 ;
  assign n6324 = ~n2247 & n6323 ;
  assign n6325 = n1996 & ~n3778 ;
  assign n6326 = n3986 ^ x61 ^ 1'b0 ;
  assign n6327 = n6326 ^ n2500 ^ n2395 ;
  assign n6328 = n6327 ^ n2050 ^ n1671 ;
  assign n6329 = n6325 & ~n6328 ;
  assign n6330 = n6329 ^ n3796 ^ 1'b0 ;
  assign n6331 = x157 | n4024 ;
  assign n6332 = n3123 ^ n2055 ^ 1'b0 ;
  assign n6333 = n1777 | n6332 ;
  assign n6334 = n5754 ^ n1093 ^ 1'b0 ;
  assign n6335 = n6243 | n6334 ;
  assign n6336 = n1387 ^ n681 ^ 1'b0 ;
  assign n6337 = n1596 & n6336 ;
  assign n6338 = n1165 & n6337 ;
  assign n6339 = n6338 ^ n4935 ^ 1'b0 ;
  assign n6340 = n4198 ^ n1793 ^ 1'b0 ;
  assign n6341 = ( ~n675 & n6339 ) | ( ~n675 & n6340 ) | ( n6339 & n6340 ) ;
  assign n6342 = ~n1976 & n2115 ;
  assign n6343 = n4569 & n6342 ;
  assign n6344 = n5492 ^ n5021 ^ 1'b0 ;
  assign n6345 = n4172 ^ n2778 ^ 1'b0 ;
  assign n6346 = n3397 & n6345 ;
  assign n6347 = n6346 ^ n2889 ^ 1'b0 ;
  assign n6348 = n904 | n6347 ;
  assign n6349 = n3790 ^ n1735 ^ 1'b0 ;
  assign n6350 = n5134 | n6349 ;
  assign n6351 = n6350 ^ n4734 ^ n3091 ;
  assign n6352 = n6351 ^ x17 ^ 1'b0 ;
  assign n6353 = ~n1785 & n6352 ;
  assign n6354 = n1643 ^ n958 ^ 1'b0 ;
  assign n6355 = ~x154 & n6354 ;
  assign n6356 = n3065 & n6355 ;
  assign n6357 = n3302 & n6356 ;
  assign n6358 = n6357 ^ n3830 ^ 1'b0 ;
  assign n6359 = n3054 & ~n6358 ;
  assign n6360 = n825 & n3175 ;
  assign n6361 = n2675 & n6360 ;
  assign n6362 = ~n1376 & n6361 ;
  assign n6363 = n566 & n5143 ;
  assign n6364 = ~n1951 & n3765 ;
  assign n6365 = ~n5139 & n6364 ;
  assign n6366 = ~n3451 & n5904 ;
  assign n6367 = n2103 & ~n4757 ;
  assign n6368 = n6367 ^ n493 ^ 1'b0 ;
  assign n6369 = n2505 ^ x1 ^ 1'b0 ;
  assign n6370 = ~n2720 & n6369 ;
  assign n6371 = ~n4579 & n6370 ;
  assign n6374 = n1727 & ~n2776 ;
  assign n6375 = n2906 & n6374 ;
  assign n6372 = n4049 ^ n2079 ^ 1'b0 ;
  assign n6373 = n6372 ^ n3928 ^ n490 ;
  assign n6376 = n6375 ^ n6373 ^ n552 ;
  assign n6377 = ~n5152 & n6376 ;
  assign n6378 = n6377 ^ n4718 ^ 1'b0 ;
  assign n6379 = x27 & n4160 ;
  assign n6380 = x145 ^ x90 ^ 1'b0 ;
  assign n6381 = n5457 & n6380 ;
  assign n6382 = n6381 ^ n3050 ^ 1'b0 ;
  assign n6383 = n5620 ^ n871 ^ 1'b0 ;
  assign n6384 = x34 & ~n3345 ;
  assign n6385 = n3223 & n6384 ;
  assign n6386 = n1903 ^ n1703 ^ 1'b0 ;
  assign n6387 = ~n6385 & n6386 ;
  assign n6388 = n1423 & n5164 ;
  assign n6389 = n6388 ^ n1548 ^ 1'b0 ;
  assign n6390 = n6389 ^ n4678 ^ 1'b0 ;
  assign n6391 = n6369 | n6390 ;
  assign n6392 = n816 & n2682 ;
  assign n6393 = n428 | n1683 ;
  assign n6394 = n6393 ^ n4158 ^ 1'b0 ;
  assign n6395 = ~n1988 & n6346 ;
  assign n6396 = ~n6394 & n6395 ;
  assign n6397 = n4238 ^ n3735 ^ 1'b0 ;
  assign n6398 = x178 & n6397 ;
  assign n6399 = n2072 & ~n3939 ;
  assign n6400 = n2387 & ~n4170 ;
  assign n6401 = n1249 & n6400 ;
  assign n6402 = n2001 & ~n5419 ;
  assign n6403 = ~n1167 & n4283 ;
  assign n6404 = n6403 ^ n1529 ^ 1'b0 ;
  assign n6405 = n2188 & ~n6404 ;
  assign n6406 = n3989 ^ n672 ^ 1'b0 ;
  assign n6407 = n1663 & n6406 ;
  assign n6408 = ~n5450 & n6407 ;
  assign n6409 = n645 | n5271 ;
  assign n6410 = n6409 ^ n5026 ^ 1'b0 ;
  assign n6411 = ~n1139 & n3073 ;
  assign n6412 = ~n666 & n6411 ;
  assign n6413 = n2340 ^ n1262 ^ 1'b0 ;
  assign n6414 = n934 ^ n663 ^ 1'b0 ;
  assign n6415 = n6414 ^ n1126 ^ 1'b0 ;
  assign n6416 = ~n4743 & n6415 ;
  assign n6417 = ~n5867 & n6416 ;
  assign n6418 = n6413 & n6417 ;
  assign n6419 = n5927 ^ n1141 ^ 1'b0 ;
  assign n6420 = n3773 ^ n795 ^ 1'b0 ;
  assign n6421 = n4026 ^ n3339 ^ 1'b0 ;
  assign n6422 = ~n2225 & n5692 ;
  assign n6423 = n399 & ~n3633 ;
  assign n6424 = n6423 ^ n3132 ^ 1'b0 ;
  assign n6425 = ~n6422 & n6424 ;
  assign n6426 = n3387 ^ n1451 ^ 1'b0 ;
  assign n6427 = n6425 & ~n6426 ;
  assign n6428 = ~n817 & n6427 ;
  assign n6429 = ~n1016 & n5076 ;
  assign n6430 = n4622 & n6429 ;
  assign n6431 = ~n2306 & n4586 ;
  assign n6432 = n3304 ^ x174 ^ 1'b0 ;
  assign n6433 = ~n3501 & n6432 ;
  assign n6434 = n2624 & n6433 ;
  assign n6435 = ~n2766 & n5110 ;
  assign n6436 = n2835 ^ x127 ^ 1'b0 ;
  assign n6437 = n2105 | n6436 ;
  assign n6438 = ~n2964 & n6437 ;
  assign n6439 = n1797 & n6438 ;
  assign n6440 = x231 & ~n2564 ;
  assign n6441 = n1601 & n2714 ;
  assign n6442 = x84 & n6441 ;
  assign n6443 = n6442 ^ n2232 ^ 1'b0 ;
  assign n6444 = n3678 & n6443 ;
  assign n6445 = n6444 ^ n3798 ^ 1'b0 ;
  assign n6446 = n6440 & ~n6445 ;
  assign n6449 = n3431 ^ n3137 ^ 1'b0 ;
  assign n6450 = n5845 & n6449 ;
  assign n6447 = n5120 ^ n4579 ^ 1'b0 ;
  assign n6448 = n3152 | n6447 ;
  assign n6451 = n6450 ^ n6448 ^ 1'b0 ;
  assign n6452 = n1620 ^ x116 ^ 1'b0 ;
  assign n6453 = n2712 & n6452 ;
  assign n6454 = n2463 & ~n5194 ;
  assign n6455 = n6454 ^ x254 ^ 1'b0 ;
  assign n6456 = x191 & n2624 ;
  assign n6457 = n1111 | n5525 ;
  assign n6458 = n6456 | n6457 ;
  assign n6459 = ~n2536 & n6458 ;
  assign n6460 = ~n6455 & n6459 ;
  assign n6461 = ~x168 & n6246 ;
  assign n6462 = n1845 ^ n1248 ^ 1'b0 ;
  assign n6463 = ~n1611 & n6462 ;
  assign n6464 = n2292 & n3759 ;
  assign n6465 = n6463 & ~n6464 ;
  assign n6466 = n6465 ^ n392 ^ 1'b0 ;
  assign n6467 = n6466 ^ n3834 ^ 1'b0 ;
  assign n6468 = ~n3993 & n6467 ;
  assign n6469 = n3466 ^ n921 ^ 1'b0 ;
  assign n6470 = n3144 & ~n6413 ;
  assign n6471 = n2895 & n6470 ;
  assign n6472 = n490 & ~n5004 ;
  assign n6473 = n440 & n6472 ;
  assign n6474 = n2684 & ~n6473 ;
  assign n6475 = n3472 & n6474 ;
  assign n6476 = n1783 ^ n1701 ^ 1'b0 ;
  assign n6477 = n5598 & ~n6476 ;
  assign n6478 = x115 & ~n2299 ;
  assign n6479 = n6478 ^ n884 ^ 1'b0 ;
  assign n6480 = ~n2343 & n2941 ;
  assign n6481 = n2720 | n3137 ;
  assign n6482 = n6480 | n6481 ;
  assign n6483 = n434 | n4002 ;
  assign n6484 = n3328 & ~n6483 ;
  assign n6486 = ~n4138 & n5358 ;
  assign n6485 = n559 & n5855 ;
  assign n6487 = n6486 ^ n6485 ^ 1'b0 ;
  assign n6488 = ~n905 & n5242 ;
  assign n6489 = ~n4904 & n6488 ;
  assign n6490 = n2725 & ~n4068 ;
  assign n6491 = n6489 & n6490 ;
  assign n6492 = ~n1126 & n3669 ;
  assign n6493 = n6492 ^ x59 ^ 1'b0 ;
  assign n6494 = n3328 ^ n1247 ^ 1'b0 ;
  assign n6495 = n1050 ^ n481 ^ 1'b0 ;
  assign n6496 = n779 & ~n6495 ;
  assign n6497 = n2867 & n6496 ;
  assign n6498 = n3115 & n6497 ;
  assign n6499 = n895 & ~n3784 ;
  assign n6500 = n1646 ^ n432 ^ 1'b0 ;
  assign n6501 = ~n2286 & n6167 ;
  assign n6502 = n6500 & n6501 ;
  assign n6503 = n3277 & n5110 ;
  assign n6504 = ~n4570 & n6503 ;
  assign n6505 = ~n4695 & n6504 ;
  assign n6506 = n1242 | n6320 ;
  assign n6507 = n6506 ^ n3845 ^ 1'b0 ;
  assign n6508 = x13 & n4256 ;
  assign n6509 = n6508 ^ x169 ^ 1'b0 ;
  assign n6510 = n956 | n5591 ;
  assign n6511 = n6097 | n6510 ;
  assign n6512 = n720 & n1829 ;
  assign n6513 = n6512 ^ x104 ^ 1'b0 ;
  assign n6514 = n3841 | n6513 ;
  assign n6515 = n6514 ^ n5588 ^ 1'b0 ;
  assign n6516 = n539 & ~n5166 ;
  assign n6517 = n6133 ^ n1453 ^ 1'b0 ;
  assign n6518 = n1642 & ~n1799 ;
  assign n6519 = ~n6203 & n6518 ;
  assign n6520 = n5164 ^ n399 ^ 1'b0 ;
  assign n6521 = ~n361 & n6520 ;
  assign n6522 = n2804 | n6521 ;
  assign n6524 = x180 & ~n2420 ;
  assign n6523 = n4397 ^ n300 ^ 1'b0 ;
  assign n6525 = n6524 ^ n6523 ^ 1'b0 ;
  assign n6526 = n5571 ^ x58 ^ 1'b0 ;
  assign n6527 = n4002 | n6526 ;
  assign n6528 = n1591 | n1974 ;
  assign n6529 = n5111 ^ n3709 ^ 1'b0 ;
  assign n6530 = n6298 | n6529 ;
  assign n6531 = n6530 ^ n434 ^ 1'b0 ;
  assign n6532 = n6531 ^ n3294 ^ 1'b0 ;
  assign n6533 = n5401 | n6502 ;
  assign n6534 = n6533 ^ n2997 ^ 1'b0 ;
  assign n6535 = n2008 & n6463 ;
  assign n6536 = ~n583 & n6535 ;
  assign n6537 = n6536 ^ n2378 ^ n2124 ;
  assign n6538 = n6537 ^ x188 ^ 1'b0 ;
  assign n6539 = ~n4166 & n6538 ;
  assign n6540 = n6539 ^ n2910 ^ 1'b0 ;
  assign n6541 = n720 & ~n1573 ;
  assign n6542 = n6541 ^ n3816 ^ 1'b0 ;
  assign n6543 = n4808 ^ n2397 ^ n1983 ;
  assign n6544 = n2827 & n4313 ;
  assign n6545 = n6544 ^ n3941 ^ 1'b0 ;
  assign n6546 = ~n6543 & n6545 ;
  assign n6547 = ~n3588 & n4289 ;
  assign n6548 = n6547 ^ n614 ^ 1'b0 ;
  assign n6549 = x87 & n6548 ;
  assign n6550 = n6549 ^ x186 ^ 1'b0 ;
  assign n6551 = n508 & n6253 ;
  assign n6552 = n1513 ^ n866 ^ 1'b0 ;
  assign n6553 = ~n2587 & n6552 ;
  assign n6554 = n2978 & n5061 ;
  assign n6555 = n2095 & n6554 ;
  assign n6556 = n3982 | n5942 ;
  assign n6557 = ( ~n955 & n1301 ) | ( ~n955 & n2480 ) | ( n1301 & n2480 ) ;
  assign n6558 = n4255 & n6557 ;
  assign n6559 = ~n1650 & n3248 ;
  assign n6560 = ~n550 & n6559 ;
  assign n6561 = n724 & n5733 ;
  assign n6562 = n6561 ^ n5781 ^ 1'b0 ;
  assign n6563 = n2011 & n4705 ;
  assign n6564 = ~n2183 & n6563 ;
  assign n6565 = n2244 & ~n6149 ;
  assign n6566 = n6565 ^ n1919 ^ 1'b0 ;
  assign n6567 = ~n1240 & n1554 ;
  assign n6568 = ~n1479 & n6567 ;
  assign n6569 = n2474 ^ n2109 ^ 1'b0 ;
  assign n6570 = n2449 | n6569 ;
  assign n6571 = ( n6566 & n6568 ) | ( n6566 & n6570 ) | ( n6568 & n6570 ) ;
  assign n6572 = n6571 ^ n432 ^ 1'b0 ;
  assign n6573 = n5090 | n6224 ;
  assign n6574 = ~n3842 & n6573 ;
  assign n6575 = n4066 | n6574 ;
  assign n6576 = n4421 | n6575 ;
  assign n6577 = n3068 ^ n1783 ^ 1'b0 ;
  assign n6578 = n3067 & n6577 ;
  assign n6579 = n2133 & ~n2455 ;
  assign n6580 = n6579 ^ n1350 ^ 1'b0 ;
  assign n6581 = ~n768 & n6580 ;
  assign n6582 = ~n1617 & n6581 ;
  assign n6583 = ~n2248 & n6582 ;
  assign n6584 = n597 & n2439 ;
  assign n6585 = ( n1544 & n2854 ) | ( n1544 & n6584 ) | ( n2854 & n6584 ) ;
  assign n6586 = n510 | n5355 ;
  assign n6587 = x21 | n1312 ;
  assign n6588 = n1438 & n1749 ;
  assign n6589 = n6588 ^ n3868 ^ 1'b0 ;
  assign n6590 = n6589 ^ n2812 ^ 1'b0 ;
  assign n6591 = ~n1505 & n6590 ;
  assign n6592 = n6584 & n6591 ;
  assign n6593 = n6587 & ~n6592 ;
  assign n6594 = x130 & ~n2849 ;
  assign n6595 = n3284 & n6594 ;
  assign n6596 = ~n6593 & n6595 ;
  assign n6597 = n6596 ^ n1328 ^ 1'b0 ;
  assign n6598 = n6586 & n6597 ;
  assign n6599 = n6598 ^ n3210 ^ 1'b0 ;
  assign n6600 = n538 & n812 ;
  assign n6601 = ~x16 & n6600 ;
  assign n6602 = n1271 | n1736 ;
  assign n6603 = n899 & n4449 ;
  assign n6611 = n5685 ^ n2623 ^ 1'b0 ;
  assign n6612 = n1808 & n6611 ;
  assign n6604 = n946 & n1286 ;
  assign n6605 = ~n1808 & n6604 ;
  assign n6607 = n2925 ^ n1611 ^ 1'b0 ;
  assign n6608 = n1633 | n6607 ;
  assign n6606 = x222 & n1961 ;
  assign n6609 = n6608 ^ n6606 ^ 1'b0 ;
  assign n6610 = ~n6605 & n6609 ;
  assign n6613 = n6612 ^ n6610 ^ 1'b0 ;
  assign n6614 = n2697 & n6613 ;
  assign n6617 = n490 | n2247 ;
  assign n6618 = n3545 & ~n6617 ;
  assign n6615 = n1553 | n5606 ;
  assign n6616 = n6615 ^ n2299 ^ 1'b0 ;
  assign n6619 = n6618 ^ n6616 ^ n6147 ;
  assign n6620 = n1517 ^ n318 ^ 1'b0 ;
  assign n6621 = n6620 ^ n1784 ^ 1'b0 ;
  assign n6622 = n6621 ^ n2861 ^ 1'b0 ;
  assign n6623 = n1974 | n6622 ;
  assign n6624 = n618 | n628 ;
  assign n6625 = n6624 ^ n2804 ^ 1'b0 ;
  assign n6626 = x127 | n6625 ;
  assign n6627 = n1675 & n1969 ;
  assign n6628 = n6627 ^ n1455 ^ 1'b0 ;
  assign n6629 = n6626 & ~n6628 ;
  assign n6630 = n465 | n2833 ;
  assign n6633 = n2704 & n2901 ;
  assign n6634 = n6192 & n6633 ;
  assign n6635 = n2682 & n6634 ;
  assign n6631 = n4545 ^ n351 ^ 1'b0 ;
  assign n6632 = ~n5490 & n6631 ;
  assign n6636 = n6635 ^ n6632 ^ 1'b0 ;
  assign n6637 = n1194 & ~n2467 ;
  assign n6638 = x200 & n1521 ;
  assign n6639 = n6638 ^ n918 ^ 1'b0 ;
  assign n6640 = n6639 ^ n4870 ^ 1'b0 ;
  assign n6641 = n6640 ^ n5586 ^ 1'b0 ;
  assign n6642 = n6637 & ~n6641 ;
  assign n6643 = x231 & n1788 ;
  assign n6644 = n6643 ^ n3043 ^ 1'b0 ;
  assign n6645 = n771 & n6342 ;
  assign n6646 = n6645 ^ n1973 ^ 1'b0 ;
  assign n6647 = n3960 ^ x191 ^ 1'b0 ;
  assign n6648 = n6647 ^ n1922 ^ 1'b0 ;
  assign n6649 = ~n6646 & n6648 ;
  assign n6650 = n1905 & ~n3234 ;
  assign n6651 = n6650 ^ n3705 ^ 1'b0 ;
  assign n6652 = n1952 & ~n6651 ;
  assign n6653 = n5136 & n6652 ;
  assign n6654 = ~n380 & n4652 ;
  assign n6655 = n6654 ^ n3768 ^ 1'b0 ;
  assign n6656 = n4812 | n6655 ;
  assign n6657 = n5357 & ~n6656 ;
  assign n6658 = n1299 ^ n286 ^ 1'b0 ;
  assign n6659 = x249 & ~n6658 ;
  assign n6660 = n1390 & ~n5642 ;
  assign n6661 = n4459 & n6660 ;
  assign n6662 = n1337 ^ n1172 ^ 1'b0 ;
  assign n6663 = n1825 | n3721 ;
  assign n6664 = n1479 & ~n6663 ;
  assign n6665 = n6664 ^ n3576 ^ 1'b0 ;
  assign n6666 = n3326 & n3368 ;
  assign n6667 = ~n3081 & n4721 ;
  assign n6668 = n971 & n4091 ;
  assign n6669 = n2097 & ~n4919 ;
  assign n6670 = ~n1047 & n6669 ;
  assign n6671 = n4638 | n6670 ;
  assign n6672 = n6671 ^ n5778 ^ 1'b0 ;
  assign n6674 = n2019 ^ x172 ^ 1'b0 ;
  assign n6673 = n4091 & n5573 ;
  assign n6675 = n6674 ^ n6673 ^ 1'b0 ;
  assign n6681 = n2416 ^ n836 ^ 1'b0 ;
  assign n6676 = n6165 ^ n3542 ^ 1'b0 ;
  assign n6677 = n2113 ^ n1914 ^ n573 ;
  assign n6678 = n6677 ^ n1732 ^ 1'b0 ;
  assign n6679 = n4268 & n6678 ;
  assign n6680 = n6676 & n6679 ;
  assign n6682 = n6681 ^ n6680 ^ 1'b0 ;
  assign n6685 = ~n2644 & n2720 ;
  assign n6683 = n644 & ~n4117 ;
  assign n6684 = n5817 & n6683 ;
  assign n6686 = n6685 ^ n6684 ^ 1'b0 ;
  assign n6687 = n288 & ~n3509 ;
  assign n6688 = ~n2536 & n2974 ;
  assign n6689 = n6688 ^ n1093 ^ 1'b0 ;
  assign n6690 = ~n2477 & n4638 ;
  assign n6691 = ~x213 & n6690 ;
  assign n6692 = n6691 ^ n929 ^ 1'b0 ;
  assign n6693 = ~n1660 & n6692 ;
  assign n6694 = ~n5047 & n6693 ;
  assign n6695 = n3489 ^ x171 ^ 1'b0 ;
  assign n6696 = x192 & ~n6695 ;
  assign n6697 = ~n1016 & n6696 ;
  assign n6698 = n6697 ^ n549 ^ 1'b0 ;
  assign n6699 = n1435 | n1623 ;
  assign n6700 = n6699 ^ n5390 ^ 1'b0 ;
  assign n6701 = n3000 | n4263 ;
  assign n6702 = n2371 & ~n6701 ;
  assign n6703 = n6702 ^ n5763 ^ 1'b0 ;
  assign n6704 = n2309 ^ n919 ^ 1'b0 ;
  assign n6705 = n855 & ~n1684 ;
  assign n6706 = ~n1639 & n6705 ;
  assign n6707 = n6704 | n6706 ;
  assign n6708 = n6412 ^ n681 ^ 1'b0 ;
  assign n6709 = ~n2289 & n5229 ;
  assign n6710 = ~n1877 & n6709 ;
  assign n6711 = n2187 ^ n1694 ^ 1'b0 ;
  assign n6712 = n446 & ~n6711 ;
  assign n6713 = n1164 & n2082 ;
  assign n6714 = n6713 ^ n2778 ^ 1'b0 ;
  assign n6715 = ~n2863 & n6679 ;
  assign n6716 = n1269 & n5598 ;
  assign n6717 = n4888 ^ n1488 ^ 1'b0 ;
  assign n6718 = n3187 ^ n426 ^ 1'b0 ;
  assign n6719 = n3862 & ~n6718 ;
  assign n6720 = n3146 ^ n1948 ^ 1'b0 ;
  assign n6721 = ~n1216 & n6720 ;
  assign n6722 = n3512 & ~n6721 ;
  assign n6723 = n3414 & n5171 ;
  assign n6724 = ~x65 & n6723 ;
  assign n6725 = n532 | n6724 ;
  assign n6726 = n6722 | n6725 ;
  assign n6727 = n761 & ~n6726 ;
  assign n6734 = n1694 | n2338 ;
  assign n6735 = n6734 ^ n4913 ^ 1'b0 ;
  assign n6736 = n994 & n2896 ;
  assign n6737 = n6735 | n6736 ;
  assign n6728 = n677 | n3043 ;
  assign n6729 = n3319 & ~n6728 ;
  assign n6730 = n647 & n2071 ;
  assign n6731 = n2336 & ~n6730 ;
  assign n6732 = n6731 ^ n2486 ^ 1'b0 ;
  assign n6733 = n6729 | n6732 ;
  assign n6738 = n6737 ^ n6733 ^ 1'b0 ;
  assign n6739 = ( ~n1614 & n2011 ) | ( ~n1614 & n2293 ) | ( n2011 & n2293 ) ;
  assign n6740 = n6739 ^ n450 ^ 1'b0 ;
  assign n6741 = ~n3576 & n6740 ;
  assign n6742 = ~n2949 & n6741 ;
  assign n6743 = n5323 ^ n3125 ^ 1'b0 ;
  assign n6744 = n6019 ^ n2857 ^ 1'b0 ;
  assign n6745 = n6744 ^ x126 ^ 1'b0 ;
  assign n6746 = n4190 & ~n6295 ;
  assign n6747 = n6746 ^ n4373 ^ 1'b0 ;
  assign n6748 = n3437 ^ n1840 ^ x112 ;
  assign n6749 = n1818 | n4862 ;
  assign n6750 = n844 | n6749 ;
  assign n6751 = ~n1539 & n2998 ;
  assign n6752 = n6751 ^ n3669 ^ 1'b0 ;
  assign n6753 = ~n2632 & n6752 ;
  assign n6754 = n1974 & n6753 ;
  assign n6755 = n6239 ^ n568 ^ 1'b0 ;
  assign n6756 = n2565 & ~n6755 ;
  assign n6757 = ~n3521 & n6756 ;
  assign n6758 = n3248 ^ n1449 ^ 1'b0 ;
  assign n6759 = n2129 & ~n6758 ;
  assign n6760 = n5849 ^ n1765 ^ 1'b0 ;
  assign n6761 = n6760 ^ x88 ^ 1'b0 ;
  assign n6762 = n538 & ~n784 ;
  assign n6763 = n6587 & n6762 ;
  assign n6764 = ( n1217 & ~n4865 ) | ( n1217 & n6763 ) | ( ~n4865 & n6763 ) ;
  assign n6765 = n3437 ^ n1419 ^ 1'b0 ;
  assign n6766 = n1021 | n6765 ;
  assign n6767 = n1073 & ~n6766 ;
  assign n6768 = n6767 ^ x146 ^ 1'b0 ;
  assign n6769 = ~n4006 & n6768 ;
  assign n6770 = n723 & ~n6386 ;
  assign n6771 = n6770 ^ n866 ^ 1'b0 ;
  assign n6772 = n3479 ^ n2606 ^ 1'b0 ;
  assign n6773 = n2420 ^ n2271 ^ 1'b0 ;
  assign n6774 = ~n3874 & n6773 ;
  assign n6775 = ~n6455 & n6774 ;
  assign n6776 = ~n2493 & n6775 ;
  assign n6777 = n6776 ^ n1832 ^ 1'b0 ;
  assign n6778 = n5958 ^ n2008 ^ 1'b0 ;
  assign n6779 = n6777 & ~n6778 ;
  assign n6780 = n6779 ^ n1635 ^ 1'b0 ;
  assign n6781 = ( ~n1314 & n1402 ) | ( ~n1314 & n1890 ) | ( n1402 & n1890 ) ;
  assign n6782 = n2035 ^ n894 ^ 1'b0 ;
  assign n6783 = n4914 | n5530 ;
  assign n6784 = n3496 ^ n1111 ^ 1'b0 ;
  assign n6785 = n6784 ^ n4334 ^ 1'b0 ;
  assign n6786 = n1429 | n3628 ;
  assign n6787 = n5100 | n6786 ;
  assign n6788 = n6787 ^ n3304 ^ 1'b0 ;
  assign n6789 = n1081 & ~n1939 ;
  assign n6790 = n6789 ^ n928 ^ 1'b0 ;
  assign n6791 = n4609 & n6790 ;
  assign n6792 = ~n1969 & n3009 ;
  assign n6793 = n3991 ^ n2885 ^ 1'b0 ;
  assign n6794 = n6792 & ~n6793 ;
  assign n6795 = n6791 | n6794 ;
  assign n6796 = n296 & ~n904 ;
  assign n6797 = n6796 ^ n669 ^ 1'b0 ;
  assign n6798 = ~n4449 & n6797 ;
  assign n6799 = ~n3322 & n6798 ;
  assign n6800 = ~n538 & n1916 ;
  assign n6801 = n3416 & n6800 ;
  assign n6802 = n5690 & ~n6801 ;
  assign n6803 = n6281 ^ x249 ^ 1'b0 ;
  assign n6804 = n365 | n2491 ;
  assign n6805 = n6804 ^ n1111 ^ 1'b0 ;
  assign n6806 = n1614 & ~n1783 ;
  assign n6807 = n6806 ^ x216 ^ 1'b0 ;
  assign n6808 = n2070 | n6807 ;
  assign n6809 = n6808 ^ n867 ^ 1'b0 ;
  assign n6810 = n4106 & n6809 ;
  assign n6811 = n913 & n6810 ;
  assign n6812 = n710 & n6744 ;
  assign n6813 = n1295 & n6812 ;
  assign n6814 = n4787 & ~n6813 ;
  assign n6815 = n6814 ^ n3908 ^ 1'b0 ;
  assign n6816 = n6815 ^ n5678 ^ 1'b0 ;
  assign n6817 = n3032 & ~n4118 ;
  assign n6818 = ~n3078 & n6817 ;
  assign n6819 = n6818 ^ n4979 ^ 1'b0 ;
  assign n6821 = n2772 ^ n1648 ^ n1111 ;
  assign n6820 = n5799 & ~n6623 ;
  assign n6822 = n6821 ^ n6820 ^ 1'b0 ;
  assign n6823 = n4868 ^ n4217 ^ 1'b0 ;
  assign n6824 = n5690 ^ n5617 ^ 1'b0 ;
  assign n6825 = n2075 & ~n6215 ;
  assign n6826 = n4409 ^ n1272 ^ x75 ;
  assign n6827 = n6608 & n6826 ;
  assign n6828 = n2048 & n6827 ;
  assign n6829 = ~n1692 & n6828 ;
  assign n6830 = n956 & n1098 ;
  assign n6831 = n876 ^ x31 ^ 1'b0 ;
  assign n6832 = n6830 & n6831 ;
  assign n6833 = n1834 | n6729 ;
  assign n6834 = n1872 & ~n6833 ;
  assign n6835 = n2276 & ~n6834 ;
  assign n6836 = n1195 & n6835 ;
  assign n6837 = n6832 & ~n6836 ;
  assign n6838 = n6837 ^ n4970 ^ 1'b0 ;
  assign n6839 = ~n4910 & n6551 ;
  assign n6840 = n6839 ^ n3816 ^ 1'b0 ;
  assign n6841 = n3436 ^ x111 ^ 1'b0 ;
  assign n6842 = n2219 | n6841 ;
  assign n6843 = n3153 | n4949 ;
  assign n6844 = ~n529 & n6843 ;
  assign n6845 = ~n2857 & n6844 ;
  assign n6846 = n5385 ^ x6 ^ 1'b0 ;
  assign n6847 = n2164 & n2593 ;
  assign n6848 = n1160 ^ x138 ^ 1'b0 ;
  assign n6849 = n6847 & n6848 ;
  assign n6853 = x150 & n2796 ;
  assign n6854 = n2427 & n6853 ;
  assign n6855 = n6310 ^ n5638 ^ 1'b0 ;
  assign n6856 = n6854 | n6855 ;
  assign n6851 = n776 | n4957 ;
  assign n6852 = n1557 | n6851 ;
  assign n6857 = n6856 ^ n6852 ^ 1'b0 ;
  assign n6850 = n2581 & ~n4054 ;
  assign n6858 = n6857 ^ n6850 ^ 1'b0 ;
  assign n6860 = n1658 | n1904 ;
  assign n6861 = n6034 | n6860 ;
  assign n6859 = n4615 ^ n3895 ^ x50 ;
  assign n6862 = n6861 ^ n6859 ^ 1'b0 ;
  assign n6863 = n5351 | n6862 ;
  assign n6864 = n6863 ^ n4079 ^ 1'b0 ;
  assign n6865 = n1912 & n6864 ;
  assign n6866 = n5581 ^ n2697 ^ n1234 ;
  assign n6867 = n2986 ^ n1083 ^ 1'b0 ;
  assign n6868 = n6866 & ~n6867 ;
  assign n6869 = n2581 ^ x182 ^ 1'b0 ;
  assign n6870 = n538 & n1572 ;
  assign n6871 = n4164 & n6870 ;
  assign n6872 = n6871 ^ x136 ^ 1'b0 ;
  assign n6873 = n6869 | n6872 ;
  assign n6874 = n6873 ^ n4933 ^ 1'b0 ;
  assign n6875 = n2129 & ~n5248 ;
  assign n6876 = n6875 ^ n5569 ^ 1'b0 ;
  assign n6877 = n1765 & n6876 ;
  assign n6878 = n1693 & n6877 ;
  assign n6879 = ~n3541 & n4461 ;
  assign n6880 = n4209 | n6879 ;
  assign n6881 = n6878 & ~n6880 ;
  assign n6882 = n4615 ^ n4307 ^ n497 ;
  assign n6883 = n6882 ^ n2141 ^ 1'b0 ;
  assign n6884 = n1792 & ~n2046 ;
  assign n6885 = n6715 | n6884 ;
  assign n6886 = n345 & ~n4787 ;
  assign n6887 = ~n6630 & n6886 ;
  assign n6888 = n6023 & n6887 ;
  assign n6890 = n1382 | n4083 ;
  assign n6891 = n4810 | n6890 ;
  assign n6889 = n798 & ~n1897 ;
  assign n6892 = n6891 ^ n6889 ^ n2973 ;
  assign n6893 = n6892 ^ x237 ^ 1'b0 ;
  assign n6894 = n633 & n1928 ;
  assign n6895 = ~n1829 & n6894 ;
  assign n6896 = ~n3386 & n5944 ;
  assign n6897 = n6895 & n6896 ;
  assign n6898 = n3239 & ~n6205 ;
  assign n6899 = n502 | n1677 ;
  assign n6900 = ~n1453 & n3810 ;
  assign n6901 = n3603 ^ n2470 ^ 1'b0 ;
  assign n6902 = ~n6900 & n6901 ;
  assign n6903 = n6902 ^ n570 ^ 1'b0 ;
  assign n6904 = n6409 ^ n6264 ^ 1'b0 ;
  assign n6911 = x197 & n337 ;
  assign n6912 = ~n337 & n6911 ;
  assign n6913 = n6912 ^ n320 ^ 1'b0 ;
  assign n6914 = n461 & n1018 ;
  assign n6915 = ~n1018 & n6914 ;
  assign n6916 = n648 & n6915 ;
  assign n6917 = x234 & n6916 ;
  assign n6918 = n1343 & n6917 ;
  assign n6919 = n325 | n6918 ;
  assign n6920 = n325 & ~n6919 ;
  assign n6921 = n6913 | n6920 ;
  assign n6922 = n6913 & ~n6921 ;
  assign n6923 = n6325 & n6922 ;
  assign n6906 = x202 & x253 ;
  assign n6907 = ~x253 & n6906 ;
  assign n6908 = x78 & ~n6907 ;
  assign n6909 = n6907 & n6908 ;
  assign n6910 = ~n1327 & n6909 ;
  assign n6905 = n3902 ^ n2164 ^ n1179 ;
  assign n6924 = n6923 ^ n6910 ^ n6905 ;
  assign n6926 = n4075 ^ n1492 ^ 1'b0 ;
  assign n6927 = x253 & ~n6926 ;
  assign n6925 = ~n2348 & n6311 ;
  assign n6928 = n6927 ^ n6925 ^ 1'b0 ;
  assign n6929 = n6928 ^ n1551 ^ 1'b0 ;
  assign n6930 = n1463 ^ n345 ^ 1'b0 ;
  assign n6931 = ~n2663 & n6930 ;
  assign n6932 = n6931 ^ n1354 ^ 1'b0 ;
  assign n6933 = n2644 ^ n2115 ^ 1'b0 ;
  assign n6934 = n6933 ^ x97 ^ 1'b0 ;
  assign n6935 = ~n1951 & n2333 ;
  assign n6936 = n3431 & n3694 ;
  assign n6937 = n2237 ^ n801 ^ 1'b0 ;
  assign n6938 = n5968 & n6937 ;
  assign n6939 = n6938 ^ n3008 ^ 1'b0 ;
  assign n6940 = n6936 & ~n6939 ;
  assign n6941 = n6271 ^ n1969 ^ 1'b0 ;
  assign n6942 = n2466 & n4797 ;
  assign n6943 = n6942 ^ n4888 ^ 1'b0 ;
  assign n6944 = n2658 & ~n6943 ;
  assign n6945 = n1646 ^ n259 ^ 1'b0 ;
  assign n6946 = n696 & ~n3479 ;
  assign n6947 = n4253 & n6946 ;
  assign n6948 = n6947 ^ n3813 ^ 1'b0 ;
  assign n6950 = ~n2939 & n5463 ;
  assign n6949 = x234 & n5445 ;
  assign n6951 = n6950 ^ n6949 ^ 1'b0 ;
  assign n6952 = n1172 ^ n415 ^ 1'b0 ;
  assign n6953 = n3656 | n6952 ;
  assign n6954 = ~n296 & n6953 ;
  assign n6955 = n6954 ^ n3947 ^ 1'b0 ;
  assign n6956 = ~n2061 & n6955 ;
  assign n6957 = n3561 ^ n1318 ^ 1'b0 ;
  assign n6958 = n3751 | n6957 ;
  assign n6959 = ~n3132 & n6798 ;
  assign n6960 = n6958 & n6959 ;
  assign n6961 = n959 & ~n1964 ;
  assign n6962 = n6961 ^ n339 ^ 1'b0 ;
  assign n6963 = n304 | n6962 ;
  assign n6964 = x252 & n3116 ;
  assign n6965 = n265 & n6964 ;
  assign n6966 = n6965 ^ n5143 ^ 1'b0 ;
  assign n6967 = n4096 & ~n5642 ;
  assign n6968 = ~n1049 & n3842 ;
  assign n6969 = ~n6967 & n6968 ;
  assign n6970 = n4461 ^ n4286 ^ 1'b0 ;
  assign n6971 = n3171 & ~n6970 ;
  assign n6972 = n6971 ^ n3376 ^ 1'b0 ;
  assign n6973 = n6972 ^ n5310 ^ 1'b0 ;
  assign n6974 = n1802 & ~n6973 ;
  assign n6975 = n4660 ^ n2013 ^ 1'b0 ;
  assign n6976 = n2652 & n6165 ;
  assign n6977 = ~n552 & n2900 ;
  assign n6978 = n766 & n923 ;
  assign n6979 = n6977 & n6978 ;
  assign n6980 = n6979 ^ n2062 ^ 1'b0 ;
  assign n6981 = n6976 & n6980 ;
  assign n6982 = n6981 ^ n6271 ^ 1'b0 ;
  assign n6983 = n1324 & n6982 ;
  assign n6984 = n354 & ~n1027 ;
  assign n6985 = n6984 ^ n1710 ^ 1'b0 ;
  assign n6986 = n354 & ~n6985 ;
  assign n6987 = n1974 & ~n6986 ;
  assign n6988 = n1021 & n6987 ;
  assign n6989 = n3569 ^ n968 ^ 1'b0 ;
  assign n6990 = n3999 ^ n2575 ^ n2303 ;
  assign n6991 = x246 & n6990 ;
  assign n6992 = n6863 & ~n6991 ;
  assign n6993 = n6989 & n6992 ;
  assign n6994 = n1065 & ~n6642 ;
  assign n6995 = ~n2179 & n3733 ;
  assign n6999 = n5205 ^ n2944 ^ 1'b0 ;
  assign n7000 = n6999 ^ n748 ^ 1'b0 ;
  assign n6996 = n4169 ^ n2274 ^ 1'b0 ;
  assign n6997 = ~n5968 & n6996 ;
  assign n6998 = n3448 | n6997 ;
  assign n7001 = n7000 ^ n6998 ^ 1'b0 ;
  assign n7002 = ~n6995 & n7001 ;
  assign n7003 = n897 | n5250 ;
  assign n7004 = n2164 & ~n3405 ;
  assign n7005 = n6040 & ~n7004 ;
  assign n7007 = ~n1873 & n5346 ;
  assign n7008 = n7007 ^ x88 ^ 1'b0 ;
  assign n7009 = n3294 & n7008 ;
  assign n7006 = x76 | n2900 ;
  assign n7010 = n7009 ^ n7006 ^ n633 ;
  assign n7011 = n1952 & ~n2737 ;
  assign n7012 = n2796 & n7011 ;
  assign n7013 = n1269 & n7012 ;
  assign n7014 = n2433 | n6702 ;
  assign n7015 = n1920 & n2633 ;
  assign n7016 = ~x226 & n1453 ;
  assign n7017 = ~n4767 & n6125 ;
  assign n7018 = n2351 ^ x105 ^ 1'b0 ;
  assign n7019 = n2893 & n7018 ;
  assign n7020 = n1258 & ~n7019 ;
  assign n7021 = n7020 ^ n5598 ^ n4456 ;
  assign n7022 = n1593 | n4532 ;
  assign n7023 = n7022 ^ n4261 ^ 1'b0 ;
  assign n7024 = n2515 | n4603 ;
  assign n7025 = n4191 & ~n6331 ;
  assign n7026 = x85 & ~n2740 ;
  assign n7027 = n5089 ^ n5045 ^ 1'b0 ;
  assign n7028 = ~n1064 & n7027 ;
  assign n7029 = n2990 & ~n3925 ;
  assign n7030 = n7029 ^ n2257 ^ 1'b0 ;
  assign n7031 = ~n1018 & n1512 ;
  assign n7032 = n6631 & n7031 ;
  assign n7033 = n6325 ^ n887 ^ 1'b0 ;
  assign n7034 = n2336 & ~n7033 ;
  assign n7035 = n7034 ^ n5079 ^ 1'b0 ;
  assign n7036 = n4065 | n7035 ;
  assign n7037 = ( x83 & n315 ) | ( x83 & ~n1111 ) | ( n315 & ~n1111 ) ;
  assign n7038 = n1249 & ~n5233 ;
  assign n7039 = n7038 ^ n5336 ^ 1'b0 ;
  assign n7040 = n6797 ^ n6677 ^ 1'b0 ;
  assign n7041 = x73 ^ x43 ^ 1'b0 ;
  assign n7042 = ~n1236 & n7041 ;
  assign n7043 = n803 & n7042 ;
  assign n7044 = ~n1447 & n7043 ;
  assign n7045 = n7044 ^ n1914 ^ 1'b0 ;
  assign n7046 = n3984 & n7045 ;
  assign n7047 = n6359 ^ n2011 ^ 1'b0 ;
  assign n7048 = n7047 ^ n4013 ^ 1'b0 ;
  assign n7049 = n7046 | n7048 ;
  assign n7050 = n4197 & n5555 ;
  assign n7051 = n4037 ^ n3891 ^ 1'b0 ;
  assign n7052 = n3212 | n6596 ;
  assign n7053 = n401 | n2172 ;
  assign n7054 = n7053 ^ n557 ^ 1'b0 ;
  assign n7055 = n7054 ^ n1291 ^ n820 ;
  assign n7056 = ~n1651 & n4027 ;
  assign n7057 = n5290 & n7056 ;
  assign n7058 = ~n987 & n4275 ;
  assign n7059 = n3008 & ~n7058 ;
  assign n7060 = n7059 ^ n761 ^ 1'b0 ;
  assign n7061 = n7060 ^ x108 ^ 1'b0 ;
  assign n7062 = n2394 | n3459 ;
  assign n7063 = n4605 ^ n1817 ^ 1'b0 ;
  assign n7064 = n6620 | n7063 ;
  assign n7065 = n6749 ^ n5864 ^ 1'b0 ;
  assign n7066 = ~n7064 & n7065 ;
  assign n7067 = n3031 & n5356 ;
  assign n7068 = ~n2624 & n7067 ;
  assign n7069 = n2627 ^ x195 ^ 1'b0 ;
  assign n7070 = n2803 ^ n2309 ^ 1'b0 ;
  assign n7071 = ~n988 & n5662 ;
  assign n7072 = n1188 & n7071 ;
  assign n7073 = n1739 | n3893 ;
  assign n7074 = n7073 ^ n1782 ^ 1'b0 ;
  assign n7075 = n673 ^ n347 ^ 1'b0 ;
  assign n7076 = x197 & n7075 ;
  assign n7077 = n7076 ^ n1249 ^ 1'b0 ;
  assign n7078 = n7077 ^ n2241 ^ 1'b0 ;
  assign n7079 = x167 & n7078 ;
  assign n7080 = n7079 ^ n667 ^ 1'b0 ;
  assign n7081 = n1856 & ~n7080 ;
  assign n7082 = n4067 & n7081 ;
  assign n7083 = n1527 & n7082 ;
  assign n7084 = x246 & ~n5093 ;
  assign n7085 = ~x246 & n7084 ;
  assign n7086 = n749 | n7085 ;
  assign n7087 = n7085 & ~n7086 ;
  assign n7088 = n318 & n1020 ;
  assign n7089 = ~n1020 & n7088 ;
  assign n7090 = n1906 & ~n7089 ;
  assign n7091 = n7087 & n7090 ;
  assign n7092 = ~n283 & n587 ;
  assign n7093 = n283 & n7092 ;
  assign n7094 = n7091 & ~n7093 ;
  assign n7095 = ~n7091 & n7094 ;
  assign n7096 = n7095 ^ n4502 ^ n3499 ;
  assign n7097 = n686 | n2555 ;
  assign n7098 = n7097 ^ n4377 ^ 1'b0 ;
  assign n7099 = n4787 & ~n5442 ;
  assign n7100 = n7098 & n7099 ;
  assign n7101 = x17 & ~n5521 ;
  assign n7102 = n3136 & n7101 ;
  assign n7103 = n1803 | n2902 ;
  assign n7104 = n5744 & n6325 ;
  assign n7105 = n440 & n7104 ;
  assign n7106 = n4625 | n7105 ;
  assign n7107 = n1535 & ~n7106 ;
  assign n7108 = n2807 ^ n1326 ^ x67 ;
  assign n7109 = n4361 ^ n4084 ^ 1'b0 ;
  assign n7110 = n415 & ~n1686 ;
  assign n7111 = n7109 & n7110 ;
  assign n7112 = n1360 & ~n5445 ;
  assign n7113 = n7112 ^ n4103 ^ 1'b0 ;
  assign n7114 = n6162 | n7113 ;
  assign n7115 = n7114 ^ n4177 ^ 1'b0 ;
  assign n7116 = n370 & n3454 ;
  assign n7117 = n7116 ^ n3721 ^ 1'b0 ;
  assign n7118 = ( n1539 & ~n7115 ) | ( n1539 & n7117 ) | ( ~n7115 & n7117 ) ;
  assign n7119 = n7118 ^ n5989 ^ 1'b0 ;
  assign n7120 = x132 & ~n7119 ;
  assign n7121 = ~n987 & n3636 ;
  assign n7122 = x184 & n2505 ;
  assign n7123 = n7122 ^ n1033 ^ 1'b0 ;
  assign n7124 = n7121 & ~n7123 ;
  assign n7125 = n5703 ^ n1977 ^ 1'b0 ;
  assign n7126 = ~n6271 & n7125 ;
  assign n7127 = n6290 ^ n1742 ^ 1'b0 ;
  assign n7128 = n7127 ^ n5396 ^ 1'b0 ;
  assign n7129 = n6700 | n7128 ;
  assign n7130 = n1390 ^ x221 ^ 1'b0 ;
  assign n7131 = n571 | n7130 ;
  assign n7132 = n4006 & ~n7131 ;
  assign n7133 = n1283 ^ n288 ^ 1'b0 ;
  assign n7134 = n3862 ^ n651 ^ 1'b0 ;
  assign n7135 = n5645 & ~n7134 ;
  assign n7136 = n2427 & ~n6194 ;
  assign n7137 = n7136 ^ n2190 ^ 1'b0 ;
  assign n7138 = n3003 & ~n5600 ;
  assign n7139 = n5004 | n5450 ;
  assign n7140 = n7138 & ~n7139 ;
  assign n7141 = n1369 | n7140 ;
  assign n7142 = n1621 | n7141 ;
  assign n7143 = n6635 ^ n4705 ^ 1'b0 ;
  assign n7144 = n7143 ^ n5384 ^ n3532 ;
  assign n7145 = x152 & ~n1739 ;
  assign n7146 = n7145 ^ x140 ^ 1'b0 ;
  assign n7147 = n4352 & ~n7146 ;
  assign n7148 = n7147 ^ x114 ^ 1'b0 ;
  assign n7149 = n7144 & ~n7148 ;
  assign n7150 = n3373 & ~n3392 ;
  assign n7151 = n7150 ^ n5495 ^ 1'b0 ;
  assign n7152 = n4822 & n6203 ;
  assign n7153 = n7152 ^ n1490 ^ 1'b0 ;
  assign n7154 = n7151 & n7153 ;
  assign n7155 = ~n376 & n2686 ;
  assign n7156 = n2576 ^ n1223 ^ x222 ;
  assign n7157 = n1535 | n7156 ;
  assign n7158 = n7155 & ~n7157 ;
  assign n7159 = n1480 | n6970 ;
  assign n7160 = n1832 | n7159 ;
  assign n7161 = ~n2076 & n4647 ;
  assign n7162 = n5493 ^ n1606 ^ 1'b0 ;
  assign n7164 = ~n1810 & n2466 ;
  assign n7165 = n7164 ^ n4515 ^ 1'b0 ;
  assign n7166 = n7165 ^ n3985 ^ 1'b0 ;
  assign n7167 = n7166 ^ n3152 ^ 1'b0 ;
  assign n7168 = n5665 & n7167 ;
  assign n7163 = n1424 & ~n1546 ;
  assign n7169 = n7168 ^ n7163 ^ 1'b0 ;
  assign n7170 = n6869 ^ n3524 ^ 1'b0 ;
  assign n7171 = n5588 ^ n5150 ^ 1'b0 ;
  assign n7172 = n4161 ^ n4031 ^ 1'b0 ;
  assign n7173 = n2615 ^ x47 ^ 1'b0 ;
  assign n7174 = n4024 ^ n2869 ^ 1'b0 ;
  assign n7175 = n1335 | n4068 ;
  assign n7176 = n7175 ^ n5071 ^ 1'b0 ;
  assign n7177 = n7174 & ~n7176 ;
  assign n7178 = n3420 ^ n347 ^ 1'b0 ;
  assign n7179 = ~n2476 & n7178 ;
  assign n7180 = x222 & n4310 ;
  assign n7181 = n5443 & n7180 ;
  assign n7182 = n4812 | n5179 ;
  assign n7183 = n2475 | n7182 ;
  assign n7184 = x227 & ~n533 ;
  assign n7185 = ~n1601 & n7184 ;
  assign n7186 = n5334 & n5961 ;
  assign n7187 = n7185 & n7186 ;
  assign n7188 = n7183 & ~n7187 ;
  assign n7189 = n7181 & n7188 ;
  assign n7190 = n6019 ^ n3043 ^ 1'b0 ;
  assign n7191 = n1301 & ~n7190 ;
  assign n7192 = n7191 ^ n3910 ^ 1'b0 ;
  assign n7193 = n1093 & n7192 ;
  assign n7194 = n318 | n7193 ;
  assign n7196 = x47 & n1325 ;
  assign n7195 = n562 | n1741 ;
  assign n7197 = n7196 ^ n7195 ^ 1'b0 ;
  assign n7198 = n7197 ^ n724 ^ 1'b0 ;
  assign n7199 = n2356 & ~n7198 ;
  assign n7200 = n4502 & ~n6195 ;
  assign n7201 = ~n1883 & n4498 ;
  assign n7202 = n956 & n7201 ;
  assign n7203 = n6484 | n7202 ;
  assign n7204 = n7203 ^ n3304 ^ 1'b0 ;
  assign n7205 = x234 & ~n4495 ;
  assign n7206 = n672 & n7205 ;
  assign n7207 = n5032 & n7206 ;
  assign n7208 = ~n628 & n2055 ;
  assign n7209 = x212 & n872 ;
  assign n7210 = ~n3144 & n7209 ;
  assign n7211 = n7210 ^ n3163 ^ 1'b0 ;
  assign n7212 = n2052 ^ n1039 ^ 1'b0 ;
  assign n7213 = ~n5759 & n7212 ;
  assign n7214 = n7213 ^ n1974 ^ 1'b0 ;
  assign n7215 = n7214 ^ n2750 ^ n1368 ;
  assign n7216 = n3043 & ~n5920 ;
  assign n7217 = n3386 ^ n1777 ^ 1'b0 ;
  assign n7218 = n553 & n2904 ;
  assign n7219 = n7218 ^ n1905 ^ n415 ;
  assign n7220 = ~n7217 & n7219 ;
  assign n7221 = n7220 ^ n7026 ^ 1'b0 ;
  assign n7222 = n6001 | n6735 ;
  assign n7223 = n7222 ^ n458 ^ 1'b0 ;
  assign n7227 = n6999 ^ n1970 ^ n1318 ;
  assign n7228 = n3571 | n7227 ;
  assign n7224 = n6892 ^ n3971 ^ 1'b0 ;
  assign n7225 = x207 & n7224 ;
  assign n7226 = ~n795 & n7225 ;
  assign n7229 = n7228 ^ n7226 ^ 1'b0 ;
  assign n7230 = n2762 | n5635 ;
  assign n7231 = x213 & ~n1149 ;
  assign n7232 = n7231 ^ n1332 ^ 1'b0 ;
  assign n7233 = ~n3339 & n7232 ;
  assign n7234 = n7230 & n7233 ;
  assign n7235 = n4389 & ~n7234 ;
  assign n7236 = n7235 ^ n807 ^ 1'b0 ;
  assign n7237 = n3599 ^ n2080 ^ 1'b0 ;
  assign n7238 = n3226 ^ x208 ^ 1'b0 ;
  assign n7239 = x80 & n7238 ;
  assign n7240 = n1073 & ~n1632 ;
  assign n7241 = ~n7239 & n7240 ;
  assign n7242 = n972 | n1805 ;
  assign n7243 = x151 | n7242 ;
  assign n7244 = n7243 ^ n5793 ^ 1'b0 ;
  assign n7247 = n2544 ^ n1391 ^ 1'b0 ;
  assign n7248 = n7247 ^ n5484 ^ 1'b0 ;
  assign n7245 = ~n637 & n6830 ;
  assign n7246 = n7245 ^ n1566 ^ 1'b0 ;
  assign n7249 = n7248 ^ n7246 ^ 1'b0 ;
  assign n7250 = ~n3703 & n7249 ;
  assign n7251 = ~n2910 & n7250 ;
  assign n7252 = n3856 ^ n505 ^ 1'b0 ;
  assign n7253 = n3158 | n7252 ;
  assign n7254 = n4867 ^ n891 ^ 1'b0 ;
  assign n7255 = n1749 & ~n7254 ;
  assign n7256 = n781 & n7255 ;
  assign n7257 = n2772 ^ n2634 ^ 1'b0 ;
  assign n7258 = ~n1999 & n4779 ;
  assign n7259 = n1593 | n3381 ;
  assign n7260 = x100 & ~n6214 ;
  assign n7261 = ~n5427 & n7260 ;
  assign n7262 = n6998 ^ x174 ^ 1'b0 ;
  assign n7263 = n2379 | n4340 ;
  assign n7264 = n7263 ^ n3528 ^ 1'b0 ;
  assign n7265 = n793 & ~n1805 ;
  assign n7266 = x200 & n1099 ;
  assign n7267 = n978 & ~n7266 ;
  assign n7268 = n7267 ^ n2087 ^ 1'b0 ;
  assign n7269 = ~n6742 & n7096 ;
  assign n7270 = n6229 & ~n7269 ;
  assign n7271 = x76 & ~n6891 ;
  assign n7272 = ~x130 & n2393 ;
  assign n7273 = n564 & n2819 ;
  assign n7274 = ~n7272 & n7273 ;
  assign n7275 = n7274 ^ n1703 ^ 1'b0 ;
  assign n7278 = n6483 ^ n3328 ^ 1'b0 ;
  assign n7277 = n302 | n3197 ;
  assign n7279 = n7278 ^ n7277 ^ 1'b0 ;
  assign n7276 = ~n498 & n6060 ;
  assign n7280 = n7279 ^ n7276 ^ 1'b0 ;
  assign n7281 = n1223 ^ x32 ^ 1'b0 ;
  assign n7282 = n288 & ~n7281 ;
  assign n7283 = n1468 & n6541 ;
  assign n7284 = ~n7282 & n7283 ;
  assign n7285 = n6511 ^ n2673 ^ 1'b0 ;
  assign n7286 = n5283 ^ n1320 ^ 1'b0 ;
  assign n7287 = n5651 & ~n7286 ;
  assign n7288 = n7287 ^ n5290 ^ n3651 ;
  assign n7289 = n7288 ^ n360 ^ 1'b0 ;
  assign n7290 = n1105 & ~n7289 ;
  assign n7291 = x63 | n1083 ;
  assign n7292 = n579 & ~n6663 ;
  assign n7293 = ~n7291 & n7292 ;
  assign n7294 = n828 | n3880 ;
  assign n7295 = n7293 & ~n7294 ;
  assign n7296 = n6702 ^ n3573 ^ 1'b0 ;
  assign n7297 = n3139 | n5134 ;
  assign n7298 = n509 & ~n7297 ;
  assign n7299 = n5476 & ~n7298 ;
  assign n7300 = ~x253 & n1226 ;
  assign n7301 = n1720 | n4347 ;
  assign n7302 = n7300 & n7301 ;
  assign n7303 = ~n3648 & n7302 ;
  assign n7304 = n5277 | n5433 ;
  assign n7305 = n7304 ^ n5752 ^ 1'b0 ;
  assign n7306 = ~x134 & n2129 ;
  assign n7307 = n5484 | n7306 ;
  assign n7308 = x98 | n7307 ;
  assign n7309 = n820 | n3405 ;
  assign n7310 = ~n4386 & n7309 ;
  assign n7311 = n790 | n7310 ;
  assign n7312 = n7311 ^ x174 ^ 1'b0 ;
  assign n7313 = ~n6751 & n7312 ;
  assign n7314 = ~n5060 & n7313 ;
  assign n7315 = n725 & ~n2266 ;
  assign n7316 = n2811 & n7315 ;
  assign n7317 = n5042 | n7316 ;
  assign n7318 = n1487 & n5235 ;
  assign n7319 = ~n4026 & n7318 ;
  assign n7320 = n4815 | n6246 ;
  assign n7321 = n3219 ^ n724 ^ 1'b0 ;
  assign n7322 = n1675 ^ n1606 ^ 1'b0 ;
  assign n7323 = n4255 | n7322 ;
  assign n7324 = n5450 | n7323 ;
  assign n7325 = n7324 ^ x126 ^ 1'b0 ;
  assign n7326 = n2384 | n7325 ;
  assign n7327 = ~n7321 & n7326 ;
  assign n7328 = n892 | n7327 ;
  assign n7329 = n508 | n7328 ;
  assign n7330 = n1539 & n1807 ;
  assign n7331 = n7330 ^ x88 ^ 1'b0 ;
  assign n7332 = n1599 ^ n1379 ^ 1'b0 ;
  assign n7333 = x167 & ~n7332 ;
  assign n7334 = n7333 ^ n3868 ^ 1'b0 ;
  assign n7335 = n1427 | n7334 ;
  assign n7336 = ~n4423 & n6241 ;
  assign n7337 = n7336 ^ n649 ^ 1'b0 ;
  assign n7338 = n4358 | n7337 ;
  assign n7339 = n2153 ^ n313 ^ 1'b0 ;
  assign n7340 = n7339 ^ n1419 ^ n1038 ;
  assign n7341 = n1843 & n1949 ;
  assign n7342 = n2358 & n4671 ;
  assign n7343 = n7342 ^ n672 ^ 1'b0 ;
  assign n7344 = n2227 ^ n1378 ^ 1'b0 ;
  assign n7345 = ~n2191 & n7344 ;
  assign n7346 = n4333 ^ x11 ^ 1'b0 ;
  assign n7347 = n2711 | n7346 ;
  assign n7348 = n5913 ^ n1829 ^ 1'b0 ;
  assign n7349 = ~n7347 & n7348 ;
  assign n7350 = n7345 & ~n7349 ;
  assign n7351 = n1293 | n2266 ;
  assign n7352 = n7351 ^ n1832 ^ 1'b0 ;
  assign n7353 = n7352 ^ n3159 ^ n1896 ;
  assign n7354 = n6737 & ~n7121 ;
  assign n7355 = n4065 & n7354 ;
  assign n7356 = x145 & n2148 ;
  assign n7357 = n7356 ^ n707 ^ 1'b0 ;
  assign n7358 = n6866 | n7357 ;
  assign n7359 = n833 & n4873 ;
  assign n7360 = ~n672 & n1992 ;
  assign n7361 = n7360 ^ n2261 ^ 1'b0 ;
  assign n7362 = n7361 ^ n5350 ^ 1'b0 ;
  assign n7363 = n4644 & n5940 ;
  assign n7364 = n7363 ^ n3850 ^ 1'b0 ;
  assign n7365 = ~n438 & n7364 ;
  assign n7366 = n1903 | n3524 ;
  assign n7367 = n3107 ^ n1260 ^ n1188 ;
  assign n7368 = n2730 & n6065 ;
  assign n7369 = n4903 & n6610 ;
  assign n7370 = ~n5266 & n7369 ;
  assign n7371 = n7368 & n7370 ;
  assign n7372 = ~x216 & n7371 ;
  assign n7373 = n5015 & n6065 ;
  assign n7374 = n3047 & n5462 ;
  assign n7375 = n2503 | n5311 ;
  assign n7376 = n7374 & ~n7375 ;
  assign n7377 = n2414 & ~n7376 ;
  assign n7378 = n7377 ^ n4009 ^ 1'b0 ;
  assign n7380 = ~n3331 & n3982 ;
  assign n7381 = n7380 ^ n5830 ^ 1'b0 ;
  assign n7379 = n5567 | n6450 ;
  assign n7382 = n7381 ^ n7379 ^ 1'b0 ;
  assign n7383 = n6022 ^ n4024 ^ 1'b0 ;
  assign n7384 = n7155 ^ n3707 ^ 1'b0 ;
  assign n7385 = n3377 ^ n292 ^ 1'b0 ;
  assign n7386 = n1158 & ~n7385 ;
  assign n7387 = n4753 ^ n1223 ^ 1'b0 ;
  assign n7388 = ~n1994 & n2008 ;
  assign n7389 = ~n366 & n7388 ;
  assign n7390 = n7389 ^ n951 ^ 1'b0 ;
  assign n7391 = n2188 & n4791 ;
  assign n7392 = ( n3725 & n5155 ) | ( n3725 & n7391 ) | ( n5155 & n7391 ) ;
  assign n7393 = n3473 | n4490 ;
  assign n7394 = n7393 ^ n2564 ^ 1'b0 ;
  assign n7395 = n1464 & ~n2165 ;
  assign n7396 = n7395 ^ n3881 ^ 1'b0 ;
  assign n7397 = n3431 & n7396 ;
  assign n7399 = n3928 ^ n1028 ^ 1'b0 ;
  assign n7400 = n2035 | n7399 ;
  assign n7398 = n7131 ^ n7108 ^ 1'b0 ;
  assign n7401 = n7400 ^ n7398 ^ 1'b0 ;
  assign n7402 = n2371 | n2441 ;
  assign n7403 = n7402 ^ n4274 ^ 1'b0 ;
  assign n7404 = n3953 ^ n817 ^ 1'b0 ;
  assign n7405 = ~n3567 & n3891 ;
  assign n7406 = n897 & n7405 ;
  assign n7407 = n3340 | n6412 ;
  assign n7408 = n1219 & ~n4162 ;
  assign n7409 = n2210 | n4217 ;
  assign n7410 = n7408 & ~n7409 ;
  assign n7411 = n2796 & n3998 ;
  assign n7412 = n6748 ^ n5328 ^ 1'b0 ;
  assign n7413 = n7411 | n7412 ;
  assign n7414 = n6025 | n7181 ;
  assign n7415 = n3694 & ~n5646 ;
  assign n7416 = n7415 ^ x42 ^ 1'b0 ;
  assign n7418 = n2358 ^ n2143 ^ 1'b0 ;
  assign n7419 = ~n2122 & n7418 ;
  assign n7417 = x202 & ~n796 ;
  assign n7420 = n7419 ^ n7417 ^ 1'b0 ;
  assign n7421 = n3626 ^ n2914 ^ n2172 ;
  assign n7422 = n4459 ^ n1537 ^ 1'b0 ;
  assign n7423 = n7421 & ~n7422 ;
  assign n7424 = x189 & n7423 ;
  assign n7425 = n7424 ^ n339 ^ 1'b0 ;
  assign n7426 = n3611 ^ x80 ^ 1'b0 ;
  assign n7427 = n6522 & n7426 ;
  assign n7428 = n1832 | n7427 ;
  assign n7429 = n7425 & ~n7428 ;
  assign n7430 = ~n1832 & n1883 ;
  assign n7433 = ~n1350 & n1757 ;
  assign n7434 = n7433 ^ n265 ^ 1'b0 ;
  assign n7435 = n3165 ^ n1081 ^ 1'b0 ;
  assign n7436 = x115 & ~n7435 ;
  assign n7437 = n7434 | n7436 ;
  assign n7431 = n2609 ^ n1106 ^ 1'b0 ;
  assign n7432 = ~n4709 & n7431 ;
  assign n7438 = n7437 ^ n7432 ^ 1'b0 ;
  assign n7439 = n1947 & n3333 ;
  assign n7440 = n7439 ^ n6950 ^ 1'b0 ;
  assign n7441 = x163 & ~n1865 ;
  assign n7442 = n7441 ^ n4509 ^ 1'b0 ;
  assign n7443 = ( n3373 & n7440 ) | ( n3373 & ~n7442 ) | ( n7440 & ~n7442 ) ;
  assign n7444 = x28 | n4715 ;
  assign n7445 = ~n2467 & n7444 ;
  assign n7446 = n7445 ^ n4840 ^ 1'b0 ;
  assign n7447 = n1791 & ~n1951 ;
  assign n7448 = n7447 ^ n655 ^ 1'b0 ;
  assign n7449 = n2686 & ~n6509 ;
  assign n7451 = n1310 & ~n2134 ;
  assign n7452 = ~n1139 & n7451 ;
  assign n7450 = ( n313 & n1967 ) | ( n313 & n2129 ) | ( n1967 & n2129 ) ;
  assign n7453 = n7452 ^ n7450 ^ 1'b0 ;
  assign n7454 = ~n4149 & n7453 ;
  assign n7455 = n1867 | n3451 ;
  assign n7456 = n7455 ^ n6768 ^ 1'b0 ;
  assign n7457 = n1521 & ~n7456 ;
  assign n7458 = n5184 & n6047 ;
  assign n7459 = n7458 ^ n3750 ^ 1'b0 ;
  assign n7460 = n1320 | n5193 ;
  assign n7461 = n7460 ^ n2681 ^ 1'b0 ;
  assign n7462 = x98 & n3270 ;
  assign n7463 = ~n7461 & n7462 ;
  assign n7464 = n988 | n7463 ;
  assign n7465 = n2629 | n7464 ;
  assign n7466 = n3799 & n7465 ;
  assign n7467 = x186 & ~n5061 ;
  assign n7468 = n2119 & n4169 ;
  assign n7469 = ~n3410 & n7468 ;
  assign n7470 = n7469 ^ n1628 ^ 1'b0 ;
  assign n7471 = n6190 & ~n7470 ;
  assign n7472 = n630 & ~n696 ;
  assign n7473 = n2293 & n7472 ;
  assign n7474 = n6537 & n7473 ;
  assign n7475 = n7474 ^ n3902 ^ 1'b0 ;
  assign n7476 = n6228 ^ n5613 ^ 1'b0 ;
  assign n7477 = n7476 ^ n747 ^ 1'b0 ;
  assign n7478 = n2476 ^ n1066 ^ 1'b0 ;
  assign n7479 = ~n543 & n7478 ;
  assign n7480 = n2908 & ~n7479 ;
  assign n7481 = n7480 ^ n6057 ^ 1'b0 ;
  assign n7482 = n1423 & n3881 ;
  assign n7483 = n7482 ^ n1035 ^ 1'b0 ;
  assign n7484 = n2487 & ~n5189 ;
  assign n7485 = n3807 | n4993 ;
  assign n7486 = n2132 ^ n760 ^ 1'b0 ;
  assign n7487 = n6473 | n7486 ;
  assign n7488 = n3585 & ~n7487 ;
  assign n7489 = x84 & ~n7488 ;
  assign n7490 = ~n705 & n1514 ;
  assign n7491 = ~n6935 & n7490 ;
  assign n7492 = n1077 | n5030 ;
  assign n7493 = n7400 & ~n7492 ;
  assign n7494 = n639 & ~n7493 ;
  assign n7495 = n2017 ^ n1780 ^ 1'b0 ;
  assign n7496 = n1861 ^ n1792 ^ 1'b0 ;
  assign n7497 = n2741 & ~n7496 ;
  assign n7498 = n5779 & n6061 ;
  assign n7500 = n3740 ^ n918 ^ 1'b0 ;
  assign n7499 = ~x115 & n7243 ;
  assign n7501 = n7500 ^ n7499 ^ 1'b0 ;
  assign n7502 = n669 | n1693 ;
  assign n7503 = n2074 & ~n4117 ;
  assign n7504 = n7502 & n7503 ;
  assign n7509 = n1483 & ~n2320 ;
  assign n7506 = ~n1619 & n6626 ;
  assign n7507 = ~x2 & n7506 ;
  assign n7505 = n647 & n1773 ;
  assign n7508 = n7507 ^ n7505 ^ 1'b0 ;
  assign n7510 = n7509 ^ n7508 ^ 1'b0 ;
  assign n7511 = n7510 ^ n4671 ^ 1'b0 ;
  assign n7512 = n7504 | n7511 ;
  assign n7513 = n3267 & n7512 ;
  assign n7514 = n946 & n2184 ;
  assign n7515 = n7514 ^ n2903 ^ 1'b0 ;
  assign n7516 = n1381 ^ n1073 ^ 1'b0 ;
  assign n7517 = n2026 ^ n1195 ^ 1'b0 ;
  assign n7518 = n641 | n7517 ;
  assign n7519 = n7518 ^ n6962 ^ 1'b0 ;
  assign n7524 = n598 | n1347 ;
  assign n7525 = ~n4718 & n7524 ;
  assign n7526 = n7525 ^ n2247 ^ 1'b0 ;
  assign n7520 = n6859 ^ n5438 ^ 1'b0 ;
  assign n7521 = n7520 ^ n7115 ^ 1'b0 ;
  assign n7522 = n2082 & ~n7521 ;
  assign n7523 = n5173 & n7522 ;
  assign n7527 = n7526 ^ n7523 ^ 1'b0 ;
  assign n7528 = n4536 ^ n2604 ^ 1'b0 ;
  assign n7529 = n3270 ^ n1031 ^ 1'b0 ;
  assign n7530 = n7529 ^ n2469 ^ 1'b0 ;
  assign n7531 = ~n7528 & n7530 ;
  assign n7532 = n5907 & ~n7117 ;
  assign n7533 = n7532 ^ n3678 ^ 1'b0 ;
  assign n7534 = n3475 ^ x233 ^ 1'b0 ;
  assign n7535 = n387 & ~n7534 ;
  assign n7536 = n7535 ^ x195 ^ 1'b0 ;
  assign n7537 = n3269 ^ n1973 ^ 1'b0 ;
  assign n7538 = n4626 | n7537 ;
  assign n7539 = n4380 & n7538 ;
  assign n7540 = n7539 ^ n3275 ^ 1'b0 ;
  assign n7541 = ~n1451 & n2820 ;
  assign n7542 = n5926 & n7541 ;
  assign n7543 = n6482 ^ n4429 ^ 1'b0 ;
  assign n7544 = n7542 | n7543 ;
  assign n7545 = n637 | n1327 ;
  assign n7546 = n7545 ^ n6189 ^ 1'b0 ;
  assign n7547 = n5023 & n7546 ;
  assign n7548 = n2740 ^ n1936 ^ x179 ;
  assign n7549 = n7548 ^ n4083 ^ 1'b0 ;
  assign n7550 = n3033 ^ n1688 ^ 1'b0 ;
  assign n7551 = n1639 & ~n4980 ;
  assign n7552 = n7551 ^ n3938 ^ 1'b0 ;
  assign n7553 = n894 & ~n1606 ;
  assign n7554 = n7553 ^ x218 ^ 1'b0 ;
  assign n7555 = n571 | n7554 ;
  assign n7556 = n4352 | n7555 ;
  assign n7557 = ~n564 & n7556 ;
  assign n7558 = n1154 | n2085 ;
  assign n7559 = ( x49 & n2500 ) | ( x49 & ~n4728 ) | ( n2500 & ~n4728 ) ;
  assign n7560 = n7558 & ~n7559 ;
  assign n7561 = ~n1419 & n1864 ;
  assign n7562 = n7561 ^ n3145 ^ 1'b0 ;
  assign n7563 = n6617 ^ n4147 ^ 1'b0 ;
  assign n7567 = n3154 & n7034 ;
  assign n7564 = ~n368 & n1195 ;
  assign n7565 = ~n4120 & n7564 ;
  assign n7566 = n1333 | n7565 ;
  assign n7568 = n7567 ^ n7566 ^ 1'b0 ;
  assign n7569 = n1955 & ~n5683 ;
  assign n7570 = n6483 & ~n7569 ;
  assign n7571 = n7570 ^ n1925 ^ 1'b0 ;
  assign n7572 = n2073 & n7571 ;
  assign n7573 = ~n6379 & n7572 ;
  assign n7574 = n4913 & ~n6469 ;
  assign n7575 = n7552 & n7574 ;
  assign n7579 = n504 | n3739 ;
  assign n7580 = n1846 | n7579 ;
  assign n7581 = ~n493 & n7580 ;
  assign n7582 = n7581 ^ n7034 ^ 1'b0 ;
  assign n7576 = n3522 ^ n3140 ^ 1'b0 ;
  assign n7577 = ~n5728 & n7576 ;
  assign n7578 = n7577 ^ n2359 ^ 1'b0 ;
  assign n7583 = n7582 ^ n7578 ^ n7512 ;
  assign n7584 = n2166 & ~n3466 ;
  assign n7585 = n4222 | n4306 ;
  assign n7586 = n502 & n7585 ;
  assign n7587 = n7586 ^ n6895 ^ 1'b0 ;
  assign n7588 = n959 & n7587 ;
  assign n7589 = x130 & n1310 ;
  assign n7590 = n6239 & n7589 ;
  assign n7591 = n417 | n7590 ;
  assign n7592 = ~n901 & n6034 ;
  assign n7593 = n7592 ^ n3960 ^ 1'b0 ;
  assign n7594 = n2896 & n4801 ;
  assign n7595 = n5552 ^ n2846 ^ 1'b0 ;
  assign n7596 = n428 | n3635 ;
  assign n7597 = n7596 ^ n1351 ^ 1'b0 ;
  assign n7598 = ~n2887 & n7597 ;
  assign n7599 = ~n2633 & n7598 ;
  assign n7600 = n703 & n3812 ;
  assign n7601 = n7599 & n7600 ;
  assign n7602 = n1183 | n4347 ;
  assign n7603 = n1382 & ~n7602 ;
  assign n7604 = n623 | n1191 ;
  assign n7605 = n7604 ^ n6460 ^ n1608 ;
  assign n7606 = n2081 & ~n2853 ;
  assign n7607 = n7606 ^ n2256 ^ 1'b0 ;
  assign n7608 = ~n6236 & n7607 ;
  assign n7609 = ~n1381 & n6117 ;
  assign n7610 = n1931 ^ n261 ^ 1'b0 ;
  assign n7611 = n6617 | n7610 ;
  assign n7612 = n7611 ^ n1953 ^ 1'b0 ;
  assign n7613 = n666 & ~n7612 ;
  assign n7614 = n3561 ^ n1160 ^ 1'b0 ;
  assign n7615 = ~n1447 & n7614 ;
  assign n7616 = ~n5527 & n7615 ;
  assign n7617 = n4590 & n7616 ;
  assign n7618 = n7617 ^ n5089 ^ 1'b0 ;
  assign n7619 = ~n1410 & n5578 ;
  assign n7620 = n4834 ^ n354 ^ 1'b0 ;
  assign n7621 = ~n3845 & n7620 ;
  assign n7622 = ~n6809 & n7621 ;
  assign n7623 = x11 & ~n3345 ;
  assign n7624 = ~n1344 & n7623 ;
  assign n7625 = n5496 & n7061 ;
  assign n7628 = n3169 ^ n2844 ^ 1'b0 ;
  assign n7626 = ~n1806 & n3452 ;
  assign n7627 = n7626 ^ n315 ^ 1'b0 ;
  assign n7629 = n7628 ^ n7627 ^ 1'b0 ;
  assign n7630 = n6442 & ~n7629 ;
  assign n7631 = n2997 & ~n5255 ;
  assign n7632 = ~n271 & n7631 ;
  assign n7633 = n4256 ^ n1974 ^ 1'b0 ;
  assign n7634 = n1513 | n5867 ;
  assign n7635 = n1305 ^ n1077 ^ 1'b0 ;
  assign n7636 = ~n3953 & n7635 ;
  assign n7637 = n7253 | n7636 ;
  assign n7638 = n5733 ^ n2581 ^ 1'b0 ;
  assign n7639 = n7638 ^ n4236 ^ 1'b0 ;
  assign n7640 = ~n1059 & n3707 ;
  assign n7641 = n7640 ^ n4822 ^ 1'b0 ;
  assign n7642 = n3611 | n3731 ;
  assign n7643 = n1243 | n4063 ;
  assign n7644 = n2839 & ~n4709 ;
  assign n7645 = ~n2869 & n7644 ;
  assign n7646 = n7645 ^ n6846 ^ 1'b0 ;
  assign n7647 = n5840 ^ n446 ^ 1'b0 ;
  assign n7648 = n4117 | n7647 ;
  assign n7649 = n3388 ^ n2789 ^ 1'b0 ;
  assign n7650 = ~n1807 & n7649 ;
  assign n7651 = n7648 | n7650 ;
  assign n7652 = x24 | n7651 ;
  assign n7653 = n3254 ^ x16 ^ 1'b0 ;
  assign n7654 = n2868 & ~n7653 ;
  assign n7655 = n4551 ^ n2565 ^ n600 ;
  assign n7656 = ~n7654 & n7655 ;
  assign n7657 = n603 & n7656 ;
  assign n7659 = n2136 & n3175 ;
  assign n7658 = n1847 & n4143 ;
  assign n7660 = n7659 ^ n7658 ^ 1'b0 ;
  assign n7661 = n4172 ^ n4122 ^ 1'b0 ;
  assign n7667 = n1134 & n1818 ;
  assign n7662 = n2075 | n3729 ;
  assign n7663 = n7662 ^ n1506 ^ 1'b0 ;
  assign n7664 = n6544 & n7663 ;
  assign n7665 = n3636 & ~n4573 ;
  assign n7666 = ~n7664 & n7665 ;
  assign n7668 = n7667 ^ n7666 ^ n4838 ;
  assign n7669 = n6825 ^ n3703 ^ 1'b0 ;
  assign n7670 = n7669 ^ n7352 ^ 1'b0 ;
  assign n7671 = n4688 & n6369 ;
  assign n7672 = ~n5796 & n7671 ;
  assign n7673 = n6033 & n7672 ;
  assign n7674 = n5124 & ~n7673 ;
  assign n7675 = n7674 ^ n381 ^ 1'b0 ;
  assign n7679 = n1451 & ~n3122 ;
  assign n7676 = x47 & ~n954 ;
  assign n7677 = n7676 ^ n4331 ^ 1'b0 ;
  assign n7678 = n2116 | n7677 ;
  assign n7680 = n7679 ^ n7678 ^ 1'b0 ;
  assign n7681 = n1646 & n7680 ;
  assign n7682 = n2850 ^ n478 ^ 1'b0 ;
  assign n7683 = n5569 ^ n3266 ^ 1'b0 ;
  assign n7684 = n6740 & n7683 ;
  assign n7685 = n3780 & ~n5205 ;
  assign n7686 = ~n1216 & n4031 ;
  assign n7687 = n1893 & n7686 ;
  assign n7688 = ( n1130 & n7548 ) | ( n1130 & n7687 ) | ( n7548 & n7687 ) ;
  assign n7689 = n4040 ^ n1904 ^ 1'b0 ;
  assign n7690 = n1576 | n6502 ;
  assign n7691 = n6328 & n7039 ;
  assign n7692 = n7461 ^ n2116 ^ 1'b0 ;
  assign n7693 = n5287 & ~n7677 ;
  assign n7694 = ( ~n1114 & n5233 ) | ( ~n1114 & n7693 ) | ( n5233 & n7693 ) ;
  assign n7695 = n4376 & ~n4806 ;
  assign n7696 = n880 & ~n7695 ;
  assign n7697 = n4742 ^ x137 ^ 1'b0 ;
  assign n7699 = n1040 & n1945 ;
  assign n7700 = n3703 & n7699 ;
  assign n7698 = ~n528 & n729 ;
  assign n7701 = n7700 ^ n7698 ^ 1'b0 ;
  assign n7702 = n5442 ^ n571 ^ 1'b0 ;
  assign n7703 = n1576 & ~n7702 ;
  assign n7704 = n5989 ^ n4091 ^ 1'b0 ;
  assign n7705 = n2521 & ~n6546 ;
  assign n7706 = n1361 & ~n4608 ;
  assign n7707 = n3725 ^ n2003 ^ 1'b0 ;
  assign n7708 = n5424 & ~n7707 ;
  assign n7709 = ~n4548 & n7708 ;
  assign n7710 = n5530 ^ n2406 ^ 1'b0 ;
  assign n7711 = n7153 ^ n1720 ^ 1'b0 ;
  assign n7712 = n1948 ^ n748 ^ 1'b0 ;
  assign n7713 = n4834 | n7712 ;
  assign n7716 = n7640 ^ n3645 ^ 1'b0 ;
  assign n7714 = n1463 & ~n4002 ;
  assign n7715 = ~n2376 & n7714 ;
  assign n7717 = n7716 ^ n7715 ^ 1'b0 ;
  assign n7718 = ~n2476 & n3346 ;
  assign n7722 = n5452 ^ n335 ^ 1'b0 ;
  assign n7723 = n1787 & ~n7722 ;
  assign n7719 = n461 & ~n4204 ;
  assign n7720 = n4709 & n7719 ;
  assign n7721 = n7720 ^ n2629 ^ 1'b0 ;
  assign n7724 = n7723 ^ n7721 ^ 1'b0 ;
  assign n7725 = n7718 & ~n7724 ;
  assign n7726 = n7725 ^ n1324 ^ 1'b0 ;
  assign n7727 = n2890 | n4709 ;
  assign n7728 = n7403 ^ n6963 ^ 1'b0 ;
  assign n7729 = ~n7727 & n7728 ;
  assign n7730 = ~n3633 & n4788 ;
  assign n7731 = n2345 & ~n2836 ;
  assign n7732 = n7731 ^ n1620 ^ 1'b0 ;
  assign n7733 = x133 | n4527 ;
  assign n7734 = n7733 ^ n872 ^ 1'b0 ;
  assign n7735 = n6083 ^ n2034 ^ 1'b0 ;
  assign n7736 = n285 | n7735 ;
  assign n7737 = n6298 ^ x202 ^ 1'b0 ;
  assign n7738 = n3772 & ~n7737 ;
  assign n7739 = ~n1507 & n7097 ;
  assign n7740 = n2129 & ~n3620 ;
  assign n7741 = ~n3399 & n7740 ;
  assign n7742 = n846 | n7741 ;
  assign n7743 = n7583 | n7742 ;
  assign n7744 = x60 & n5132 ;
  assign n7745 = n7744 ^ n4176 ^ 1'b0 ;
  assign n7746 = n566 & n6026 ;
  assign n7747 = ~n1236 & n6141 ;
  assign n7748 = n5282 & n7747 ;
  assign n7749 = n7748 ^ x151 ^ 1'b0 ;
  assign n7750 = n7220 ^ n869 ^ 1'b0 ;
  assign n7752 = n3345 ^ n1035 ^ 1'b0 ;
  assign n7753 = n4502 & ~n7752 ;
  assign n7751 = n6228 & ~n7131 ;
  assign n7754 = n7753 ^ n7751 ^ 1'b0 ;
  assign n7755 = n5478 ^ n4658 ^ 1'b0 ;
  assign n7756 = n384 | n5770 ;
  assign n7759 = n1677 ^ n1190 ^ 1'b0 ;
  assign n7760 = n3481 & n7759 ;
  assign n7757 = x169 & n3015 ;
  assign n7758 = n6524 & n7757 ;
  assign n7761 = n7760 ^ n7758 ^ 1'b0 ;
  assign n7762 = n6548 & ~n7278 ;
  assign n7763 = ~x204 & n7762 ;
  assign n7764 = n7763 ^ n4701 ^ 1'b0 ;
  assign n7768 = ~n2286 & n3197 ;
  assign n7765 = x123 & n7325 ;
  assign n7766 = n7765 ^ n1999 ^ 1'b0 ;
  assign n7767 = x182 & n7766 ;
  assign n7769 = n7768 ^ n7767 ^ 1'b0 ;
  assign n7770 = n3349 ^ x160 ^ 1'b0 ;
  assign n7771 = n3267 & n7770 ;
  assign n7772 = n6019 ^ n1176 ^ 1'b0 ;
  assign n7773 = n7771 & ~n7772 ;
  assign n7774 = n3648 & n7773 ;
  assign n7775 = n2964 & n7774 ;
  assign n7776 = n545 | n7775 ;
  assign n7777 = n7776 ^ n6933 ^ 1'b0 ;
  assign n7778 = n2949 ^ n456 ^ 1'b0 ;
  assign n7779 = n4664 ^ n3221 ^ 1'b0 ;
  assign n7780 = ~n4035 & n7779 ;
  assign n7781 = n7780 ^ n7706 ^ 1'b0 ;
  assign n7782 = n1762 & ~n7381 ;
  assign n7783 = n6749 & n7782 ;
  assign n7784 = n2019 | n3659 ;
  assign n7785 = n7784 ^ n4850 ^ 1'b0 ;
  assign n7786 = n546 & ~n4873 ;
  assign n7787 = n832 & n7786 ;
  assign n7788 = ( n4400 & ~n5378 ) | ( n4400 & n7199 ) | ( ~n5378 & n7199 ) ;
  assign n7789 = n1453 & n6882 ;
  assign n7790 = n3214 ^ n2526 ^ 1'b0 ;
  assign n7791 = n2891 & n7790 ;
  assign n7792 = n1337 & ~n6127 ;
  assign n7793 = n325 | n2207 ;
  assign n7794 = n7793 ^ n2186 ^ 1'b0 ;
  assign n7795 = ~n2799 & n7794 ;
  assign n7796 = n7795 ^ n821 ^ 1'b0 ;
  assign n7797 = ~n1324 & n3288 ;
  assign n7798 = ~n6355 & n7797 ;
  assign n7799 = ~n1689 & n6935 ;
  assign n7800 = n7798 & n7799 ;
  assign n7801 = n2097 ^ n644 ^ 1'b0 ;
  assign n7802 = n1791 & n7801 ;
  assign n7803 = n7132 & n7802 ;
  assign n7804 = n7803 ^ n2024 ^ 1'b0 ;
  assign n7805 = n901 | n5444 ;
  assign n7806 = n4222 & ~n7805 ;
  assign n7807 = n7806 ^ n3417 ^ 1'b0 ;
  assign n7808 = n2194 & n6320 ;
  assign n7809 = n7808 ^ n7644 ^ 1'b0 ;
  assign n7810 = n4432 | n5915 ;
  assign n7812 = n279 | n4051 ;
  assign n7813 = n2402 & ~n7812 ;
  assign n7811 = x22 & n1014 ;
  assign n7814 = n7813 ^ n7811 ^ 1'b0 ;
  assign n7815 = n788 | n2301 ;
  assign n7816 = n7815 ^ n4541 ^ 1'b0 ;
  assign n7817 = n7816 ^ n7257 ^ 1'b0 ;
  assign n7818 = n3181 & n7817 ;
  assign n7819 = n5129 ^ n3068 ^ 1'b0 ;
  assign n7820 = n2517 & ~n7819 ;
  assign n7821 = n1383 | n7820 ;
  assign n7822 = ~x147 & n795 ;
  assign n7823 = ~n1667 & n2672 ;
  assign n7824 = n7823 ^ n685 ^ 1'b0 ;
  assign n7825 = ~n2677 & n6285 ;
  assign n7826 = ~n7824 & n7825 ;
  assign n7827 = n7826 ^ n1909 ^ n1644 ;
  assign n7828 = ( ~n1139 & n3081 ) | ( ~n1139 & n4229 ) | ( n3081 & n4229 ) ;
  assign n7829 = n2243 & ~n5179 ;
  assign n7830 = x0 & x3 ;
  assign n7831 = n2035 | n7830 ;
  assign n7832 = n7831 ^ n921 ^ 1'b0 ;
  assign n7833 = n4810 & n7832 ;
  assign n7834 = n7829 | n7833 ;
  assign n7835 = n7834 ^ n3714 ^ 1'b0 ;
  assign n7836 = n4518 ^ n3487 ^ 1'b0 ;
  assign n7837 = n4018 ^ x23 ^ 1'b0 ;
  assign n7838 = n7836 & n7837 ;
  assign n7839 = ~n1483 & n7838 ;
  assign n7840 = n1324 & ~n7839 ;
  assign n7841 = ~x114 & n7840 ;
  assign n7845 = ~n2322 & n4671 ;
  assign n7842 = n1718 | n4445 ;
  assign n7843 = n4972 & n7842 ;
  assign n7844 = n3331 & n7843 ;
  assign n7846 = n7845 ^ n7844 ^ 1'b0 ;
  assign n7847 = n445 ^ x67 ^ 1'b0 ;
  assign n7848 = n5761 ^ n2652 ^ 1'b0 ;
  assign n7849 = n7442 | n7848 ;
  assign n7850 = x205 & n7627 ;
  assign n7851 = n7850 ^ n3955 ^ 1'b0 ;
  assign n7852 = n6133 | n7851 ;
  assign n7853 = n7852 ^ n503 ^ 1'b0 ;
  assign n7854 = n5512 & ~n7853 ;
  assign n7855 = n4964 & n7854 ;
  assign n7856 = x15 & n1228 ;
  assign n7857 = n1819 & n7856 ;
  assign n7858 = n4134 & n7857 ;
  assign n7868 = n470 | n2722 ;
  assign n7867 = n3823 ^ n3681 ^ 1'b0 ;
  assign n7869 = n7868 ^ n7867 ^ 1'b0 ;
  assign n7863 = ~n2179 & n7357 ;
  assign n7859 = n1010 & ~n1729 ;
  assign n7860 = ~n2531 & n7859 ;
  assign n7861 = n1616 & ~n7860 ;
  assign n7862 = n7861 ^ n5155 ^ 1'b0 ;
  assign n7864 = n7863 ^ n7862 ^ 1'b0 ;
  assign n7865 = n6506 ^ n1808 ^ 1'b0 ;
  assign n7866 = n7864 & ~n7865 ;
  assign n7870 = n7869 ^ n7866 ^ 1'b0 ;
  assign n7871 = n934 | n2519 ;
  assign n7872 = n1952 & ~n7871 ;
  assign n7873 = n3858 ^ n1867 ^ 1'b0 ;
  assign n7874 = n3326 & n7873 ;
  assign n7875 = ~n7872 & n7874 ;
  assign n7876 = n7875 ^ n1644 ^ 1'b0 ;
  assign n7877 = n7876 ^ n7391 ^ 1'b0 ;
  assign n7878 = n6416 & n7877 ;
  assign n7879 = n5468 ^ n3901 ^ 1'b0 ;
  assign n7880 = n7878 & ~n7879 ;
  assign n7881 = ~n2709 & n6328 ;
  assign n7882 = n7881 ^ n1622 ^ 1'b0 ;
  assign n7883 = x80 & ~x92 ;
  assign n7884 = n4063 ^ n3489 ^ 1'b0 ;
  assign n7885 = ~n1288 & n7884 ;
  assign n7886 = n1678 & ~n5923 ;
  assign n7887 = n7886 ^ n1337 ^ 1'b0 ;
  assign n7888 = n7887 ^ n2357 ^ 1'b0 ;
  assign n7889 = n4631 | n7888 ;
  assign n7890 = n7757 | n7889 ;
  assign n7891 = ~n1783 & n7890 ;
  assign n7892 = ~n7007 & n7891 ;
  assign n7893 = n3574 & n6719 ;
  assign n7894 = n768 ^ x85 ^ 1'b0 ;
  assign n7895 = n7679 ^ n5366 ^ 1'b0 ;
  assign n7896 = n285 | n6564 ;
  assign n7897 = n6493 | n7896 ;
  assign n7898 = n1622 ^ x27 ^ 1'b0 ;
  assign n7899 = n7898 ^ n1440 ^ 1'b0 ;
  assign n7900 = ~n623 & n4258 ;
  assign n7901 = ~n7124 & n7900 ;
  assign n7902 = n1204 ^ n610 ^ x247 ;
  assign n7903 = n7902 ^ n1523 ^ 1'b0 ;
  assign n7904 = n7903 ^ n2750 ^ 1'b0 ;
  assign n7905 = n623 & n7904 ;
  assign n7906 = n1239 ^ n553 ^ 1'b0 ;
  assign n7907 = ~n1546 & n7906 ;
  assign n7908 = ( n4376 & ~n7005 ) | ( n4376 & n7907 ) | ( ~n7005 & n7907 ) ;
  assign n7909 = n728 & n1112 ;
  assign n7910 = n7909 ^ n1521 ^ 1'b0 ;
  assign n7911 = n7910 ^ n2185 ^ 1'b0 ;
  assign n7912 = n1920 & n7911 ;
  assign n7914 = n3187 | n3801 ;
  assign n7913 = n2867 & ~n3436 ;
  assign n7915 = n7914 ^ n7913 ^ 1'b0 ;
  assign n7916 = x199 & ~n3321 ;
  assign n7917 = n2770 | n7916 ;
  assign n7918 = n2704 & ~n3462 ;
  assign n7919 = n6772 ^ n6278 ^ 1'b0 ;
  assign n7920 = n1814 & ~n7919 ;
  assign n7921 = n1089 & ~n5691 ;
  assign n7922 = ~n6902 & n7921 ;
  assign n7923 = n7922 ^ n4061 ^ 1'b0 ;
  assign n7924 = n7920 & ~n7923 ;
  assign n7925 = n623 | n7924 ;
  assign n7926 = n4009 ^ n3580 ^ 1'b0 ;
  assign n7927 = n7926 ^ n3144 ^ 1'b0 ;
  assign n7928 = n426 & ~n7927 ;
  assign n7929 = n5079 & n6043 ;
  assign n7930 = ~n6160 & n7562 ;
  assign n7931 = n7930 ^ n5193 ^ 1'b0 ;
  assign n7932 = n3855 | n5612 ;
  assign n7933 = n2019 & ~n7932 ;
  assign n7934 = n1836 ^ n994 ^ 1'b0 ;
  assign n7935 = ~n3337 & n7934 ;
  assign n7936 = ~n2143 & n7935 ;
  assign n7937 = n3017 | n7936 ;
  assign n7938 = n3763 ^ n2731 ^ 1'b0 ;
  assign n7939 = n6274 ^ n3385 ^ 1'b0 ;
  assign n7940 = n1380 & n7939 ;
  assign n7941 = n7940 ^ n6179 ^ 1'b0 ;
  assign n7942 = n7938 | n7941 ;
  assign n7943 = n6593 ^ n5372 ^ 1'b0 ;
  assign n7944 = x211 & ~n7943 ;
  assign n7945 = x29 & ~n7928 ;
  assign n7946 = ~n1805 & n7112 ;
  assign n7947 = ~n5703 & n7946 ;
  assign n7948 = n5877 ^ n1335 ^ 1'b0 ;
  assign n7949 = n1857 & ~n7948 ;
  assign n7950 = n1114 & n7415 ;
  assign n7951 = n2572 ^ x41 ^ 1'b0 ;
  assign n7952 = n7951 ^ n2796 ^ 1'b0 ;
  assign n7953 = n5610 & ~n7952 ;
  assign n7954 = n3049 & n5275 ;
  assign n7955 = n2289 | n2384 ;
  assign n7956 = n7955 ^ n796 ^ 1'b0 ;
  assign n7957 = n6564 | n7956 ;
  assign n7959 = n2665 ^ n996 ^ 1'b0 ;
  assign n7958 = ~n1835 & n2629 ;
  assign n7960 = n7959 ^ n7958 ^ 1'b0 ;
  assign n7963 = n1252 & ~n1391 ;
  assign n7964 = ~n3073 & n7963 ;
  assign n7961 = n2550 ^ x185 ^ 1'b0 ;
  assign n7962 = x231 & n7961 ;
  assign n7965 = n7964 ^ n7962 ^ 1'b0 ;
  assign n7966 = n7960 & ~n7965 ;
  assign n7967 = n3283 ^ n2089 ^ 1'b0 ;
  assign n7968 = ~n562 & n979 ;
  assign n7969 = n7968 ^ n1814 ^ 1'b0 ;
  assign n7970 = n7967 & ~n7969 ;
  assign n7971 = ( x193 & n1556 ) | ( x193 & n1914 ) | ( n1556 & n1914 ) ;
  assign n7972 = n7971 ^ n3031 ^ 1'b0 ;
  assign n7973 = ~n3446 & n7972 ;
  assign n7974 = n3548 & ~n7590 ;
  assign n7975 = ~n1588 & n2303 ;
  assign n7976 = n7975 ^ n4602 ^ 1'b0 ;
  assign n7977 = n1146 | n7976 ;
  assign n7978 = n1846 & n4783 ;
  assign n7979 = n4310 & n7978 ;
  assign n7980 = n7979 ^ n4611 ^ 1'b0 ;
  assign n7981 = n3493 & n7980 ;
  assign n7982 = n892 | n4671 ;
  assign n7983 = n5569 ^ n946 ^ 1'b0 ;
  assign n7984 = n7982 | n7983 ;
  assign n7985 = n3199 & ~n6584 ;
  assign n7986 = n7984 & n7985 ;
  assign n7987 = n7986 ^ n3255 ^ 1'b0 ;
  assign n7988 = n2437 & ~n7987 ;
  assign n7989 = n3158 ^ n2063 ^ n602 ;
  assign n7990 = n5645 & n7723 ;
  assign n7991 = n7990 ^ n1130 ^ 1'b0 ;
  assign n7992 = n7991 ^ n6681 ^ n3823 ;
  assign n7993 = n7989 & ~n7992 ;
  assign n7994 = ~n3675 & n5079 ;
  assign n7995 = n7994 ^ n3487 ^ 1'b0 ;
  assign n7996 = n1356 ^ x198 ^ 1'b0 ;
  assign n7997 = n4919 ^ n3250 ^ 1'b0 ;
  assign n7998 = ~n7996 & n7997 ;
  assign n7999 = n6325 ^ n2342 ^ 1'b0 ;
  assign n8000 = n5672 & n7999 ;
  assign n8001 = n1158 & ~n8000 ;
  assign n8002 = n1814 ^ n1540 ^ n349 ;
  assign n8003 = ~n1440 & n8002 ;
  assign n8004 = n8003 ^ n3577 ^ 1'b0 ;
  assign n8005 = n5574 & ~n6327 ;
  assign n8006 = ~n2334 & n2549 ;
  assign n8007 = n1576 ^ n813 ^ 1'b0 ;
  assign n8008 = n3801 & ~n8007 ;
  assign n8009 = n2319 ^ n756 ^ 1'b0 ;
  assign n8010 = n1249 & n8009 ;
  assign n8011 = n3430 & n8010 ;
  assign n8012 = n8008 & ~n8011 ;
  assign n8013 = n1646 ^ x33 ^ 1'b0 ;
  assign n8014 = n4295 & n8013 ;
  assign n8015 = n2698 & ~n6084 ;
  assign n8016 = n8015 ^ n3676 ^ 1'b0 ;
  assign n8017 = ( ~n288 & n8014 ) | ( ~n288 & n8016 ) | ( n8014 & n8016 ) ;
  assign n8018 = x20 | n5196 ;
  assign n8019 = n4688 & n8018 ;
  assign n8020 = n5285 ^ n2591 ^ 1'b0 ;
  assign n8021 = n5879 ^ n830 ^ 1'b0 ;
  assign n8022 = n3314 & ~n8021 ;
  assign n8023 = n2639 & ~n8022 ;
  assign n8024 = n2334 | n4341 ;
  assign n8025 = n1689 ^ n357 ^ 1'b0 ;
  assign n8026 = ~n6595 & n7395 ;
  assign n8027 = n8026 ^ n5213 ^ 1'b0 ;
  assign n8028 = ( n488 & n633 ) | ( n488 & ~n3014 ) | ( n633 & ~n3014 ) ;
  assign n8029 = n4756 ^ n3362 ^ 1'b0 ;
  assign n8030 = n8029 ^ n2938 ^ 1'b0 ;
  assign n8031 = n2527 & n8030 ;
  assign n8032 = n8031 ^ n2672 ^ 1'b0 ;
  assign n8033 = n1947 & n8032 ;
  assign n8034 = n415 & n4389 ;
  assign n8035 = ~n8033 & n8034 ;
  assign n8036 = ~n512 & n4617 ;
  assign n8037 = ~n1255 & n6478 ;
  assign n8038 = ~n8036 & n8037 ;
  assign n8039 = n3842 ^ n1988 ^ 1'b0 ;
  assign n8040 = n1710 & ~n2643 ;
  assign n8041 = n8040 ^ n3040 ^ 1'b0 ;
  assign n8042 = x107 & ~n4992 ;
  assign n8043 = n8042 ^ n5952 ^ 1'b0 ;
  assign n8044 = n8043 ^ n3888 ^ 1'b0 ;
  assign n8045 = ~n2055 & n8044 ;
  assign n8046 = n4753 ^ n2055 ^ 1'b0 ;
  assign n8047 = x228 & ~n8046 ;
  assign n8048 = n7982 & n8047 ;
  assign n8049 = n5134 ^ n2012 ^ 1'b0 ;
  assign n8050 = n836 & n8049 ;
  assign n8051 = n8050 ^ n7195 ^ 1'b0 ;
  assign n8052 = n6486 ^ n808 ^ 1'b0 ;
  assign n8053 = n8051 & ~n8052 ;
  assign n8054 = n726 & n8053 ;
  assign n8055 = n3377 & n8054 ;
  assign n8056 = ~n816 & n4290 ;
  assign n8057 = n2080 & n3756 ;
  assign n8058 = n1326 & n8057 ;
  assign n8059 = n7507 ^ x7 ^ 1'b0 ;
  assign n8060 = n5278 | n6635 ;
  assign n8061 = ~n647 & n1405 ;
  assign n8062 = n8061 ^ n5578 ^ 1'b0 ;
  assign n8063 = n3171 & ~n8062 ;
  assign n8064 = n3226 ^ n1981 ^ 1'b0 ;
  assign n8065 = ~n456 & n1604 ;
  assign n8066 = n2099 | n8065 ;
  assign n8067 = n8066 ^ n3884 ^ 1'b0 ;
  assign n8068 = ~x254 & n8067 ;
  assign n8069 = n8068 ^ n1361 ^ 1'b0 ;
  assign n8070 = n2462 | n8069 ;
  assign n8071 = n4283 ^ n1792 ^ 1'b0 ;
  assign n8072 = ~n1441 & n8071 ;
  assign n8073 = n4207 ^ n1709 ^ 1'b0 ;
  assign n8074 = n4804 & ~n8073 ;
  assign n8075 = n6295 | n8074 ;
  assign n8076 = n8072 | n8075 ;
  assign n8077 = n3758 ^ n2893 ^ 1'b0 ;
  assign n8078 = n6953 ^ n5243 ^ 1'b0 ;
  assign n8079 = ~n8077 & n8078 ;
  assign n8080 = n1056 & ~n1969 ;
  assign n8081 = n6548 & n8080 ;
  assign n8082 = n3522 | n5768 ;
  assign n8083 = n6214 & n7258 ;
  assign n8084 = n2938 | n5564 ;
  assign n8086 = n3385 | n3896 ;
  assign n8087 = n2578 & ~n8086 ;
  assign n8088 = ~n3473 & n8087 ;
  assign n8085 = n1385 & ~n7320 ;
  assign n8089 = n8088 ^ n8085 ^ 1'b0 ;
  assign n8090 = n3632 ^ n610 ^ 1'b0 ;
  assign n8091 = n2870 & ~n8090 ;
  assign n8092 = ~n1661 & n5167 ;
  assign n8093 = n8092 ^ n7654 ^ n1741 ;
  assign n8094 = n675 | n4613 ;
  assign n8095 = n2181 & ~n8094 ;
  assign n8097 = n747 & n3543 ;
  assign n8098 = n1803 ^ n580 ^ 1'b0 ;
  assign n8099 = n8097 & n8098 ;
  assign n8096 = n4061 | n4775 ;
  assign n8100 = n8099 ^ n8096 ^ 1'b0 ;
  assign n8101 = x25 | n8100 ;
  assign n8102 = n2103 ^ n1087 ^ 1'b0 ;
  assign n8103 = n8102 ^ n3634 ^ 1'b0 ;
  assign n8104 = n8103 ^ x4 ^ 1'b0 ;
  assign n8105 = n4907 & ~n5679 ;
  assign n8106 = n4627 & n8105 ;
  assign n8107 = n3774 ^ n1395 ^ 1'b0 ;
  assign n8108 = n1751 | n3172 ;
  assign n8109 = n2896 & ~n4485 ;
  assign n8110 = n8109 ^ n4681 ^ 1'b0 ;
  assign n8111 = ~n611 & n8110 ;
  assign n8112 = n6582 | n7807 ;
  assign n8113 = n663 ^ n374 ^ 1'b0 ;
  assign n8114 = n7173 ^ n6626 ^ 1'b0 ;
  assign n8115 = n3083 | n8114 ;
  assign n8116 = n5529 & n7326 ;
  assign n8117 = n6423 ^ n4107 ^ 1'b0 ;
  assign n8118 = n1291 | n8117 ;
  assign n8120 = n4276 ^ x213 ^ 1'b0 ;
  assign n8119 = n2565 & ~n5150 ;
  assign n8121 = n8120 ^ n8119 ^ 1'b0 ;
  assign n8125 = n566 & ~n1865 ;
  assign n8126 = n8125 ^ n1391 ^ 1'b0 ;
  assign n8122 = ~x199 & n4140 ;
  assign n8123 = ~n2921 & n8122 ;
  assign n8124 = n3614 | n8123 ;
  assign n8127 = n8126 ^ n8124 ^ 1'b0 ;
  assign n8128 = ( n3328 & ~n6665 ) | ( n3328 & n7706 ) | ( ~n6665 & n7706 ) ;
  assign n8129 = n5200 ^ n3854 ^ 1'b0 ;
  assign n8130 = n8129 ^ n860 ^ 1'b0 ;
  assign n8131 = ( ~n1014 & n3040 ) | ( ~n1014 & n7138 ) | ( n3040 & n7138 ) ;
  assign n8132 = n8131 ^ n5737 ^ 1'b0 ;
  assign n8133 = n2675 & n8132 ;
  assign n8134 = ~n3115 & n3476 ;
  assign n8135 = n8134 ^ n1832 ^ 1'b0 ;
  assign n8136 = n8135 ^ n5056 ^ 1'b0 ;
  assign n8137 = n2665 & ~n8136 ;
  assign n8138 = n1783 & n8137 ;
  assign n8139 = n1899 ^ n994 ^ 1'b0 ;
  assign n8140 = n987 & n3619 ;
  assign n8141 = n8140 ^ x232 ^ 1'b0 ;
  assign n8142 = n705 & n8029 ;
  assign n8143 = ~n8141 & n8142 ;
  assign n8144 = ~n2378 & n8143 ;
  assign n8145 = n4501 & ~n5682 ;
  assign n8146 = n7374 ^ n6620 ^ 1'b0 ;
  assign n8147 = n7050 ^ n4485 ^ 1'b0 ;
  assign n8148 = n8006 & n8147 ;
  assign n8149 = n3308 | n4718 ;
  assign n8150 = n8149 ^ n2655 ^ 1'b0 ;
  assign n8151 = x24 & ~n7132 ;
  assign n8152 = n2183 ^ n1513 ^ 1'b0 ;
  assign n8153 = ~n6327 & n8152 ;
  assign n8154 = n3798 | n8153 ;
  assign n8155 = n8024 & n8154 ;
  assign n8159 = x161 & ~n2254 ;
  assign n8160 = n8159 ^ n4705 ^ 1'b0 ;
  assign n8156 = n5062 ^ n4569 ^ 1'b0 ;
  assign n8157 = n7127 & ~n8156 ;
  assign n8158 = ~n6087 & n8157 ;
  assign n8161 = n8160 ^ n8158 ^ 1'b0 ;
  assign n8162 = n1354 | n1657 ;
  assign n8163 = n1111 | n2696 ;
  assign n8164 = n1896 & ~n8163 ;
  assign n8165 = n3468 & ~n8164 ;
  assign n8166 = ~n5864 & n7196 ;
  assign n8167 = ~n8165 & n8166 ;
  assign n8168 = n6780 & n8167 ;
  assign n8169 = n2223 ^ n1087 ^ 1'b0 ;
  assign n8170 = n5928 ^ n3529 ^ 1'b0 ;
  assign n8172 = n3807 & n5292 ;
  assign n8173 = n1181 & n8172 ;
  assign n8171 = ~n1490 & n3694 ;
  assign n8174 = n8173 ^ n8171 ^ 1'b0 ;
  assign n8175 = n1783 & ~n5288 ;
  assign n8176 = n4051 | n6870 ;
  assign n8178 = n480 | n534 ;
  assign n8179 = n8178 ^ n5277 ^ 1'b0 ;
  assign n8177 = x210 & n397 ;
  assign n8180 = n8179 ^ n8177 ^ 1'b0 ;
  assign n8181 = n7281 ^ n1843 ^ 1'b0 ;
  assign n8182 = n1772 | n1787 ;
  assign n8183 = n1680 | n6878 ;
  assign n8184 = n8183 ^ n3950 ^ 1'b0 ;
  assign n8185 = n3723 ^ n903 ^ 1'b0 ;
  assign n8186 = ~n2516 & n8185 ;
  assign n8187 = n4449 & ~n8186 ;
  assign n8188 = n311 | n8187 ;
  assign n8189 = n8188 ^ n5207 ^ 1'b0 ;
  assign n8190 = n8184 & ~n8189 ;
  assign n8191 = n8182 & ~n8190 ;
  assign n8192 = n456 & n1814 ;
  assign n8193 = ~n315 & n6340 ;
  assign n8194 = n8192 & n8193 ;
  assign n8195 = ~n4586 & n8194 ;
  assign n8196 = ~n2485 & n5535 ;
  assign n8201 = ~n1753 & n1953 ;
  assign n8199 = n2119 & ~n3683 ;
  assign n8200 = n8199 ^ n3270 ^ 1'b0 ;
  assign n8197 = n405 | n6813 ;
  assign n8198 = n4209 & ~n8197 ;
  assign n8202 = n8201 ^ n8200 ^ n8198 ;
  assign n8203 = n2764 | n3796 ;
  assign n8204 = ~n723 & n4065 ;
  assign n8205 = n8204 ^ n6511 ^ 1'b0 ;
  assign n8206 = n4432 & n7368 ;
  assign n8207 = n8206 ^ x196 ^ 1'b0 ;
  assign n8208 = n2304 & n8207 ;
  assign n8209 = n1395 & ~n7822 ;
  assign n8210 = n3057 ^ n988 ^ 1'b0 ;
  assign n8211 = ~n2997 & n8210 ;
  assign n8212 = n1333 | n2648 ;
  assign n8213 = n8212 ^ n1411 ^ 1'b0 ;
  assign n8214 = n8211 & ~n8213 ;
  assign n8215 = n2014 & ~n3081 ;
  assign n8216 = n7484 ^ n2089 ^ 1'b0 ;
  assign n8217 = x64 & ~n2295 ;
  assign n8218 = n3624 ^ n883 ^ 1'b0 ;
  assign n8219 = n1749 & ~n4711 ;
  assign n8220 = ~n8218 & n8219 ;
  assign n8221 = ~n5989 & n8220 ;
  assign n8222 = n5804 ^ x159 ^ 1'b0 ;
  assign n8223 = n3358 & n8222 ;
  assign n8224 = n8223 ^ n3667 ^ 1'b0 ;
  assign n8225 = n7288 & ~n8224 ;
  assign n8226 = n6190 & n8225 ;
  assign n8228 = n6407 ^ n2026 ^ 1'b0 ;
  assign n8227 = ~n1339 & n1682 ;
  assign n8229 = n8228 ^ n8227 ^ 1'b0 ;
  assign n8230 = ( n587 & ~n2973 ) | ( n587 & n4734 ) | ( ~n2973 & n4734 ) ;
  assign n8231 = n1682 ^ n1474 ^ 1'b0 ;
  assign n8232 = ~n4037 & n4796 ;
  assign n8233 = n4063 ^ n3759 ^ 1'b0 ;
  assign n8234 = n1801 ^ x4 ^ 1'b0 ;
  assign n8235 = n3361 & n7248 ;
  assign n8236 = ~n8234 & n8235 ;
  assign n8237 = n1920 & n2003 ;
  assign n8239 = n4680 ^ n2159 ^ 1'b0 ;
  assign n8240 = ~n3577 & n8239 ;
  assign n8238 = n468 | n6840 ;
  assign n8241 = n8240 ^ n8238 ^ 1'b0 ;
  assign n8242 = n5748 ^ n2632 ^ x250 ;
  assign n8243 = ( n1116 & n1849 ) | ( n1116 & ~n5909 ) | ( n1849 & ~n5909 ) ;
  assign n8244 = n8243 ^ n5535 ^ 1'b0 ;
  assign n8245 = n653 & n6324 ;
  assign n8246 = n8245 ^ n4378 ^ 1'b0 ;
  assign n8247 = x20 & n6586 ;
  assign n8248 = n4879 & n8247 ;
  assign n8249 = n5898 | n7563 ;
  assign n8250 = n2165 ^ x60 ^ 1'b0 ;
  assign n8253 = ~x5 & n3065 ;
  assign n8251 = n2013 & ~n5004 ;
  assign n8252 = n7469 | n8251 ;
  assign n8254 = n8253 ^ n8252 ^ 1'b0 ;
  assign n8258 = n7964 ^ n4406 ^ 1'b0 ;
  assign n8255 = n3762 | n4104 ;
  assign n8256 = n8255 ^ n3939 ^ 1'b0 ;
  assign n8257 = n8256 ^ n6196 ^ 1'b0 ;
  assign n8259 = n8258 ^ n8257 ^ 1'b0 ;
  assign n8260 = n2152 | n8259 ;
  assign n8261 = n3297 | n8260 ;
  assign n8262 = n4750 | n4979 ;
  assign n8263 = n7054 & ~n8262 ;
  assign n8264 = n5328 | n6312 ;
  assign n8265 = n6312 & ~n8264 ;
  assign n8266 = n3548 | n3571 ;
  assign n8267 = n3548 & ~n8266 ;
  assign n8268 = n3880 & ~n5702 ;
  assign n8269 = n8267 | n8268 ;
  assign n8270 = n8267 & ~n8269 ;
  assign n8271 = n8265 | n8270 ;
  assign n8272 = n2990 ^ n2316 ^ 1'b0 ;
  assign n8273 = n8271 | n8272 ;
  assign n8274 = n1849 | n6499 ;
  assign n8275 = n8274 ^ n4188 ^ 1'b0 ;
  assign n8276 = ~n4076 & n8275 ;
  assign n8277 = n2219 & n2241 ;
  assign n8278 = n8277 ^ n1194 ^ 1'b0 ;
  assign n8279 = x151 & ~n6974 ;
  assign n8280 = x148 & n5650 ;
  assign n8283 = n1970 | n7518 ;
  assign n8281 = n1724 ^ n1269 ^ 1'b0 ;
  assign n8282 = n1159 & n8281 ;
  assign n8284 = n8283 ^ n8282 ^ 1'b0 ;
  assign n8285 = n1417 | n8284 ;
  assign n8286 = x5 & n1897 ;
  assign n8287 = n7498 & ~n8286 ;
  assign n8288 = n3569 | n6020 ;
  assign n8289 = ~n3549 & n4393 ;
  assign n8290 = n3468 ^ x64 ^ 1'b0 ;
  assign n8291 = n4615 | n8290 ;
  assign n8292 = ~n5210 & n6055 ;
  assign n8293 = n8292 ^ n3115 ^ 1'b0 ;
  assign n8294 = n3212 & ~n7876 ;
  assign n8295 = n7507 ^ n4988 ^ x161 ;
  assign n8296 = n7977 ^ n288 ^ 1'b0 ;
  assign n8297 = n8127 & ~n8296 ;
  assign n8298 = n4641 | n6400 ;
  assign n8299 = ~n1027 & n8298 ;
  assign n8300 = x115 | n2689 ;
  assign n8301 = n1787 & n8300 ;
  assign n8302 = n1682 ^ x44 ^ 1'b0 ;
  assign n8303 = ~n4205 & n8302 ;
  assign n8304 = n8303 ^ n1182 ^ 1'b0 ;
  assign n8305 = n4168 | n8304 ;
  assign n8306 = n3091 | n6123 ;
  assign n8307 = n8306 ^ n950 ^ 1'b0 ;
  assign n8308 = n1732 & n3402 ;
  assign n8309 = n8308 ^ n6637 ^ 1'b0 ;
  assign n8310 = n8309 ^ n6788 ^ 1'b0 ;
  assign n8311 = n8307 | n8310 ;
  assign n8312 = ~n948 & n2624 ;
  assign n8313 = x92 & n8312 ;
  assign n8314 = n8311 & n8313 ;
  assign n8315 = n3672 & n6768 ;
  assign n8316 = ~n6988 & n8315 ;
  assign n8317 = n7316 & n8316 ;
  assign n8318 = n2581 | n8317 ;
  assign n8319 = n8318 ^ n3242 ^ 1'b0 ;
  assign n8320 = n2510 ^ n978 ^ 1'b0 ;
  assign n8321 = n5021 ^ n3998 ^ 1'b0 ;
  assign n8322 = n8320 | n8321 ;
  assign n8324 = ~n4257 & n4580 ;
  assign n8325 = n1048 & n4507 ;
  assign n8326 = n5514 & n8325 ;
  assign n8327 = n8324 & ~n8326 ;
  assign n8328 = n1212 & n8327 ;
  assign n8323 = n1208 & ~n3819 ;
  assign n8329 = n8328 ^ n8323 ^ 1'b0 ;
  assign n8330 = n8099 ^ n5521 ^ 1'b0 ;
  assign n8331 = ~n4048 & n8330 ;
  assign n8332 = ~n5215 & n8115 ;
  assign n8333 = x25 & ~n1021 ;
  assign n8334 = n956 | n8333 ;
  assign n8335 = n820 | n3000 ;
  assign n8336 = n8335 ^ x145 ^ 1'b0 ;
  assign n8337 = n3158 | n3313 ;
  assign n8338 = n8336 | n8337 ;
  assign n8339 = ~n5360 & n8338 ;
  assign n8340 = ~n4991 & n8339 ;
  assign n8341 = n7739 & ~n8340 ;
  assign n8348 = n3511 ^ n2173 ^ 1'b0 ;
  assign n8342 = n2373 & n5665 ;
  assign n8343 = ~n8201 & n8342 ;
  assign n8344 = n1368 & ~n2534 ;
  assign n8345 = ~n2607 & n8344 ;
  assign n8346 = n1117 | n8345 ;
  assign n8347 = n8343 & ~n8346 ;
  assign n8349 = n8348 ^ n8347 ^ n4565 ;
  assign n8350 = n6489 ^ n3624 ^ 1'b0 ;
  assign n8351 = ~n3790 & n8350 ;
  assign n8352 = n2779 & ~n6939 ;
  assign n8353 = n1704 | n8352 ;
  assign n8354 = n8353 ^ n766 ^ 1'b0 ;
  assign n8355 = n8354 ^ x200 ^ 1'b0 ;
  assign n8356 = n2487 | n8355 ;
  assign n8358 = n6373 ^ n3812 ^ 1'b0 ;
  assign n8359 = n4083 & n8358 ;
  assign n8357 = n4329 & ~n6970 ;
  assign n8360 = n8359 ^ n8357 ^ 1'b0 ;
  assign n8361 = x15 & ~n1893 ;
  assign n8362 = ~n1850 & n8361 ;
  assign n8363 = n8362 ^ n8070 ^ 1'b0 ;
  assign n8364 = x141 & ~n4728 ;
  assign n8365 = n7137 ^ n1360 ^ 1'b0 ;
  assign n8366 = ~n2596 & n4668 ;
  assign n8367 = ~n4481 & n8366 ;
  assign n8368 = x221 & n2746 ;
  assign n8369 = n538 & n8368 ;
  assign n8370 = n1841 & ~n4862 ;
  assign n8371 = n8370 ^ n3198 ^ 1'b0 ;
  assign n8372 = ~n1814 & n8371 ;
  assign n8373 = n2916 & n8372 ;
  assign n8374 = n1380 | n1718 ;
  assign n8375 = n1810 & ~n3790 ;
  assign n8376 = n5791 & n8375 ;
  assign n8377 = ( ~n6004 & n8374 ) | ( ~n6004 & n8376 ) | ( n8374 & n8376 ) ;
  assign n8378 = n397 | n6892 ;
  assign n8379 = ~n2115 & n6290 ;
  assign n8380 = ~n8378 & n8379 ;
  assign n8381 = n8380 ^ n2591 ^ 1'b0 ;
  assign n8382 = n2149 & ~n2561 ;
  assign n8383 = n2962 ^ n859 ^ 1'b0 ;
  assign n8384 = n3182 & n3928 ;
  assign n8385 = n2027 ^ n1546 ^ 1'b0 ;
  assign n8386 = ~n3770 & n8385 ;
  assign n8387 = ~n2704 & n8386 ;
  assign n8388 = n825 & ~n8387 ;
  assign n8389 = n6756 ^ n3939 ^ 1'b0 ;
  assign n8394 = n1442 ^ n452 ^ 1'b0 ;
  assign n8395 = ~n323 & n8394 ;
  assign n8390 = n822 & ~n6768 ;
  assign n8391 = n8390 ^ n4222 ^ 1'b0 ;
  assign n8392 = ~n7826 & n8391 ;
  assign n8393 = ~n1481 & n8392 ;
  assign n8396 = n8395 ^ n8393 ^ 1'b0 ;
  assign n8397 = n1973 ^ n575 ^ 1'b0 ;
  assign n8398 = n8397 ^ n1451 ^ 1'b0 ;
  assign n8399 = n8396 | n8398 ;
  assign n8400 = n957 & ~n8399 ;
  assign n8401 = ~n1148 & n8400 ;
  assign n8402 = n458 | n3413 ;
  assign n8403 = n8402 ^ x184 ^ 1'b0 ;
  assign n8404 = n8403 ^ n529 ^ 1'b0 ;
  assign n8405 = n2175 & n5444 ;
  assign n8406 = ~n3878 & n8405 ;
  assign n8407 = n2098 | n6350 ;
  assign n8408 = n8407 ^ n2846 ^ 1'b0 ;
  assign n8409 = n825 & ~n1330 ;
  assign n8410 = n2964 | n8409 ;
  assign n8411 = n633 ^ x81 ^ 1'b0 ;
  assign n8413 = n2158 & ~n7138 ;
  assign n8414 = n2626 & n8413 ;
  assign n8412 = n281 & ~n2723 ;
  assign n8415 = n8414 ^ n8412 ^ 1'b0 ;
  assign n8416 = n7031 | n8231 ;
  assign n8417 = n6006 & ~n7504 ;
  assign n8418 = n2432 ^ x17 ^ 1'b0 ;
  assign n8419 = n6762 | n8418 ;
  assign n8420 = n2248 | n8419 ;
  assign n8421 = x33 & ~n8420 ;
  assign n8422 = n8421 ^ n3376 ^ 1'b0 ;
  assign n8423 = n5112 & n8422 ;
  assign n8424 = n6298 & n8423 ;
  assign n8425 = ~n3521 & n4720 ;
  assign n8426 = n8425 ^ n4797 ^ 1'b0 ;
  assign n8427 = n8424 | n8426 ;
  assign n8428 = ~n895 & n5587 ;
  assign n8429 = n2697 & n3250 ;
  assign n8430 = n8429 ^ n3212 ^ 1'b0 ;
  assign n8431 = n8430 ^ n1495 ^ 1'b0 ;
  assign n8432 = n2542 & ~n8431 ;
  assign n8433 = n8432 ^ n7555 ^ n2910 ;
  assign n8434 = n3630 & n4976 ;
  assign n8435 = ~n1521 & n8434 ;
  assign n8436 = n5793 | n8435 ;
  assign n8437 = n1566 & n5926 ;
  assign n8438 = n3825 ^ n790 ^ 1'b0 ;
  assign n8439 = n4661 ^ n521 ^ 1'b0 ;
  assign n8440 = ~n548 & n8439 ;
  assign n8441 = n6618 ^ n2244 ^ 1'b0 ;
  assign n8442 = n8440 & ~n8441 ;
  assign n8443 = n8442 ^ n959 ^ 1'b0 ;
  assign n8444 = n8352 ^ n1405 ^ 1'b0 ;
  assign n8445 = n7476 ^ n2575 ^ 1'b0 ;
  assign n8446 = n8445 ^ n8301 ^ 1'b0 ;
  assign n8447 = n903 | n3986 ;
  assign n8448 = n4791 | n8447 ;
  assign n8450 = x155 & n866 ;
  assign n8451 = n8450 ^ n1822 ^ 1'b0 ;
  assign n8449 = ~n930 & n1969 ;
  assign n8452 = n8451 ^ n8449 ^ 1'b0 ;
  assign n8453 = x191 & ~n8452 ;
  assign n8454 = n2076 | n2630 ;
  assign n8455 = x252 & n1990 ;
  assign n8456 = ~n3995 & n8455 ;
  assign n8457 = ~x115 & n8456 ;
  assign n8458 = n747 | n4532 ;
  assign n8459 = n8458 ^ n6584 ^ 1'b0 ;
  assign n8460 = n387 & ~n8459 ;
  assign n8461 = n2336 & ~n5890 ;
  assign n8462 = n458 | n1689 ;
  assign n8463 = n6162 ^ n3290 ^ 1'b0 ;
  assign n8464 = n2247 | n5656 ;
  assign n8465 = ( x172 & ~n1930 ) | ( x172 & n3834 ) | ( ~n1930 & n3834 ) ;
  assign n8466 = ~n5920 & n8465 ;
  assign n8467 = n4538 & n8466 ;
  assign n8468 = n2966 & ~n5231 ;
  assign n8469 = n8319 & ~n8468 ;
  assign n8470 = n1635 & ~n3606 ;
  assign n8471 = n3270 & n3611 ;
  assign n8472 = n6023 & n8471 ;
  assign n8473 = n6389 ^ x151 ^ 1'b0 ;
  assign n8474 = n8473 ^ n4777 ^ 1'b0 ;
  assign n8475 = n331 & n8049 ;
  assign n8476 = ~n623 & n3239 ;
  assign n8477 = n8476 ^ n2165 ^ 1'b0 ;
  assign n8478 = n987 & n1658 ;
  assign n8479 = n3751 | n8478 ;
  assign n8480 = n8479 ^ n8010 ^ 1'b0 ;
  assign n8481 = n5984 ^ n1085 ^ 1'b0 ;
  assign n8483 = n818 & ~n2760 ;
  assign n8484 = ~x3 & n8483 ;
  assign n8482 = n7272 & n8324 ;
  assign n8485 = n8484 ^ n8482 ^ 1'b0 ;
  assign n8486 = n8485 ^ n3533 ^ 1'b0 ;
  assign n8487 = n8481 & n8486 ;
  assign n8488 = n4118 ^ n1826 ^ 1'b0 ;
  assign n8489 = n4327 | n8488 ;
  assign n8490 = n754 & ~n3854 ;
  assign n8491 = ~n1321 & n8490 ;
  assign n8492 = n1619 | n8491 ;
  assign n8493 = ~n8489 & n8492 ;
  assign n8494 = n8493 ^ n1803 ^ 1'b0 ;
  assign n8495 = n2269 & n8494 ;
  assign n8496 = n8495 ^ n2486 ^ 1'b0 ;
  assign n8497 = n2807 & n8496 ;
  assign n8498 = n4788 ^ n436 ^ 1'b0 ;
  assign n8499 = n1536 | n8498 ;
  assign n8500 = n3224 & n8499 ;
  assign n8501 = n5076 ^ n3477 ^ 1'b0 ;
  assign n8502 = n1261 & n1464 ;
  assign n8503 = n950 & n8502 ;
  assign n8504 = x181 & n8503 ;
  assign n8505 = ~n1354 & n8504 ;
  assign n8506 = n7128 & n8505 ;
  assign n8507 = n3020 & n4168 ;
  assign n8508 = ~n4373 & n5932 ;
  assign n8509 = n2177 ^ n934 ^ 1'b0 ;
  assign n8510 = n8509 ^ n6032 ^ 1'b0 ;
  assign n8511 = n2477 | n8510 ;
  assign n8512 = n5232 ^ n571 ^ 1'b0 ;
  assign n8513 = n8512 ^ n2197 ^ 1'b0 ;
  assign n8515 = n3446 ^ n633 ^ 1'b0 ;
  assign n8514 = x147 | n3042 ;
  assign n8516 = n8515 ^ n8514 ^ 1'b0 ;
  assign n8517 = ~n1339 & n1397 ;
  assign n8518 = n8517 ^ n5494 ^ 1'b0 ;
  assign n8519 = ~n8516 & n8518 ;
  assign n8520 = ~n5758 & n8519 ;
  assign n8521 = x229 & ~n2936 ;
  assign n8522 = n1068 & n8521 ;
  assign n8523 = n2582 & n4941 ;
  assign n8524 = n8523 ^ n7720 ^ 1'b0 ;
  assign n8525 = n1105 ^ n793 ^ 1'b0 ;
  assign n8526 = ~n7554 & n7559 ;
  assign n8527 = ~n808 & n1760 ;
  assign n8528 = n895 | n8527 ;
  assign n8529 = x154 | n1770 ;
  assign n8530 = n3641 ^ n2217 ^ 1'b0 ;
  assign n8531 = ~n894 & n8530 ;
  assign n8532 = ( n6136 & ~n8529 ) | ( n6136 & n8531 ) | ( ~n8529 & n8531 ) ;
  assign n8533 = n4010 ^ n1277 ^ 1'b0 ;
  assign n8534 = x30 & ~n8533 ;
  assign n8535 = n8534 ^ n4426 ^ 1'b0 ;
  assign n8536 = ~n8532 & n8535 ;
  assign n8537 = n1093 | n7206 ;
  assign n8538 = n4203 & ~n8537 ;
  assign n8539 = n975 & ~n4063 ;
  assign n8540 = n8538 & n8539 ;
  assign n8541 = n4173 & n6797 ;
  assign n8542 = n2414 & n8541 ;
  assign n8543 = n8540 & n8542 ;
  assign n8544 = n703 | n1843 ;
  assign n8545 = ( n1096 & n5170 ) | ( n1096 & ~n8544 ) | ( n5170 & ~n8544 ) ;
  assign n8546 = x106 & n1354 ;
  assign n8547 = n4617 & ~n5505 ;
  assign n8548 = ~n2029 & n4615 ;
  assign n8549 = x236 & ~n8548 ;
  assign n8550 = n8547 & n8549 ;
  assign n8551 = x145 & n796 ;
  assign n8552 = n666 & ~n8551 ;
  assign n8553 = n8552 ^ n4995 ^ 1'b0 ;
  assign n8554 = n8553 ^ n7407 ^ 1'b0 ;
  assign n8555 = ~n671 & n776 ;
  assign n8556 = n1717 | n7321 ;
  assign n8557 = n2387 ^ n1553 ^ 1'b0 ;
  assign n8558 = n8556 & n8557 ;
  assign n8559 = n8558 ^ n6537 ^ 1'b0 ;
  assign n8560 = n4354 ^ n3473 ^ 1'b0 ;
  assign n8561 = n4684 | n8560 ;
  assign n8562 = n3854 & ~n8561 ;
  assign n8563 = ~n2114 & n5700 ;
  assign n8564 = n8563 ^ n2987 ^ 1'b0 ;
  assign n8565 = ( n492 & n3449 ) | ( n492 & ~n4385 ) | ( n3449 & ~n4385 ) ;
  assign n8566 = n3760 & n4324 ;
  assign n8567 = n8566 ^ n2232 ^ 1'b0 ;
  assign n8568 = ~n8565 & n8567 ;
  assign n8569 = n1419 | n5023 ;
  assign n8570 = n1738 | n8569 ;
  assign n8571 = n6288 & n8570 ;
  assign n8572 = n8571 ^ n8137 ^ 1'b0 ;
  assign n8573 = n390 | n3590 ;
  assign n8574 = n1787 ^ n1757 ^ 1'b0 ;
  assign n8575 = n787 & ~n8574 ;
  assign n8576 = n1859 & n8575 ;
  assign n8577 = n5398 ^ n1949 ^ 1'b0 ;
  assign n8578 = n3963 | n8577 ;
  assign n8579 = x67 & ~n4653 ;
  assign n8580 = n8579 ^ n2152 ^ 1'b0 ;
  assign n8581 = ~n3055 & n8580 ;
  assign n8582 = ~x173 & n8581 ;
  assign n8583 = n920 | n4100 ;
  assign n8584 = n8583 ^ n2804 ^ 1'b0 ;
  assign n8585 = n956 | n8584 ;
  assign n8586 = x218 & ~n8585 ;
  assign n8587 = n8582 | n8586 ;
  assign n8588 = n8578 & ~n8587 ;
  assign n8589 = n470 & n2184 ;
  assign n8590 = n3403 | n8589 ;
  assign n8591 = n8590 ^ n5043 ^ 1'b0 ;
  assign n8592 = n1417 | n3625 ;
  assign n8593 = n8497 ^ n6781 ^ 1'b0 ;
  assign n8594 = ~n8592 & n8593 ;
  assign n8595 = n2219 | n3067 ;
  assign n8596 = n8595 ^ n1987 ^ 1'b0 ;
  assign n8597 = n8596 ^ n3565 ^ 1'b0 ;
  assign n8598 = n6030 ^ n5056 ^ 1'b0 ;
  assign n8599 = n540 & n8598 ;
  assign n8600 = n8599 ^ x2 ^ 1'b0 ;
  assign n8601 = n1825 & n4447 ;
  assign n8602 = ~n4198 & n8601 ;
  assign n8603 = n7284 ^ n4298 ^ 1'b0 ;
  assign n8604 = n4726 & n8603 ;
  assign n8605 = n710 & n1819 ;
  assign n8606 = ~n2082 & n8605 ;
  assign n8607 = n8606 ^ n1814 ^ 1'b0 ;
  assign n8608 = n955 & n8607 ;
  assign n8609 = n4340 ^ n3323 ^ 1'b0 ;
  assign n8610 = n5974 ^ n1037 ^ 1'b0 ;
  assign n8611 = ~n7558 & n8610 ;
  assign n8612 = ( n1897 & ~n2505 ) | ( n1897 & n8611 ) | ( ~n2505 & n8611 ) ;
  assign n8613 = n655 | n8612 ;
  assign n8614 = ~n1802 & n2779 ;
  assign n8615 = n1379 & ~n8614 ;
  assign n8616 = n1159 ^ n1002 ^ 1'b0 ;
  assign n8617 = n8615 & n8616 ;
  assign n8618 = n1776 ^ n1146 ^ 1'b0 ;
  assign n8619 = n3847 & n8618 ;
  assign n8620 = n3410 ^ n1444 ^ 1'b0 ;
  assign n8621 = n8619 & n8620 ;
  assign n8622 = n3181 ^ n2600 ^ 1'b0 ;
  assign n8623 = n1031 | n8622 ;
  assign n8624 = n2072 & ~n8623 ;
  assign n8625 = n8624 ^ n1859 ^ 1'b0 ;
  assign n8626 = ( n1159 & n2414 ) | ( n1159 & ~n3065 ) | ( n2414 & ~n3065 ) ;
  assign n8627 = n8626 ^ n5217 ^ 1'b0 ;
  assign n8628 = n8625 & n8627 ;
  assign n8629 = n8628 ^ n2526 ^ 1'b0 ;
  assign n8630 = n8621 & n8629 ;
  assign n8631 = n3536 ^ n1378 ^ 1'b0 ;
  assign n8632 = n3328 ^ n2476 ^ 1'b0 ;
  assign n8633 = n8632 ^ n4313 ^ 1'b0 ;
  assign n8634 = n4246 & ~n7343 ;
  assign n8635 = ~n3265 & n8634 ;
  assign n8638 = ~n1979 & n7212 ;
  assign n8636 = x254 | n1409 ;
  assign n8637 = n2806 | n8636 ;
  assign n8639 = n8638 ^ n8637 ^ 1'b0 ;
  assign n8640 = ~n4336 & n8639 ;
  assign n8641 = ~n3812 & n5765 ;
  assign n8642 = n8641 ^ n5255 ^ 1'b0 ;
  assign n8643 = ~n2861 & n4469 ;
  assign n8644 = ~n1815 & n8643 ;
  assign n8645 = x233 & ~n8644 ;
  assign n8646 = n895 & ~n5568 ;
  assign n8647 = ~n552 & n2042 ;
  assign n8648 = n6071 ^ n1987 ^ 1'b0 ;
  assign n8649 = ~n8647 & n8648 ;
  assign n8650 = n1727 & n8108 ;
  assign n8651 = n2004 & n8650 ;
  assign n8654 = n1438 | n3624 ;
  assign n8652 = n2298 | n3337 ;
  assign n8653 = n2561 & ~n8652 ;
  assign n8655 = n8654 ^ n8653 ^ 1'b0 ;
  assign n8656 = ~n5110 & n8655 ;
  assign n8657 = n600 & ~n4502 ;
  assign n8658 = n4903 ^ n4521 ^ 1'b0 ;
  assign n8659 = n8658 ^ n5776 ^ n4021 ;
  assign n8660 = n956 | n2083 ;
  assign n8661 = ~n6450 & n8660 ;
  assign n8662 = ~n1835 & n4671 ;
  assign n8663 = ~n8661 & n8662 ;
  assign n8664 = n694 | n2146 ;
  assign n8665 = n1105 | n8664 ;
  assign n8666 = n1042 & n4712 ;
  assign n8667 = ~n7994 & n8666 ;
  assign n8668 = ~n2541 & n6790 ;
  assign n8669 = n691 & n8668 ;
  assign n8672 = n3373 & n6121 ;
  assign n8673 = n546 & n8672 ;
  assign n8670 = n4032 & n6954 ;
  assign n8671 = n2517 & ~n8670 ;
  assign n8674 = n8673 ^ n8671 ^ 1'b0 ;
  assign n8675 = x122 | n856 ;
  assign n8676 = n1701 & n8334 ;
  assign n8677 = n8676 ^ n7196 ^ 1'b0 ;
  assign n8678 = n1370 & ~n6500 ;
  assign n8679 = n8678 ^ n7117 ^ 1'b0 ;
  assign n8680 = n7060 & n8534 ;
  assign n8681 = n8680 ^ n4251 ^ 1'b0 ;
  assign n8682 = n8681 ^ n7945 ^ 1'b0 ;
  assign n8683 = n1219 | n8682 ;
  assign n8684 = n4671 ^ n725 ^ 1'b0 ;
  assign n8685 = x118 & x171 ;
  assign n8686 = ~n972 & n1573 ;
  assign n8687 = n8686 ^ n1606 ^ 1'b0 ;
  assign n8688 = n8687 ^ n6278 ^ 1'b0 ;
  assign n8689 = n8685 & ~n8688 ;
  assign n8691 = n4385 & ~n5288 ;
  assign n8690 = x216 & ~n7570 ;
  assign n8692 = n8691 ^ n8690 ^ 1'b0 ;
  assign n8693 = n4720 ^ n3593 ^ 1'b0 ;
  assign n8694 = n728 & n2698 ;
  assign n8695 = n8694 ^ n6327 ^ 1'b0 ;
  assign n8696 = n8695 ^ n2856 ^ 1'b0 ;
  assign n8697 = n5970 ^ n3879 ^ 1'b0 ;
  assign n8698 = n5929 & ~n6851 ;
  assign n8699 = x26 | n1216 ;
  assign n8700 = n8699 ^ x4 ^ 1'b0 ;
  assign n8701 = ~n1188 & n1372 ;
  assign n8702 = n8701 ^ n1006 ^ 1'b0 ;
  assign n8703 = ~n1037 & n8406 ;
  assign n8704 = ~n903 & n8295 ;
  assign n8705 = n1023 ^ x214 ^ 1'b0 ;
  assign n8706 = n2475 & n8705 ;
  assign n8707 = n3255 & n8706 ;
  assign n8708 = n5105 ^ n3616 ^ 1'b0 ;
  assign n8709 = ~n580 & n8708 ;
  assign n8710 = n7907 ^ n858 ^ 1'b0 ;
  assign n8711 = n4112 | n7325 ;
  assign n8712 = n5751 & n8711 ;
  assign n8713 = n8712 ^ n7536 ^ 1'b0 ;
  assign n8714 = n3456 ^ n3042 ^ 1'b0 ;
  assign n8715 = n2498 & ~n8714 ;
  assign n8716 = ~n744 & n8715 ;
  assign n8717 = n1757 & ~n1806 ;
  assign n8718 = ~n2412 & n8717 ;
  assign n8719 = n8718 ^ n897 ^ 1'b0 ;
  assign n8720 = n2861 | n8719 ;
  assign n8721 = n4578 | n8720 ;
  assign n8722 = n6625 ^ n1048 ^ 1'b0 ;
  assign n8723 = n6885 ^ n4313 ^ 1'b0 ;
  assign n8724 = n8722 | n8723 ;
  assign n8726 = n4995 ^ n456 ^ 1'b0 ;
  assign n8727 = n1045 & n8726 ;
  assign n8725 = n4708 ^ n4442 ^ 1'b0 ;
  assign n8728 = n8727 ^ n8725 ^ 1'b0 ;
  assign n8729 = n8728 ^ n7193 ^ 1'b0 ;
  assign n8730 = n830 ^ n708 ^ 1'b0 ;
  assign n8731 = n3700 | n8730 ;
  assign n8732 = n4378 ^ n1689 ^ 1'b0 ;
  assign n8733 = n302 & ~n8732 ;
  assign n8734 = x228 & n8733 ;
  assign n8735 = n4338 & n5435 ;
  assign n8736 = n1671 ^ n629 ^ 1'b0 ;
  assign n8737 = ~n1383 & n8736 ;
  assign n8738 = n2141 & n8737 ;
  assign n8739 = n8738 ^ n1856 ^ 1'b0 ;
  assign n8740 = n720 & n8739 ;
  assign n8741 = n5337 ^ n2672 ^ 1'b0 ;
  assign n8742 = n6423 | n8741 ;
  assign n8743 = n2714 & n8742 ;
  assign n8744 = n4834 ^ n987 ^ 1'b0 ;
  assign n8745 = ~n7408 & n8744 ;
  assign n8746 = n8745 ^ n2698 ^ 1'b0 ;
  assign n8747 = ~n6365 & n8746 ;
  assign n8748 = n1775 & ~n7097 ;
  assign n8749 = n985 | n8748 ;
  assign n8750 = n8749 ^ n2218 ^ 1'b0 ;
  assign n8751 = ~n2852 & n6998 ;
  assign n8752 = n8352 & n8751 ;
  assign n8755 = n4015 ^ n1330 ^ 1'b0 ;
  assign n8756 = ~n701 & n8755 ;
  assign n8757 = n6886 ^ n4989 ^ 1'b0 ;
  assign n8758 = n8756 & n8757 ;
  assign n8753 = n4406 ^ n2476 ^ 1'b0 ;
  assign n8754 = n3288 | n8753 ;
  assign n8759 = n8758 ^ n8754 ^ 1'b0 ;
  assign n8760 = n8409 ^ n8223 ^ 1'b0 ;
  assign n8761 = n2527 & ~n8760 ;
  assign n8762 = ~n2796 & n3353 ;
  assign n8763 = ~n8097 & n8762 ;
  assign n8764 = n7997 & n8763 ;
  assign n8765 = n749 ^ n718 ^ 1'b0 ;
  assign n8766 = n6288 & ~n8765 ;
  assign n8767 = n8766 ^ n8307 ^ 1'b0 ;
  assign n8768 = n5253 ^ x241 ^ 1'b0 ;
  assign n8769 = n7528 ^ x246 ^ 1'b0 ;
  assign n8770 = n3791 & ~n8769 ;
  assign n8771 = ~n6951 & n8770 ;
  assign n8772 = n4388 & ~n4871 ;
  assign n8773 = x104 & x143 ;
  assign n8774 = ~n8772 & n8773 ;
  assign n8775 = ~n4021 & n6178 ;
  assign n8776 = n8775 ^ n3336 ^ 1'b0 ;
  assign n8777 = ~n339 & n575 ;
  assign n8778 = ~n575 & n8777 ;
  assign n8779 = n4246 & ~n8778 ;
  assign n8780 = n8778 & n8779 ;
  assign n8781 = n423 & ~n440 ;
  assign n8782 = n440 & n8781 ;
  assign n8783 = x94 & x223 ;
  assign n8784 = ~x94 & n8783 ;
  assign n8785 = n2040 & ~n8784 ;
  assign n8786 = ~n8782 & n8785 ;
  assign n8787 = n8780 & n8786 ;
  assign n8788 = n8776 & ~n8787 ;
  assign n8789 = ~n8776 & n8788 ;
  assign n8790 = n5784 & ~n8789 ;
  assign n8791 = ~n5784 & n8790 ;
  assign n8792 = n5945 ^ n5400 ^ 1'b0 ;
  assign n8793 = n4333 & n8767 ;
  assign n8794 = x21 & n4865 ;
  assign n8795 = n8794 ^ n7117 ^ 1'b0 ;
  assign n8796 = n8721 & ~n8795 ;
  assign n8797 = n3024 | n7881 ;
  assign n8798 = ~n4995 & n8797 ;
  assign n8799 = ~n7321 & n8798 ;
  assign n8800 = n1997 ^ x156 ^ 1'b0 ;
  assign n8801 = ~n2162 & n8800 ;
  assign n8802 = ~n418 & n8801 ;
  assign n8803 = n8802 ^ n994 ^ 1'b0 ;
  assign n8804 = n8803 ^ n6059 ^ 1'b0 ;
  assign n8805 = x95 & ~n2187 ;
  assign n8806 = ~n1604 & n8805 ;
  assign n8807 = n8806 ^ n1938 ^ 1'b0 ;
  assign n8808 = x137 & ~n8807 ;
  assign n8809 = n8808 ^ n3807 ^ 1'b0 ;
  assign n8810 = n3053 ^ n1333 ^ 1'b0 ;
  assign n8811 = x99 & n8810 ;
  assign n8812 = n8811 ^ n5286 ^ 1'b0 ;
  assign n8813 = n6580 & ~n8812 ;
  assign n8814 = ~n2463 & n8813 ;
  assign n8815 = n8307 ^ n6014 ^ 1'b0 ;
  assign n8816 = n8200 | n8815 ;
  assign n8817 = n1749 & ~n2895 ;
  assign n8818 = n8817 ^ n7376 ^ 1'b0 ;
  assign n8819 = n6446 & n8818 ;
  assign n8820 = n3410 | n3845 ;
  assign n8821 = n6721 ^ n703 ^ 1'b0 ;
  assign n8822 = n8821 ^ n2423 ^ 1'b0 ;
  assign n8823 = n7039 & n8822 ;
  assign n8824 = n8503 & ~n8765 ;
  assign n8825 = ~n8823 & n8824 ;
  assign n8826 = ~n3195 & n3322 ;
  assign n8827 = ~n2466 & n8826 ;
  assign n8828 = n7771 ^ n1472 ^ 1'b0 ;
  assign n8829 = n8827 | n8828 ;
  assign n8830 = n8829 ^ n7570 ^ x187 ;
  assign n8831 = n754 & n4278 ;
  assign n8832 = ~n4645 & n8831 ;
  assign n8833 = x92 & ~n527 ;
  assign n8834 = ~n4671 & n8833 ;
  assign n8835 = n5673 & ~n5739 ;
  assign n8836 = n1857 & ~n7118 ;
  assign n8837 = ( n593 & ~n1004 ) | ( n593 & n8836 ) | ( ~n1004 & n8836 ) ;
  assign n8839 = n3528 | n4173 ;
  assign n8840 = n354 | n8839 ;
  assign n8838 = n1400 & ~n3624 ;
  assign n8841 = n8840 ^ n8838 ^ 1'b0 ;
  assign n8842 = n1701 & n5792 ;
  assign n8843 = n6433 ^ n5091 ^ 1'b0 ;
  assign n8844 = n6807 ^ n1503 ^ 1'b0 ;
  assign n8845 = n8843 & n8844 ;
  assign n8846 = n985 & n8845 ;
  assign n8849 = ~n514 & n607 ;
  assign n8847 = n5849 ^ n1125 ^ 1'b0 ;
  assign n8848 = n2476 & ~n8847 ;
  assign n8850 = n8849 ^ n8848 ^ 1'b0 ;
  assign n8851 = ~n3688 & n4680 ;
  assign n8853 = ( n2274 & n4230 ) | ( n2274 & n4580 ) | ( n4230 & n4580 ) ;
  assign n8854 = ~n4625 & n8853 ;
  assign n8852 = n1643 & n2498 ;
  assign n8855 = n8854 ^ n8852 ^ 1'b0 ;
  assign n8856 = x207 & n4664 ;
  assign n8857 = n2031 | n3580 ;
  assign n8858 = n2031 & ~n8857 ;
  assign n8859 = n791 & ~n8858 ;
  assign n8860 = ~n791 & n8859 ;
  assign n8861 = ~n1102 & n4283 ;
  assign n8862 = n8860 & n8861 ;
  assign n8863 = n608 | n685 ;
  assign n8864 = n685 & ~n8863 ;
  assign n8865 = n625 | n8864 ;
  assign n8866 = n8864 & ~n8865 ;
  assign n8867 = n6744 & ~n8866 ;
  assign n8868 = n8866 & n8867 ;
  assign n8869 = n8862 | n8868 ;
  assign n8870 = n8862 & ~n8869 ;
  assign n8875 = n707 & n6116 ;
  assign n8876 = n2120 & ~n8875 ;
  assign n8871 = n1738 & ~n4267 ;
  assign n8872 = ~n2755 & n8871 ;
  assign n8873 = ~n5826 & n8872 ;
  assign n8874 = x7 & ~n8873 ;
  assign n8877 = n8876 ^ n8874 ^ n6202 ;
  assign n8878 = n8303 ^ n1628 ^ 1'b0 ;
  assign n8879 = n4756 & n8878 ;
  assign n8880 = n1156 ^ n468 ^ 1'b0 ;
  assign n8881 = ~n5163 & n8880 ;
  assign n8887 = n1243 & ~n2543 ;
  assign n8882 = n7321 ^ x151 ^ 1'b0 ;
  assign n8883 = n3833 & n8882 ;
  assign n8884 = n3524 ^ n3247 ^ 1'b0 ;
  assign n8885 = ~n4063 & n8884 ;
  assign n8886 = n8883 & n8885 ;
  assign n8888 = n8887 ^ n8886 ^ 1'b0 ;
  assign n8889 = n4063 & ~n7496 ;
  assign n8890 = n6015 ^ n4731 ^ 1'b0 ;
  assign n8891 = n8890 ^ n1038 ^ 1'b0 ;
  assign n8892 = x177 & ~n8891 ;
  assign n8893 = ~n6267 & n6464 ;
  assign n8894 = n2066 & n5284 ;
  assign n8895 = n1926 ^ n357 ^ 1'b0 ;
  assign n8896 = ~n8894 & n8895 ;
  assign n8897 = n7023 ^ n4169 ^ 1'b0 ;
  assign n8898 = n2437 & ~n4751 ;
  assign n8899 = n8898 ^ n1184 ^ 1'b0 ;
  assign n8900 = n8899 ^ n2784 ^ 1'b0 ;
  assign n8901 = n3983 | n8900 ;
  assign n8902 = n3558 ^ x175 ^ 1'b0 ;
  assign n8903 = n8801 & ~n8902 ;
  assign n8904 = n800 & ~n5150 ;
  assign n8905 = ~n8903 & n8904 ;
  assign n8906 = n7982 ^ n5723 ^ 1'b0 ;
  assign n8907 = n5585 & ~n8906 ;
  assign n8908 = n2844 ^ n1447 ^ 1'b0 ;
  assign n8909 = n8908 ^ n6768 ^ 1'b0 ;
  assign n8910 = n3869 & n6635 ;
  assign n8911 = n3825 ^ n322 ^ 1'b0 ;
  assign n8912 = n1899 & n8911 ;
  assign n8913 = n8453 ^ n7984 ^ 1'b0 ;
  assign n8914 = n5357 ^ n954 ^ 1'b0 ;
  assign n8915 = ~n8328 & n8914 ;
  assign n8916 = n8915 ^ n5833 ^ 1'b0 ;
  assign n8917 = n4644 & ~n6252 ;
  assign n8918 = n8917 ^ n8305 ^ 1'b0 ;
  assign n8919 = ~n2143 & n2827 ;
  assign n8922 = n4140 ^ n3901 ^ 1'b0 ;
  assign n8920 = ~n6160 & n6521 ;
  assign n8921 = n7411 & n8920 ;
  assign n8923 = n8922 ^ n8921 ^ n8389 ;
  assign n8924 = n7497 & n8219 ;
  assign n8925 = ~n1529 & n8924 ;
  assign n8926 = x141 & n5125 ;
  assign n8927 = n3606 & n8926 ;
  assign n8928 = n8927 ^ n7741 ^ 1'b0 ;
  assign n8929 = n8928 ^ n5261 ^ n3323 ;
  assign n8930 = n6583 ^ n421 ^ 1'b0 ;
  assign n8931 = n8309 ^ n1264 ^ n1075 ;
  assign n8932 = n8930 | n8931 ;
  assign n8933 = ( n1914 & ~n5296 ) | ( n1914 & n6482 ) | ( ~n5296 & n6482 ) ;
  assign n8934 = n3974 & n4905 ;
  assign n8935 = n8934 ^ n6938 ^ 1'b0 ;
  assign n8936 = n4780 | n8935 ;
  assign n8937 = n8936 ^ n1896 ^ 1'b0 ;
  assign n8938 = n3715 ^ n1658 ^ 1'b0 ;
  assign n8939 = ~n3850 & n8938 ;
  assign n8940 = n1593 ^ n309 ^ 1'b0 ;
  assign n8941 = n1738 | n8940 ;
  assign n8942 = n3862 & n8941 ;
  assign n8943 = x132 & n3737 ;
  assign n8944 = n8943 ^ n4955 ^ 1'b0 ;
  assign n8945 = ( ~n1339 & n2074 ) | ( ~n1339 & n8944 ) | ( n2074 & n8944 ) ;
  assign n8948 = n3137 & ~n4111 ;
  assign n8947 = n452 ^ n370 ^ 1'b0 ;
  assign n8949 = n8948 ^ n8947 ^ 1'b0 ;
  assign n8950 = x184 & n8949 ;
  assign n8946 = n6587 & n7301 ;
  assign n8951 = n8950 ^ n8946 ^ 1'b0 ;
  assign n8952 = n8108 & ~n8951 ;
  assign n8953 = n3549 & n8952 ;
  assign n8954 = ~n1754 & n4737 ;
  assign n8955 = n8954 ^ n4094 ^ 1'b0 ;
  assign n8956 = n4094 & n8955 ;
  assign n8957 = ~n3736 & n8956 ;
  assign n8958 = n1831 & ~n3411 ;
  assign n8959 = n8958 ^ n2613 ^ 1'b0 ;
  assign n8960 = n1709 & ~n2903 ;
  assign n8963 = n7408 ^ n3855 ^ 1'b0 ;
  assign n8961 = n4978 & n6490 ;
  assign n8962 = n8961 ^ n5223 ^ 1'b0 ;
  assign n8964 = n8963 ^ n8962 ^ 1'b0 ;
  assign n8965 = ~n2861 & n3727 ;
  assign n8966 = n8965 ^ n6791 ^ 1'b0 ;
  assign n8967 = n7200 | n8966 ;
  assign n8968 = n1671 & ~n3729 ;
  assign n8969 = n8968 ^ n4534 ^ 1'b0 ;
  assign n8970 = n1169 & ~n8969 ;
  assign n8971 = n2074 & ~n8970 ;
  assign n8972 = n8971 ^ n969 ^ 1'b0 ;
  assign n8973 = n2065 ^ n1697 ^ 1'b0 ;
  assign n8974 = n2395 & ~n8973 ;
  assign n8975 = n8974 ^ n4027 ^ 1'b0 ;
  assign n8976 = ~n320 & n8975 ;
  assign n8986 = ~n1239 & n1540 ;
  assign n8987 = ~n1540 & n8986 ;
  assign n8988 = n8987 ^ n5026 ^ 1'b0 ;
  assign n8977 = n3620 ^ x148 ^ 1'b0 ;
  assign n8978 = n1704 & n3794 ;
  assign n8979 = n8977 | n8978 ;
  assign n8980 = n8977 & ~n8979 ;
  assign n8981 = n1663 & ~n3657 ;
  assign n8982 = n8980 & n8981 ;
  assign n8983 = n4949 | n7217 ;
  assign n8984 = n7217 & ~n8983 ;
  assign n8985 = n8982 | n8984 ;
  assign n8989 = n8988 ^ n8985 ^ 1'b0 ;
  assign n8990 = n3255 & n8602 ;
  assign n8991 = n1325 ^ n974 ^ 1'b0 ;
  assign n8992 = n1094 & ~n8991 ;
  assign n8993 = n8329 & ~n8992 ;
  assign n8994 = n7029 & n7243 ;
  assign n8995 = n8994 ^ n4314 ^ 1'b0 ;
  assign n8996 = n8995 ^ n4300 ^ 1'b0 ;
  assign n8997 = n3184 | n8996 ;
  assign n8999 = ~n994 & n2753 ;
  assign n9000 = n8999 ^ n3067 ^ 1'b0 ;
  assign n8998 = ~x223 & n4857 ;
  assign n9001 = n9000 ^ n8998 ^ 1'b0 ;
  assign n9002 = n1867 ^ n1073 ^ 1'b0 ;
  assign n9003 = n6071 | n9002 ;
  assign n9004 = n6757 ^ n5401 ^ n4652 ;
  assign n9005 = x22 | n707 ;
  assign n9006 = n2761 ^ x34 ^ 1'b0 ;
  assign n9007 = n9006 ^ n7497 ^ 1'b0 ;
  assign n9008 = n1931 | n3736 ;
  assign n9009 = n9008 ^ n686 ^ 1'b0 ;
  assign n9010 = n9007 & ~n9009 ;
  assign n9011 = n1779 & n4176 ;
  assign n9012 = n8309 ^ n6408 ^ 1'b0 ;
  assign n9013 = n4764 ^ n3687 ^ 1'b0 ;
  assign n9014 = n9013 ^ n4164 ^ 1'b0 ;
  assign n9015 = n9012 & n9014 ;
  assign n9016 = n3499 ^ n942 ^ 1'b0 ;
  assign n9017 = n6560 ^ n6399 ^ 1'b0 ;
  assign n9018 = n9016 & ~n9017 ;
  assign n9019 = n891 | n8930 ;
  assign n9023 = n4775 ^ n4005 ^ 1'b0 ;
  assign n9024 = n723 & ~n9023 ;
  assign n9025 = n4397 & ~n9024 ;
  assign n9020 = n4491 & ~n7098 ;
  assign n9021 = n9020 ^ n1657 ^ 1'b0 ;
  assign n9022 = ~n2006 & n9021 ;
  assign n9026 = n9025 ^ n9022 ^ 1'b0 ;
  assign n9027 = n887 & ~n2776 ;
  assign n9033 = n4694 ^ n725 ^ 1'b0 ;
  assign n9031 = ~n2632 & n6566 ;
  assign n9032 = n9031 ^ n331 ^ 1'b0 ;
  assign n9034 = n9033 ^ n9032 ^ 1'b0 ;
  assign n9028 = n2124 & n6985 ;
  assign n9029 = n9028 ^ n2324 ^ 1'b0 ;
  assign n9030 = n5269 & ~n9029 ;
  assign n9035 = n9034 ^ n9030 ^ 1'b0 ;
  assign n9037 = n6199 ^ n2082 ^ 1'b0 ;
  assign n9038 = n2485 | n9037 ;
  assign n9039 = n4003 & ~n9038 ;
  assign n9036 = n1825 & n4833 ;
  assign n9040 = n9039 ^ n9036 ^ 1'b0 ;
  assign n9041 = ( n4152 & n6325 ) | ( n4152 & ~n9040 ) | ( n6325 & ~n9040 ) ;
  assign n9042 = ~n641 & n1033 ;
  assign n9043 = n623 & n9042 ;
  assign n9044 = n9043 ^ n8025 ^ 1'b0 ;
  assign n9045 = ~n7257 & n9044 ;
  assign n9046 = n643 & n2018 ;
  assign n9047 = n9046 ^ n957 ^ 1'b0 ;
  assign n9048 = n3209 & ~n9047 ;
  assign n9049 = n9048 ^ n6548 ^ 1'b0 ;
  assign n9050 = n8345 ^ n1969 ^ 1'b0 ;
  assign n9051 = n6355 ^ n561 ^ 1'b0 ;
  assign n9052 = n3995 & n9051 ;
  assign n9053 = n5457 | n9052 ;
  assign n9054 = ~n9050 & n9053 ;
  assign n9055 = ~n1854 & n9054 ;
  assign n9056 = n1293 | n4771 ;
  assign n9057 = n9056 ^ n5557 ^ 1'b0 ;
  assign n9058 = n760 & ~n1871 ;
  assign n9059 = ~n4253 & n9058 ;
  assign n9060 = n1893 & ~n2146 ;
  assign n9061 = n1991 | n6169 ;
  assign n9062 = n1979 & n4144 ;
  assign n9063 = n1139 ^ n1056 ^ n749 ;
  assign n9064 = n4455 ^ n1740 ^ 1'b0 ;
  assign n9065 = n5587 & ~n9064 ;
  assign n9068 = n1395 | n3386 ;
  assign n9069 = n9068 ^ n4327 ^ 1'b0 ;
  assign n9070 = n9069 ^ n1459 ^ 1'b0 ;
  assign n9071 = n827 & n9070 ;
  assign n9066 = n836 ^ x169 ^ 1'b0 ;
  assign n9067 = n6840 | n9066 ;
  assign n9072 = n9071 ^ n9067 ^ 1'b0 ;
  assign n9073 = n5361 ^ n1944 ^ 1'b0 ;
  assign n9074 = n9073 ^ n2865 ^ 1'b0 ;
  assign n9075 = n4376 & ~n8572 ;
  assign n9076 = x225 | n2219 ;
  assign n9077 = n376 & ~n1366 ;
  assign n9078 = ~n3074 & n9077 ;
  assign n9079 = n2099 ^ n1617 ^ 1'b0 ;
  assign n9080 = n3599 | n9079 ;
  assign n9081 = n2972 ^ n552 ^ 1'b0 ;
  assign n9082 = ~n1453 & n6752 ;
  assign n9083 = ~n7037 & n9082 ;
  assign n9084 = n4430 & ~n7416 ;
  assign n9085 = ( n281 & n6620 ) | ( n281 & n6772 ) | ( n6620 & n6772 ) ;
  assign n9086 = ~n3198 & n3672 ;
  assign n9087 = ( ~n2443 & n3601 ) | ( ~n2443 & n4301 ) | ( n3601 & n4301 ) ;
  assign n9088 = n7395 ^ n2863 ^ 1'b0 ;
  assign n9089 = n9087 & ~n9088 ;
  assign n9090 = n3603 ^ n2482 ^ 1'b0 ;
  assign n9091 = n8645 & ~n9090 ;
  assign n9092 = ~n9089 & n9091 ;
  assign n9093 = x100 & ~n7123 ;
  assign n9094 = n9093 ^ n4416 ^ 1'b0 ;
  assign n9095 = n3999 & ~n9094 ;
  assign n9096 = n6311 ^ n5551 ^ 1'b0 ;
  assign n9097 = n3033 & n9096 ;
  assign n9098 = n7362 & n8440 ;
  assign n9099 = n9098 ^ n3305 ^ 1'b0 ;
  assign n9100 = n7255 ^ n930 ^ 1'b0 ;
  assign n9101 = ~n2072 & n6715 ;
  assign n9102 = n6655 ^ n901 ^ 1'b0 ;
  assign n9103 = ~n1344 & n9102 ;
  assign n9104 = ( ~n2889 & n3068 ) | ( ~n2889 & n7622 ) | ( n3068 & n7622 ) ;
  assign n9105 = n3027 ^ n1843 ^ 1'b0 ;
  assign n9106 = n4108 ^ n1143 ^ 1'b0 ;
  assign n9107 = n9106 ^ n5492 ^ 1'b0 ;
  assign n9108 = n8776 & ~n9107 ;
  assign n9109 = n4764 ^ n2495 ^ 1'b0 ;
  assign n9110 = n6032 ^ n2075 ^ 1'b0 ;
  assign n9111 = n3711 | n9110 ;
  assign n9112 = n4686 | n9111 ;
  assign n9113 = n1541 | n9112 ;
  assign n9114 = n9113 ^ n1380 ^ 1'b0 ;
  assign n9115 = n4399 ^ n854 ^ 1'b0 ;
  assign n9116 = ~n8491 & n9115 ;
  assign n9117 = ~x186 & n9116 ;
  assign n9118 = n478 | n4546 ;
  assign n9119 = ~n5030 & n5141 ;
  assign n9120 = n722 & n1779 ;
  assign n9121 = ~n4068 & n9120 ;
  assign n9122 = n4169 & n9121 ;
  assign n9123 = n4982 & n5900 ;
  assign n9124 = ~n9122 & n9123 ;
  assign n9125 = ~n9119 & n9124 ;
  assign n9126 = x67 | n6169 ;
  assign n9127 = n2933 | n3860 ;
  assign n9128 = n5869 | n9127 ;
  assign n9129 = n5622 ^ n2938 ^ n1299 ;
  assign n9130 = n6039 ^ n2307 ^ 1'b0 ;
  assign n9131 = n3480 & n9130 ;
  assign n9132 = n9131 ^ n3855 ^ 1'b0 ;
  assign n9133 = ~n3466 & n7367 ;
  assign n9134 = n776 & n1385 ;
  assign n9135 = n3403 & n9134 ;
  assign n9136 = n4849 | n9135 ;
  assign n9137 = n9133 & ~n9136 ;
  assign n9138 = n6759 & ~n9137 ;
  assign n9139 = ~n5392 & n9138 ;
  assign n9140 = n1533 ^ n1271 ^ 1'b0 ;
  assign n9141 = n7248 & ~n9140 ;
  assign n9142 = n267 & n7115 ;
  assign n9143 = n9142 ^ n1820 ^ 1'b0 ;
  assign n9144 = n3578 & n9143 ;
  assign n9145 = x104 & n6416 ;
  assign n9146 = n9145 ^ n7591 ^ 1'b0 ;
  assign n9147 = ~n3184 & n4031 ;
  assign n9148 = n7271 & n9147 ;
  assign n9149 = n8419 ^ n3537 ^ 1'b0 ;
  assign n9150 = n5566 ^ n854 ^ 1'b0 ;
  assign n9151 = n9150 ^ n1479 ^ 1'b0 ;
  assign n9152 = n9149 & ~n9151 ;
  assign n9153 = n5639 & n6993 ;
  assign n9154 = n2609 & ~n6195 ;
  assign n9155 = n3083 & ~n4568 ;
  assign n9156 = n9155 ^ n3780 ^ 1'b0 ;
  assign n9157 = n1537 | n9156 ;
  assign n9158 = n9157 ^ n1910 ^ 1'b0 ;
  assign n9159 = n3295 & ~n9158 ;
  assign n9160 = n9159 ^ n3856 ^ 1'b0 ;
  assign n9161 = n1080 & n5146 ;
  assign n9162 = ~n2119 & n9161 ;
  assign n9163 = n8722 ^ n2681 ^ 1'b0 ;
  assign n9164 = n2517 & n9163 ;
  assign n9165 = ~n5645 & n9164 ;
  assign n9166 = n691 | n9165 ;
  assign n9167 = ( n5579 & n9162 ) | ( n5579 & n9166 ) | ( n9162 & n9166 ) ;
  assign n9168 = ~n1926 & n5036 ;
  assign n9169 = ~n8317 & n9168 ;
  assign n9170 = n9169 ^ n7692 ^ 1'b0 ;
  assign n9171 = n2286 & n5379 ;
  assign n9172 = n9171 ^ n5519 ^ 1'b0 ;
  assign n9173 = x235 & n9172 ;
  assign n9174 = x249 | n3336 ;
  assign n9175 = n9174 ^ n2331 ^ 1'b0 ;
  assign n9176 = n844 & n3216 ;
  assign n9177 = ~n3047 & n5356 ;
  assign n9178 = n7079 ^ n3093 ^ n2997 ;
  assign n9179 = n9178 ^ n965 ^ 1'b0 ;
  assign n9180 = n9177 | n9179 ;
  assign n9181 = n9152 | n9180 ;
  assign n9182 = x206 & n5950 ;
  assign n9183 = ~n3057 & n9182 ;
  assign n9184 = ( n4502 & ~n4678 ) | ( n4502 & n9183 ) | ( ~n4678 & n9183 ) ;
  assign n9185 = ~n651 & n1159 ;
  assign n9186 = ~n840 & n9185 ;
  assign n9187 = x181 & ~n3336 ;
  assign n9188 = n9187 ^ n1562 ^ 1'b0 ;
  assign n9189 = ~n1124 & n9188 ;
  assign n9190 = ~n4289 & n9189 ;
  assign n9191 = n5922 ^ x73 ^ 1'b0 ;
  assign n9192 = ~n1395 & n9191 ;
  assign n9193 = n9192 ^ n2001 ^ 1'b0 ;
  assign n9194 = n9193 ^ n1810 ^ 1'b0 ;
  assign n9195 = n3984 ^ n349 ^ 1'b0 ;
  assign n9196 = n1630 & ~n2070 ;
  assign n9197 = n8708 ^ n6951 ^ 1'b0 ;
  assign n9198 = ~n1192 & n4888 ;
  assign n9199 = n9198 ^ x214 ^ 1'b0 ;
  assign n9200 = n5235 & ~n9199 ;
  assign n9201 = ~n1094 & n9200 ;
  assign n9202 = n4576 | n9201 ;
  assign n9203 = n4448 | n9202 ;
  assign n9204 = ~n965 & n4954 ;
  assign n9205 = ~n4521 & n9204 ;
  assign n9206 = x226 | n7300 ;
  assign n9207 = n1912 & n9206 ;
  assign n9208 = n4075 ^ n2035 ^ 1'b0 ;
  assign n9209 = x87 & ~n4225 ;
  assign n9210 = n3540 & n9209 ;
  assign n9211 = n9208 | n9210 ;
  assign n9212 = ~n354 & n5229 ;
  assign n9213 = n3735 & ~n7109 ;
  assign n9214 = n1260 ^ x142 ^ 1'b0 ;
  assign n9215 = n1575 | n7169 ;
  assign n9216 = n9215 ^ n1255 ^ 1'b0 ;
  assign n9217 = x92 & n9216 ;
  assign n9218 = n3073 & ~n3195 ;
  assign n9219 = n7015 & n9218 ;
  assign n9220 = n7836 ^ x182 ^ 1'b0 ;
  assign n9221 = n4804 | n9220 ;
  assign n9222 = ~n9219 & n9221 ;
  assign n9223 = n341 ^ x217 ^ 1'b0 ;
  assign n9224 = n4318 | n9223 ;
  assign n9225 = x17 | n9224 ;
  assign n9226 = x233 & ~n4803 ;
  assign n9227 = n9226 ^ n6676 ^ 1'b0 ;
  assign n9228 = ~n7674 & n8693 ;
  assign n9229 = n9228 ^ n2281 ^ 1'b0 ;
  assign n9230 = n9229 ^ n5662 ^ 1'b0 ;
  assign n9231 = n1864 & n9230 ;
  assign n9232 = n2951 ^ n1324 ^ 1'b0 ;
  assign n9233 = n4691 ^ n1156 ^ 1'b0 ;
  assign n9234 = n2014 & n3687 ;
  assign n9235 = n1423 & n8738 ;
  assign n9236 = n9235 ^ n4142 ^ 1'b0 ;
  assign n9237 = n9236 ^ n3112 ^ 1'b0 ;
  assign n9238 = ~n9234 & n9237 ;
  assign n9243 = n2158 ^ n574 ^ 1'b0 ;
  assign n9239 = n1237 ^ n1176 ^ 1'b0 ;
  assign n9240 = n9239 ^ n5519 ^ 1'b0 ;
  assign n9241 = n6058 & n9240 ;
  assign n9242 = n9241 ^ n3678 ^ 1'b0 ;
  assign n9244 = n9243 ^ n9242 ^ 1'b0 ;
  assign n9245 = n3780 ^ n3628 ^ 1'b0 ;
  assign n9246 = n6246 & n9245 ;
  assign n9247 = n9246 ^ n3419 ^ 1'b0 ;
  assign n9248 = n2158 | n9247 ;
  assign n9249 = n7681 ^ n4971 ^ 1'b0 ;
  assign n9250 = n5896 | n9249 ;
  assign n9251 = n504 & ~n6739 ;
  assign n9252 = n3501 | n9251 ;
  assign n9254 = n2715 ^ n1625 ^ n694 ;
  assign n9255 = n1728 ^ n1075 ^ 1'b0 ;
  assign n9256 = n9254 & ~n9255 ;
  assign n9253 = ~n2333 & n5559 ;
  assign n9257 = n9256 ^ n9253 ^ 1'b0 ;
  assign n9258 = ~n623 & n9257 ;
  assign n9259 = n9258 ^ n2078 ^ 1'b0 ;
  assign n9260 = n394 | n4579 ;
  assign n9261 = ~n1102 & n9260 ;
  assign n9262 = n8795 & ~n9261 ;
  assign n9263 = ~n9259 & n9262 ;
  assign n9264 = n7608 ^ n4605 ^ 1'b0 ;
  assign n9265 = n707 & ~n6074 ;
  assign n9266 = n9265 ^ n2018 ^ 1'b0 ;
  assign n9267 = n9266 ^ n2474 ^ 1'b0 ;
  assign n9270 = ~x226 & n1249 ;
  assign n9268 = n3454 & ~n3991 ;
  assign n9269 = n9268 ^ n7793 ^ 1'b0 ;
  assign n9271 = n9270 ^ n9269 ^ 1'b0 ;
  assign n9272 = n791 & n9271 ;
  assign n9275 = n1236 | n3822 ;
  assign n9276 = n9275 ^ n1159 ^ 1'b0 ;
  assign n9273 = n3741 & n8523 ;
  assign n9274 = n1496 & n9273 ;
  assign n9277 = n9276 ^ n9274 ^ 1'b0 ;
  assign n9278 = ~n1290 & n1527 ;
  assign n9279 = ( n1563 & n7164 ) | ( n1563 & ~n9278 ) | ( n7164 & ~n9278 ) ;
  assign n9280 = n633 | n7314 ;
  assign n9281 = n9280 ^ n2089 ^ 1'b0 ;
  assign n9283 = ~n1156 & n1867 ;
  assign n9284 = n9283 ^ n7902 ^ n1154 ;
  assign n9282 = n1304 | n2001 ;
  assign n9285 = n9284 ^ n9282 ^ 1'b0 ;
  assign n9286 = ~n6647 & n9285 ;
  assign n9287 = n9286 ^ n8110 ^ 1'b0 ;
  assign n9288 = n1228 & n7627 ;
  assign n9289 = n9288 ^ n2333 ^ 1'b0 ;
  assign n9290 = n3976 & n9289 ;
  assign n9291 = n6065 ^ n3139 ^ 1'b0 ;
  assign n9294 = n4204 ^ n2364 ^ 1'b0 ;
  assign n9292 = n6568 ^ n2566 ^ 1'b0 ;
  assign n9293 = n4430 & ~n9292 ;
  assign n9295 = n9294 ^ n9293 ^ 1'b0 ;
  assign n9296 = n9295 ^ n8733 ^ n1328 ;
  assign n9298 = n5244 | n5779 ;
  assign n9299 = n9298 ^ n2820 ^ 1'b0 ;
  assign n9297 = n1854 & n6885 ;
  assign n9300 = n9299 ^ n9297 ^ 1'b0 ;
  assign n9301 = n4772 ^ n4180 ^ 1'b0 ;
  assign n9302 = n968 & ~n9301 ;
  assign n9303 = n5031 & n9302 ;
  assign n9304 = n6900 ^ n1080 ^ 1'b0 ;
  assign n9305 = n9304 ^ n5242 ^ 1'b0 ;
  assign n9306 = ( ~n814 & n7654 ) | ( ~n814 & n8076 ) | ( n7654 & n8076 ) ;
  assign n9307 = n3678 ^ n2587 ^ 1'b0 ;
  assign n9308 = n9307 ^ n8309 ^ 1'b0 ;
  assign n9309 = n5188 ^ n4476 ^ 1'b0 ;
  assign n9310 = ~n395 & n9309 ;
  assign n9311 = n8833 ^ n2315 ^ 1'b0 ;
  assign n9312 = n628 | n5985 ;
  assign n9313 = n9312 ^ n9018 ^ 1'b0 ;
  assign n9314 = n385 & ~n8836 ;
  assign n9315 = n9226 ^ n3073 ^ 1'b0 ;
  assign n9317 = n361 | n3145 ;
  assign n9318 = n1754 | n9317 ;
  assign n9319 = n9318 ^ n3995 ^ 1'b0 ;
  assign n9320 = n1653 & ~n9319 ;
  assign n9316 = n1399 | n4575 ;
  assign n9321 = n9320 ^ n9316 ^ 1'b0 ;
  assign n9322 = ~n573 & n5882 ;
  assign n9323 = n9322 ^ n5419 ^ 1'b0 ;
  assign n9324 = n9323 ^ n6106 ^ 1'b0 ;
  assign n9325 = n1241 | n6392 ;
  assign n9326 = n9325 ^ n7860 ^ 1'b0 ;
  assign n9327 = n426 & ~n3622 ;
  assign n9328 = n498 & ~n3308 ;
  assign n9329 = n864 & n9328 ;
  assign n9330 = ~n3532 & n5196 ;
  assign n9331 = ~n1264 & n9330 ;
  assign n9332 = n9329 | n9331 ;
  assign n9333 = n9332 ^ n1894 ^ 1'b0 ;
  assign n9334 = n9101 ^ n6838 ^ 1'b0 ;
  assign n9335 = n9333 & ~n9334 ;
  assign n9336 = n6606 ^ n2750 ^ 1'b0 ;
  assign n9337 = n3902 & n9336 ;
  assign n9338 = n4580 ^ n3234 ^ 1'b0 ;
  assign n9339 = ~n5445 & n9338 ;
  assign n9340 = n2384 | n9339 ;
  assign n9341 = n9340 ^ n8381 ^ 1'b0 ;
  assign n9342 = n2693 ^ n1773 ^ 1'b0 ;
  assign n9343 = ~n4211 & n9342 ;
  assign n9344 = n3795 | n5850 ;
  assign n9345 = n6456 & ~n7451 ;
  assign n9346 = n4652 & ~n9345 ;
  assign n9347 = n9346 ^ n3961 ^ 1'b0 ;
  assign n9348 = n3062 & n7126 ;
  assign n9349 = ~n9347 & n9348 ;
  assign n9350 = n7882 ^ n7190 ^ n3822 ;
  assign n9351 = n568 ^ n405 ^ 1'b0 ;
  assign n9352 = ~n1271 & n9351 ;
  assign n9354 = n2107 ^ n1451 ^ 1'b0 ;
  assign n9355 = x183 & ~n5984 ;
  assign n9356 = n9354 & n9355 ;
  assign n9357 = n1635 & ~n3165 ;
  assign n9358 = n3329 & n9357 ;
  assign n9359 = n9356 | n9358 ;
  assign n9360 = n907 & ~n9359 ;
  assign n9353 = ~n4203 & n7397 ;
  assign n9361 = n9360 ^ n9353 ^ n2660 ;
  assign n9362 = n9353 ^ n6400 ^ 1'b0 ;
  assign n9363 = ~n3226 & n9163 ;
  assign n9364 = ~n1334 & n3599 ;
  assign n9365 = n9364 ^ n8808 ^ 1'b0 ;
  assign n9366 = n6358 | n9365 ;
  assign n9367 = n6138 & ~n9366 ;
  assign n9368 = n8730 ^ n7421 ^ 1'b0 ;
  assign n9369 = x27 & n8369 ;
  assign n9370 = ~n6313 & n6562 ;
  assign n9371 = n7519 & n9370 ;
  assign n9372 = n3781 | n6200 ;
  assign n9373 = n9372 ^ n2591 ^ 1'b0 ;
  assign n9374 = n6885 ^ n820 ^ 1'b0 ;
  assign n9375 = n791 & n6617 ;
  assign n9376 = n9375 ^ n5348 ^ 1'b0 ;
  assign n9377 = n4372 & ~n5924 ;
  assign n9378 = ~n611 & n5837 ;
  assign n9379 = n967 & n1052 ;
  assign n9380 = ~n1850 & n9379 ;
  assign n9381 = n4972 | n9380 ;
  assign n9382 = ( n1404 & ~n5896 ) | ( n1404 & n8211 ) | ( ~n5896 & n8211 ) ;
  assign n9383 = n4459 ^ x66 ^ 1'b0 ;
  assign n9384 = n5835 | n9383 ;
  assign n9385 = n2180 | n9384 ;
  assign n9386 = n9385 ^ n4490 ^ 1'b0 ;
  assign n9387 = ~n2757 & n8065 ;
  assign n9388 = n3107 & n9387 ;
  assign n9389 = ~n3206 & n4351 ;
  assign n9390 = n9389 ^ n4701 ^ 1'b0 ;
  assign n9391 = n7542 | n9390 ;
  assign n9392 = n2928 & ~n4263 ;
  assign n9393 = n3931 & n9392 ;
  assign n9394 = ~n4603 & n4892 ;
  assign n9395 = n9313 ^ n6670 ^ 1'b0 ;
  assign n9396 = ~n1368 & n7029 ;
  assign n9397 = n3381 | n8728 ;
  assign n9398 = n9397 ^ n9375 ^ x27 ;
  assign n9399 = n2790 | n7648 ;
  assign n9400 = n1683 & ~n1694 ;
  assign n9401 = n5983 | n9400 ;
  assign n9402 = n2212 | n9401 ;
  assign n9406 = ~n1654 & n3405 ;
  assign n9407 = ~n5255 & n9406 ;
  assign n9403 = n6111 & n6716 ;
  assign n9404 = n9403 ^ n4488 ^ 1'b0 ;
  assign n9405 = n5955 & n9404 ;
  assign n9408 = n9407 ^ n9405 ^ 1'b0 ;
  assign n9409 = n7434 ^ n1334 ^ 1'b0 ;
  assign n9410 = ~n440 & n9409 ;
  assign n9411 = n9410 ^ n5152 ^ 1'b0 ;
  assign n9412 = n9408 & ~n9411 ;
  assign n9413 = n5902 | n7839 ;
  assign n9414 = n7326 ^ n1810 ^ 1'b0 ;
  assign n9415 = n1593 & n9414 ;
  assign n9416 = n315 | n2112 ;
  assign n9417 = n8733 & ~n9416 ;
  assign n9418 = ~n4493 & n5146 ;
  assign n9420 = n5672 ^ n3162 ^ 1'b0 ;
  assign n9419 = x196 & n3707 ;
  assign n9421 = n9420 ^ n9419 ^ 1'b0 ;
  assign n9422 = n8343 ^ n7057 ^ 1'b0 ;
  assign n9423 = n9421 & n9422 ;
  assign n9424 = ~n9418 & n9423 ;
  assign n9425 = n9424 ^ n6003 ^ 1'b0 ;
  assign n9426 = n3735 ^ n343 ^ 1'b0 ;
  assign n9427 = ~n341 & n9426 ;
  assign n9428 = n7611 ^ n4191 ^ 1'b0 ;
  assign n9429 = ~n3520 & n9428 ;
  assign n9430 = ~n3071 & n9429 ;
  assign n9431 = n7221 ^ n928 ^ 1'b0 ;
  assign n9432 = n8877 ^ n3458 ^ 1'b0 ;
  assign n9435 = x215 & n6882 ;
  assign n9436 = n9435 ^ n1345 ^ 1'b0 ;
  assign n9437 = n9436 ^ n7043 ^ n4393 ;
  assign n9433 = n1049 & n1622 ;
  assign n9434 = ~n5929 & n9433 ;
  assign n9438 = n9437 ^ n9434 ^ 1'b0 ;
  assign n9439 = n8612 ^ n3016 ^ 1'b0 ;
  assign n9440 = n2632 ^ n2314 ^ n2061 ;
  assign n9441 = n929 | n9440 ;
  assign n9442 = n9441 ^ n3862 ^ 1'b0 ;
  assign n9443 = ~n623 & n2871 ;
  assign n9444 = n9443 ^ n5360 ^ 1'b0 ;
  assign n9445 = n5343 & ~n9444 ;
  assign n9446 = n1850 & n7108 ;
  assign n9447 = ~n934 & n9446 ;
  assign n9448 = n3825 & n9447 ;
  assign n9449 = n1885 & ~n2004 ;
  assign n9450 = n9449 ^ n2972 ^ 1'b0 ;
  assign n9451 = ~n7058 & n9450 ;
  assign n9452 = n1648 & ~n3411 ;
  assign n9453 = ~x76 & n9452 ;
  assign n9454 = n8118 & n9453 ;
  assign n9455 = n840 | n1814 ;
  assign n9457 = n568 & ~n1769 ;
  assign n9458 = ~n1841 & n9457 ;
  assign n9459 = n2597 ^ n705 ^ 1'b0 ;
  assign n9460 = n2642 | n9459 ;
  assign n9461 = n3577 & ~n9460 ;
  assign n9462 = n9458 | n9461 ;
  assign n9463 = n9462 ^ n4734 ^ 1'b0 ;
  assign n9456 = n1825 & ~n3778 ;
  assign n9464 = n9463 ^ n9456 ^ 1'b0 ;
  assign n9465 = n9455 | n9464 ;
  assign n9466 = n6944 ^ n4440 ^ n1350 ;
  assign n9467 = n6241 & ~n9466 ;
  assign n9468 = n8127 & n9467 ;
  assign n9469 = n9371 ^ n5588 ^ 1'b0 ;
  assign n9470 = n1242 & n9469 ;
  assign n9471 = n7508 ^ n675 ^ 1'b0 ;
  assign n9472 = n9471 ^ n4195 ^ 1'b0 ;
  assign n9473 = n6927 | n9472 ;
  assign n9474 = n7933 | n8635 ;
  assign n9475 = n9474 ^ n5478 ^ 1'b0 ;
  assign n9476 = ~n2590 & n5629 ;
  assign n9477 = ~x195 & n9476 ;
  assign n9478 = n6702 | n9477 ;
  assign n9479 = n9478 ^ n2966 ^ 1'b0 ;
  assign n9480 = n6975 & ~n8237 ;
  assign n9481 = n9480 ^ n8047 ^ 1'b0 ;
  assign n9482 = ~n9301 & n9481 ;
  assign n9483 = x118 & ~n2987 ;
  assign n9484 = n2482 & ~n9483 ;
  assign n9485 = n5331 ^ n903 ^ 1'b0 ;
  assign n9486 = n9485 ^ n7507 ^ 1'b0 ;
  assign n9487 = ~n1510 & n9486 ;
  assign n9488 = n3495 & n5993 ;
  assign n9489 = ~x143 & n9488 ;
  assign n9490 = n9487 & ~n9489 ;
  assign n9491 = n7111 & n9490 ;
  assign n9492 = n927 | n9156 ;
  assign n9493 = ~x174 & n2149 ;
  assign n9494 = n6612 ^ n6229 ^ 1'b0 ;
  assign n9495 = n9493 & ~n9494 ;
  assign n9496 = n1835 ^ n1181 ^ 1'b0 ;
  assign n9497 = n2875 & n9496 ;
  assign n9498 = n7172 ^ n4133 ^ 1'b0 ;
  assign n9499 = n1275 & ~n9233 ;
  assign n9500 = n832 | n5525 ;
  assign n9501 = n7103 | n9500 ;
  assign n9502 = n9501 ^ n1164 ^ 1'b0 ;
  assign n9503 = n744 ^ n585 ^ 1'b0 ;
  assign n9504 = n1797 & n9503 ;
  assign n9505 = ~n1797 & n9504 ;
  assign n9506 = n7431 & ~n9505 ;
  assign n9507 = n9505 & n9506 ;
  assign n9508 = n3765 ^ x19 ^ 1'b0 ;
  assign n9509 = ~n9507 & n9508 ;
  assign n9510 = ~n1686 & n1977 ;
  assign n9511 = ~n1977 & n9510 ;
  assign n9512 = n4605 | n9511 ;
  assign n9513 = n8051 & ~n9512 ;
  assign n9514 = ~n9509 & n9513 ;
  assign n9515 = n1409 & ~n1897 ;
  assign n9516 = n1361 & n9515 ;
  assign n9517 = ( n3603 & n7345 ) | ( n3603 & ~n8298 ) | ( n7345 & ~n8298 ) ;
  assign n9521 = n3820 ^ n1370 ^ 1'b0 ;
  assign n9522 = n3373 & n9521 ;
  assign n9518 = n4934 ^ n2712 ^ 1'b0 ;
  assign n9519 = ~n4495 & n9518 ;
  assign n9520 = n1068 & n9519 ;
  assign n9523 = n9522 ^ n9520 ^ 1'b0 ;
  assign n9526 = n1360 & n5038 ;
  assign n9527 = n9526 ^ n1983 ^ 1'b0 ;
  assign n9524 = n7278 ^ n4594 ^ 1'b0 ;
  assign n9525 = n3175 | n9524 ;
  assign n9528 = n9527 ^ n9525 ^ 1'b0 ;
  assign n9529 = x99 & n2244 ;
  assign n9530 = n9529 ^ n1105 ^ 1'b0 ;
  assign n9531 = n5384 ^ n4416 ^ 1'b0 ;
  assign n9532 = n9530 | n9531 ;
  assign n9533 = n863 | n1694 ;
  assign n9534 = n928 | n9533 ;
  assign n9535 = n9534 ^ n4932 ^ n2715 ;
  assign n9536 = n1429 ^ x155 ^ 1'b0 ;
  assign n9537 = n6580 & n9536 ;
  assign n9538 = ~n729 & n1105 ;
  assign n9539 = n9538 ^ n4645 ^ 1'b0 ;
  assign n9540 = n9537 | n9539 ;
  assign n9541 = n1974 ^ n927 ^ 1'b0 ;
  assign n9542 = ~n493 & n859 ;
  assign n9543 = n2806 | n9542 ;
  assign n9544 = ~n877 & n1736 ;
  assign n9545 = n848 & n9544 ;
  assign n9546 = n9545 ^ n394 ^ 1'b0 ;
  assign n9547 = n9543 & ~n9546 ;
  assign n9548 = n1818 & n7712 ;
  assign n9549 = ~n307 & n4867 ;
  assign n9550 = ~n927 & n9549 ;
  assign n9551 = n9550 ^ n7571 ^ 1'b0 ;
  assign n9552 = n9548 & n9551 ;
  assign n9553 = ~n5454 & n9552 ;
  assign n9554 = ~n703 & n2868 ;
  assign n9555 = ~n448 & n7960 ;
  assign n9556 = ~n1397 & n7451 ;
  assign n9557 = n3123 ^ n1663 ^ 1'b0 ;
  assign n9558 = n3115 | n9557 ;
  assign n9559 = n9558 ^ n7457 ^ 1'b0 ;
  assign n9560 = ~n3181 & n6167 ;
  assign n9561 = ~n740 & n2590 ;
  assign n9562 = n9561 ^ n3552 ^ 1'b0 ;
  assign n9563 = n623 | n2343 ;
  assign n9564 = ~n9562 & n9563 ;
  assign n9565 = n1255 & n4047 ;
  assign n9566 = n4175 ^ n944 ^ 1'b0 ;
  assign n9567 = n3839 | n9566 ;
  assign n9568 = n9567 ^ n5242 ^ 1'b0 ;
  assign n9569 = ( ~x14 & x206 ) | ( ~x14 & n897 ) | ( x206 & n897 ) ;
  assign n9570 = n1252 & ~n9569 ;
  assign n9571 = ~n2351 & n9570 ;
  assign n9572 = n1945 & n9053 ;
  assign n9573 = ~n3670 & n9572 ;
  assign n9574 = n9269 & ~n9573 ;
  assign n9575 = ~x249 & n9574 ;
  assign n9576 = n955 | n9575 ;
  assign n9577 = n7518 ^ n7508 ^ 1'b0 ;
  assign n9578 = n4596 & ~n9577 ;
  assign n9579 = n4741 ^ n1591 ^ 1'b0 ;
  assign n9580 = n6967 & n9579 ;
  assign n9584 = ~x245 & n2106 ;
  assign n9581 = n6964 & n7535 ;
  assign n9582 = n6972 & n9581 ;
  assign n9583 = ~n9234 & n9582 ;
  assign n9585 = n9584 ^ n9583 ^ 1'b0 ;
  assign n9586 = n7220 ^ x83 ^ 1'b0 ;
  assign n9587 = n9493 & n9586 ;
  assign n9588 = ( n401 & ~n5826 ) | ( n401 & n8099 ) | ( ~n5826 & n8099 ) ;
  assign n9590 = n482 ^ n277 ^ 1'b0 ;
  assign n9591 = n1264 & ~n9590 ;
  assign n9592 = n9591 ^ n5703 ^ 1'b0 ;
  assign n9589 = n8908 ^ n1846 ^ 1'b0 ;
  assign n9593 = n9592 ^ n9589 ^ 1'b0 ;
  assign n9594 = n4273 ^ n985 ^ 1'b0 ;
  assign n9595 = n9594 ^ n3756 ^ 1'b0 ;
  assign n9596 = x113 & n9595 ;
  assign n9597 = n3637 & ~n9596 ;
  assign n9598 = n1777 | n3239 ;
  assign n9599 = n5346 & n6999 ;
  assign n9600 = n6702 & n9599 ;
  assign n9601 = ~n1907 & n3277 ;
  assign n9602 = n9601 ^ n1968 ^ 1'b0 ;
  assign n9603 = x39 & n9602 ;
  assign n9604 = n9603 ^ n6414 ^ 1'b0 ;
  assign n9605 = n9604 ^ n3743 ^ 1'b0 ;
  assign n9606 = n2356 & n9605 ;
  assign n9607 = n8931 ^ n1720 ^ 1'b0 ;
  assign n9608 = ~n9394 & n9607 ;
  assign n9609 = n5188 & ~n7303 ;
  assign n9610 = n6856 ^ n1863 ^ 1'b0 ;
  assign n9611 = ~n2426 & n9610 ;
  assign n9612 = n5382 | n9611 ;
  assign n9613 = ~n9609 & n9612 ;
  assign n9614 = n1805 & n4195 ;
  assign n9615 = n9614 ^ n6874 ^ 1'b0 ;
  assign n9616 = ~n9613 & n9615 ;
  assign n9617 = x144 & n3683 ;
  assign n9621 = n1840 | n8644 ;
  assign n9618 = x54 & ~n1760 ;
  assign n9619 = n9618 ^ n9256 ^ 1'b0 ;
  assign n9620 = ~n1926 & n9619 ;
  assign n9622 = n9621 ^ n9620 ^ 1'b0 ;
  assign n9623 = ~x84 & n3558 ;
  assign n9624 = ~n7910 & n9623 ;
  assign n9625 = n4321 & ~n9624 ;
  assign n9626 = n7411 & n9625 ;
  assign n9627 = n3071 & n5000 ;
  assign n9630 = n2437 ^ n968 ^ 1'b0 ;
  assign n9628 = n2362 | n5121 ;
  assign n9629 = x114 | n9628 ;
  assign n9631 = n9630 ^ n9629 ^ 1'b0 ;
  assign n9632 = ~n4520 & n9631 ;
  assign n9633 = n2507 & ~n4366 ;
  assign n9634 = n9633 ^ n1899 ^ 1'b0 ;
  assign n9635 = n9634 ^ n5310 ^ 1'b0 ;
  assign n9636 = ~n1928 & n9635 ;
  assign n9642 = n1522 ^ n903 ^ 1'b0 ;
  assign n9643 = ~n832 & n9642 ;
  assign n9644 = n4791 & n9643 ;
  assign n9645 = ~n9643 & n9644 ;
  assign n9641 = ~n5370 & n6866 ;
  assign n9646 = n9645 ^ n9641 ^ 1'b0 ;
  assign n9647 = n7730 ^ n2105 ^ 1'b0 ;
  assign n9648 = n9646 & n9647 ;
  assign n9637 = x98 & x239 ;
  assign n9638 = n9637 ^ n1291 ^ 1'b0 ;
  assign n9639 = ~n4849 & n9638 ;
  assign n9640 = ~n2006 & n9639 ;
  assign n9649 = n9648 ^ n9640 ^ 1'b0 ;
  assign n9650 = n472 | n3284 ;
  assign n9651 = n683 & ~n9650 ;
  assign n9652 = ( n1608 & n3323 ) | ( n1608 & n9651 ) | ( n3323 & n9651 ) ;
  assign n9653 = n9652 ^ n2510 ^ 1'b0 ;
  assign n9654 = ( ~n1286 & n6033 ) | ( ~n1286 & n9653 ) | ( n6033 & n9653 ) ;
  assign n9655 = n9654 ^ n3413 ^ 1'b0 ;
  assign n9660 = x248 & n3152 ;
  assign n9656 = ~n3430 & n5296 ;
  assign n9657 = n9656 ^ n3444 ^ 1'b0 ;
  assign n9658 = n1360 & ~n9657 ;
  assign n9659 = n9658 ^ n7423 ^ 1'b0 ;
  assign n9661 = n9660 ^ n9659 ^ 1'b0 ;
  assign n9662 = n9055 ^ n8108 ^ 1'b0 ;
  assign n9663 = n3880 | n9662 ;
  assign n9664 = n492 & n4793 ;
  assign n9665 = ~n2597 & n9664 ;
  assign n9666 = n1441 | n7089 ;
  assign n9667 = n1441 & ~n9666 ;
  assign n9671 = x145 & x220 ;
  assign n9672 = ~x145 & n9671 ;
  assign n9668 = ~n3324 & n4385 ;
  assign n9669 = n3324 & n9668 ;
  assign n9670 = n546 & ~n9669 ;
  assign n9673 = n9672 ^ n9670 ^ 1'b0 ;
  assign n9674 = n5417 & n9673 ;
  assign n9675 = n9667 & n9674 ;
  assign n9676 = x0 & ~n9675 ;
  assign n9677 = ~x0 & n9676 ;
  assign n9678 = n2357 ^ n1596 ^ 1'b0 ;
  assign n9679 = ~n3679 & n9678 ;
  assign n9680 = n3655 & ~n6851 ;
  assign n9681 = n9680 ^ n3186 ^ 1'b0 ;
  assign n9682 = n1223 & ~n9681 ;
  assign n9683 = n9682 ^ n9000 ^ 1'b0 ;
  assign n9684 = n9679 & n9683 ;
  assign n9685 = n4251 ^ n3531 ^ x235 ;
  assign n9686 = n1361 & ~n1782 ;
  assign n9687 = n2841 & n9686 ;
  assign n9688 = n2951 ^ n1693 ^ 1'b0 ;
  assign n9689 = n4719 & ~n8933 ;
  assign n9690 = ~n9688 & n9689 ;
  assign n9691 = n361 & n4826 ;
  assign n9692 = n9691 ^ n3269 ^ 1'b0 ;
  assign n9693 = n2083 & ~n4520 ;
  assign n9694 = n6262 ^ n3016 ^ 1'b0 ;
  assign n9695 = n9693 | n9694 ;
  assign n9696 = ( n4143 & ~n9692 ) | ( n4143 & n9695 ) | ( ~n9692 & n9695 ) ;
  assign n9697 = n4727 ^ n4615 ^ 1'b0 ;
  assign n9698 = n681 & n3366 ;
  assign n9699 = n9697 & ~n9698 ;
  assign n9700 = n9699 ^ n608 ^ 1'b0 ;
  assign n9701 = x14 & ~n628 ;
  assign n9702 = n9701 ^ n1685 ^ 1'b0 ;
  assign n9703 = n4860 & n9702 ;
  assign n9707 = n3576 & n4481 ;
  assign n9704 = n500 & ~n514 ;
  assign n9705 = n9704 ^ n4190 ^ 1'b0 ;
  assign n9706 = n9705 ^ n1593 ^ 1'b0 ;
  assign n9708 = n9707 ^ n9706 ^ 1'b0 ;
  assign n9709 = n337 & ~n5199 ;
  assign n9710 = n9709 ^ n3053 ^ 1'b0 ;
  assign n9711 = n8371 ^ n7560 ^ 1'b0 ;
  assign n9712 = ~n985 & n5346 ;
  assign n9713 = ~n9711 & n9712 ;
  assign n9714 = n9713 ^ n1427 ^ 1'b0 ;
  assign n9715 = n707 & ~n708 ;
  assign n9716 = n9715 ^ x82 ^ 1'b0 ;
  assign n9717 = n4067 | n9716 ;
  assign n9718 = n1413 & n6111 ;
  assign n9719 = n9718 ^ n760 ^ 1'b0 ;
  assign n9720 = n8456 & ~n9719 ;
  assign n9721 = n3381 ^ n840 ^ 1'b0 ;
  assign n9722 = ~n4054 & n9721 ;
  assign n9723 = n9722 ^ n4613 ^ 1'b0 ;
  assign n9724 = n9723 ^ n4731 ^ 1'b0 ;
  assign n9725 = n6566 | n9724 ;
  assign n9726 = n9725 ^ n2737 ^ 1'b0 ;
  assign n9727 = n7961 ^ n4009 ^ 1'b0 ;
  assign n9728 = n6111 & ~n9727 ;
  assign n9729 = n1638 | n2208 ;
  assign n9730 = n9728 | n9729 ;
  assign n9731 = n9133 ^ n7239 ^ 1'b0 ;
  assign n9732 = n3379 | n3865 ;
  assign n9733 = x3 & ~n4766 ;
  assign n9734 = n9733 ^ n2861 ^ 1'b0 ;
  assign n9735 = ~n1071 & n9734 ;
  assign n9736 = n9735 ^ n8691 ^ 1'b0 ;
  assign n9737 = n485 & ~n2735 ;
  assign n9738 = n9737 ^ n566 ^ 1'b0 ;
  assign n9739 = n9736 | n9738 ;
  assign n9740 = ~n8842 & n9022 ;
  assign n9741 = n9740 ^ n8324 ^ 1'b0 ;
  assign n9744 = n5823 ^ n2768 ^ 1'b0 ;
  assign n9743 = n3614 | n4505 ;
  assign n9745 = n9744 ^ n9743 ^ 1'b0 ;
  assign n9746 = ~n1893 & n9745 ;
  assign n9747 = ~n786 & n9746 ;
  assign n9748 = n3989 ^ n887 ^ 1'b0 ;
  assign n9749 = n9747 | n9748 ;
  assign n9750 = n7339 | n9749 ;
  assign n9751 = n9750 ^ n6493 ^ 1'b0 ;
  assign n9742 = ~n858 & n8094 ;
  assign n9752 = n9751 ^ n9742 ^ 1'b0 ;
  assign n9753 = ~n3043 & n7077 ;
  assign n9754 = ~x117 & n9753 ;
  assign n9755 = n9333 | n9754 ;
  assign n9759 = n3082 | n6421 ;
  assign n9756 = n1044 & ~n1280 ;
  assign n9757 = n9756 ^ n5791 ^ 1'b0 ;
  assign n9758 = ~n4874 & n9757 ;
  assign n9760 = n9759 ^ n9758 ^ 1'b0 ;
  assign n9761 = n3499 & ~n3632 ;
  assign n9762 = n2310 | n5151 ;
  assign n9763 = n9762 ^ n4540 ^ 1'b0 ;
  assign n9764 = n9761 & ~n9763 ;
  assign n9765 = n8065 ^ n3813 ^ 1'b0 ;
  assign n9766 = n9765 ^ n8377 ^ 1'b0 ;
  assign n9767 = n8813 ^ n2962 ^ 1'b0 ;
  assign n9768 = ~n6333 & n9767 ;
  assign n9769 = ~x197 & n9768 ;
  assign n9770 = n9769 ^ n1361 ^ 1'b0 ;
  assign n9771 = n7353 & n9770 ;
  assign n9772 = n4630 ^ x172 ^ 1'b0 ;
  assign n9773 = n1894 & n9772 ;
  assign n9774 = n9773 ^ n3408 ^ 1'b0 ;
  assign n9775 = n3669 & n9774 ;
  assign n9776 = n440 ^ n339 ^ 1'b0 ;
  assign n9777 = n9776 ^ x123 ^ 1'b0 ;
  assign n9778 = n4553 & ~n9777 ;
  assign n9779 = n8122 ^ n4120 ^ 1'b0 ;
  assign n9780 = n9778 & ~n9779 ;
  assign n9781 = ~n9775 & n9780 ;
  assign n9782 = n5932 ^ n5424 ^ 1'b0 ;
  assign n9783 = ~n3091 & n9782 ;
  assign n9784 = n1383 & ~n3561 ;
  assign n9785 = ~n4236 & n9784 ;
  assign n9786 = n9783 & ~n9785 ;
  assign n9787 = n434 & n5356 ;
  assign n9788 = n1588 | n9787 ;
  assign n9789 = n833 | n1427 ;
  assign n9790 = ~n3078 & n3842 ;
  assign n9791 = ~n6902 & n9790 ;
  assign n9792 = n461 ^ n366 ^ 1'b0 ;
  assign n9793 = n1255 | n9792 ;
  assign n9794 = n1568 | n2589 ;
  assign n9795 = n2011 & n6516 ;
  assign n9796 = n5004 ^ n2962 ^ 1'b0 ;
  assign n9797 = n6586 ^ n4623 ^ 1'b0 ;
  assign n9798 = n6703 ^ n6647 ^ 1'b0 ;
  assign n9799 = n7248 & ~n9798 ;
  assign n9800 = n9799 ^ n1424 ^ 1'b0 ;
  assign n9801 = ~n9797 & n9800 ;
  assign n9802 = n9801 ^ n3882 ^ 1'b0 ;
  assign n9803 = n2129 & ~n2215 ;
  assign n9804 = x20 & ~n3651 ;
  assign n9805 = ~n2076 & n7725 ;
  assign n9806 = n9804 & n9805 ;
  assign n9810 = n6192 ^ n4233 ^ 1'b0 ;
  assign n9808 = ( ~x151 & n715 ) | ( ~x151 & n923 ) | ( n715 & n923 ) ;
  assign n9807 = n2590 | n6573 ;
  assign n9809 = n9808 ^ n9807 ^ 1'b0 ;
  assign n9811 = n9810 ^ n9809 ^ 1'b0 ;
  assign n9814 = ~n1510 & n3189 ;
  assign n9815 = n9814 ^ n2066 ^ 1'b0 ;
  assign n9813 = ~n2855 & n5714 ;
  assign n9816 = n9815 ^ n9813 ^ 1'b0 ;
  assign n9812 = ~n3331 & n7778 ;
  assign n9817 = n9816 ^ n9812 ^ 1'b0 ;
  assign n9818 = ~n3187 & n6612 ;
  assign n9819 = n1356 & n9818 ;
  assign n9820 = ~n1318 & n5207 ;
  assign n9821 = n2129 | n2581 ;
  assign n9822 = n265 & ~n283 ;
  assign n9823 = n1480 & n9822 ;
  assign n9824 = n2279 & n9823 ;
  assign n9825 = n9824 ^ n4822 ^ 1'b0 ;
  assign n9826 = n3939 | n9825 ;
  assign n9827 = n3459 | n9826 ;
  assign n9829 = ~n1361 & n3210 ;
  assign n9830 = n2853 & n9829 ;
  assign n9828 = n1696 & ~n8241 ;
  assign n9831 = n9830 ^ n9828 ^ 1'b0 ;
  assign n9832 = n1052 & ~n4158 ;
  assign n9833 = n9832 ^ n5853 ^ 1'b0 ;
  assign n9834 = ~n2135 & n9833 ;
  assign n9835 = n4106 | n9690 ;
  assign n9836 = n8731 ^ n6290 ^ 1'b0 ;
  assign n9837 = ~n4130 & n5199 ;
  assign n9838 = x254 & n1426 ;
  assign n9839 = ~n1426 & n9838 ;
  assign n9840 = n2185 & n9839 ;
  assign n9841 = x85 & ~n848 ;
  assign n9842 = n848 & n9841 ;
  assign n9843 = x241 & ~n2467 ;
  assign n9844 = n2467 & n9843 ;
  assign n9845 = n1521 & ~n9844 ;
  assign n9846 = n9844 & n9845 ;
  assign n9847 = n9842 | n9846 ;
  assign n9848 = n9842 & ~n9847 ;
  assign n9849 = n566 & n1249 ;
  assign n9850 = n9848 & n9849 ;
  assign n9851 = n9840 | n9850 ;
  assign n9852 = n1644 & ~n9851 ;
  assign n9853 = n1635 & ~n7045 ;
  assign n9854 = n9853 ^ n5846 ^ 1'b0 ;
  assign n9855 = ~n1866 & n2865 ;
  assign n9856 = n5137 & n9855 ;
  assign n9857 = ~n7531 & n9856 ;
  assign n9859 = n6570 ^ n2136 ^ 1'b0 ;
  assign n9860 = n3884 | n9859 ;
  assign n9858 = n1351 & ~n4661 ;
  assign n9861 = n9860 ^ n9858 ^ 1'b0 ;
  assign n9862 = n9861 ^ n4899 ^ 1'b0 ;
  assign n9863 = n6891 ^ n2491 ^ 1'b0 ;
  assign n9864 = n886 & ~n7130 ;
  assign n9865 = n3976 & n9864 ;
  assign n9866 = n2589 ^ n1345 ^ 1'b0 ;
  assign n9867 = n673 | n6551 ;
  assign n9868 = n9867 ^ n2190 ^ 1'b0 ;
  assign n9869 = n5796 & n9868 ;
  assign n9870 = n5042 ^ n2909 ^ x98 ;
  assign n9871 = n2274 & ~n6174 ;
  assign n9872 = n9870 & n9871 ;
  assign n9873 = ( ~n444 & n2358 ) | ( ~n444 & n9872 ) | ( n2358 & n9872 ) ;
  assign n9874 = ~n2247 & n2451 ;
  assign n9875 = x117 & n2935 ;
  assign n9876 = n9875 ^ n8556 ^ 1'b0 ;
  assign n9877 = n2318 & ~n8462 ;
  assign n9878 = n4791 & ~n5891 ;
  assign n9879 = n9878 ^ n5125 ^ 1'b0 ;
  assign n9880 = n2080 & n4997 ;
  assign n9881 = ~n1893 & n9880 ;
  assign n9886 = n4157 ^ n363 ^ 1'b0 ;
  assign n9882 = n5587 | n7050 ;
  assign n9883 = n5730 | n9882 ;
  assign n9884 = n8922 ^ n5824 ^ 1'b0 ;
  assign n9885 = n9883 & n9884 ;
  assign n9887 = n9886 ^ n9885 ^ 1'b0 ;
  assign n9888 = n7305 | n9887 ;
  assign n9889 = ~x71 & n1850 ;
  assign n9890 = ~n5535 & n9889 ;
  assign n9891 = n756 ^ n486 ^ 1'b0 ;
  assign n9895 = n4840 ^ x156 ^ 1'b0 ;
  assign n9892 = n3637 & ~n6032 ;
  assign n9893 = n9892 ^ n884 ^ 1'b0 ;
  assign n9894 = n9893 ^ n8963 ^ 1'b0 ;
  assign n9896 = n9895 ^ n9894 ^ n8633 ;
  assign n9897 = n9525 ^ n1117 ^ 1'b0 ;
  assign n9898 = n1548 ^ n504 ^ 1'b0 ;
  assign n9899 = n9898 ^ n6774 ^ 1'b0 ;
  assign n9900 = n2361 & ~n9899 ;
  assign n9901 = n8312 ^ n6463 ^ 1'b0 ;
  assign n9902 = n880 & n9901 ;
  assign n9903 = n8836 ^ n2920 ^ 1'b0 ;
  assign n9904 = n9902 & ~n9903 ;
  assign n9905 = ~n9900 & n9904 ;
  assign n9906 = n1642 ^ x241 ^ 1'b0 ;
  assign n9907 = n397 & ~n9906 ;
  assign n9908 = n2768 & n8718 ;
  assign n9909 = n9908 ^ n7821 ^ 1'b0 ;
  assign n9910 = ~n1814 & n3197 ;
  assign n9911 = n9910 ^ n2787 ^ x34 ;
  assign n9912 = n9911 ^ n3546 ^ 1'b0 ;
  assign n9913 = n1780 & ~n2263 ;
  assign n9914 = ~n6749 & n9913 ;
  assign n9915 = n9914 ^ n2004 ^ 1'b0 ;
  assign n9916 = n9915 ^ n3432 ^ 1'b0 ;
  assign n9917 = n9205 ^ n1488 ^ 1'b0 ;
  assign n9918 = n3441 | n9917 ;
  assign n9919 = n9916 & ~n9918 ;
  assign n9920 = n9912 & ~n9919 ;
  assign n9921 = ~n3678 & n9920 ;
  assign n9922 = n6989 ^ n6225 ^ n5846 ;
  assign n9923 = n887 & n1641 ;
  assign n9924 = n2629 ^ n1156 ^ 1'b0 ;
  assign n9925 = n1376 & n9924 ;
  assign n9926 = n9925 ^ n8582 ^ 1'b0 ;
  assign n9927 = n4939 & ~n7117 ;
  assign n9928 = n3235 & n9927 ;
  assign n9929 = n685 | n4787 ;
  assign n9930 = n3575 | n6729 ;
  assign n9931 = n3911 & n9930 ;
  assign n9932 = n9929 & n9931 ;
  assign n9933 = n9932 ^ n941 ^ 1'b0 ;
  assign n9934 = n3906 ^ n1117 ^ 1'b0 ;
  assign n9935 = n9122 ^ n903 ^ 1'b0 ;
  assign n9936 = n2269 & n9935 ;
  assign n9937 = n9936 ^ n2409 ^ 1'b0 ;
  assign n9938 = n9530 ^ n972 ^ 1'b0 ;
  assign n9939 = ~n1383 & n9938 ;
  assign n9940 = n9939 ^ n399 ^ 1'b0 ;
  assign n9941 = ~x9 & n2786 ;
  assign n9942 = n9941 ^ n2318 ^ 1'b0 ;
  assign n9943 = n2881 & ~n4707 ;
  assign n9944 = n9943 ^ n2190 ^ 1'b0 ;
  assign n9945 = n9944 ^ n1810 ^ 1'b0 ;
  assign n9946 = n9942 & ~n9945 ;
  assign n9947 = ~n9940 & n9946 ;
  assign n9948 = n4310 ^ n589 ^ 1'b0 ;
  assign n9949 = n9905 & n9948 ;
  assign n9950 = ~n9947 & n9949 ;
  assign n9951 = n9069 ^ n5137 ^ 1'b0 ;
  assign n9952 = n2837 ^ n892 ^ 1'b0 ;
  assign n9953 = n6437 | n9952 ;
  assign n9954 = n9951 & ~n9953 ;
  assign n9955 = n9954 ^ n2247 ^ 1'b0 ;
  assign n9956 = n2026 & ~n2315 ;
  assign n9957 = n6169 ^ n4198 ^ 1'b0 ;
  assign n9958 = ~n3511 & n8211 ;
  assign n9959 = n2761 & n9958 ;
  assign n9960 = n2073 ^ n1064 ^ 1'b0 ;
  assign n9961 = n9959 | n9960 ;
  assign n9962 = n9961 ^ n932 ^ 1'b0 ;
  assign n9963 = n9957 | n9962 ;
  assign n9964 = n8728 ^ n2426 ^ 1'b0 ;
  assign n9965 = n2087 & ~n8139 ;
  assign n9966 = ~n647 & n1262 ;
  assign n9967 = n9966 ^ n1501 ^ 1'b0 ;
  assign n9968 = n5196 ^ n1740 ^ 1'b0 ;
  assign n9969 = n9967 & n9968 ;
  assign n9970 = ~n2235 & n4328 ;
  assign n9971 = ~n1736 & n9970 ;
  assign n9972 = n9971 ^ n8765 ^ 1'b0 ;
  assign n9973 = n2098 ^ n1678 ^ 1'b0 ;
  assign n9974 = n9307 & ~n9973 ;
  assign n9975 = n9974 ^ n1991 ^ 1'b0 ;
  assign n9976 = n9972 & ~n9975 ;
  assign n9977 = n1736 & n3071 ;
  assign n9978 = ~n8646 & n9977 ;
  assign n9979 = n1239 ^ n1031 ^ 1'b0 ;
  assign n9980 = n5989 & n9979 ;
  assign n9983 = n4888 ^ n354 ^ 1'b0 ;
  assign n9984 = ~n1435 & n9983 ;
  assign n9985 = n9984 ^ n3030 ^ 1'b0 ;
  assign n9986 = n9985 ^ n4106 ^ 1'b0 ;
  assign n9981 = n6889 ^ n6464 ^ n4417 ;
  assign n9982 = ~n7671 & n9981 ;
  assign n9987 = n9986 ^ n9982 ^ 1'b0 ;
  assign n9988 = n9980 & n9987 ;
  assign n9989 = n1898 & ~n3045 ;
  assign n9990 = ( n4304 & n5767 ) | ( n4304 & n8244 ) | ( n5767 & n8244 ) ;
  assign n9991 = n9990 ^ n7552 ^ 1'b0 ;
  assign n9992 = n749 | n6179 ;
  assign n9993 = n2886 | n3926 ;
  assign n9994 = n6394 ^ n2554 ^ 1'b0 ;
  assign n9995 = n9824 | n9994 ;
  assign n9996 = n1429 & n9995 ;
  assign n9997 = n6325 ^ n977 ^ 1'b0 ;
  assign n9998 = x28 & ~n9997 ;
  assign n9999 = n9998 ^ n4395 ^ 1'b0 ;
  assign n10000 = ~n5194 & n9999 ;
  assign n10001 = n6649 & n10000 ;
  assign n10002 = n10001 ^ n9402 ^ 1'b0 ;
  assign n10003 = n1062 & ~n3950 ;
  assign n10004 = n5814 & n10003 ;
  assign n10005 = n3511 | n10004 ;
  assign n10006 = n3336 | n7133 ;
  assign n10007 = n5723 & n9415 ;
  assign n10008 = n10007 ^ x253 ^ 1'b0 ;
  assign n10009 = n3221 ^ n1657 ^ 1'b0 ;
  assign n10010 = ~n3549 & n10009 ;
  assign n10011 = n4205 | n7244 ;
  assign n10012 = n7524 | n10011 ;
  assign n10013 = ~x154 & n3288 ;
  assign n10014 = ~n10012 & n10013 ;
  assign n10015 = n10014 ^ n8257 ^ 1'b0 ;
  assign n10016 = n10010 & n10015 ;
  assign n10017 = n5440 ^ x59 ^ 1'b0 ;
  assign n10018 = n5354 ^ n4227 ^ 1'b0 ;
  assign n10019 = ~n3035 & n10018 ;
  assign n10020 = ~n5867 & n7621 ;
  assign n10021 = n1499 & n10020 ;
  assign n10022 = n2150 & ~n10021 ;
  assign n10023 = n1004 & ~n10022 ;
  assign n10024 = n4677 | n5389 ;
  assign n10025 = n3483 & n10024 ;
  assign n10026 = n1334 | n3112 ;
  assign n10027 = n6885 & n9463 ;
  assign n10028 = n2575 & ~n3545 ;
  assign n10029 = n3239 & n9947 ;
  assign n10030 = ~n10028 & n10029 ;
  assign n10031 = n4945 ^ n4208 ^ n1849 ;
  assign n10032 = n5446 & ~n10031 ;
  assign n10033 = n1980 & n10032 ;
  assign n10034 = n4813 ^ n2500 ^ 1'b0 ;
  assign n10035 = n2825 & n10034 ;
  assign n10036 = ~n5152 & n10035 ;
  assign n10037 = n9737 & n10036 ;
  assign n10038 = n2658 | n3389 ;
  assign n10039 = x158 | n414 ;
  assign n10040 = n10039 ^ n2287 ^ 1'b0 ;
  assign n10041 = ~n4075 & n10040 ;
  assign n10042 = ~n10038 & n10041 ;
  assign n10043 = n6546 & ~n10042 ;
  assign n10044 = n10043 ^ n7642 ^ 1'b0 ;
  assign n10045 = n800 & ~n4063 ;
  assign n10046 = n6858 & n10045 ;
  assign n10047 = n3152 ^ n2925 ^ 1'b0 ;
  assign n10048 = n6990 & ~n10047 ;
  assign n10049 = n6900 ^ n2345 ^ 1'b0 ;
  assign n10050 = n10049 ^ n3414 ^ 1'b0 ;
  assign n10051 = n366 & n10050 ;
  assign n10052 = x81 & ~n9074 ;
  assign n10053 = n6413 ^ n533 ^ 1'b0 ;
  assign n10054 = ~n1411 & n10053 ;
  assign n10055 = ~n6813 & n10054 ;
  assign n10056 = n10055 ^ n4154 ^ 1'b0 ;
  assign n10057 = n5788 ^ n1996 ^ 1'b0 ;
  assign n10058 = n2129 & ~n10057 ;
  assign n10059 = n5154 & ~n10058 ;
  assign n10060 = n6966 ^ n1271 ^ 1'b0 ;
  assign n10061 = n10059 | n10060 ;
  assign n10062 = n8442 ^ n1075 ^ 1'b0 ;
  assign n10063 = n4140 & n10062 ;
  assign n10064 = n2704 ^ n762 ^ 1'b0 ;
  assign n10065 = n10064 ^ n1945 ^ 1'b0 ;
  assign n10066 = n7395 & ~n10065 ;
  assign n10067 = n10066 ^ n2423 ^ 1'b0 ;
  assign n10068 = ~n9219 & n10067 ;
  assign n10069 = n522 & n3803 ;
  assign n10070 = n10069 ^ x191 ^ 1'b0 ;
  assign n10071 = n1814 & ~n10070 ;
  assign n10072 = n10071 ^ n2402 ^ 1'b0 ;
  assign n10074 = n2725 & ~n4961 ;
  assign n10075 = n10074 ^ n2457 ^ 1'b0 ;
  assign n10073 = n4433 & ~n8212 ;
  assign n10076 = n10075 ^ n10073 ^ 1'b0 ;
  assign n10077 = n966 & n1801 ;
  assign n10078 = ~n10076 & n10077 ;
  assign n10080 = n4658 ^ n3275 ^ 1'b0 ;
  assign n10079 = n2320 & n2752 ;
  assign n10081 = n10080 ^ n10079 ^ 1'b0 ;
  assign n10082 = n7047 ^ n4116 ^ 1'b0 ;
  assign n10083 = n1646 & n6817 ;
  assign n10084 = n10083 ^ n10027 ^ 1'b0 ;
  assign n10085 = n8872 ^ n5045 ^ 1'b0 ;
  assign n10086 = n4047 & ~n10085 ;
  assign n10087 = n3690 & ~n7630 ;
  assign n10088 = n1100 ^ n965 ^ 1'b0 ;
  assign n10089 = n1499 | n10088 ;
  assign n10090 = n3879 & n5929 ;
  assign n10091 = ~n895 & n2989 ;
  assign n10092 = n10091 ^ n1643 ^ 1'b0 ;
  assign n10093 = n7563 | n10092 ;
  assign n10094 = n10090 & ~n10093 ;
  assign n10095 = n10089 | n10094 ;
  assign n10097 = n358 | n3059 ;
  assign n10096 = n3258 & n4395 ;
  assign n10098 = n10097 ^ n10096 ^ 1'b0 ;
  assign n10099 = n747 & ~n6233 ;
  assign n10100 = n10099 ^ n4615 ^ 1'b0 ;
  assign n10101 = n4053 & ~n10100 ;
  assign n10102 = n942 & n8480 ;
  assign n10105 = n1643 & ~n3882 ;
  assign n10103 = n4341 | n5890 ;
  assign n10104 = n2042 & ~n10103 ;
  assign n10106 = n10105 ^ n10104 ^ 1'b0 ;
  assign n10107 = n2248 & n2587 ;
  assign n10108 = n1883 & n10107 ;
  assign n10111 = n959 | n3328 ;
  assign n10112 = ~n869 & n10111 ;
  assign n10109 = ~n2936 & n3428 ;
  assign n10110 = n1527 & n10109 ;
  assign n10113 = n10112 ^ n10110 ^ 1'b0 ;
  assign n10114 = n3128 & n10113 ;
  assign n10115 = n3516 | n4896 ;
  assign n10116 = x232 | n10115 ;
  assign n10117 = n10116 ^ n2143 ^ 1'b0 ;
  assign n10118 = n9875 & n10117 ;
  assign n10119 = n6974 ^ n415 ^ 1'b0 ;
  assign n10120 = n10118 & ~n10119 ;
  assign n10121 = n5496 & ~n8324 ;
  assign n10122 = n7630 ^ n2089 ^ 1'b0 ;
  assign n10123 = n1302 & ~n9116 ;
  assign n10124 = n10123 ^ n1321 ^ 1'b0 ;
  assign n10125 = x60 | n4910 ;
  assign n10126 = n10125 ^ n3903 ^ 1'b0 ;
  assign n10127 = x140 & ~n6473 ;
  assign n10128 = n10127 ^ x200 ^ 1'b0 ;
  assign n10129 = n5619 ^ n2246 ^ 1'b0 ;
  assign n10130 = n2463 & ~n10129 ;
  assign n10131 = ~n10128 & n10130 ;
  assign n10132 = n10131 ^ n7855 ^ 1'b0 ;
  assign n10133 = n10126 & ~n10132 ;
  assign n10134 = n2678 & ~n3896 ;
  assign n10135 = n3834 & n10134 ;
  assign n10136 = ~n3477 & n10135 ;
  assign n10137 = n552 | n1059 ;
  assign n10138 = n7109 & ~n10137 ;
  assign n10139 = n3891 | n4189 ;
  assign n10140 = n2979 | n10139 ;
  assign n10141 = ~n3902 & n10140 ;
  assign n10142 = n10138 | n10141 ;
  assign n10143 = n10142 ^ n4026 ^ 1'b0 ;
  assign n10144 = n2150 | n9170 ;
  assign n10145 = n9001 & n10144 ;
  assign n10146 = n4263 ^ n1391 ^ 1'b0 ;
  assign n10147 = n10146 ^ n9068 ^ 1'b0 ;
  assign n10148 = n1743 | n3122 ;
  assign n10149 = n6847 | n10148 ;
  assign n10150 = n1443 | n10149 ;
  assign n10151 = n3128 & n6506 ;
  assign n10153 = n1419 & n9630 ;
  assign n10152 = n5262 ^ n4743 ^ n4328 ;
  assign n10154 = n10153 ^ n10152 ^ n1441 ;
  assign n10155 = n7168 | n10154 ;
  assign n10156 = n10151 | n10155 ;
  assign n10157 = n10089 & ~n10156 ;
  assign n10158 = n6295 | n10157 ;
  assign n10159 = x112 & ~n4314 ;
  assign n10160 = n1820 & n10159 ;
  assign n10161 = n3105 & n7655 ;
  assign n10162 = n5471 & n10161 ;
  assign n10163 = n6213 & ~n10162 ;
  assign n10164 = n1562 | n6667 ;
  assign n10165 = n8956 ^ n3558 ^ 1'b0 ;
  assign n10166 = n1777 | n10165 ;
  assign n10167 = n864 | n6060 ;
  assign n10168 = n2536 & ~n7689 ;
  assign n10169 = n2549 & n8236 ;
  assign n10170 = n5639 & n7661 ;
  assign n10171 = n10170 ^ n6446 ^ 1'b0 ;
  assign n10173 = n3910 ^ n2537 ^ 1'b0 ;
  assign n10174 = n1488 | n10173 ;
  assign n10172 = ~n2949 & n8899 ;
  assign n10175 = n10174 ^ n10172 ^ 1'b0 ;
  assign n10176 = x203 & n10175 ;
  assign n10177 = ~n1646 & n10176 ;
  assign n10178 = n9223 ^ x249 ^ 1'b0 ;
  assign n10179 = ( x89 & ~n4776 ) | ( x89 & n10178 ) | ( ~n4776 & n10178 ) ;
  assign n10180 = n8995 ^ n3336 ^ 1'b0 ;
  assign n10181 = n10179 & ~n10180 ;
  assign n10182 = n1143 ^ x253 ^ 1'b0 ;
  assign n10183 = n2489 | n2870 ;
  assign n10184 = n4625 | n10183 ;
  assign n10185 = n10182 & ~n10184 ;
  assign n10186 = n9651 ^ n2393 ^ 1'b0 ;
  assign n10187 = ~n4370 & n10186 ;
  assign n10188 = n1740 | n10187 ;
  assign n10189 = n1260 & ~n9053 ;
  assign n10191 = n4630 ^ n602 ^ 1'b0 ;
  assign n10192 = ~n3365 & n10191 ;
  assign n10193 = n10192 ^ n7124 ^ 1'b0 ;
  assign n10194 = n7061 & ~n10193 ;
  assign n10190 = ~n1449 & n5207 ;
  assign n10195 = n10194 ^ n10190 ^ 1'b0 ;
  assign n10196 = n736 ^ n337 ^ 1'b0 ;
  assign n10197 = n6879 | n10196 ;
  assign n10198 = x101 | n10197 ;
  assign n10199 = x64 & ~n9939 ;
  assign n10200 = n4473 & ~n10199 ;
  assign n10201 = n2660 & n10200 ;
  assign n10202 = n833 & n9445 ;
  assign n10203 = n10202 ^ n5928 ^ 1'b0 ;
  assign n10204 = ~n351 & n1133 ;
  assign n10205 = n10204 ^ n8604 ^ 1'b0 ;
  assign n10206 = n6325 ^ n6017 ^ n4745 ;
  assign n10207 = n9655 | n10206 ;
  assign n10208 = n10206 & ~n10207 ;
  assign n10209 = n2035 & ~n4256 ;
  assign n10210 = n3673 & n10209 ;
  assign n10211 = n643 | n6123 ;
  assign n10216 = n6757 & n9525 ;
  assign n10217 = n10216 ^ n1790 ^ 1'b0 ;
  assign n10212 = n420 & ~n2385 ;
  assign n10213 = n10212 ^ n1118 ^ 1'b0 ;
  assign n10214 = n10213 ^ n1473 ^ 1'b0 ;
  assign n10215 = n1164 & n10214 ;
  assign n10218 = n10217 ^ n10215 ^ 1'b0 ;
  assign n10219 = n860 & n7290 ;
  assign n10220 = n10219 ^ n9678 ^ 1'b0 ;
  assign n10221 = n2868 ^ n492 ^ 1'b0 ;
  assign n10222 = n10221 ^ n2557 ^ 1'b0 ;
  assign n10223 = n4099 & ~n5232 ;
  assign n10224 = n10223 ^ n2018 ^ 1'b0 ;
  assign n10225 = n1499 | n10224 ;
  assign n10226 = n3274 & n3524 ;
  assign n10231 = ~n2944 & n5177 ;
  assign n10232 = ~x61 & n10231 ;
  assign n10233 = n2936 & ~n10232 ;
  assign n10227 = n456 | n7867 ;
  assign n10228 = n694 & ~n10227 ;
  assign n10229 = n2366 & ~n10228 ;
  assign n10230 = n4193 & ~n10229 ;
  assign n10234 = n10233 ^ n10230 ^ 1'b0 ;
  assign n10235 = n1173 & n2184 ;
  assign n10236 = n10235 ^ n1148 ^ 1'b0 ;
  assign n10237 = n4539 & n10236 ;
  assign n10238 = n6104 ^ n3219 ^ n1672 ;
  assign n10239 = ~n5593 & n10087 ;
  assign n10240 = n7195 ^ n4851 ^ 1'b0 ;
  assign n10241 = n7901 ^ n5495 ^ 1'b0 ;
  assign n10248 = n915 & n941 ;
  assign n10249 = ~n915 & n10248 ;
  assign n10250 = x208 & x252 ;
  assign n10251 = n10249 & n10250 ;
  assign n10252 = x216 & n5060 ;
  assign n10253 = ~x216 & n10252 ;
  assign n10254 = n10253 ^ n3125 ^ 1'b0 ;
  assign n10255 = n10251 & ~n10254 ;
  assign n10256 = n10255 ^ n3855 ^ 1'b0 ;
  assign n10242 = ~n1732 & n1985 ;
  assign n10243 = n1732 & n10242 ;
  assign n10244 = x7 & ~n1729 ;
  assign n10245 = n10243 & n10244 ;
  assign n10246 = ~n4203 & n10245 ;
  assign n10247 = n10222 | n10246 ;
  assign n10257 = n10256 ^ n10247 ^ 1'b0 ;
  assign n10258 = n10257 ^ n436 ^ 1'b0 ;
  assign n10259 = n1630 | n3656 ;
  assign n10260 = n10259 ^ n2392 ^ 1'b0 ;
  assign n10261 = n10126 & n10260 ;
  assign n10262 = n3264 & ~n7148 ;
  assign n10263 = ~n1554 & n3493 ;
  assign n10264 = n5945 & ~n6667 ;
  assign n10265 = n7496 & n10264 ;
  assign n10266 = ~n1922 & n7836 ;
  assign n10267 = n10266 ^ n3836 ^ 1'b0 ;
  assign n10268 = n9356 ^ n2957 ^ 1'b0 ;
  assign n10269 = n3936 & n10268 ;
  assign n10270 = n3387 & n10269 ;
  assign n10271 = n2722 & n4498 ;
  assign n10272 = n7287 ^ n1468 ^ 1'b0 ;
  assign n10273 = n9731 & n10272 ;
  assign n10274 = n856 & n5715 ;
  assign n10275 = n4209 & n10274 ;
  assign n10276 = n10275 ^ n5835 ^ n3026 ;
  assign n10277 = n1049 | n9055 ;
  assign n10278 = n4938 | n10277 ;
  assign n10279 = n8263 & n10278 ;
  assign n10280 = n4560 ^ x85 ^ 1'b0 ;
  assign n10281 = n6012 & n6403 ;
  assign n10282 = ~n651 & n4324 ;
  assign n10283 = n10282 ^ n4796 ^ 1'b0 ;
  assign n10284 = n5000 ^ n3212 ^ 1'b0 ;
  assign n10285 = n10284 ^ n6205 ^ 1'b0 ;
  assign n10286 = n3551 & n10285 ;
  assign n10287 = ( ~n2409 & n4001 ) | ( ~n2409 & n4523 ) | ( n4001 & n4523 ) ;
  assign n10288 = n797 | n1012 ;
  assign n10289 = n7723 ^ n3370 ^ 1'b0 ;
  assign n10290 = n10288 & n10289 ;
  assign n10291 = ~n10287 & n10290 ;
  assign n10292 = ~n3307 & n10291 ;
  assign n10293 = n10292 ^ n4338 ^ 1'b0 ;
  assign n10294 = n10286 & ~n10293 ;
  assign n10295 = n9974 ^ x125 ^ 1'b0 ;
  assign n10296 = n4058 & n10295 ;
  assign n10297 = ~n5312 & n10296 ;
  assign n10298 = x128 & ~n6661 ;
  assign n10300 = ~n2644 & n3524 ;
  assign n10301 = n3933 ^ n1130 ^ 1'b0 ;
  assign n10302 = n10300 & n10301 ;
  assign n10299 = n4154 | n10150 ;
  assign n10303 = n10302 ^ n10299 ^ 1'b0 ;
  assign n10304 = x166 & n6595 ;
  assign n10305 = n6524 | n10304 ;
  assign n10306 = ~n2632 & n3521 ;
  assign n10307 = n10306 ^ n2373 ^ 1'b0 ;
  assign n10308 = ~n8586 & n10307 ;
  assign n10309 = n3493 ^ n2976 ^ 1'b0 ;
  assign n10310 = ~n5307 & n10309 ;
  assign n10311 = n10310 ^ n4166 ^ 1'b0 ;
  assign n10312 = n2472 & ~n3182 ;
  assign n10313 = n10312 ^ n2057 ^ 1'b0 ;
  assign n10314 = n8215 | n10313 ;
  assign n10320 = n2892 | n6231 ;
  assign n10321 = n4669 & ~n10320 ;
  assign n10316 = ~x24 & n1831 ;
  assign n10317 = n10316 ^ n5704 ^ 1'b0 ;
  assign n10318 = n10317 ^ n4467 ^ 1'b0 ;
  assign n10319 = n1639 & n10318 ;
  assign n10322 = n10321 ^ n10319 ^ 1'b0 ;
  assign n10315 = ~n4063 & n6371 ;
  assign n10323 = n10322 ^ n10315 ^ 1'b0 ;
  assign n10324 = n2536 | n5170 ;
  assign n10325 = n2569 | n10324 ;
  assign n10331 = n4992 ^ n1018 ^ 1'b0 ;
  assign n10326 = n3300 & n7733 ;
  assign n10327 = n384 & n10326 ;
  assign n10328 = ~n3360 & n7217 ;
  assign n10329 = n10327 & n10328 ;
  assign n10330 = n495 | n10329 ;
  assign n10332 = n10331 ^ n10330 ^ 1'b0 ;
  assign n10333 = x123 & n6171 ;
  assign n10334 = n4143 & n10333 ;
  assign n10335 = n1639 & ~n3413 ;
  assign n10336 = n10335 ^ n2293 ^ 1'b0 ;
  assign n10337 = ~n2352 & n10336 ;
  assign n10338 = n3039 & n10337 ;
  assign n10339 = n6583 & ~n7997 ;
  assign n10340 = n10338 & n10339 ;
  assign n10341 = n5530 | n10340 ;
  assign n10342 = n2026 | n10341 ;
  assign n10343 = n5409 | n10342 ;
  assign n10344 = n10334 & ~n10343 ;
  assign n10345 = n9034 ^ n4773 ^ 1'b0 ;
  assign n10346 = n5385 ^ n3480 ^ 1'b0 ;
  assign n10347 = n10346 ^ x222 ^ 1'b0 ;
  assign n10348 = n6214 ^ n637 ^ 1'b0 ;
  assign n10349 = n5709 | n10348 ;
  assign n10350 = n10349 ^ n9451 ^ 1'b0 ;
  assign n10351 = n4431 ^ n1568 ^ 1'b0 ;
  assign n10352 = n9345 | n10351 ;
  assign n10354 = n2723 & n7741 ;
  assign n10353 = x101 & ~n468 ;
  assign n10355 = n10354 ^ n10353 ^ 1'b0 ;
  assign n10356 = ~n10352 & n10355 ;
  assign n10357 = ~n5422 & n6322 ;
  assign n10358 = n10357 ^ n8957 ^ 1'b0 ;
  assign n10359 = x160 | n1124 ;
  assign n10360 = ~n6158 & n8083 ;
  assign n10373 = n3310 ^ n3076 ^ 1'b0 ;
  assign n10369 = n1706 | n3197 ;
  assign n10370 = n7337 & ~n10369 ;
  assign n10366 = n577 & n5168 ;
  assign n10367 = n5918 & ~n10366 ;
  assign n10368 = ~n2219 & n10367 ;
  assign n10371 = n10370 ^ n10368 ^ 1'b0 ;
  assign n10372 = ~n4083 & n10371 ;
  assign n10374 = n10373 ^ n10372 ^ 1'b0 ;
  assign n10361 = n3343 & n7961 ;
  assign n10362 = ~n3423 & n4287 ;
  assign n10363 = n10362 ^ n3639 ^ 1'b0 ;
  assign n10364 = n1605 | n10363 ;
  assign n10365 = n10361 & n10364 ;
  assign n10375 = n10374 ^ n10365 ^ 1'b0 ;
  assign n10376 = x239 & ~n816 ;
  assign n10377 = n3694 ^ n669 ^ 1'b0 ;
  assign n10378 = n4092 & n10377 ;
  assign n10379 = n10378 ^ n1450 ^ 1'b0 ;
  assign n10380 = n6735 | n10379 ;
  assign n10381 = n10380 ^ n3181 ^ 1'b0 ;
  assign n10382 = ~n2047 & n3988 ;
  assign n10383 = n1515 & ~n3745 ;
  assign n10386 = n1083 | n6473 ;
  assign n10387 = n1873 | n10386 ;
  assign n10384 = x8 & ~x131 ;
  assign n10385 = x47 & n10384 ;
  assign n10388 = n10387 ^ n10385 ^ 1'b0 ;
  assign n10389 = ~n4694 & n10388 ;
  assign n10390 = n7971 ^ n5015 ^ 1'b0 ;
  assign n10391 = n5414 & ~n10390 ;
  assign n10392 = n10391 ^ x163 ^ 1'b0 ;
  assign n10394 = n2883 & ~n4538 ;
  assign n10393 = n5237 & n6792 ;
  assign n10395 = n10394 ^ n10393 ^ n2115 ;
  assign n10397 = n1628 & n4190 ;
  assign n10396 = n1223 ^ n616 ^ 1'b0 ;
  assign n10398 = n10397 ^ n10396 ^ n1969 ;
  assign n10399 = n10398 ^ n2569 ^ 1'b0 ;
  assign n10401 = n2436 ^ n1337 ^ 1'b0 ;
  assign n10400 = n2668 | n3694 ;
  assign n10402 = n10401 ^ n10400 ^ 1'b0 ;
  assign n10403 = n1159 | n1784 ;
  assign n10404 = n10403 ^ n5111 ^ 1'b0 ;
  assign n10405 = n5956 ^ n3501 ^ 1'b0 ;
  assign n10406 = n10404 | n10405 ;
  assign n10407 = ~n6813 & n8655 ;
  assign n10408 = n7323 & n10407 ;
  assign n10409 = n5756 ^ n5664 ^ 1'b0 ;
  assign n10410 = ~n1207 & n10409 ;
  assign n10412 = x180 & n7625 ;
  assign n10413 = ~n8485 & n10412 ;
  assign n10411 = x166 & ~n4159 ;
  assign n10414 = n10413 ^ n10411 ^ 1'b0 ;
  assign n10415 = n2728 & ~n9418 ;
  assign n10416 = ~n2134 & n10415 ;
  assign n10417 = n2731 ^ n904 ^ 1'b0 ;
  assign n10418 = ~n9190 & n10417 ;
  assign n10419 = n2143 ^ n452 ^ 1'b0 ;
  assign n10420 = ~n8107 & n10419 ;
  assign n10421 = n4656 ^ n3368 ^ 1'b0 ;
  assign n10422 = n7565 | n10421 ;
  assign n10423 = n10422 ^ n3946 ^ n1654 ;
  assign n10429 = x214 & n4031 ;
  assign n10430 = ~x15 & n10429 ;
  assign n10431 = n10430 ^ n3531 ^ 1'b0 ;
  assign n10432 = n913 | n10431 ;
  assign n10428 = n461 & n3610 ;
  assign n10433 = n10432 ^ n10428 ^ 1'b0 ;
  assign n10424 = n2367 & ~n4720 ;
  assign n10425 = ~x182 & n10424 ;
  assign n10426 = n6774 | n10425 ;
  assign n10427 = n662 & ~n10426 ;
  assign n10434 = n10433 ^ n10427 ^ 1'b0 ;
  assign n10435 = n3529 | n10434 ;
  assign n10436 = n7989 | n10435 ;
  assign n10437 = ( x58 & ~n1096 ) | ( x58 & n3767 ) | ( ~n1096 & n3767 ) ;
  assign n10438 = n2577 & n10437 ;
  assign n10439 = n10111 | n10438 ;
  assign n10440 = n1537 | n10439 ;
  assign n10441 = n10440 ^ n1066 ^ 1'b0 ;
  assign n10442 = n722 & ~n10441 ;
  assign n10443 = n5928 & n10442 ;
  assign n10444 = n5189 ^ x239 ^ 1'b0 ;
  assign n10445 = n9480 & ~n10444 ;
  assign n10447 = n3224 ^ n2241 ^ 1'b0 ;
  assign n10448 = n331 & ~n10447 ;
  assign n10446 = n9254 ^ n5000 ^ 1'b0 ;
  assign n10449 = n10448 ^ n10446 ^ 1'b0 ;
  assign n10450 = n3707 | n10449 ;
  assign n10451 = n10450 ^ n1910 ^ 1'b0 ;
  assign n10452 = ( ~n903 & n3403 ) | ( ~n903 & n10399 ) | ( n3403 & n10399 ) ;
  assign n10453 = ~n2191 & n2467 ;
  assign n10454 = n10453 ^ x213 ^ 1'b0 ;
  assign n10455 = n4936 ^ n304 ^ 1'b0 ;
  assign n10456 = n4286 & ~n10455 ;
  assign n10457 = ( ~n381 & n8058 ) | ( ~n381 & n10456 ) | ( n8058 & n10456 ) ;
  assign n10458 = n703 ^ x3 ^ 1'b0 ;
  assign n10459 = n1010 & n4363 ;
  assign n10460 = n6811 ^ n2482 ^ 1'b0 ;
  assign n10461 = n10460 ^ n672 ^ 1'b0 ;
  assign n10462 = n10459 & ~n10461 ;
  assign n10463 = n7262 & ~n10325 ;
  assign n10464 = n10463 ^ n8504 ^ 1'b0 ;
  assign n10465 = n8572 ^ n4625 ^ 1'b0 ;
  assign n10466 = n4625 ^ x253 ^ 1'b0 ;
  assign n10467 = n6075 | n10466 ;
  assign n10468 = n10467 ^ n1668 ^ n1352 ;
  assign n10469 = ~n6846 & n8716 ;
  assign n10470 = n2844 | n5023 ;
  assign n10471 = n8493 | n10470 ;
  assign n10472 = n4290 ^ n2306 ^ 1'b0 ;
  assign n10473 = n4373 ^ n1016 ^ 1'b0 ;
  assign n10474 = x226 & ~n2168 ;
  assign n10475 = n2168 & n10474 ;
  assign n10476 = n10039 & ~n10475 ;
  assign n10478 = ~n290 & n1653 ;
  assign n10479 = ~n1653 & n10478 ;
  assign n10477 = n1570 & n4432 ;
  assign n10480 = n10479 ^ n10477 ^ 1'b0 ;
  assign n10481 = n7725 & ~n10480 ;
  assign n10482 = ~n10476 & n10481 ;
  assign n10483 = ~n3860 & n5017 ;
  assign n10484 = ~n5026 & n10483 ;
  assign n10485 = n4181 & n10484 ;
  assign n10486 = n552 ^ n493 ^ 1'b0 ;
  assign n10487 = n8765 | n10486 ;
  assign n10488 = n3022 | n4071 ;
  assign n10489 = n10487 | n10488 ;
  assign n10490 = n810 & ~n10489 ;
  assign n10491 = x81 & n5398 ;
  assign n10492 = n3633 & ~n10491 ;
  assign n10494 = ~n4281 & n4729 ;
  assign n10495 = n10494 ^ n5031 ^ 1'b0 ;
  assign n10493 = n5112 & n7914 ;
  assign n10496 = n10495 ^ n10493 ^ 1'b0 ;
  assign n10497 = ~n2849 & n2925 ;
  assign n10498 = n10497 ^ n2997 ^ 1'b0 ;
  assign n10499 = n277 & ~n5124 ;
  assign n10500 = n10499 ^ n3687 ^ 1'b0 ;
  assign n10501 = n4652 | n10500 ;
  assign n10502 = n10501 ^ n1141 ^ 1'b0 ;
  assign n10503 = n10498 & ~n10502 ;
  assign n10504 = n3251 ^ n1361 ^ 1'b0 ;
  assign n10505 = n3331 | n4014 ;
  assign n10506 = ~n821 & n3543 ;
  assign n10507 = ~n2737 & n10506 ;
  assign n10508 = n3325 | n4149 ;
  assign n10509 = n7628 & ~n10508 ;
  assign n10510 = n10509 ^ n825 ^ 1'b0 ;
  assign n10511 = n8347 | n10510 ;
  assign n10512 = ~n3187 & n3985 ;
  assign n10513 = n10512 ^ n1385 ^ 1'b0 ;
  assign n10514 = n1701 | n10513 ;
  assign n10515 = ~n1021 & n1120 ;
  assign n10516 = n2841 & n10515 ;
  assign n10517 = n3371 | n5354 ;
  assign n10518 = n10517 ^ x228 ^ 1'b0 ;
  assign n10519 = ~n10516 & n10518 ;
  assign n10520 = ~n1697 & n5373 ;
  assign n10521 = n3112 & n10520 ;
  assign n10522 = n10521 ^ n8604 ^ 1'b0 ;
  assign n10523 = n4529 ^ n1085 ^ 1'b0 ;
  assign n10524 = n10523 ^ n781 ^ 1'b0 ;
  assign n10525 = n10140 & n10524 ;
  assign n10526 = n8118 | n10525 ;
  assign n10527 = n9003 ^ n2827 ^ 1'b0 ;
  assign n10528 = n2013 & n9102 ;
  assign n10529 = n6700 & n10528 ;
  assign n10530 = n1159 & n10529 ;
  assign n10531 = n3373 & n10530 ;
  assign n10532 = n1207 | n9068 ;
  assign n10533 = n10532 ^ n6812 ^ 1'b0 ;
  assign n10534 = n1594 & n10533 ;
  assign n10535 = ~n10531 & n10534 ;
  assign n10536 = n1857 & n4164 ;
  assign n10537 = n3197 & n10536 ;
  assign n10538 = n1950 & n2011 ;
  assign n10539 = ~n3552 & n10538 ;
  assign n10540 = ~n10537 & n10539 ;
  assign n10541 = n3599 ^ n2021 ^ 1'b0 ;
  assign n10542 = n895 | n4336 ;
  assign n10543 = n10541 & ~n10542 ;
  assign n10544 = ~x25 & n2846 ;
  assign n10545 = n10543 & n10544 ;
  assign n10550 = ~n623 & n1560 ;
  assign n10546 = x197 & ~n1717 ;
  assign n10547 = ~n987 & n5025 ;
  assign n10548 = n10546 & ~n10547 ;
  assign n10549 = n5876 & n10548 ;
  assign n10551 = n10550 ^ n10549 ^ 1'b0 ;
  assign n10552 = n760 | n5132 ;
  assign n10553 = n10552 ^ n2213 ^ 1'b0 ;
  assign n10554 = n10495 ^ n1016 ^ 1'b0 ;
  assign n10555 = n3331 | n10554 ;
  assign n10556 = n6293 & ~n10555 ;
  assign n10557 = ( n723 & n4242 ) | ( n723 & ~n7212 ) | ( n4242 & ~n7212 ) ;
  assign n10558 = n2918 & ~n5527 ;
  assign n10559 = ~n987 & n8201 ;
  assign n10560 = ~x44 & n593 ;
  assign n10561 = n10559 | n10560 ;
  assign n10562 = ~n3181 & n9837 ;
  assign n10563 = n10562 ^ n1621 ^ 1'b0 ;
  assign n10564 = n1535 | n3032 ;
  assign n10570 = n4499 ^ n1059 ^ 1'b0 ;
  assign n10571 = n8538 | n10570 ;
  assign n10566 = n5059 ^ x91 ^ 1'b0 ;
  assign n10565 = ~n456 & n6999 ;
  assign n10567 = n10566 ^ n10565 ^ 1'b0 ;
  assign n10568 = n6253 & n10567 ;
  assign n10569 = ~n2711 & n10568 ;
  assign n10572 = n10571 ^ n10569 ^ 1'b0 ;
  assign n10573 = ~n10564 & n10572 ;
  assign n10574 = n9487 ^ n8921 ^ 1'b0 ;
  assign n10575 = n3768 & ~n10574 ;
  assign n10576 = ~n3633 & n10575 ;
  assign n10577 = ( n2188 & n7232 ) | ( n2188 & n10149 ) | ( n7232 & n10149 ) ;
  assign n10578 = n442 | n920 ;
  assign n10579 = n10578 ^ n1646 ^ 1'b0 ;
  assign n10580 = n655 & ~n10579 ;
  assign n10581 = ~n1877 & n10580 ;
  assign n10582 = n10581 ^ n862 ^ 1'b0 ;
  assign n10583 = n10582 ^ n3739 ^ 1'b0 ;
  assign n10584 = ~n5262 & n7262 ;
  assign n10585 = n7905 ^ n562 ^ 1'b0 ;
  assign n10586 = n7436 ^ n3480 ^ 1'b0 ;
  assign n10587 = ~n10585 & n10586 ;
  assign n10588 = n1079 & n10354 ;
  assign n10589 = ~n535 & n4772 ;
  assign n10590 = n3618 & n10589 ;
  assign n10591 = n618 & n3364 ;
  assign n10592 = n10591 ^ n514 ^ 1'b0 ;
  assign n10593 = n10590 | n10592 ;
  assign n10594 = n2022 | n6504 ;
  assign n10595 = n10594 ^ n7284 ^ 1'b0 ;
  assign n10596 = x190 & ~n1210 ;
  assign n10597 = n2769 | n7140 ;
  assign n10598 = n7681 | n10597 ;
  assign n10599 = n10596 | n10598 ;
  assign n10600 = x44 & ~n10259 ;
  assign n10601 = n10600 ^ n1736 ^ 1'b0 ;
  assign n10602 = n6990 ^ n1967 ^ 1'b0 ;
  assign n10603 = n4363 ^ n3405 ^ 1'b0 ;
  assign n10604 = ~n6082 & n10603 ;
  assign n10605 = n5610 & ~n6715 ;
  assign n10606 = n1158 | n1904 ;
  assign n10607 = n1446 & ~n3359 ;
  assign n10608 = n791 | n10607 ;
  assign n10609 = n10606 | n10608 ;
  assign n10610 = n10609 ^ n4982 ^ 1'b0 ;
  assign n10611 = n3950 ^ n3755 ^ 1'b0 ;
  assign n10612 = ~n7272 & n10611 ;
  assign n10613 = n3428 | n5105 ;
  assign n10614 = ~n896 & n10613 ;
  assign n10615 = n4306 ^ n971 ^ n808 ;
  assign n10616 = n10615 ^ n10603 ^ n1056 ;
  assign n10617 = n498 & ~n1361 ;
  assign n10618 = n3561 ^ n1070 ^ 1'b0 ;
  assign n10619 = n6215 & n10618 ;
  assign n10620 = ~n8611 & n10619 ;
  assign n10621 = n4485 | n10620 ;
  assign n10622 = n10621 ^ n3484 ^ 1'b0 ;
  assign n10623 = n2966 ^ n1646 ^ 1'b0 ;
  assign n10624 = n7520 ^ n472 ^ 1'b0 ;
  assign n10625 = ~n1903 & n2542 ;
  assign n10626 = n8538 & n10625 ;
  assign n10627 = ~n2731 & n10626 ;
  assign n10628 = x65 & ~n7343 ;
  assign n10629 = ~n1793 & n10628 ;
  assign n10630 = ~n1512 & n2531 ;
  assign n10631 = n2252 ^ n1467 ^ 1'b0 ;
  assign n10632 = n10630 | n10631 ;
  assign n10636 = ~n2770 & n7325 ;
  assign n10637 = n10636 ^ n2070 ^ 1'b0 ;
  assign n10638 = n10637 ^ n1207 ^ 1'b0 ;
  assign n10639 = n1529 & n9149 ;
  assign n10640 = n10638 & n10639 ;
  assign n10633 = n4473 ^ x128 ^ 1'b0 ;
  assign n10634 = n10633 ^ n7929 ^ 1'b0 ;
  assign n10635 = n2736 & n10634 ;
  assign n10641 = n10640 ^ n10635 ^ 1'b0 ;
  assign n10642 = n3239 & ~n10641 ;
  assign n10643 = n2188 & ~n3545 ;
  assign n10644 = n3405 ^ n800 ^ 1'b0 ;
  assign n10645 = ~n4932 & n10644 ;
  assign n10646 = n10645 ^ n7768 ^ 1'b0 ;
  assign n10647 = n1427 | n5535 ;
  assign n10648 = n10370 | n10647 ;
  assign n10649 = n996 | n10648 ;
  assign n10650 = n3153 ^ n633 ^ 1'b0 ;
  assign n10651 = n4497 & n10650 ;
  assign n10652 = n10651 ^ n4534 ^ 1'b0 ;
  assign n10653 = n2420 & ~n10652 ;
  assign n10654 = ~n294 & n8209 ;
  assign n10655 = n10654 ^ n7153 ^ 1'b0 ;
  assign n10657 = n5442 ^ x12 ^ 1'b0 ;
  assign n10658 = n2352 & n10657 ;
  assign n10656 = n2429 & ~n2712 ;
  assign n10659 = n10658 ^ n10656 ^ 1'b0 ;
  assign n10660 = n545 | n3828 ;
  assign n10661 = n333 | n10660 ;
  assign n10662 = n1635 & n2816 ;
  assign n10663 = ~n3976 & n10662 ;
  assign n10664 = n7312 & ~n10663 ;
  assign n10665 = ~n10661 & n10664 ;
  assign n10666 = n7370 & n8737 ;
  assign n10667 = n1249 & n2998 ;
  assign n10668 = n2858 & n10667 ;
  assign n10669 = n566 & n10668 ;
  assign n10671 = n2065 ^ n1783 ^ 1'b0 ;
  assign n10670 = ~n683 & n1589 ;
  assign n10672 = n10671 ^ n10670 ^ 1'b0 ;
  assign n10673 = n3554 ^ n812 ^ 1'b0 ;
  assign n10674 = n7137 & ~n10673 ;
  assign n10677 = n1290 | n3931 ;
  assign n10676 = n3610 & ~n5124 ;
  assign n10678 = n10677 ^ n10676 ^ 1'b0 ;
  assign n10675 = n7648 ^ n4538 ^ 1'b0 ;
  assign n10679 = n10678 ^ n10675 ^ 1'b0 ;
  assign n10680 = n6171 & n8628 ;
  assign n10681 = n4848 & n10680 ;
  assign n10682 = n10541 ^ x41 ^ 1'b0 ;
  assign n10683 = ~x178 & n10682 ;
  assign n10684 = n5504 & n10683 ;
  assign n10685 = n2423 & ~n3750 ;
  assign n10686 = n5531 & ~n10685 ;
  assign n10687 = n10686 ^ n7384 ^ 1'b0 ;
  assign n10688 = n354 & ~n4766 ;
  assign n10689 = n10688 ^ n6433 ^ 1'b0 ;
  assign n10690 = n7149 & ~n10689 ;
  assign n10691 = n9487 ^ n9417 ^ 1'b0 ;
  assign n10692 = ( n3750 & ~n4112 ) | ( n3750 & n10691 ) | ( ~n4112 & n10691 ) ;
  assign n10693 = x235 & ~n4884 ;
  assign n10694 = ~x29 & n10693 ;
  assign n10695 = n10375 | n10694 ;
  assign n10696 = n4382 | n8160 ;
  assign n10697 = n10696 ^ n1328 ^ 1'b0 ;
  assign n10698 = n820 & ~n6511 ;
  assign n10699 = ~n3903 & n5452 ;
  assign n10700 = ~n5358 & n10699 ;
  assign n10701 = n5167 ^ n1321 ^ 1'b0 ;
  assign n10702 = n4764 ^ n4260 ^ 1'b0 ;
  assign n10703 = ~n3112 & n5618 ;
  assign n10704 = n6121 & n6368 ;
  assign n10705 = n10704 ^ n9714 ^ 1'b0 ;
  assign n10706 = n6991 | n9678 ;
  assign n10707 = n2672 ^ n522 ^ 1'b0 ;
  assign n10708 = n10706 & n10707 ;
  assign n10709 = n4755 ^ n3533 ^ 1'b0 ;
  assign n10710 = n6050 ^ n4220 ^ 1'b0 ;
  assign n10711 = n2912 | n10710 ;
  assign n10712 = n10711 ^ n655 ^ 1'b0 ;
  assign n10713 = n2439 & ~n9220 ;
  assign n10714 = n10713 ^ n6821 ^ 1'b0 ;
  assign n10715 = n10714 ^ n5401 ^ 1'b0 ;
  assign n10716 = n8212 | n10715 ;
  assign n10717 = n3729 ^ n1991 ^ 1'b0 ;
  assign n10718 = n10717 ^ n7667 ^ 1'b0 ;
  assign n10719 = n5170 ^ n4345 ^ 1'b0 ;
  assign n10720 = n10719 ^ n3639 ^ 1'b0 ;
  assign n10721 = n2239 & n10720 ;
  assign n10722 = n9449 ^ n5140 ^ 1'b0 ;
  assign n10723 = ~n1728 & n10722 ;
  assign n10724 = n9254 | n10281 ;
  assign n10725 = n2700 & n4065 ;
  assign n10726 = ~x67 & n611 ;
  assign n10727 = n4562 & n10726 ;
  assign n10728 = n10226 & n10727 ;
  assign n10729 = n1234 | n10728 ;
  assign n10730 = n7760 & n9977 ;
  assign n10731 = n10730 ^ n4013 ^ 1'b0 ;
  assign n10732 = ~n875 & n10731 ;
  assign n10733 = n10729 & n10732 ;
  assign n10738 = n3814 ^ n1910 ^ 1'b0 ;
  assign n10739 = n3748 & n10738 ;
  assign n10737 = n2322 | n7387 ;
  assign n10740 = n10739 ^ n10737 ^ 1'b0 ;
  assign n10734 = n1703 | n1863 ;
  assign n10735 = n430 & ~n10734 ;
  assign n10736 = n4733 | n10735 ;
  assign n10741 = n10740 ^ n10736 ^ 1'b0 ;
  assign n10742 = ( n6253 & n6698 ) | ( n6253 & ~n10615 ) | ( n6698 & ~n10615 ) ;
  assign n10743 = n8087 ^ n1351 ^ 1'b0 ;
  assign n10744 = n708 | n10743 ;
  assign n10745 = n6491 ^ n5905 ^ 1'b0 ;
  assign n10746 = ~n10744 & n10745 ;
  assign n10747 = n8501 & n10746 ;
  assign n10748 = n8481 & ~n10747 ;
  assign n10749 = n10546 ^ n1710 ^ 1'b0 ;
  assign n10750 = n361 & ~n10749 ;
  assign n10751 = ~n3740 & n10750 ;
  assign n10752 = n7679 ^ n1677 ^ 1'b0 ;
  assign n10753 = n1402 & ~n10752 ;
  assign n10754 = n5023 & n10038 ;
  assign n10755 = n2555 | n10754 ;
  assign n10756 = n10755 ^ n7274 ^ 1'b0 ;
  assign n10757 = n7736 | n10756 ;
  assign n10758 = n4119 & n4278 ;
  assign n10759 = n4223 ^ n3436 ^ 1'b0 ;
  assign n10760 = n6990 & n10759 ;
  assign n10762 = ~n488 & n5261 ;
  assign n10763 = n10762 ^ x57 ^ 1'b0 ;
  assign n10761 = n5026 & n7028 ;
  assign n10764 = n10763 ^ n10761 ^ 1'b0 ;
  assign n10765 = n8796 ^ n3899 ^ 1'b0 ;
  assign n10766 = ~n9713 & n10765 ;
  assign n10767 = n2678 & ~n3324 ;
  assign n10768 = n8460 ^ n858 ^ 1'b0 ;
  assign n10769 = n10430 ^ n4698 ^ 1'b0 ;
  assign n10770 = x25 & n10769 ;
  assign n10771 = n8625 ^ n3153 ^ 1'b0 ;
  assign n10772 = ~n3641 & n6665 ;
  assign n10773 = n8263 & n10772 ;
  assign n10774 = n6479 & n8165 ;
  assign n10775 = n10313 ^ n7526 ^ 1'b0 ;
  assign n10776 = n6373 | n10775 ;
  assign n10777 = n8444 ^ n4660 ^ 1'b0 ;
  assign n10778 = n7844 & n9163 ;
  assign n10779 = n5761 ^ n5341 ^ n4129 ;
  assign n10780 = n2517 & ~n10779 ;
  assign n10781 = ~n9239 & n9692 ;
  assign n10782 = n8833 ^ n1775 ^ 1'b0 ;
  assign n10783 = x28 & x111 ;
  assign n10784 = n8170 & ~n9802 ;
  assign n10785 = ~n8823 & n10784 ;
  assign n10786 = n1671 & ~n2536 ;
  assign n10787 = n10786 ^ n6830 ^ 1'b0 ;
  assign n10788 = n1436 | n2870 ;
  assign n10789 = n5634 ^ n2492 ^ 1'b0 ;
  assign n10790 = n8885 & ~n10789 ;
  assign n10791 = ~n10788 & n10790 ;
  assign n10792 = n10787 & n10791 ;
  assign n10794 = n2578 & ~n4695 ;
  assign n10793 = n3670 & n9040 ;
  assign n10795 = n10794 ^ n10793 ^ 1'b0 ;
  assign n10796 = x67 & ~n1680 ;
  assign n10797 = ~n6020 & n10796 ;
  assign n10798 = n3240 | n10797 ;
  assign n10799 = x97 & ~n2938 ;
  assign n10800 = n10799 ^ n3917 ^ 1'b0 ;
  assign n10801 = n5271 | n6942 ;
  assign n10802 = n10800 & n10801 ;
  assign n10803 = n10802 ^ n8888 ^ 1'b0 ;
  assign n10806 = ~n1646 & n2001 ;
  assign n10807 = n10806 ^ n4103 ^ 1'b0 ;
  assign n10808 = n698 | n10807 ;
  assign n10804 = ~x213 & n4195 ;
  assign n10805 = ~n2402 & n10804 ;
  assign n10809 = n10808 ^ n10805 ^ 1'b0 ;
  assign n10813 = n1173 & ~n3132 ;
  assign n10810 = n958 & n2148 ;
  assign n10811 = ~n5562 & n10810 ;
  assign n10812 = n6200 | n10811 ;
  assign n10814 = n10813 ^ n10812 ^ 1'b0 ;
  assign n10815 = n10814 ^ n4601 ^ 1'b0 ;
  assign n10816 = n10815 ^ n3537 ^ 1'b0 ;
  assign n10817 = n9470 ^ n673 ^ 1'b0 ;
  assign n10818 = n8087 ^ n2400 ^ 1'b0 ;
  assign n10820 = n557 & n1972 ;
  assign n10819 = x68 & n7249 ;
  assign n10821 = n10820 ^ n10819 ^ 1'b0 ;
  assign n10822 = n1981 ^ n323 ^ 1'b0 ;
  assign n10823 = n1937 | n7601 ;
  assign n10824 = n10823 ^ n4295 ^ 1'b0 ;
  assign n10825 = ~n562 & n6576 ;
  assign n10826 = ~n2812 & n10825 ;
  assign n10827 = n7230 ^ n5385 ^ 1'b0 ;
  assign n10828 = n10827 ^ n1111 ^ 1'b0 ;
  assign n10829 = ~n10826 & n10828 ;
  assign n10830 = n809 & n10829 ;
  assign n10831 = n3540 & n10830 ;
  assign n10832 = n4734 ^ n2283 ^ 1'b0 ;
  assign n10833 = x245 & n10832 ;
  assign n10834 = n3484 & ~n10833 ;
  assign n10835 = n2591 & n8995 ;
  assign n10836 = n10834 & ~n10835 ;
  assign n10837 = n1620 | n8998 ;
  assign n10838 = n10837 ^ n2528 ^ 1'b0 ;
  assign n10839 = ~n539 & n1892 ;
  assign n10840 = ~n1738 & n10839 ;
  assign n10841 = n1935 & ~n10840 ;
  assign n10842 = n10841 ^ n10158 ^ 1'b0 ;
  assign n10843 = n10540 ^ n10141 ^ 1'b0 ;
  assign n10844 = n3130 ^ n2001 ^ 1'b0 ;
  assign n10845 = n7668 ^ n5484 ^ 1'b0 ;
  assign n10846 = n7303 | n10845 ;
  assign n10847 = n1330 & ~n10846 ;
  assign n10848 = ~n696 & n1793 ;
  assign n10849 = n10848 ^ n294 ^ 1'b0 ;
  assign n10850 = ~n3175 & n10849 ;
  assign n10851 = n9719 & n10850 ;
  assign n10852 = n3020 & n3845 ;
  assign n10853 = ~n4366 & n10852 ;
  assign n10854 = n3091 & n10853 ;
  assign n10855 = n1742 & n6425 ;
  assign n10856 = n736 | n6856 ;
  assign n10857 = n5152 ^ n3334 ^ 1'b0 ;
  assign n10858 = n10857 ^ n5125 ^ n1007 ;
  assign n10859 = n8768 | n8908 ;
  assign n10860 = n5828 & n10859 ;
  assign n10861 = n1879 ^ n1563 ^ 1'b0 ;
  assign n10862 = n3714 ^ n1262 ^ 1'b0 ;
  assign n10863 = ~n10861 & n10862 ;
  assign n10864 = n10082 ^ n5804 ^ n1029 ;
  assign n10865 = n2197 ^ n527 ^ 1'b0 ;
  assign n10866 = n6195 | n10865 ;
  assign n10867 = n6458 | n10866 ;
  assign n10868 = ~n480 & n1549 ;
  assign n10869 = n3953 ^ n3171 ^ 1'b0 ;
  assign n10870 = n10869 ^ n2148 ^ 1'b0 ;
  assign n10871 = n10868 & n10870 ;
  assign n10872 = n9302 & n10140 ;
  assign n10873 = n10872 ^ n4579 ^ 1'b0 ;
  assign n10875 = n3951 ^ n2491 ^ 1'b0 ;
  assign n10876 = n10875 ^ n493 ^ 1'b0 ;
  assign n10877 = n4962 | n10876 ;
  assign n10874 = n3191 & ~n9371 ;
  assign n10878 = n10877 ^ n10874 ^ 1'b0 ;
  assign n10879 = n5492 ^ n1181 ^ 1'b0 ;
  assign n10880 = ~n4010 & n10879 ;
  assign n10881 = n10880 ^ n4579 ^ 1'b0 ;
  assign n10882 = n9445 & n10881 ;
  assign n10883 = n10882 ^ n4290 ^ 1'b0 ;
  assign n10884 = n1450 & ~n10883 ;
  assign n10885 = ~n2440 & n10884 ;
  assign n10886 = n7146 ^ n5692 ^ 1'b0 ;
  assign n10887 = ~n360 & n1947 ;
  assign n10888 = n10887 ^ x174 ^ x128 ;
  assign n10889 = ~n2576 & n8655 ;
  assign n10890 = ~n5356 & n10889 ;
  assign n10891 = n2565 & n2733 ;
  assign n10892 = n10891 ^ n1882 ^ 1'b0 ;
  assign n10893 = n5259 & ~n10892 ;
  assign n10894 = ~n2392 & n9913 ;
  assign n10895 = n10894 ^ n6317 ^ 1'b0 ;
  assign n10896 = n7483 ^ n4627 ^ 1'b0 ;
  assign n10897 = n10188 & n10896 ;
  assign n10898 = n10897 ^ n3670 ^ 1'b0 ;
  assign n10899 = n4209 ^ n3419 ^ 1'b0 ;
  assign n10900 = n8538 | n10899 ;
  assign n10901 = ~n7884 & n9071 ;
  assign n10902 = n10901 ^ n4548 ^ 1'b0 ;
  assign n10903 = ~n10900 & n10902 ;
  assign n10904 = n10903 ^ n10056 ^ 1'b0 ;
  assign n10905 = x112 | n1917 ;
  assign n10906 = n7890 | n10905 ;
  assign n10907 = n5050 | n6491 ;
  assign n10908 = n10907 ^ n2019 ^ 1'b0 ;
  assign n10909 = n10908 ^ n3621 ^ 1'b0 ;
  assign n10910 = x194 & n859 ;
  assign n10911 = ~n2698 & n10910 ;
  assign n10912 = n7494 ^ n3499 ^ 1'b0 ;
  assign n10913 = n3503 & n4291 ;
  assign n10914 = n4328 & n5726 ;
  assign n10915 = n6522 & ~n6794 ;
  assign n10916 = n4431 & ~n10348 ;
  assign n10917 = ~n4617 & n10916 ;
  assign n10918 = n10917 ^ n7611 ^ 1'b0 ;
  assign n10919 = n2735 ^ n1379 ^ 1'b0 ;
  assign n10920 = x141 & ~n6431 ;
  assign n10921 = n10920 ^ n3240 ^ 1'b0 ;
  assign n10922 = n2423 & ~n10921 ;
  assign n10923 = n1977 & ~n5849 ;
  assign n10924 = ~n2438 & n10923 ;
  assign n10925 = n3727 | n10924 ;
  assign n10926 = n7148 & ~n10925 ;
  assign n10927 = n3433 ^ n1027 ^ 1'b0 ;
  assign n10928 = ~n10926 & n10927 ;
  assign n10929 = x137 & n1883 ;
  assign n10930 = n3847 & n8727 ;
  assign n10931 = ~n4719 & n10930 ;
  assign n10932 = n9558 ^ n5913 ^ 1'b0 ;
  assign n10933 = ( ~n8237 & n10931 ) | ( ~n8237 & n10932 ) | ( n10931 & n10932 ) ;
  assign n10934 = n6456 & n9238 ;
  assign n10935 = n4300 & n10934 ;
  assign n10936 = n3235 & ~n10935 ;
  assign n10937 = x113 | n3204 ;
  assign n10938 = n1429 & ~n3006 ;
  assign n10939 = n4846 & n10938 ;
  assign n10940 = n10937 & ~n10939 ;
  assign n10941 = n10940 ^ n2216 ^ 1'b0 ;
  assign n10942 = n607 | n10941 ;
  assign n10943 = ~n521 & n8611 ;
  assign n10944 = n10943 ^ x174 ^ 1'b0 ;
  assign n10945 = n10944 ^ n911 ^ 1'b0 ;
  assign n10946 = x149 & ~n10945 ;
  assign n10947 = ~n1980 & n6372 ;
  assign n10948 = ~n8713 & n10947 ;
  assign n10949 = n1682 & n7043 ;
  assign n10950 = n10949 ^ n1683 ^ 1'b0 ;
  assign n10951 = n7443 & ~n9086 ;
  assign n10952 = n3695 ^ n2136 ^ 1'b0 ;
  assign n10953 = n1488 & ~n10952 ;
  assign n10954 = n8329 ^ n1569 ^ 1'b0 ;
  assign n10955 = n859 & ~n4130 ;
  assign n10956 = n1736 & n4954 ;
  assign n10957 = n10956 ^ n5535 ^ 1'b0 ;
  assign n10958 = ~n412 & n5698 ;
  assign n10959 = n7888 | n8406 ;
  assign n10960 = n10959 ^ n2757 ^ 1'b0 ;
  assign n10961 = n3145 ^ n1018 ^ 1'b0 ;
  assign n10962 = ~n9094 & n10961 ;
  assign n10963 = n4107 & n5879 ;
  assign n10964 = x184 & n10963 ;
  assign n10965 = ~n8727 & n10964 ;
  assign n10969 = n4555 ^ n3016 ^ 1'b0 ;
  assign n10966 = n1379 & n1670 ;
  assign n10967 = ~n8281 & n10966 ;
  assign n10968 = n10967 ^ n3049 ^ 1'b0 ;
  assign n10970 = n10969 ^ n10968 ^ 1'b0 ;
  assign n10971 = n4705 ^ n733 ^ 1'b0 ;
  assign n10972 = n4416 & n10971 ;
  assign n10973 = n7451 ^ n3678 ^ 1'b0 ;
  assign n10974 = n10972 & ~n10973 ;
  assign n10975 = n956 | n10877 ;
  assign n10976 = n10975 ^ n6809 ^ 1'b0 ;
  assign n10977 = n10976 ^ n6541 ^ 1'b0 ;
  assign n10978 = ~n10352 & n10977 ;
  assign n10979 = n10974 & ~n10978 ;
  assign n10980 = n286 & n7627 ;
  assign n10981 = x133 | n300 ;
  assign n10982 = n5730 & n9951 ;
  assign n10983 = ~n9935 & n10982 ;
  assign n10984 = n3893 ^ n1442 ^ 1'b0 ;
  assign n10985 = n2877 & ~n10984 ;
  assign n10986 = n2292 & n10985 ;
  assign n10987 = n8283 & ~n8829 ;
  assign n10988 = n1291 & n10987 ;
  assign n10989 = n5280 | n6585 ;
  assign n10990 = n5686 | n10989 ;
  assign n10991 = n10990 ^ n9083 ^ 1'b0 ;
  assign n10992 = n3040 | n5690 ;
  assign n10993 = n10992 ^ n4886 ^ 1'b0 ;
  assign n10994 = ( n8512 & ~n9639 ) | ( n8512 & n10993 ) | ( ~n9639 & n10993 ) ;
  assign n10995 = n1795 & ~n7466 ;
  assign n10996 = n10995 ^ n10888 ^ 1'b0 ;
  assign n10997 = ~n2142 & n2281 ;
  assign n10998 = n7362 & ~n10997 ;
  assign n10999 = n8609 & n10998 ;
  assign n11000 = n2037 ^ n803 ^ 1'b0 ;
  assign n11001 = x181 & n11000 ;
  assign n11002 = n1075 & n7597 ;
  assign n11003 = ~n11001 & n11002 ;
  assign n11004 = ~n4803 & n5945 ;
  assign n11005 = n11004 ^ n7942 ^ n5696 ;
  assign n11006 = n6768 | n10744 ;
  assign n11007 = n423 | n11006 ;
  assign n11008 = n1745 | n5450 ;
  assign n11009 = n11008 ^ n10887 ^ 1'b0 ;
  assign n11010 = n11007 & ~n11009 ;
  assign n11011 = n1252 & ~n2700 ;
  assign n11012 = n11011 ^ n538 ^ 1'b0 ;
  assign n11013 = n1337 & n11012 ;
  assign n11014 = n10187 ^ n3855 ^ 1'b0 ;
  assign n11015 = n11014 ^ n2180 ^ 1'b0 ;
  assign n11016 = n11013 & ~n11015 ;
  assign n11017 = n2644 | n6663 ;
  assign n11018 = n2644 & ~n11017 ;
  assign n11028 = ~n4267 & n7451 ;
  assign n11029 = n4267 & n11028 ;
  assign n11030 = ~n1910 & n11029 ;
  assign n11019 = x71 & x90 ;
  assign n11020 = ~x71 & n11019 ;
  assign n11021 = x223 & ~n11020 ;
  assign n11022 = ~x223 & n11021 ;
  assign n11023 = n4124 & ~n11022 ;
  assign n11024 = ~n4124 & n11023 ;
  assign n11025 = n623 | n11024 ;
  assign n11026 = n623 & ~n11025 ;
  assign n11027 = n4913 | n11026 ;
  assign n11031 = n11030 ^ n11027 ^ 1'b0 ;
  assign n11032 = ~n11018 & n11031 ;
  assign n11033 = x218 & ~n3943 ;
  assign n11034 = n11033 ^ n4484 ^ 1'b0 ;
  assign n11035 = ~n9345 & n11034 ;
  assign n11036 = n9345 & n11035 ;
  assign n11037 = n9296 ^ n8509 ^ x82 ;
  assign n11038 = n8879 ^ n1031 ^ 1'b0 ;
  assign n11039 = n8461 & ~n10002 ;
  assign n11040 = n4554 & n11039 ;
  assign n11041 = n5444 ^ n3862 ^ 1'b0 ;
  assign n11042 = n9569 | n11041 ;
  assign n11043 = n11042 ^ n7109 ^ 1'b0 ;
  assign n11044 = n10762 & n11043 ;
  assign n11045 = ~n7458 & n11044 ;
  assign n11046 = ~x68 & n3368 ;
  assign n11047 = n3591 & n9188 ;
  assign n11048 = n2931 & n11047 ;
  assign n11049 = n1977 & n5175 ;
  assign n11050 = n11049 ^ n2021 ^ 1'b0 ;
  assign n11051 = ~n2047 & n11050 ;
  assign n11052 = n2892 & n11051 ;
  assign n11053 = ~n407 & n6975 ;
  assign n11054 = n11052 & n11053 ;
  assign n11055 = n11054 ^ n10944 ^ 1'b0 ;
  assign n11056 = n2576 ^ n1614 ^ 1'b0 ;
  assign n11057 = n2715 | n11056 ;
  assign n11058 = n11057 ^ n5510 ^ 1'b0 ;
  assign n11059 = ( ~x222 & n2642 ) | ( ~x222 & n8489 ) | ( n2642 & n8489 ) ;
  assign n11060 = n4689 ^ x190 ^ 1'b0 ;
  assign n11061 = n11059 | n11060 ;
  assign n11062 = ~n8201 & n9682 ;
  assign n11063 = n11062 ^ n6049 ^ 1'b0 ;
  assign n11064 = n8947 ^ n4931 ^ 1'b0 ;
  assign n11065 = n11063 & ~n11064 ;
  assign n11066 = ~n2256 & n8479 ;
  assign n11067 = ~n476 & n8596 ;
  assign n11068 = x106 | n11067 ;
  assign n11069 = n7868 ^ n2837 ^ n2715 ;
  assign n11070 = n6123 | n11069 ;
  assign n11071 = n11070 ^ n3143 ^ 1'b0 ;
  assign n11072 = ( n1111 & n3591 ) | ( n1111 & ~n8773 ) | ( n3591 & ~n8773 ) ;
  assign n11073 = n11072 ^ x27 ^ 1'b0 ;
  assign n11074 = n5285 ^ n985 ^ 1'b0 ;
  assign n11075 = n4753 & ~n4804 ;
  assign n11076 = n11075 ^ n540 ^ 1'b0 ;
  assign n11077 = n4366 & n11076 ;
  assign n11078 = n7621 | n10747 ;
  assign n11079 = n4617 & ~n11078 ;
  assign n11080 = n11079 ^ n5261 ^ 1'b0 ;
  assign n11081 = n7901 ^ n7809 ^ 1'b0 ;
  assign n11082 = n10423 ^ x155 ^ 1'b0 ;
  assign n11083 = n4276 & n8014 ;
  assign n11084 = n10559 | n11083 ;
  assign n11085 = n11084 ^ n7076 ^ 1'b0 ;
  assign n11086 = n2415 & n11085 ;
  assign n11087 = n6751 & n11086 ;
  assign n11088 = n1772 | n2142 ;
  assign n11089 = n11088 ^ n10120 ^ 1'b0 ;
  assign n11090 = x141 & n3356 ;
  assign n11091 = n11090 ^ n8703 ^ 1'b0 ;
  assign n11092 = x100 & ~n598 ;
  assign n11093 = n11092 ^ x3 ^ 1'b0 ;
  assign n11094 = n8090 & n10150 ;
  assign n11095 = n11094 ^ n5464 ^ 1'b0 ;
  assign n11096 = n11093 & ~n11095 ;
  assign n11097 = ( n296 & ~n1839 ) | ( n296 & n6573 ) | ( ~n1839 & n6573 ) ;
  assign n11098 = ~n3854 & n4851 ;
  assign n11099 = ~n11097 & n11098 ;
  assign n11100 = ~n1483 & n1485 ;
  assign n11101 = n11100 ^ n4930 ^ 1'b0 ;
  assign n11102 = n10762 ^ n3179 ^ 1'b0 ;
  assign n11103 = n3022 | n11102 ;
  assign n11104 = ~n11101 & n11103 ;
  assign n11105 = n593 & n1226 ;
  assign n11106 = n3130 | n3298 ;
  assign n11107 = n11105 | n11106 ;
  assign n11108 = ~n1849 & n11107 ;
  assign n11109 = ~n4376 & n9203 ;
  assign n11110 = n6932 ^ n1318 ^ 1'b0 ;
  assign n11111 = n10540 ^ n3226 ^ 1'b0 ;
  assign n11112 = n11111 ^ n2660 ^ 1'b0 ;
  assign n11113 = ~n11110 & n11112 ;
  assign n11115 = n5920 ^ n2571 ^ 1'b0 ;
  assign n11114 = n7769 & n8715 ;
  assign n11116 = n11115 ^ n11114 ^ 1'b0 ;
  assign n11117 = n8497 ^ n3204 ^ x52 ;
  assign n11118 = ~n749 & n11117 ;
  assign n11119 = n11118 ^ n9955 ^ 1'b0 ;
  assign n11120 = n430 & n1787 ;
  assign n11121 = n1818 ^ x132 ^ 1'b0 ;
  assign n11122 = ~n4743 & n11121 ;
  assign n11123 = n832 & ~n11122 ;
  assign n11124 = n781 & ~n7434 ;
  assign n11125 = n11124 ^ n2643 ^ n2487 ;
  assign n11126 = n10733 ^ n5703 ^ 1'b0 ;
  assign n11127 = n4283 & ~n11126 ;
  assign n11128 = n8200 ^ n1141 ^ 1'b0 ;
  assign n11129 = n11128 ^ n9877 ^ 1'b0 ;
  assign n11130 = n3593 & ~n6438 ;
  assign n11131 = ~n9697 & n11130 ;
  assign n11133 = n2112 ^ n2001 ^ 1'b0 ;
  assign n11134 = n11133 ^ n3772 ^ 1'b0 ;
  assign n11132 = n5381 & n7390 ;
  assign n11135 = n11134 ^ n11132 ^ 1'b0 ;
  assign n11136 = n11135 ^ n2942 ^ 1'b0 ;
  assign n11137 = n1854 & n7263 ;
  assign n11138 = n1696 | n7387 ;
  assign n11139 = n1696 & ~n11138 ;
  assign n11140 = n4122 ^ n1723 ^ 1'b0 ;
  assign n11141 = n538 & n11140 ;
  assign n11142 = n708 & n11141 ;
  assign n11143 = n6031 & ~n11142 ;
  assign n11145 = ~n2577 & n4543 ;
  assign n11146 = n2782 & n11145 ;
  assign n11147 = n11146 ^ n6146 ^ 1'b0 ;
  assign n11144 = n5755 ^ n5575 ^ n951 ;
  assign n11148 = n11147 ^ n11144 ^ 1'b0 ;
  assign n11149 = n4721 & ~n7374 ;
  assign n11150 = n3026 ^ x106 ^ 1'b0 ;
  assign n11151 = n5447 ^ n3181 ^ 1'b0 ;
  assign n11152 = n6587 & ~n11151 ;
  assign n11153 = n5812 ^ n1775 ^ 1'b0 ;
  assign n11154 = n11152 & n11153 ;
  assign n11155 = n3441 | n4360 ;
  assign n11156 = n11155 ^ n1228 ^ 1'b0 ;
  assign n11157 = n1083 & ~n11156 ;
  assign n11158 = ~n6311 & n11157 ;
  assign n11159 = n4680 & ~n10381 ;
  assign n11160 = n1579 ^ n932 ^ 1'b0 ;
  assign n11161 = ~n8328 & n11160 ;
  assign n11162 = ~n3545 & n10197 ;
  assign n11163 = n1825 & ~n5880 ;
  assign n11164 = ~x244 & n11163 ;
  assign n11165 = n1917 & ~n11164 ;
  assign n11166 = n825 | n1354 ;
  assign n11172 = ~x115 & x190 ;
  assign n11167 = n661 & n9183 ;
  assign n11168 = n2629 & ~n11167 ;
  assign n11169 = n11168 ^ n2526 ^ 1'b0 ;
  assign n11170 = n11169 ^ n6038 ^ 1'b0 ;
  assign n11171 = x152 & ~n11170 ;
  assign n11173 = n11172 ^ n11171 ^ 1'b0 ;
  assign n11175 = n833 & n2762 ;
  assign n11174 = n904 | n9693 ;
  assign n11176 = n11175 ^ n11174 ^ 1'b0 ;
  assign n11177 = n10460 ^ n10322 ^ 1'b0 ;
  assign n11179 = n3495 ^ n3239 ^ 1'b0 ;
  assign n11180 = n4723 & n11179 ;
  assign n11178 = n3862 & ~n4133 ;
  assign n11181 = n11180 ^ n11178 ^ 1'b0 ;
  assign n11182 = n11181 ^ n8635 ^ 1'b0 ;
  assign n11183 = n8280 & n11182 ;
  assign n11184 = ~n8638 & n11183 ;
  assign n11185 = n756 & n3765 ;
  assign n11186 = ~n2855 & n8303 ;
  assign n11187 = n11185 & n11186 ;
  assign n11188 = ~n7023 & n7248 ;
  assign n11189 = ~n4385 & n11188 ;
  assign n11190 = n4720 | n5439 ;
  assign n11191 = n482 | n11190 ;
  assign n11192 = n417 & ~n1553 ;
  assign n11193 = n11192 ^ n820 ^ 1'b0 ;
  assign n11194 = n5089 & ~n11193 ;
  assign n11195 = n5530 ^ n1634 ^ 1'b0 ;
  assign n11196 = n5413 & n11195 ;
  assign n11197 = n1630 | n2908 ;
  assign n11198 = n5407 ^ n3700 ^ 1'b0 ;
  assign n11199 = ~n1772 & n11198 ;
  assign n11200 = n5012 | n6735 ;
  assign n11201 = n11200 ^ n349 ^ 1'b0 ;
  assign n11202 = n566 | n11201 ;
  assign n11203 = ~n1125 & n11202 ;
  assign n11204 = n5378 & ~n11203 ;
  assign n11205 = n7862 & ~n11204 ;
  assign n11206 = n4179 ^ n2489 ^ 1'b0 ;
  assign n11207 = ( n4686 & ~n6551 ) | ( n4686 & n11206 ) | ( ~n6551 & n11206 ) ;
  assign n11209 = n872 & ~n1111 ;
  assign n11210 = n5909 & ~n11209 ;
  assign n11208 = n1914 & n9211 ;
  assign n11211 = n11210 ^ n11208 ^ 1'b0 ;
  assign n11212 = x226 & n979 ;
  assign n11213 = n2066 & n11212 ;
  assign n11214 = n3880 | n4238 ;
  assign n11215 = n11214 ^ n10198 ^ 1'b0 ;
  assign n11216 = n11213 | n11215 ;
  assign n11217 = n10606 ^ n3886 ^ n809 ;
  assign n11218 = n11217 ^ n2766 ^ 1'b0 ;
  assign n11219 = n10640 & n11218 ;
  assign n11220 = n7054 ^ n561 ^ x81 ;
  assign n11221 = n10021 | n10327 ;
  assign n11222 = n11221 ^ n7778 ^ 1'b0 ;
  assign n11223 = n11220 & ~n11222 ;
  assign n11224 = ~x178 & n11223 ;
  assign n11225 = n6110 ^ n2590 ^ 1'b0 ;
  assign n11226 = n269 | n11225 ;
  assign n11227 = n1277 ^ x57 ^ 1'b0 ;
  assign n11228 = ~n2510 & n11227 ;
  assign n11229 = n11228 ^ n5755 ^ 1'b0 ;
  assign n11230 = n2423 & ~n11229 ;
  assign n11231 = ~n11226 & n11230 ;
  assign n11232 = ~n2528 & n3616 ;
  assign n11233 = n11232 ^ n6972 ^ 1'b0 ;
  assign n11234 = n956 ^ n930 ^ 1'b0 ;
  assign n11235 = n8509 ^ x67 ^ 1'b0 ;
  assign n11236 = n11234 & n11235 ;
  assign n11237 = ~n1772 & n11236 ;
  assign n11238 = n11237 ^ n4076 ^ 1'b0 ;
  assign n11239 = n11233 | n11238 ;
  assign n11240 = n2076 | n8586 ;
  assign n11241 = n2502 & ~n3333 ;
  assign n11242 = n2760 & ~n11241 ;
  assign n11243 = n6502 | n11242 ;
  assign n11244 = n2527 & n2954 ;
  assign n11245 = n11244 ^ n5151 ^ 1'b0 ;
  assign n11246 = ~n4501 & n8234 ;
  assign n11247 = ( n876 & n8363 ) | ( n876 & ~n10265 ) | ( n8363 & ~n10265 ) ;
  assign n11248 = n8512 ^ n8232 ^ 1'b0 ;
  assign n11249 = n5509 | n11248 ;
  assign n11250 = n11249 ^ n2155 ^ 1'b0 ;
  assign n11251 = n3657 | n10321 ;
  assign n11252 = n11251 ^ n3541 ^ 1'b0 ;
  assign n11253 = ~n3069 & n8442 ;
  assign n11254 = n3666 & n11253 ;
  assign n11255 = n5493 ^ n649 ^ 1'b0 ;
  assign n11256 = n9356 | n11255 ;
  assign n11257 = x73 & n343 ;
  assign n11258 = n1291 & n11257 ;
  assign n11259 = n1501 & ~n3001 ;
  assign n11260 = n2460 | n11259 ;
  assign n11261 = n7830 & ~n11260 ;
  assign n11262 = n6307 & ~n11261 ;
  assign n11263 = n994 & n11262 ;
  assign n11264 = n11258 & n11263 ;
  assign n11265 = n793 & n1935 ;
  assign n11266 = ~n8883 & n11265 ;
  assign n11267 = n6717 ^ n4300 ^ 1'b0 ;
  assign n11268 = ~n11266 & n11267 ;
  assign n11269 = n1738 & n4586 ;
  assign n11270 = n5686 ^ n4418 ^ 1'b0 ;
  assign n11271 = n11269 | n11270 ;
  assign n11272 = n8011 ^ n4676 ^ 1'b0 ;
  assign n11273 = n7613 ^ n5185 ^ n5135 ;
  assign n11274 = n6884 ^ n939 ^ 1'b0 ;
  assign n11275 = ~n6647 & n7135 ;
  assign n11276 = ~n11274 & n11275 ;
  assign n11277 = n1383 | n11276 ;
  assign n11278 = n11277 ^ n4047 ^ 1'b0 ;
  assign n11281 = ~n3750 & n7900 ;
  assign n11279 = n2602 ^ n1919 ^ 1'b0 ;
  assign n11280 = x33 | n11279 ;
  assign n11282 = n11281 ^ n11280 ^ n4598 ;
  assign n11283 = n1900 & n1953 ;
  assign n11284 = n11283 ^ n1818 ^ 1'b0 ;
  assign n11285 = n470 & ~n1513 ;
  assign n11286 = n11285 ^ n5435 ^ 1'b0 ;
  assign n11287 = ~n11284 & n11286 ;
  assign n11290 = n808 | n9440 ;
  assign n11291 = n11290 ^ n4040 ^ 1'b0 ;
  assign n11288 = n6762 ^ n2816 ^ 1'b0 ;
  assign n11289 = ~n5879 & n11288 ;
  assign n11292 = n11291 ^ n11289 ^ 1'b0 ;
  assign n11293 = n11292 ^ x128 ^ 1'b0 ;
  assign n11294 = n8409 ^ n7179 ^ x93 ;
  assign n11295 = n1905 & ~n11294 ;
  assign n11296 = n11295 ^ n3171 ^ 1'b0 ;
  assign n11297 = n4971 & n11296 ;
  assign n11298 = n11297 ^ n3265 ^ 1'b0 ;
  assign n11299 = ~n4480 & n11298 ;
  assign n11300 = n1285 & n11299 ;
  assign n11301 = n11300 ^ n849 ^ 1'b0 ;
  assign n11302 = n4398 & ~n11301 ;
  assign n11303 = n9464 ^ n5579 ^ 1'b0 ;
  assign n11304 = n11302 & n11303 ;
  assign n11305 = n1264 | n6164 ;
  assign n11306 = n1926 | n11305 ;
  assign n11307 = x248 & n11306 ;
  assign n11308 = ~n9955 & n11307 ;
  assign n11309 = n8962 & ~n9695 ;
  assign n11310 = ~n8844 & n11309 ;
  assign n11311 = n8635 ^ n7775 ^ 1'b0 ;
  assign n11312 = ~n4133 & n11311 ;
  assign n11313 = n6771 | n9940 ;
  assign n11314 = n6771 & ~n11313 ;
  assign n11315 = n4251 & ~n11314 ;
  assign n11316 = ~n4251 & n11315 ;
  assign n11317 = n10340 | n11316 ;
  assign n11318 = n2011 & n11317 ;
  assign n11319 = ~n5898 & n11318 ;
  assign n11320 = n895 & ~n1447 ;
  assign n11321 = n11320 ^ n7290 ^ 1'b0 ;
  assign n11322 = n10330 | n11321 ;
  assign n11323 = n1240 & ~n6189 ;
  assign n11324 = n942 & ~n9375 ;
  assign n11325 = n8412 & n11324 ;
  assign n11326 = ~n2093 & n7732 ;
  assign n11327 = n11326 ^ n7097 ^ 1'b0 ;
  assign n11328 = n11327 ^ n3093 ^ 1'b0 ;
  assign n11329 = n9249 ^ n4524 ^ 1'b0 ;
  assign n11330 = n1018 & n1467 ;
  assign n11331 = n5135 & n11330 ;
  assign n11332 = n11331 ^ n5752 ^ n3436 ;
  assign n11333 = n6498 & n9616 ;
  assign n11334 = n3759 | n10349 ;
  assign n11335 = n11334 ^ n5562 ^ 1'b0 ;
  assign n11336 = n6639 ^ x134 ^ 1'b0 ;
  assign n11337 = n725 & n11336 ;
  assign n11338 = n11337 ^ n4538 ^ 1'b0 ;
  assign n11339 = ~n3415 & n11338 ;
  assign n11340 = n4911 & ~n6766 ;
  assign n11341 = ~n1402 & n11340 ;
  assign n11342 = ~n428 & n11341 ;
  assign n11343 = n2338 & ~n7124 ;
  assign n11344 = n11343 ^ n10996 ^ 1'b0 ;
  assign n11345 = n5207 | n10471 ;
  assign n11346 = n6956 ^ n5021 ^ n294 ;
  assign n11347 = ~n2863 & n7572 ;
  assign n11348 = n11347 ^ n10169 ^ 1'b0 ;
  assign n11349 = n6903 ^ n2177 ^ 1'b0 ;
  assign n11350 = n4225 & ~n11349 ;
  assign n11353 = x63 & n3974 ;
  assign n11352 = n2529 | n5411 ;
  assign n11354 = n11353 ^ n11352 ^ 1'b0 ;
  assign n11351 = n4788 & ~n6189 ;
  assign n11355 = n11354 ^ n11351 ^ 1'b0 ;
  assign n11356 = n9071 ^ n5026 ^ 1'b0 ;
  assign n11357 = n4911 & ~n11356 ;
  assign n11358 = n381 & n11357 ;
  assign n11359 = ( n1822 & n3561 ) | ( n1822 & n11358 ) | ( n3561 & n11358 ) ;
  assign n11360 = n5495 & ~n7648 ;
  assign n11361 = n790 & n11360 ;
  assign n11362 = n778 ^ x224 ^ 1'b0 ;
  assign n11363 = ~n869 & n11362 ;
  assign n11364 = ~n7256 & n11363 ;
  assign n11365 = n11364 ^ n3102 ^ 1'b0 ;
  assign n11366 = n10875 & n11365 ;
  assign n11367 = ~n2293 & n11366 ;
  assign n11368 = n11361 & n11367 ;
  assign n11369 = n10318 ^ n8993 ^ 1'b0 ;
  assign n11370 = x27 & ~n11369 ;
  assign n11371 = n4647 ^ x21 ^ 1'b0 ;
  assign n11372 = n11371 ^ x244 ^ 1'b0 ;
  assign n11373 = n305 & n11372 ;
  assign n11374 = n11301 ^ n8879 ^ 1'b0 ;
  assign n11375 = n3162 | n9199 ;
  assign n11376 = n11375 ^ n8223 ^ 1'b0 ;
  assign n11377 = n7560 | n9415 ;
  assign n11378 = n6870 ^ n4372 ^ 1'b0 ;
  assign n11379 = n10008 ^ n6437 ^ 1'b0 ;
  assign n11380 = ~n9785 & n11379 ;
  assign n11381 = x214 & n5323 ;
  assign n11382 = n9407 ^ n4986 ^ 1'b0 ;
  assign n11383 = n4562 | n9485 ;
  assign n11387 = x231 & n2261 ;
  assign n11384 = x5 & ~n1021 ;
  assign n11385 = n7878 & ~n11384 ;
  assign n11386 = n5351 | n11385 ;
  assign n11388 = n11387 ^ n11386 ^ 1'b0 ;
  assign n11389 = n7290 & ~n7800 ;
  assign n11390 = ~n6140 & n11389 ;
  assign n11394 = n6735 ^ n4027 ^ 1'b0 ;
  assign n11391 = n1916 & n2918 ;
  assign n11392 = ~n3226 & n11391 ;
  assign n11393 = n6519 | n11392 ;
  assign n11395 = n11394 ^ n11393 ^ 1'b0 ;
  assign n11396 = n7108 & ~n11395 ;
  assign n11397 = n11396 ^ n5236 ^ 1'b0 ;
  assign n11398 = n10555 ^ n876 ^ 1'b0 ;
  assign n11399 = n8574 ^ x234 ^ 1'b0 ;
  assign n11400 = n5398 & ~n11399 ;
  assign n11401 = n11400 ^ n2046 ^ 1'b0 ;
  assign n11402 = x232 & n11401 ;
  assign n11403 = n6396 ^ n779 ^ 1'b0 ;
  assign n11407 = n430 | n557 ;
  assign n11408 = n430 & ~n11407 ;
  assign n11409 = n639 & ~n11408 ;
  assign n11410 = n11408 & n11409 ;
  assign n11404 = n1762 & ~n7206 ;
  assign n11405 = n7206 & n11404 ;
  assign n11406 = n4398 & ~n11405 ;
  assign n11411 = n11410 ^ n11406 ^ 1'b0 ;
  assign n11412 = n923 & n11411 ;
  assign n11413 = ~n923 & n11412 ;
  assign n11414 = n3303 | n6335 ;
  assign n11415 = x23 & ~n11414 ;
  assign n11416 = n4190 & ~n4382 ;
  assign n11417 = n3789 | n7364 ;
  assign n11418 = ~n9714 & n11417 ;
  assign n11419 = n11418 ^ n10728 ^ 1'b0 ;
  assign n11420 = n11416 & n11419 ;
  assign n11421 = ~n6721 & n11420 ;
  assign n11422 = x51 & ~n4613 ;
  assign n11423 = n11422 ^ n6162 ^ 1'b0 ;
  assign n11424 = n11423 ^ n5265 ^ 1'b0 ;
  assign n11425 = n6747 & n11424 ;
  assign n11426 = n11425 ^ n6255 ^ 1'b0 ;
  assign n11427 = n11426 ^ n6763 ^ 1'b0 ;
  assign n11428 = n3533 | n7785 ;
  assign n11429 = n5821 ^ n2970 ^ 1'b0 ;
  assign n11430 = n1252 & n4872 ;
  assign n11431 = n11430 ^ n5016 ^ 1'b0 ;
  assign n11432 = n11431 ^ n1785 ^ 1'b0 ;
  assign n11436 = n317 | n1929 ;
  assign n11433 = n1390 ^ n956 ^ 1'b0 ;
  assign n11434 = n11433 ^ n1853 ^ 1'b0 ;
  assign n11435 = n1684 & ~n11434 ;
  assign n11437 = n11436 ^ n11435 ^ 1'b0 ;
  assign n11438 = n5398 & ~n11437 ;
  assign n11439 = ~n5200 & n5343 ;
  assign n11440 = n866 & n11439 ;
  assign n11441 = ~n4094 & n11440 ;
  assign n11442 = n1239 | n6884 ;
  assign n11443 = n7345 ^ n3540 ^ 1'b0 ;
  assign n11444 = ~n6068 & n11443 ;
  assign n11445 = n9215 ^ n1415 ^ 1'b0 ;
  assign n11451 = x112 & n1580 ;
  assign n11446 = ~n920 & n7680 ;
  assign n11447 = n920 & n11446 ;
  assign n11448 = n3071 ^ n2017 ^ 1'b0 ;
  assign n11449 = n11448 ^ n4116 ^ 1'b0 ;
  assign n11450 = n11447 | n11449 ;
  assign n11452 = n11451 ^ n11450 ^ 1'b0 ;
  assign n11453 = ~n2315 & n7164 ;
  assign n11454 = ~n1169 & n11374 ;
  assign n11455 = n9053 ^ n8087 ^ 1'b0 ;
  assign n11456 = n2711 | n5562 ;
  assign n11457 = ~n405 & n626 ;
  assign n11458 = n11456 & ~n11457 ;
  assign n11459 = n4189 & n11458 ;
  assign n11460 = ~n3126 & n6525 ;
  assign n11461 = n11460 ^ n10042 ^ 1'b0 ;
  assign n11462 = n10620 ^ n5126 ^ 1'b0 ;
  assign n11463 = n5928 ^ n5390 ^ 1'b0 ;
  assign n11464 = n4872 ^ n2776 ^ 1'b0 ;
  assign n11465 = n390 | n11464 ;
  assign n11466 = n5494 & ~n11465 ;
  assign n11467 = ~x47 & n11466 ;
  assign n11468 = x229 & ~n259 ;
  assign n11469 = n11468 ^ n1399 ^ 1'b0 ;
  assign n11470 = n11469 ^ n11384 ^ 1'b0 ;
  assign n11471 = n1415 & n11470 ;
  assign n11472 = n3649 & n11471 ;
  assign n11473 = n6619 & ~n11472 ;
  assign n11474 = n990 | n2510 ;
  assign n11475 = ~n3943 & n5793 ;
  assign n11476 = ~n3707 & n11475 ;
  assign n11477 = n10325 & ~n11476 ;
  assign n11478 = n11477 ^ n7691 ^ n3899 ;
  assign n11479 = n1002 ^ x23 ^ 1'b0 ;
  assign n11481 = ~n4389 & n5940 ;
  assign n11480 = n2314 & n10873 ;
  assign n11482 = n11481 ^ n11480 ^ 1'b0 ;
  assign n11483 = n8626 ^ n7811 ^ 1'b0 ;
  assign n11484 = n3514 & n11483 ;
  assign n11485 = n5207 & n10414 ;
  assign n11486 = n518 & n11485 ;
  assign n11487 = ~n3331 & n7544 ;
  assign n11488 = ~n1052 & n3941 ;
  assign n11490 = ( ~x228 & n445 ) | ( ~x228 & n3509 ) | ( n445 & n3509 ) ;
  assign n11489 = n7009 & ~n10630 ;
  assign n11491 = n11490 ^ n11489 ^ 1'b0 ;
  assign n11492 = n6382 & ~n9073 ;
  assign n11493 = ~n5093 & n10852 ;
  assign n11494 = ~n2058 & n11493 ;
  assign n11495 = ~x109 & n9643 ;
  assign n11496 = n1557 | n9121 ;
  assign n11497 = n11495 | n11496 ;
  assign n11498 = n11497 ^ n7214 ^ 1'b0 ;
  assign n11499 = n5269 & n7928 ;
  assign n11500 = n11498 & n11499 ;
  assign n11501 = n3200 ^ n1025 ^ 1'b0 ;
  assign n11502 = n9086 ^ n4663 ^ 1'b0 ;
  assign n11503 = n11501 & n11502 ;
  assign n11504 = n11503 ^ n4894 ^ 1'b0 ;
  assign n11505 = ~x22 & n3088 ;
  assign n11506 = n11505 ^ n370 ^ 1'b0 ;
  assign n11507 = n7448 | n9705 ;
  assign n11508 = n1345 & ~n1761 ;
  assign n11509 = n7465 ^ n2190 ^ 1'b0 ;
  assign n11510 = ~n956 & n11509 ;
  assign n11511 = n11508 & n11510 ;
  assign n11512 = n8574 ^ n3206 ^ 1'b0 ;
  assign n11513 = n1787 & ~n5832 ;
  assign n11514 = n11513 ^ n5948 ^ 1'b0 ;
  assign n11515 = n2827 & ~n11514 ;
  assign n11516 = ~x28 & n11515 ;
  assign n11517 = n1551 | n11516 ;
  assign n11518 = n8223 ^ n6343 ^ 1'b0 ;
  assign n11519 = n3707 ^ n1926 ^ 1'b0 ;
  assign n11520 = n11519 ^ n2006 ^ 1'b0 ;
  assign n11521 = ~n573 & n3099 ;
  assign n11522 = n10883 | n11521 ;
  assign n11523 = ~n4699 & n7878 ;
  assign n11524 = n8913 | n11523 ;
  assign n11525 = n3714 & ~n8068 ;
  assign n11526 = ~n10766 & n11525 ;
  assign n11527 = n2908 & ~n6213 ;
  assign n11528 = n11527 ^ n6785 ^ 1'b0 ;
  assign n11532 = n5946 & ~n7181 ;
  assign n11533 = n11532 ^ n1133 ^ 1'b0 ;
  assign n11534 = n10790 & n11533 ;
  assign n11535 = n11534 ^ n2117 ^ 1'b0 ;
  assign n11529 = n3111 & n8002 ;
  assign n11530 = ~n1507 & n11529 ;
  assign n11531 = n4775 | n11530 ;
  assign n11536 = n11535 ^ n11531 ^ 1'b0 ;
  assign n11541 = ~n2080 & n4124 ;
  assign n11542 = n11541 ^ n10441 ^ 1'b0 ;
  assign n11543 = n990 | n11542 ;
  assign n11537 = n9407 ^ n1899 ^ 1'b0 ;
  assign n11538 = n7310 | n11537 ;
  assign n11539 = n11538 ^ n8099 ^ 1'b0 ;
  assign n11540 = n7255 & n11539 ;
  assign n11544 = n11543 ^ n11540 ^ 1'b0 ;
  assign n11545 = n329 | n2316 ;
  assign n11546 = n2316 & ~n11545 ;
  assign n11547 = n1922 & ~n6473 ;
  assign n11548 = n11546 & n11547 ;
  assign n11549 = n11548 ^ n3346 ^ 1'b0 ;
  assign n11550 = ~n430 & n3957 ;
  assign n11551 = n430 & n11550 ;
  assign n11552 = n267 & ~n1510 ;
  assign n11553 = n11551 & n11552 ;
  assign n11554 = ~n3137 & n4928 ;
  assign n11555 = n11553 & n11554 ;
  assign n11556 = x226 & n3765 ;
  assign n11557 = ~x226 & n11556 ;
  assign n11558 = n816 & n1511 ;
  assign n11559 = ~n1511 & n11558 ;
  assign n11560 = n11557 | n11559 ;
  assign n11561 = n11555 & ~n11560 ;
  assign n11562 = n11549 | n11561 ;
  assign n11563 = n11562 ^ n3284 ^ 1'b0 ;
  assign n11564 = n1832 & n9097 ;
  assign n11565 = ~n11105 & n11564 ;
  assign n11566 = n11565 ^ n4625 ^ 1'b0 ;
  assign n11567 = n5645 ^ n3088 ^ 1'b0 ;
  assign n11568 = n6425 | n11567 ;
  assign n11569 = ~n1499 & n4716 ;
  assign n11570 = ~n3065 & n11569 ;
  assign n11571 = n11570 ^ n2212 ^ 1'b0 ;
  assign n11572 = n2835 | n10833 ;
  assign n11573 = n2219 & n11572 ;
  assign n11574 = n1245 & ~n7413 ;
  assign n11575 = ~n3420 & n10514 ;
  assign n11576 = n11575 ^ n11219 ^ 1'b0 ;
  assign n11577 = n438 ^ x76 ^ 1'b0 ;
  assign n11578 = x19 & n415 ;
  assign n11579 = n5074 & ~n11578 ;
  assign n11580 = n10553 & n11579 ;
  assign n11581 = n1334 | n1799 ;
  assign n11582 = n11581 ^ n2527 ^ 1'b0 ;
  assign n11583 = ~n5077 & n11582 ;
  assign n11584 = n11583 ^ n446 ^ 1'b0 ;
  assign n11585 = n7723 & ~n11584 ;
  assign n11586 = n11585 ^ n6523 ^ 1'b0 ;
  assign n11587 = ~n1380 & n1666 ;
  assign n11588 = n11587 ^ n2122 ^ 1'b0 ;
  assign n11589 = x165 & n11588 ;
  assign n11590 = ~n5290 & n7345 ;
  assign n11591 = n11590 ^ n616 ^ 1'b0 ;
  assign n11592 = x190 & ~n6900 ;
  assign n11593 = ~n1817 & n11592 ;
  assign n11594 = n11591 & n11593 ;
  assign n11595 = ~n11589 & n11594 ;
  assign n11596 = n7898 ^ n7189 ^ 1'b0 ;
  assign n11597 = n9208 ^ n1566 ^ 1'b0 ;
  assign n11598 = n9361 & ~n11597 ;
  assign n11599 = n11598 ^ n10183 ^ 1'b0 ;
  assign n11600 = x193 & n8672 ;
  assign n11601 = ~n8672 & n11600 ;
  assign n11602 = n5613 & ~n11601 ;
  assign n11603 = n3437 & ~n11602 ;
  assign n11604 = n11603 ^ n2982 ^ 1'b0 ;
  assign n11606 = n2627 & ~n4143 ;
  assign n11607 = n11606 ^ n552 ^ 1'b0 ;
  assign n11605 = ~n1693 & n2082 ;
  assign n11608 = n11607 ^ n11605 ^ 1'b0 ;
  assign n11609 = ~n6032 & n11608 ;
  assign n11610 = n11609 ^ n4284 ^ 1'b0 ;
  assign n11612 = ~n4545 & n8654 ;
  assign n11611 = n3476 ^ n1751 ^ 1'b0 ;
  assign n11613 = n11612 ^ n11611 ^ 1'b0 ;
  assign n11614 = ~n5110 & n8773 ;
  assign n11615 = ~n4370 & n7964 ;
  assign n11618 = ~n1663 & n2345 ;
  assign n11616 = n987 ^ x129 ^ 1'b0 ;
  assign n11617 = n4456 & ~n11616 ;
  assign n11619 = n11618 ^ n11617 ^ 1'b0 ;
  assign n11620 = n6335 | n11619 ;
  assign n11621 = n8897 | n11620 ;
  assign n11622 = x222 & n11338 ;
  assign n11623 = n9261 & n11622 ;
  assign n11624 = n5646 ^ n647 ^ 1'b0 ;
  assign n11625 = ~n363 & n11624 ;
  assign n11626 = n11625 ^ n10236 ^ 1'b0 ;
  assign n11627 = n11154 ^ n4251 ^ 1'b0 ;
  assign n11628 = n3866 & ~n3970 ;
  assign n11629 = n671 | n11628 ;
  assign n11630 = n4783 | n11629 ;
  assign n11631 = ~n7688 & n11630 ;
  assign n11632 = n11631 ^ n1368 ^ 1'b0 ;
  assign n11633 = n1675 & n4917 ;
  assign n11634 = n11633 ^ n1817 ^ 1'b0 ;
  assign n11635 = ~n4595 & n11634 ;
  assign n11636 = n956 | n11635 ;
  assign n11639 = n987 & n1809 ;
  assign n11640 = ~n302 & n11639 ;
  assign n11637 = n4147 ^ n533 ^ 1'b0 ;
  assign n11638 = ( n10222 & n11246 ) | ( n10222 & n11637 ) | ( n11246 & n11637 ) ;
  assign n11641 = n11640 ^ n11638 ^ 1'b0 ;
  assign n11642 = n3776 & n11641 ;
  assign n11645 = n2105 & ~n6536 ;
  assign n11646 = n11645 ^ n1556 ^ 1'b0 ;
  assign n11647 = n2340 | n11646 ;
  assign n11644 = ~n1626 & n8192 ;
  assign n11648 = n11647 ^ n11644 ^ 1'b0 ;
  assign n11643 = n3833 & n10731 ;
  assign n11649 = n11648 ^ n11643 ^ 1'b0 ;
  assign n11650 = ~n512 & n8395 ;
  assign n11651 = n11650 ^ n5308 ^ 1'b0 ;
  assign n11652 = n1297 & n2725 ;
  assign n11653 = n11652 ^ n3399 ^ 1'b0 ;
  assign n11654 = n4298 & ~n11653 ;
  assign n11655 = n575 & ~n11654 ;
  assign n11656 = ~n6313 & n11655 ;
  assign n11657 = n1202 | n6200 ;
  assign n11658 = n10709 & ~n11657 ;
  assign n11659 = ~n6513 & n9749 ;
  assign n11660 = n7593 & n11140 ;
  assign n11661 = ~n1666 & n11660 ;
  assign n11662 = n5495 ^ n1050 ^ 1'b0 ;
  assign n11663 = n1324 & ~n11662 ;
  assign n11664 = n987 & ~n11663 ;
  assign n11665 = ~n987 & n11664 ;
  assign n11666 = n5971 & ~n11665 ;
  assign n11667 = n3454 & n7524 ;
  assign n11668 = n11667 ^ n4530 ^ 1'b0 ;
  assign n11669 = n10891 & ~n11668 ;
  assign n11670 = n8478 & n11669 ;
  assign n11671 = n11670 ^ n10181 ^ 1'b0 ;
  assign n11672 = n11666 & ~n11671 ;
  assign n11673 = n5489 ^ n749 ^ 1'b0 ;
  assign n11674 = n11673 ^ n2055 ^ 1'b0 ;
  assign n11675 = ~n589 & n11674 ;
  assign n11676 = n6205 ^ n3336 ^ 1'b0 ;
  assign n11677 = n3140 & n11676 ;
  assign n11678 = ~n11675 & n11677 ;
  assign n11679 = n6468 ^ x64 ^ 1'b0 ;
  assign n11680 = ~n7398 & n11679 ;
  assign n11681 = n5343 & ~n6102 ;
  assign n11682 = x112 & n11681 ;
  assign n11683 = n5923 ^ n4438 ^ 1'b0 ;
  assign n11684 = n2698 & ~n7098 ;
  assign n11685 = n11684 ^ n894 ^ 1'b0 ;
  assign n11686 = n4173 | n11685 ;
  assign n11687 = n11683 & ~n11686 ;
  assign n11688 = ~n1271 & n11242 ;
  assign n11689 = ~n858 & n7693 ;
  assign n11690 = n11689 ^ n4051 ^ 1'b0 ;
  assign n11691 = n11688 | n11690 ;
  assign n11692 = n11691 ^ n6493 ^ 1'b0 ;
  assign n11693 = n11692 ^ n456 ^ 1'b0 ;
  assign n11694 = n6151 & ~n11693 ;
  assign n11695 = x3 & n5665 ;
  assign n11696 = n4331 & n11695 ;
  assign n11697 = n7434 | n8225 ;
  assign n11698 = n9749 ^ n4325 ^ 1'b0 ;
  assign n11699 = ~n2926 & n11698 ;
  assign n11700 = n11699 ^ x182 ^ 1'b0 ;
  assign n11701 = x91 & n11700 ;
  assign n11702 = n1638 | n9254 ;
  assign n11703 = n1380 & n2370 ;
  assign n11704 = n1920 & n11703 ;
  assign n11705 = n1883 | n4258 ;
  assign n11706 = n3694 ^ n3349 ^ 1'b0 ;
  assign n11707 = n11705 & n11706 ;
  assign n11708 = n323 & ~n4685 ;
  assign n11709 = n3698 & n11708 ;
  assign n11710 = n1421 & n11709 ;
  assign n11711 = n3195 ^ n3018 ^ 1'b0 ;
  assign n11712 = n11224 ^ n1834 ^ 1'b0 ;
  assign n11713 = n10232 ^ n5531 ^ 1'b0 ;
  assign n11714 = n8747 | n11713 ;
  assign n11715 = n9092 | n10189 ;
  assign n11716 = n5435 | n11715 ;
  assign n11717 = n6021 ^ n4720 ^ 1'b0 ;
  assign n11718 = ~n6483 & n11717 ;
  assign n11719 = ( n1128 & n3358 ) | ( n1128 & n11718 ) | ( n3358 & n11718 ) ;
  assign n11720 = n10140 & ~n11719 ;
  assign n11721 = ~n4536 & n5902 ;
  assign n11722 = n11721 ^ n3759 ^ 1'b0 ;
  assign n11723 = n1324 | n11722 ;
  assign n11724 = n11057 ^ n1421 ^ 1'b0 ;
  assign n11725 = n11724 ^ x88 ^ 1'b0 ;
  assign n11726 = ~n5729 & n11725 ;
  assign n11727 = n11726 ^ n4179 ^ 1'b0 ;
  assign n11728 = n10233 ^ n4222 ^ 1'b0 ;
  assign n11729 = ~n7828 & n11728 ;
  assign n11730 = n8108 & n11291 ;
  assign n11731 = n11730 ^ n2427 ^ 1'b0 ;
  assign n11732 = ~n8795 & n11731 ;
  assign n11733 = n11732 ^ n10122 ^ 1'b0 ;
  assign n11734 = n4656 ^ n3918 ^ 1'b0 ;
  assign n11735 = n1360 & ~n2661 ;
  assign n11736 = n11735 ^ n876 ^ 1'b0 ;
  assign n11737 = n11736 ^ n1111 ^ 1'b0 ;
  assign n11738 = n7761 | n11737 ;
  assign n11739 = x77 & ~n10854 ;
  assign n11740 = n11739 ^ n8232 ^ 1'b0 ;
  assign n11741 = n8762 ^ n1745 ^ 1'b0 ;
  assign n11742 = n2310 & ~n11741 ;
  assign n11743 = ~n1175 & n11742 ;
  assign n11744 = ~n1405 & n11102 ;
  assign n11745 = x206 & ~n7953 ;
  assign n11746 = n7431 ^ n3976 ^ 1'b0 ;
  assign n11747 = x127 & n442 ;
  assign n11748 = n7112 & ~n11747 ;
  assign n11749 = ~n4948 & n11748 ;
  assign n11750 = n4916 | n6123 ;
  assign n11751 = n7883 & ~n11750 ;
  assign n11752 = n7359 | n11751 ;
  assign n11753 = n1701 & ~n8706 ;
  assign n11754 = n11753 ^ n3711 ^ 1'b0 ;
  assign n11755 = n9019 ^ n5754 ^ 1'b0 ;
  assign n11756 = n8234 & ~n11755 ;
  assign n11757 = n10823 ^ n5215 ^ 1'b0 ;
  assign n11758 = x130 & ~n10345 ;
  assign n11759 = ~n4575 & n10017 ;
  assign n11760 = n11759 ^ n5765 ^ 1'b0 ;
  assign n11761 = n7256 ^ n1981 ^ 1'b0 ;
  assign n11762 = n11761 ^ x89 ^ 1'b0 ;
  assign n11763 = n1826 & n11762 ;
  assign n11764 = n9611 ^ n6969 ^ 1'b0 ;
  assign n11765 = n3431 & ~n11764 ;
  assign n11766 = n11765 ^ n1489 ^ 1'b0 ;
  assign n11767 = ~n8522 & n11483 ;
  assign n11768 = n11767 ^ n2466 ^ 1'b0 ;
  assign n11769 = n1938 & ~n11768 ;
  assign n11770 = ~n5799 & n11769 ;
  assign n11771 = n5728 ^ n734 ^ 1'b0 ;
  assign n11772 = n10344 ^ n4598 ^ 1'b0 ;
  assign n11773 = n3179 & n11772 ;
  assign n11774 = ~n2819 & n4400 ;
  assign n11775 = n7894 ^ n4213 ^ 1'b0 ;
  assign n11776 = n5277 | n7703 ;
  assign n11777 = n7591 & n11776 ;
  assign n11778 = n3850 | n4133 ;
  assign n11779 = n3765 & ~n5138 ;
  assign n11780 = ( ~n3480 & n3585 ) | ( ~n3480 & n9946 ) | ( n3585 & n9946 ) ;
  assign n11783 = n4039 & n4104 ;
  assign n11781 = n969 & ~n2890 ;
  assign n11782 = n11781 ^ n1071 ^ 1'b0 ;
  assign n11784 = n11783 ^ n11782 ^ 1'b0 ;
  assign n11785 = n1855 | n11784 ;
  assign n11786 = n4551 ^ n2757 ^ 1'b0 ;
  assign n11787 = n1501 & ~n11786 ;
  assign n11788 = x20 & ~n7133 ;
  assign n11789 = ~n8137 & n11788 ;
  assign n11790 = n11749 ^ n5323 ^ 1'b0 ;
  assign n11791 = n7444 ^ n2853 ^ 1'b0 ;
  assign n11792 = n5394 | n11791 ;
  assign n11793 = n11792 ^ x143 ^ 1'b0 ;
  assign n11794 = x197 & ~n4349 ;
  assign n11795 = n8256 ^ n7630 ^ 1'b0 ;
  assign n11796 = n11794 | n11795 ;
  assign n11797 = n3726 | n6039 ;
  assign n11798 = n5466 & n11797 ;
  assign n11799 = n11798 ^ n10824 ^ 1'b0 ;
  assign n11800 = n3842 & ~n11799 ;
  assign n11801 = n5563 | n6194 ;
  assign n11802 = x151 & ~n11801 ;
  assign n11803 = n1513 ^ n641 ^ 1'b0 ;
  assign n11804 = n10189 & ~n11803 ;
  assign n11805 = n3591 & ~n6475 ;
  assign n11806 = ~n10965 & n11805 ;
  assign n11807 = n11806 ^ n8017 ^ 1'b0 ;
  assign n11808 = n3507 & ~n11807 ;
  assign n11809 = n2188 & ~n5865 ;
  assign n11810 = ~n8710 & n11809 ;
  assign n11811 = n2693 & ~n6061 ;
  assign n11812 = n11811 ^ n3711 ^ 1'b0 ;
  assign n11816 = n4272 ^ n1195 ^ 1'b0 ;
  assign n11814 = n418 | n3191 ;
  assign n11813 = n2464 & ~n10840 ;
  assign n11815 = n11814 ^ n11813 ^ 1'b0 ;
  assign n11817 = n11816 ^ n11815 ^ 1'b0 ;
  assign n11818 = n5604 ^ n4096 ^ 1'b0 ;
  assign n11819 = n7732 ^ n1544 ^ 1'b0 ;
  assign n11820 = n10048 ^ n1506 ^ 1'b0 ;
  assign n11821 = n10721 & ~n11820 ;
  assign n11822 = n703 & n987 ;
  assign n11823 = ~n987 & n11822 ;
  assign n11824 = ~n672 & n11823 ;
  assign n11825 = n1201 & n2639 ;
  assign n11826 = ~n1201 & n11825 ;
  assign n11827 = n11824 & ~n11826 ;
  assign n11833 = n420 & ~n770 ;
  assign n11834 = ~n420 & n11833 ;
  assign n11835 = x145 & ~n3258 ;
  assign n11836 = n11834 & n11835 ;
  assign n11837 = ~n2493 & n3097 ;
  assign n11838 = ~n3097 & n11837 ;
  assign n11839 = n5791 | n11838 ;
  assign n11840 = n11836 & ~n11839 ;
  assign n11841 = ~n5681 & n11840 ;
  assign n11828 = n1525 & n3040 ;
  assign n11829 = n11828 ^ n824 ^ 1'b0 ;
  assign n11830 = n583 & n11829 ;
  assign n11831 = ~n583 & n11830 ;
  assign n11832 = n6162 & ~n11831 ;
  assign n11842 = n11841 ^ n11832 ^ 1'b0 ;
  assign n11843 = n11827 & n11842 ;
  assign n11844 = n3709 ^ n787 ^ 1'b0 ;
  assign n11845 = n11843 | n11844 ;
  assign n11846 = n1230 ^ n1158 ^ 1'b0 ;
  assign n11847 = n504 | n11846 ;
  assign n11848 = n11847 ^ n10744 ^ 1'b0 ;
  assign n11849 = ~n4145 & n11848 ;
  assign n11850 = n4145 & n11849 ;
  assign n11851 = n1751 | n1994 ;
  assign n11852 = n11851 ^ n2685 ^ 1'b0 ;
  assign n11853 = ~n11850 & n11852 ;
  assign n11854 = n5838 & ~n11368 ;
  assign n11855 = n2190 | n10790 ;
  assign n11856 = n1512 & n1724 ;
  assign n11857 = n11856 ^ n9653 ^ 1'b0 ;
  assign n11858 = n11857 ^ n5122 ^ n3774 ;
  assign n11859 = n3217 & ~n11858 ;
  assign n11860 = n2420 ^ x30 ^ 1'b0 ;
  assign n11861 = n806 & ~n11860 ;
  assign n11862 = n11861 ^ n9266 ^ 1'b0 ;
  assign n11863 = n11862 ^ n8456 ^ 1'b0 ;
  assign n11864 = ~n623 & n11863 ;
  assign n11865 = n10395 ^ n1801 ^ 1'b0 ;
  assign n11866 = ~n6635 & n9898 ;
  assign n11867 = n6974 ^ n5137 ^ 1'b0 ;
  assign n11868 = ~n1857 & n11867 ;
  assign n11869 = n7542 ^ n3473 ^ 1'b0 ;
  assign n11870 = ( n11364 & ~n11868 ) | ( n11364 & n11869 ) | ( ~n11868 & n11869 ) ;
  assign n11871 = n5244 ^ n1688 ^ 1'b0 ;
  assign n11872 = n3102 & ~n11871 ;
  assign n11873 = n9530 & n11872 ;
  assign n11874 = n5758 & ~n11873 ;
  assign n11875 = n11873 & n11874 ;
  assign n11876 = x195 & ~n1677 ;
  assign n11877 = ~x195 & n11876 ;
  assign n11878 = x93 & ~n6592 ;
  assign n11879 = n6592 & n11878 ;
  assign n11880 = n2038 | n11879 ;
  assign n11881 = n2038 & ~n11880 ;
  assign n11882 = n11877 | n11881 ;
  assign n11883 = n11875 & ~n11882 ;
  assign n11884 = n3145 ^ x183 ^ 1'b0 ;
  assign n11885 = n6993 & n11214 ;
  assign n11886 = n2254 & ~n7555 ;
  assign n11887 = n11886 ^ n6985 ^ 1'b0 ;
  assign n11888 = n373 & n968 ;
  assign n11889 = n2768 & ~n6156 ;
  assign n11890 = n11889 ^ n6698 ^ 1'b0 ;
  assign n11891 = n6566 ^ n2039 ^ n1614 ;
  assign n11892 = n11891 ^ n2809 ^ 1'b0 ;
  assign n11893 = n9363 & ~n11892 ;
  assign n11894 = n9584 ^ n9301 ^ 1'b0 ;
  assign n11895 = x250 | n2302 ;
  assign n11896 = ~n8748 & n11895 ;
  assign n11897 = n11896 ^ n11331 ^ 1'b0 ;
  assign n11898 = n4409 ^ n3924 ^ 1'b0 ;
  assign n11899 = n4500 & n4804 ;
  assign n11900 = n5357 | n11899 ;
  assign n11901 = n11900 ^ n8902 ^ 1'b0 ;
  assign n11902 = ~n11898 & n11901 ;
  assign n11903 = n10077 ^ n10037 ^ 1'b0 ;
  assign n11904 = ( ~n830 & n946 ) | ( ~n830 & n3549 ) | ( n946 & n3549 ) ;
  assign n11905 = n11904 ^ n11584 ^ 1'b0 ;
  assign n11906 = ~n4846 & n11905 ;
  assign n11907 = n4502 & n11906 ;
  assign n11908 = n11907 ^ n7535 ^ 1'b0 ;
  assign n11909 = n4238 ^ n647 ^ 1'b0 ;
  assign n11910 = n5042 | n11909 ;
  assign n11911 = n9734 ^ n2417 ^ 1'b0 ;
  assign n11912 = n8874 ^ n3673 ^ 1'b0 ;
  assign n11913 = ~n5681 & n8627 ;
  assign n11914 = n11912 & n11913 ;
  assign n11916 = n509 ^ x128 ^ 1'b0 ;
  assign n11917 = n11916 ^ n8523 ^ 1'b0 ;
  assign n11918 = n4177 & ~n11917 ;
  assign n11915 = n6189 ^ x175 ^ 1'b0 ;
  assign n11919 = n11918 ^ n11915 ^ 1'b0 ;
  assign n11920 = ~x101 & n6524 ;
  assign n11921 = n1623 & n11434 ;
  assign n11922 = n11920 & n11921 ;
  assign n11923 = n508 & ~n11922 ;
  assign n11924 = n11923 ^ n9726 ^ 1'b0 ;
  assign n11925 = n1806 | n5768 ;
  assign n11926 = n11925 ^ n3670 ^ 1'b0 ;
  assign n11927 = ~n10546 & n11926 ;
  assign n11928 = ~n2380 & n5823 ;
  assign n11929 = n8495 & ~n11928 ;
  assign n11930 = n11929 ^ x77 ^ 1'b0 ;
  assign n11931 = x4 & n11930 ;
  assign n11932 = n2762 & n9068 ;
  assign n11933 = n3172 ^ n349 ^ 1'b0 ;
  assign n11934 = ~n11272 & n11933 ;
  assign n11935 = n10726 ^ n709 ^ 1'b0 ;
  assign n11936 = n1850 & ~n5279 ;
  assign n11937 = x25 & n11936 ;
  assign n11938 = n644 & ~n11937 ;
  assign n11939 = x68 & ~n2951 ;
  assign n11940 = n5293 & n11939 ;
  assign n11941 = n3546 | n6068 ;
  assign n11942 = n11941 ^ n11532 ^ 1'b0 ;
  assign n11943 = ~x67 & n6403 ;
  assign n11944 = n11943 ^ n2042 ^ 1'b0 ;
  assign n11947 = n7628 ^ n3430 ^ 1'b0 ;
  assign n11945 = n9068 ^ n5408 ^ n2536 ;
  assign n11946 = n5297 & n11945 ;
  assign n11948 = n11947 ^ n11946 ^ 1'b0 ;
  assign n11949 = n11348 ^ n1073 ^ 1'b0 ;
  assign n11950 = n747 & ~n2887 ;
  assign n11951 = x24 | n7030 ;
  assign n11952 = n1252 ^ n618 ^ 1'b0 ;
  assign n11953 = n7839 ^ n3740 ^ 1'b0 ;
  assign n11954 = n11953 ^ n11284 ^ n2693 ;
  assign n11955 = n8410 | n11954 ;
  assign n11956 = n4822 | n11955 ;
  assign n11957 = n1634 ^ n1117 ^ 1'b0 ;
  assign n11958 = n11956 & ~n11957 ;
  assign n11959 = n5819 & ~n8111 ;
  assign n11960 = n8677 & n11959 ;
  assign n11961 = n1826 ^ n1381 ^ 1'b0 ;
  assign n11962 = n7194 ^ n5443 ^ 1'b0 ;
  assign n11963 = n7637 & n11962 ;
  assign n11964 = ~n1016 & n3736 ;
  assign n11965 = n11964 ^ n7762 ^ 1'b0 ;
  assign n11966 = n1920 | n8514 ;
  assign n11967 = n11965 | n11966 ;
  assign n11968 = n3917 & ~n5489 ;
  assign n11969 = n1512 & ~n5327 ;
  assign n11970 = ~n1736 & n11969 ;
  assign n11971 = n10340 & ~n11970 ;
  assign n11972 = ~n946 & n2807 ;
  assign n11973 = n10778 & ~n11972 ;
  assign n11974 = n8258 & n10567 ;
  assign n11975 = n5350 ^ n3479 ^ 1'b0 ;
  assign n11976 = n3922 | n11975 ;
  assign n11977 = n4940 | n11976 ;
  assign n11978 = n1116 & ~n4189 ;
  assign n11979 = n5412 & n11978 ;
  assign n11980 = n855 & ~n8935 ;
  assign n11981 = n7204 & n11980 ;
  assign n11982 = n5417 ^ n2872 ^ 1'b0 ;
  assign n11983 = n4398 & ~n11982 ;
  assign n11984 = n3359 & n11983 ;
  assign n11985 = n11984 ^ n9972 ^ 1'b0 ;
  assign n11986 = n9706 ^ n8619 ^ 1'b0 ;
  assign n11987 = n8378 & ~n11986 ;
  assign n11988 = n5218 & ~n5714 ;
  assign n11989 = ~n5493 & n11988 ;
  assign n11990 = ~n361 & n6184 ;
  assign n11991 = n8367 ^ n2785 ^ 1'b0 ;
  assign n11992 = n7475 ^ n2478 ^ 1'b0 ;
  assign n11993 = n5310 | n5376 ;
  assign n11994 = n5376 & ~n11993 ;
  assign n11995 = n774 | n11994 ;
  assign n11996 = n11994 & ~n11995 ;
  assign n11997 = n3278 & ~n11996 ;
  assign n11998 = n11996 & n11997 ;
  assign n11999 = n4810 & ~n11469 ;
  assign n12000 = n11999 ^ n2921 ^ x81 ;
  assign n12001 = n4290 & n6663 ;
  assign n12002 = n9709 ^ n8513 ^ 1'b0 ;
  assign n12003 = n12002 ^ n2786 ^ 1'b0 ;
  assign n12004 = n12001 | n12003 ;
  assign n12005 = x38 & n880 ;
  assign n12006 = n12005 ^ n1961 ^ 1'b0 ;
  assign n12007 = n10267 ^ n2027 ^ 1'b0 ;
  assign n12008 = n12006 | n12007 ;
  assign n12009 = ( ~n2001 & n2039 ) | ( ~n2001 & n2289 ) | ( n2039 & n2289 ) ;
  assign n12010 = n1890 & ~n12009 ;
  assign n12011 = n12010 ^ n8025 ^ 1'b0 ;
  assign n12012 = ( n4589 & n8881 ) | ( n4589 & ~n12011 ) | ( n8881 & ~n12011 ) ;
  assign n12013 = n3872 ^ n1926 ^ 1'b0 ;
  assign n12014 = n12013 ^ n803 ^ 1'b0 ;
  assign n12015 = n5643 | n9992 ;
  assign n12016 = n4099 | n6165 ;
  assign n12017 = n3154 & ~n12016 ;
  assign n12018 = ~n1028 & n12017 ;
  assign n12019 = n11714 ^ n9503 ^ 1'b0 ;
  assign n12020 = n6477 & n7838 ;
  assign n12021 = n3569 & ~n3635 ;
  assign n12022 = ( n6119 & ~n12020 ) | ( n6119 & n12021 ) | ( ~n12020 & n12021 ) ;
  assign n12023 = n1537 | n11042 ;
  assign n12024 = ~n598 & n10168 ;
  assign n12025 = n7410 & ~n8182 ;
  assign n12026 = n11964 ^ n2970 ^ n1810 ;
  assign n12027 = n7177 & n9205 ;
  assign n12028 = n12027 ^ n4473 ^ 1'b0 ;
  assign n12029 = n1616 & n5494 ;
  assign n12030 = ~n2807 & n12029 ;
  assign n12031 = n12030 ^ n7573 ^ 1'b0 ;
  assign n12032 = n812 & n3043 ;
  assign n12034 = n2423 & ~n2785 ;
  assign n12035 = n12034 ^ n2328 ^ 1'b0 ;
  assign n12033 = x41 | n7713 ;
  assign n12036 = n12035 ^ n12033 ^ 1'b0 ;
  assign n12037 = ~n271 & n1252 ;
  assign n12038 = n1877 & n3933 ;
  assign n12039 = ~n12037 & n12038 ;
  assign n12040 = n12039 ^ n888 ^ 1'b0 ;
  assign n12041 = ~n557 & n666 ;
  assign n12042 = ~n691 & n3995 ;
  assign n12043 = ~n8002 & n12042 ;
  assign n12044 = n12043 ^ n8142 ^ 1'b0 ;
  assign n12045 = n521 ^ x190 ^ 1'b0 ;
  assign n12046 = x250 | n8588 ;
  assign n12047 = n3437 ^ n1245 ^ 1'b0 ;
  assign n12048 = n6328 | n12047 ;
  assign n12049 = n1311 & n12048 ;
  assign n12050 = ~n3784 & n6999 ;
  assign n12051 = n12050 ^ n5203 ^ 1'b0 ;
  assign n12052 = n12049 | n12051 ;
  assign n12053 = x242 & ~n6421 ;
  assign n12054 = n12053 ^ n2741 ^ 1'b0 ;
  assign n12055 = n9061 & n9861 ;
  assign n12056 = n7476 ^ x44 ^ 1'b0 ;
  assign n12057 = n6057 ^ n1694 ^ 1'b0 ;
  assign n12058 = ~n4967 & n12057 ;
  assign n12059 = n10379 ^ n849 ^ 1'b0 ;
  assign n12060 = n1385 & ~n12059 ;
  assign n12061 = n12060 ^ n3509 ^ 1'b0 ;
  assign n12062 = n3740 & ~n5162 ;
  assign n12063 = n1415 & n1762 ;
  assign n12064 = n12063 ^ n2948 ^ 1'b0 ;
  assign n12065 = ( n6881 & n11358 ) | ( n6881 & ~n12064 ) | ( n11358 & ~n12064 ) ;
  assign n12066 = ~n5880 & n9117 ;
  assign n12067 = n1295 & n7255 ;
  assign n12068 = ~n3249 & n9130 ;
  assign n12069 = n4002 & n12068 ;
  assign n12070 = ( n2095 & ~n2582 ) | ( n2095 & n2982 ) | ( ~n2582 & n2982 ) ;
  assign n12071 = n12070 ^ n9551 ^ 1'b0 ;
  assign n12072 = n2452 ^ n587 ^ 1'b0 ;
  assign n12073 = n8198 ^ n5862 ^ 1'b0 ;
  assign n12074 = n12072 | n12073 ;
  assign n12075 = n6502 ^ n5114 ^ 1'b0 ;
  assign n12076 = n10937 ^ n7397 ^ 1'b0 ;
  assign n12077 = ~n11567 & n12076 ;
  assign n12078 = ~n1239 & n12077 ;
  assign n12079 = n12078 ^ n1514 ^ 1'b0 ;
  assign n12080 = ~n988 & n12079 ;
  assign n12081 = n3404 | n5268 ;
  assign n12082 = ( x153 & x235 ) | ( x153 & ~n2901 ) | ( x235 & ~n2901 ) ;
  assign n12083 = x158 & n2186 ;
  assign n12084 = n12083 ^ n1160 ^ 1'b0 ;
  assign n12085 = n6246 ^ n3171 ^ 1'b0 ;
  assign n12086 = n12084 & n12085 ;
  assign n12087 = n5675 & ~n6637 ;
  assign n12088 = n12087 ^ n3324 ^ 1'b0 ;
  assign n12089 = n1853 & n3585 ;
  assign n12090 = n2475 & ~n12089 ;
  assign n12091 = n12089 & n12090 ;
  assign n12092 = n6162 ^ n3383 ^ 1'b0 ;
  assign n12093 = n2633 & n12092 ;
  assign n12094 = ~n5444 & n12093 ;
  assign n12104 = x105 & ~n331 ;
  assign n12105 = ~x105 & n12104 ;
  assign n12106 = x57 & n700 ;
  assign n12107 = n12105 & n12106 ;
  assign n12108 = n715 | n12107 ;
  assign n12109 = n12107 & ~n12108 ;
  assign n12110 = n1819 & ~n12109 ;
  assign n12111 = ~n1819 & n12110 ;
  assign n12112 = n1449 | n12111 ;
  assign n12113 = n1449 & ~n12112 ;
  assign n12095 = n8584 & n9799 ;
  assign n12096 = n1497 | n1658 ;
  assign n12097 = n1497 & ~n12096 ;
  assign n12098 = n2660 | n12097 ;
  assign n12099 = n2660 & ~n12098 ;
  assign n12100 = n4647 | n12099 ;
  assign n12101 = n4647 & ~n12100 ;
  assign n12102 = ~n10647 & n12101 ;
  assign n12103 = n12095 & n12102 ;
  assign n12114 = n12113 ^ n12103 ^ 1'b0 ;
  assign n12115 = n4943 & n5639 ;
  assign n12116 = n11702 ^ x190 ^ 1'b0 ;
  assign n12117 = n12116 ^ n7401 ^ 1'b0 ;
  assign n12118 = n5041 & n12117 ;
  assign n12119 = n7605 & ~n11284 ;
  assign n12120 = ~n10885 & n12119 ;
  assign n12121 = ~n1435 & n1802 ;
  assign n12122 = n12121 ^ n3511 ^ 1'b0 ;
  assign n12123 = n12087 | n12122 ;
  assign n12124 = n10888 ^ n392 ^ 1'b0 ;
  assign n12125 = n3635 | n4758 ;
  assign n12126 = n12125 ^ n7448 ^ 1'b0 ;
  assign n12127 = n1395 | n12126 ;
  assign n12128 = n8725 & ~n12127 ;
  assign n12129 = n12128 ^ n5191 ^ 1'b0 ;
  assign n12130 = n11065 & n12129 ;
  assign n12131 = n1783 & ~n5442 ;
  assign n12132 = n12131 ^ x222 ^ x31 ;
  assign n12133 = n1977 & n5266 ;
  assign n12134 = n12133 ^ n3859 ^ 1'b0 ;
  assign n12135 = ~n594 & n12134 ;
  assign n12136 = n1681 & n12135 ;
  assign n12137 = ~n3480 & n12136 ;
  assign n12138 = n9299 ^ n4734 ^ n1139 ;
  assign n12140 = n708 & n9723 ;
  assign n12139 = ~n5681 & n11154 ;
  assign n12141 = n12140 ^ n12139 ^ 1'b0 ;
  assign n12142 = n2786 & n7320 ;
  assign n12143 = n1795 & ~n12142 ;
  assign n12144 = n12143 ^ n3441 ^ 1'b0 ;
  assign n12145 = n5265 ^ n3210 ^ 1'b0 ;
  assign n12146 = n12145 ^ n1056 ^ 1'b0 ;
  assign n12147 = n7444 & n12146 ;
  assign n12148 = n12147 ^ n11725 ^ 1'b0 ;
  assign n12149 = n5070 | n8322 ;
  assign n12150 = x169 & n1605 ;
  assign n12151 = ~n1643 & n12150 ;
  assign n12152 = n1513 & n4617 ;
  assign n12153 = n1146 | n2946 ;
  assign n12154 = n12153 ^ n5207 ^ 1'b0 ;
  assign n12155 = n1137 & n12154 ;
  assign n12156 = n3419 & n4077 ;
  assign n12157 = n2432 & n12156 ;
  assign n12158 = n1365 ^ n911 ^ 1'b0 ;
  assign n12159 = n7507 | n12158 ;
  assign n12160 = n9713 | n12159 ;
  assign n12161 = n12160 ^ n786 ^ 1'b0 ;
  assign n12162 = ~n12157 & n12161 ;
  assign n12163 = n8351 & n11803 ;
  assign n12164 = n11949 & ~n12163 ;
  assign n12165 = n2006 ^ n705 ^ 1'b0 ;
  assign n12166 = n4931 ^ n4529 ^ 1'b0 ;
  assign n12167 = n12165 | n12166 ;
  assign n12168 = x100 & n1905 ;
  assign n12169 = n8328 & n12168 ;
  assign n12170 = n1339 | n7034 ;
  assign n12171 = n12170 ^ n1701 ^ 1'b0 ;
  assign n12172 = ~n1059 & n12171 ;
  assign n12173 = n10893 & n12172 ;
  assign n12174 = n9379 ^ n2017 ^ 1'b0 ;
  assign n12175 = n3181 ^ n1324 ^ 1'b0 ;
  assign n12176 = n8241 | n12175 ;
  assign n12177 = n3361 & ~n12176 ;
  assign n12178 = n3820 & n11048 ;
  assign n12179 = ~n10496 & n11377 ;
  assign n12180 = n12179 ^ n5081 ^ 1'b0 ;
  assign n12181 = n3558 | n8816 ;
  assign n12182 = n8165 | n12181 ;
  assign n12187 = n10932 ^ n2824 ^ 1'b0 ;
  assign n12188 = n7986 | n9363 ;
  assign n12189 = n12187 & ~n12188 ;
  assign n12183 = n655 & n5624 ;
  assign n12184 = n12183 ^ n932 ^ 1'b0 ;
  assign n12185 = n1441 & n2784 ;
  assign n12186 = ~n12184 & n12185 ;
  assign n12190 = n12189 ^ n12186 ^ 1'b0 ;
  assign n12191 = n11649 ^ n8287 ^ 1'b0 ;
  assign n12192 = n3616 & ~n12191 ;
  assign n12193 = ~n713 & n1909 ;
  assign n12194 = n1271 | n12193 ;
  assign n12195 = n376 | n5256 ;
  assign n12196 = n12195 ^ n6540 ^ 1'b0 ;
  assign n12197 = x245 & ~n2230 ;
  assign n12198 = ~n5510 & n12197 ;
  assign n12199 = ~n754 & n12198 ;
  assign n12200 = n5286 & ~n6900 ;
  assign n12201 = n3049 & n12200 ;
  assign n12202 = ~n8722 & n12201 ;
  assign n12203 = n12202 ^ n6960 ^ 1'b0 ;
  assign n12204 = n8638 & n12203 ;
  assign n12205 = n11524 ^ n5307 ^ 1'b0 ;
  assign n12206 = n11488 ^ n10166 ^ 1'b0 ;
  assign n12207 = n1216 | n10692 ;
  assign n12208 = n8715 | n12207 ;
  assign n12209 = n709 | n1126 ;
  assign n12210 = n12209 ^ n6466 ^ 1'b0 ;
  assign n12211 = n10488 ^ n10064 ^ 1'b0 ;
  assign n12212 = ~n4661 & n4959 ;
  assign n12213 = n10840 & n12212 ;
  assign n12214 = n1233 & ~n11870 ;
  assign n12215 = n10374 ^ n9530 ^ n7667 ;
  assign n12216 = ~n5069 & n12215 ;
  assign n12217 = ~n9162 & n10950 ;
  assign n12218 = n12217 ^ n5748 ^ 1'b0 ;
  assign n12219 = n12218 ^ n492 ^ 1'b0 ;
  assign n12220 = n2671 & ~n12219 ;
  assign n12221 = n1208 & ~n2564 ;
  assign n12222 = n12220 & ~n12221 ;
  assign n12223 = ~n4338 & n12222 ;
  assign n12224 = n12223 ^ n9205 ^ 1'b0 ;
  assign n12225 = n4233 & n12224 ;
  assign n12226 = n12225 ^ n6311 ^ 1'b0 ;
  assign n12227 = n12216 | n12226 ;
  assign n12235 = n5913 ^ n5076 ^ 1'b0 ;
  assign n12236 = n12235 ^ n4493 ^ 1'b0 ;
  assign n12228 = n3143 ^ x253 ^ x250 ;
  assign n12229 = n476 | n2581 ;
  assign n12230 = n12229 ^ n1972 ^ 1'b0 ;
  assign n12231 = x55 & n12230 ;
  assign n12232 = n12231 ^ n5700 ^ 1'b0 ;
  assign n12233 = ( n3221 & n12228 ) | ( n3221 & ~n12232 ) | ( n12228 & ~n12232 ) ;
  assign n12234 = n10708 | n12233 ;
  assign n12237 = n12236 ^ n12234 ^ 1'b0 ;
  assign n12238 = n9461 ^ n4623 ^ 1'b0 ;
  assign n12239 = n4298 | n5996 ;
  assign n12240 = n784 | n814 ;
  assign n12241 = x240 | n12240 ;
  assign n12242 = n1632 | n1685 ;
  assign n12243 = n12241 | n12242 ;
  assign n12246 = n2102 ^ n2082 ^ 1'b0 ;
  assign n12247 = n1832 & ~n12246 ;
  assign n12244 = ~n3065 & n9707 ;
  assign n12245 = n292 & n12244 ;
  assign n12248 = n12247 ^ n12245 ^ 1'b0 ;
  assign n12249 = n11702 ^ n1955 ^ 1'b0 ;
  assign n12250 = ~n2042 & n5056 ;
  assign n12251 = n12250 ^ n5457 ^ 1'b0 ;
  assign n12252 = n3076 & ~n4327 ;
  assign n12253 = n6413 & ~n11382 ;
  assign n12254 = n1372 | n2021 ;
  assign n12255 = n12254 ^ n1028 ^ 1'b0 ;
  assign n12256 = n2672 | n12255 ;
  assign n12257 = n1909 | n9539 ;
  assign n12259 = ~x103 & n285 ;
  assign n12258 = n6326 & ~n9150 ;
  assign n12260 = n12259 ^ n12258 ^ 1'b0 ;
  assign n12261 = n12081 ^ n583 ^ 1'b0 ;
  assign n12262 = ~n2559 & n12261 ;
  assign n12263 = n827 | n6080 ;
  assign n12264 = n5190 & n12075 ;
  assign n12265 = n8617 & n12264 ;
  assign n12266 = n2042 ^ n729 ^ 1'b0 ;
  assign n12267 = n4775 ^ n4420 ^ 1'b0 ;
  assign n12268 = n12267 ^ n3899 ^ 1'b0 ;
  assign n12269 = n486 ^ x93 ^ 1'b0 ;
  assign n12270 = x74 & n2928 ;
  assign n12271 = n7179 ^ n4742 ^ 1'b0 ;
  assign n12272 = ~n7323 & n12271 ;
  assign n12275 = n313 | n2065 ;
  assign n12276 = n2065 & ~n12275 ;
  assign n12273 = n4203 | n4603 ;
  assign n12274 = n1082 | n12273 ;
  assign n12277 = n12276 ^ n12274 ^ 1'b0 ;
  assign n12280 = n610 & ~n1212 ;
  assign n12281 = n1212 & n12280 ;
  assign n12282 = n7093 | n12281 ;
  assign n12283 = n7093 & ~n12282 ;
  assign n12278 = n3940 & n10869 ;
  assign n12279 = n9566 & n12278 ;
  assign n12284 = n12283 ^ n12279 ^ 1'b0 ;
  assign n12285 = ~n12277 & n12284 ;
  assign n12286 = n3860 | n9624 ;
  assign n12287 = n3743 | n12286 ;
  assign n12288 = ~n7397 & n12287 ;
  assign n12290 = ~n1633 & n6614 ;
  assign n12291 = n12290 ^ n2953 ^ 1'b0 ;
  assign n12289 = n5824 & ~n7915 ;
  assign n12292 = n12291 ^ n12289 ^ 1'b0 ;
  assign n12293 = n5399 ^ n3823 ^ 1'b0 ;
  assign n12294 = n3687 & n10813 ;
  assign n12295 = n12294 ^ n929 ^ 1'b0 ;
  assign n12296 = n8014 ^ n5508 ^ 1'b0 ;
  assign n12297 = ~n6060 & n12296 ;
  assign n12298 = ~n4086 & n12297 ;
  assign n12299 = n1291 | n11072 ;
  assign n12300 = n6886 & ~n11662 ;
  assign n12301 = n12300 ^ n5667 ^ 1'b0 ;
  assign n12302 = n12165 ^ n3810 ^ 1'b0 ;
  assign n12303 = n610 & ~n8816 ;
  assign n12304 = n12303 ^ n6205 ^ 1'b0 ;
  assign n12305 = n8041 & ~n12304 ;
  assign n12306 = n2183 & n10348 ;
  assign n12307 = n1920 & n11608 ;
  assign n12308 = n583 & ~n7155 ;
  assign n12309 = n12308 ^ x201 ^ 1'b0 ;
  assign n12310 = n6703 & n9740 ;
  assign n12311 = ~x206 & n4875 ;
  assign n12312 = ~x253 & n305 ;
  assign n12313 = n12236 | n12312 ;
  assign n12314 = n1847 | n12313 ;
  assign n12315 = ~n8600 & n12314 ;
  assign n12316 = n12315 ^ n2129 ^ 1'b0 ;
  assign n12317 = n5357 ^ n535 ^ 1'b0 ;
  assign n12318 = n957 & ~n3683 ;
  assign n12319 = n3683 & n12318 ;
  assign n12320 = ~n2568 & n12319 ;
  assign n12321 = ~n10006 & n12320 ;
  assign n12322 = n11224 & n12321 ;
  assign n12323 = n2466 ^ x28 ^ 1'b0 ;
  assign n12324 = n4978 & ~n12323 ;
  assign n12325 = n4091 & n12324 ;
  assign n12326 = n12322 & n12325 ;
  assign n12327 = n6945 ^ n6437 ^ 1'b0 ;
  assign n12328 = n3569 | n11462 ;
  assign n12329 = n3879 | n12328 ;
  assign n12330 = n12329 ^ n3979 ^ 1'b0 ;
  assign n12331 = n8329 & ~n9606 ;
  assign n12332 = n5982 ^ n3294 ^ 1'b0 ;
  assign n12333 = n816 & ~n2591 ;
  assign n12334 = n12333 ^ n1490 ^ 1'b0 ;
  assign n12335 = n2782 & ~n9771 ;
  assign n12336 = n12334 & ~n12335 ;
  assign n12337 = n12163 & n12336 ;
  assign n12338 = n12307 & ~n12337 ;
  assign n12339 = n6597 ^ n3187 ^ 1'b0 ;
  assign n12340 = x12 & n12339 ;
  assign n12341 = n1459 & ~n2470 ;
  assign n12342 = n2384 & n12341 ;
  assign n12343 = n5932 | n12342 ;
  assign n12344 = n412 & n2518 ;
  assign n12345 = ~n10817 & n12344 ;
  assign n12346 = n3107 & ~n6087 ;
  assign n12349 = n9024 ^ x253 ^ 1'b0 ;
  assign n12350 = n1423 & n5381 ;
  assign n12351 = n12349 & n12350 ;
  assign n12347 = ( n1919 & n2689 ) | ( n1919 & n9875 ) | ( n2689 & n9875 ) ;
  assign n12348 = ~n432 & n12347 ;
  assign n12352 = n12351 ^ n12348 ^ 1'b0 ;
  assign n12353 = ~n2935 & n11259 ;
  assign n12354 = n12353 ^ n2636 ^ 1'b0 ;
  assign n12355 = n7266 | n12354 ;
  assign n12356 = ~n1974 & n2465 ;
  assign n12364 = ~n9737 & n12134 ;
  assign n12357 = n1333 | n6700 ;
  assign n12360 = n4892 ^ n3402 ^ 1'b0 ;
  assign n12358 = n10413 ^ n1596 ^ 1'b0 ;
  assign n12359 = n6205 & n12358 ;
  assign n12361 = n12360 ^ n12359 ^ 1'b0 ;
  assign n12362 = ~n8160 & n12361 ;
  assign n12363 = n12357 & n12362 ;
  assign n12365 = n12364 ^ n12363 ^ 1'b0 ;
  assign n12369 = n1938 | n5608 ;
  assign n12366 = n1693 | n7936 ;
  assign n12367 = n12366 ^ n6158 ^ 1'b0 ;
  assign n12368 = n9177 & ~n12367 ;
  assign n12370 = n12369 ^ n12368 ^ 1'b0 ;
  assign n12371 = ( n2423 & ~n4726 ) | ( n2423 & n6721 ) | ( ~n4726 & n6721 ) ;
  assign n12372 = n1152 ^ n267 ^ 1'b0 ;
  assign n12373 = n12371 & ~n12372 ;
  assign n12374 = n12373 ^ n7436 ^ 1'b0 ;
  assign n12375 = n5896 ^ n2650 ^ 1'b0 ;
  assign n12376 = n12375 ^ n6433 ^ 1'b0 ;
  assign n12377 = n9977 & ~n12376 ;
  assign n12378 = n2768 & ~n4389 ;
  assign n12379 = n7813 ^ n1684 ^ 1'b0 ;
  assign n12380 = n12378 & ~n12379 ;
  assign n12381 = ~n2495 & n4395 ;
  assign n12382 = n8095 | n9592 ;
  assign n12383 = n12382 ^ n1967 ^ 1'b0 ;
  assign n12384 = n4952 ^ n1449 ^ 1'b0 ;
  assign n12385 = n4513 & n12384 ;
  assign n12386 = ( n2765 & ~n3651 ) | ( n2765 & n12385 ) | ( ~n3651 & n12385 ) ;
  assign n12387 = n12386 ^ n11336 ^ 1'b0 ;
  assign n12388 = n2562 ^ n825 ^ 1'b0 ;
  assign n12389 = n5779 | n12388 ;
  assign n12390 = n12389 ^ n5942 ^ n5597 ;
  assign n12392 = n1985 & ~n5369 ;
  assign n12391 = n2433 & ~n10201 ;
  assign n12393 = n12392 ^ n12391 ^ 1'b0 ;
  assign n12394 = ( n4249 & n7988 ) | ( n4249 & n12165 ) | ( n7988 & n12165 ) ;
  assign n12395 = n7718 ^ n4985 ^ 1'b0 ;
  assign n12396 = n12395 ^ n11395 ^ n3880 ;
  assign n12397 = n1494 & n11869 ;
  assign n12398 = n12397 ^ n10261 ^ 1'b0 ;
  assign n12399 = n407 & n6516 ;
  assign n12400 = n12399 ^ n5205 ^ 1'b0 ;
  assign n12401 = n2450 & ~n5821 ;
  assign n12402 = n12401 ^ n2190 ^ 1'b0 ;
  assign n12403 = n11915 & ~n12402 ;
  assign n12404 = n12403 ^ n3366 ^ 1'b0 ;
  assign n12405 = n519 ^ n445 ^ 1'b0 ;
  assign n12406 = n9923 ^ n2486 ^ 1'b0 ;
  assign n12407 = n9041 & ~n12406 ;
  assign n12408 = n12405 & n12407 ;
  assign n12409 = n7535 ^ n5324 ^ 1'b0 ;
  assign n12410 = n12163 | n12409 ;
  assign n12412 = n1046 & n4040 ;
  assign n12413 = n12412 ^ n4022 ^ 1'b0 ;
  assign n12414 = n1508 & n12413 ;
  assign n12415 = n12414 ^ n6131 ^ 1'b0 ;
  assign n12416 = n1307 | n12415 ;
  assign n12411 = n4191 & ~n4815 ;
  assign n12417 = n12416 ^ n12411 ^ 1'b0 ;
  assign n12418 = ~n12410 & n12417 ;
  assign n12419 = n12418 ^ n5965 ^ 1'b0 ;
  assign n12420 = n6834 ^ n5498 ^ 1'b0 ;
  assign n12421 = ( n3458 & n7293 ) | ( n3458 & n12420 ) | ( n7293 & n12420 ) ;
  assign n12422 = n3592 ^ n2414 ^ 1'b0 ;
  assign n12423 = ~n8491 & n12422 ;
  assign n12424 = n2794 ^ x204 ^ 1'b0 ;
  assign n12425 = ~n901 & n12424 ;
  assign n12426 = ~n846 & n12425 ;
  assign n12427 = ~n12423 & n12426 ;
  assign n12428 = n1594 & ~n3043 ;
  assign n12429 = n12428 ^ n394 ^ 1'b0 ;
  assign n12430 = n4814 ^ n3127 ^ 1'b0 ;
  assign n12431 = ~n12429 & n12430 ;
  assign n12432 = n12431 ^ n2143 ^ 1'b0 ;
  assign n12433 = ~n631 & n12432 ;
  assign n12434 = ~n1204 & n12433 ;
  assign n12435 = n2716 & ~n12434 ;
  assign n12436 = n12427 & n12435 ;
  assign n12437 = ~n4366 & n7914 ;
  assign n12438 = n12437 ^ n6196 ^ 1'b0 ;
  assign n12439 = n1415 & n7421 ;
  assign n12440 = n548 & n12439 ;
  assign n12441 = n12440 ^ n430 ^ 1'b0 ;
  assign n12442 = x104 & n2408 ;
  assign n12443 = ~n12441 & n12442 ;
  assign n12444 = n12443 ^ n1976 ^ 1'b0 ;
  assign n12445 = n718 & n4129 ;
  assign n12446 = n4297 & ~n7594 ;
  assign n12447 = n12446 ^ n7757 ^ 1'b0 ;
  assign n12448 = n5073 ^ n5041 ^ 1'b0 ;
  assign n12449 = n7443 ^ x70 ^ 1'b0 ;
  assign n12450 = n11285 ^ n5665 ^ 1'b0 ;
  assign n12451 = ~n12449 & n12450 ;
  assign n12452 = ~n2065 & n12451 ;
  assign n12453 = n9460 ^ n2304 ^ 1'b0 ;
  assign n12454 = n747 | n12453 ;
  assign n12455 = n9755 & ~n12454 ;
  assign n12456 = n3020 | n5029 ;
  assign n12457 = n11608 ^ n2760 ^ 1'b0 ;
  assign n12458 = n733 | n12457 ;
  assign n12459 = n1156 | n9222 ;
  assign n12460 = n9354 & ~n12459 ;
  assign n12461 = ~n5287 & n5733 ;
  assign n12466 = n1658 & n11145 ;
  assign n12467 = n5928 & n12466 ;
  assign n12462 = n2099 | n3979 ;
  assign n12463 = n11668 & ~n12462 ;
  assign n12464 = n2887 ^ n2417 ^ 1'b0 ;
  assign n12465 = ~n12463 & n12464 ;
  assign n12468 = n12467 ^ n12465 ^ 1'b0 ;
  assign n12469 = n8216 ^ n7845 ^ 1'b0 ;
  assign n12470 = n6401 | n12469 ;
  assign n12471 = n1536 & ~n12470 ;
  assign n12472 = n7949 ^ n518 ^ 1'b0 ;
  assign n12473 = n2477 | n12472 ;
  assign n12474 = n2685 ^ x222 ^ 1'b0 ;
  assign n12475 = n6790 | n12474 ;
  assign n12476 = n2900 & n4959 ;
  assign n12477 = ~n3118 & n12476 ;
  assign n12478 = n4347 & ~n12477 ;
  assign n12479 = n5990 & n9299 ;
  assign n12490 = n931 | n934 ;
  assign n12491 = n12490 ^ n669 ^ 1'b0 ;
  assign n12480 = x48 & ~n877 ;
  assign n12481 = ~x48 & n12480 ;
  assign n12482 = x59 & ~n1407 ;
  assign n12483 = n1407 & n12482 ;
  assign n12484 = n2661 | n12483 ;
  assign n12485 = n12483 & ~n12484 ;
  assign n12486 = n12485 ^ n1302 ^ 1'b0 ;
  assign n12487 = n655 & n12486 ;
  assign n12488 = n12481 & n12487 ;
  assign n12489 = n12488 ^ n3484 ^ 1'b0 ;
  assign n12492 = n12491 ^ n12489 ^ n2704 ;
  assign n12493 = n766 | n11083 ;
  assign n12494 = n3842 | n12493 ;
  assign n12495 = n12494 ^ n6022 ^ 1'b0 ;
  assign n12496 = n1890 | n9244 ;
  assign n12497 = n3842 & ~n5201 ;
  assign n12498 = n12497 ^ n8512 ^ 1'b0 ;
  assign n12499 = ~n6125 & n10580 ;
  assign n12500 = n12499 ^ n10309 ^ 1'b0 ;
  assign n12501 = n3748 ^ n1438 ^ 1'b0 ;
  assign n12502 = ~n11392 & n12501 ;
  assign n12503 = n879 | n7427 ;
  assign n12504 = ~n7190 & n10763 ;
  assign n12505 = n12503 & ~n12504 ;
  assign n12506 = n1447 ^ n1251 ^ 1'b0 ;
  assign n12507 = n3143 & ~n5384 ;
  assign n12508 = ~n11938 & n12507 ;
  assign n12509 = x41 | n1117 ;
  assign n12510 = n6370 ^ n2803 ^ 1'b0 ;
  assign n12511 = ~n12509 & n12510 ;
  assign n12512 = n12511 ^ n6741 ^ 1'b0 ;
  assign n12516 = n8345 ^ n1293 ^ 1'b0 ;
  assign n12517 = n12516 ^ n5860 ^ 1'b0 ;
  assign n12518 = n3069 | n12517 ;
  assign n12513 = ~n2794 & n4602 ;
  assign n12514 = ~n812 & n12513 ;
  assign n12515 = n12514 ^ n4343 ^ 1'b0 ;
  assign n12519 = n12518 ^ n12515 ^ 1'b0 ;
  assign n12520 = n512 | n9375 ;
  assign n12521 = n3033 & n12028 ;
  assign n12522 = n10857 ^ n5870 ^ 1'b0 ;
  assign n12523 = n7855 ^ n7813 ^ 1'b0 ;
  assign n12524 = n2159 & n12523 ;
  assign n12525 = n9957 ^ n5000 ^ 1'b0 ;
  assign n12526 = n465 ^ x123 ^ 1'b0 ;
  assign n12527 = n956 ^ n514 ^ 1'b0 ;
  assign n12528 = n5275 ^ n1181 ^ 1'b0 ;
  assign n12529 = n1880 & n12528 ;
  assign n12530 = ~n9706 & n12529 ;
  assign n12531 = n12530 ^ n7126 ^ 1'b0 ;
  assign n12532 = n12531 ^ n5176 ^ 1'b0 ;
  assign n12533 = n12527 & n12532 ;
  assign n12534 = x235 & n1634 ;
  assign n12535 = n12534 ^ n2311 ^ 1'b0 ;
  assign n12536 = ~n535 & n12535 ;
  assign n12537 = n2955 & n8223 ;
  assign n12538 = n2812 & ~n4515 ;
  assign n12539 = n12537 & n12538 ;
  assign n12540 = n10488 ^ n1152 ^ 1'b0 ;
  assign n12541 = ~n2493 & n12540 ;
  assign n12542 = n3263 ^ n2179 ^ 1'b0 ;
  assign n12543 = n1202 & ~n12542 ;
  assign n12544 = n3918 & n12543 ;
  assign n12545 = ~n12543 & n12544 ;
  assign n12546 = n5007 ^ n1886 ^ 1'b0 ;
  assign n12547 = n3713 & ~n9716 ;
  assign n12548 = n12547 ^ n6897 ^ 1'b0 ;
  assign n12549 = ~n12546 & n12548 ;
  assign n12550 = n12545 & n12549 ;
  assign n12551 = ~n2746 & n5914 ;
  assign n12552 = ~n1404 & n12551 ;
  assign n12553 = n1893 & n12552 ;
  assign n12554 = n12553 ^ n461 ^ 1'b0 ;
  assign n12555 = n4928 & n5412 ;
  assign n12556 = ~n644 & n11046 ;
  assign n12559 = n611 | n4162 ;
  assign n12557 = n1219 | n3950 ;
  assign n12558 = n2860 & ~n12557 ;
  assign n12560 = n12559 ^ n12558 ^ 1'b0 ;
  assign n12561 = n11653 | n12560 ;
  assign n12562 = n4455 & ~n5324 ;
  assign n12563 = n8089 & n11451 ;
  assign n12564 = n6998 ^ n5379 ^ 1'b0 ;
  assign n12565 = ~n6350 & n12564 ;
  assign n12568 = n4350 | n7030 ;
  assign n12566 = n7712 & ~n7882 ;
  assign n12567 = n1511 & n12566 ;
  assign n12569 = n12568 ^ n12567 ^ 1'b0 ;
  assign n12570 = n3562 ^ n2013 ^ 1'b0 ;
  assign n12571 = n5658 | n7971 ;
  assign n12572 = n12571 ^ n1817 ^ 1'b0 ;
  assign n12573 = n12572 ^ n10295 ^ n285 ;
  assign n12574 = n12573 ^ n3071 ^ 1'b0 ;
  assign n12575 = n12227 ^ n2528 ^ 1'b0 ;
  assign n12576 = n6407 ^ n3809 ^ 1'b0 ;
  assign n12577 = n12576 ^ n3423 ^ 1'b0 ;
  assign n12578 = n6348 & ~n7828 ;
  assign n12579 = n1267 & n2223 ;
  assign n12580 = n271 & n4080 ;
  assign n12581 = n12580 ^ n3989 ^ 1'b0 ;
  assign n12582 = n5755 ^ n4658 ^ 1'b0 ;
  assign n12583 = n1546 | n10272 ;
  assign n12584 = n10605 & n12583 ;
  assign n12585 = n1646 & ~n5393 ;
  assign n12586 = n795 | n2769 ;
  assign n12587 = n12586 ^ n5784 ^ n1701 ;
  assign n12588 = n3611 & ~n12587 ;
  assign n12589 = n10875 ^ n903 ^ 1'b0 ;
  assign n12590 = n2925 & ~n12589 ;
  assign n12591 = n9446 ^ n1214 ^ 1'b0 ;
  assign n12592 = n9421 & n12591 ;
  assign n12593 = n5622 & n6741 ;
  assign n12594 = ~n1130 & n12593 ;
  assign n12595 = ( n8088 & ~n12592 ) | ( n8088 & n12594 ) | ( ~n12592 & n12594 ) ;
  assign n12596 = ~n12590 & n12595 ;
  assign n12597 = n2735 & ~n3097 ;
  assign n12598 = n12597 ^ x179 ^ 1'b0 ;
  assign n12599 = n4516 & ~n5759 ;
  assign n12600 = ~n6578 & n12599 ;
  assign n12603 = n7711 ^ x101 ^ 1'b0 ;
  assign n12604 = n6446 & n12603 ;
  assign n12601 = ~n2185 & n3337 ;
  assign n12602 = n5937 | n12601 ;
  assign n12605 = n12604 ^ n12602 ^ 1'b0 ;
  assign n12606 = ~n1948 & n12423 ;
  assign n12607 = n12606 ^ n6307 ^ 1'b0 ;
  assign n12608 = n12607 ^ n6254 ^ 1'b0 ;
  assign n12609 = n12608 ^ n11299 ^ 1'b0 ;
  assign n12610 = n8823 & n12609 ;
  assign n12611 = n8151 ^ x253 ^ 1'b0 ;
  assign n12612 = n2826 | n7756 ;
  assign n12613 = ~n6315 & n11125 ;
  assign n12614 = n2376 & n6881 ;
  assign n12615 = n6003 | n10553 ;
  assign n12616 = n4032 ^ n1085 ^ 1'b0 ;
  assign n12617 = n2689 | n12616 ;
  assign n12618 = ~x155 & n6022 ;
  assign n12619 = n3477 & n7668 ;
  assign n12620 = x244 & n12619 ;
  assign n12621 = n4709 & n12620 ;
  assign n12622 = x29 & ~n12621 ;
  assign n12623 = ~n9618 & n12622 ;
  assign n12624 = n2131 & n2658 ;
  assign n12625 = n5337 & n12624 ;
  assign n12626 = n5056 ^ n4091 ^ 1'b0 ;
  assign n12627 = n12625 | n12626 ;
  assign n12628 = x3 | n8241 ;
  assign n12629 = n3142 & ~n12628 ;
  assign n12630 = n10352 ^ n8036 ^ 1'b0 ;
  assign n12631 = n7421 & ~n12630 ;
  assign n12632 = n8382 ^ n7243 ^ 1'b0 ;
  assign n12633 = ~n7800 & n12632 ;
  assign n12634 = n8090 & n12633 ;
  assign n12635 = n12634 ^ n10374 ^ 1'b0 ;
  assign n12636 = ~n6703 & n12635 ;
  assign n12637 = ~n5030 & n6442 ;
  assign n12638 = ~n6442 & n12637 ;
  assign n12639 = n1414 | n2548 ;
  assign n12640 = n12638 & ~n12639 ;
  assign n12641 = n2861 | n12640 ;
  assign n12642 = n4267 | n10327 ;
  assign n12643 = n4267 & ~n12642 ;
  assign n12644 = n1684 | n3449 ;
  assign n12645 = n12644 ^ n263 ^ 1'b0 ;
  assign n12646 = ~n12643 & n12645 ;
  assign n12647 = n12643 & n12646 ;
  assign n12648 = n6059 | n12647 ;
  assign n12649 = ~n12641 & n12648 ;
  assign n12650 = n12649 ^ n11839 ^ 1'b0 ;
  assign n12651 = ~n4627 & n8512 ;
  assign n12652 = n12651 ^ n8094 ^ 1'b0 ;
  assign n12653 = n12652 ^ n3221 ^ 1'b0 ;
  assign n12654 = n6817 & n12653 ;
  assign n12655 = n1969 | n3720 ;
  assign n12656 = n946 & ~n8960 ;
  assign n12657 = n12656 ^ x157 ^ 1'b0 ;
  assign n12658 = ~n1857 & n3328 ;
  assign n12659 = ~n278 & n12658 ;
  assign n12660 = n1414 & n12659 ;
  assign n12661 = n2465 & ~n4488 ;
  assign n12662 = ~n2465 & n12661 ;
  assign n12663 = n4118 | n12662 ;
  assign n12664 = n9698 | n12663 ;
  assign n12665 = n9698 & ~n12664 ;
  assign n12666 = ~n6286 & n11814 ;
  assign n12667 = ( n519 & n4251 ) | ( n519 & ~n12666 ) | ( n4251 & ~n12666 ) ;
  assign n12668 = ~n4380 & n4564 ;
  assign n12672 = n956 | n2366 ;
  assign n12673 = n4862 & ~n12672 ;
  assign n12674 = n2022 | n12673 ;
  assign n12675 = n700 | n12674 ;
  assign n12676 = n3772 & ~n12675 ;
  assign n12677 = n12676 ^ n4874 ^ 1'b0 ;
  assign n12670 = n6049 & ~n10666 ;
  assign n12671 = n12670 ^ n4173 ^ 1'b0 ;
  assign n12669 = n4532 ^ n3536 ^ 1'b0 ;
  assign n12678 = n12677 ^ n12671 ^ n12669 ;
  assign n12679 = n12009 ^ n9052 ^ 1'b0 ;
  assign n12680 = n12679 ^ n772 ^ 1'b0 ;
  assign n12681 = n969 & n3793 ;
  assign n12682 = n1361 & n12681 ;
  assign n12683 = n2272 | n10803 ;
  assign n12684 = n12683 ^ n1173 ^ 1'b0 ;
  assign n12685 = n4884 & n10354 ;
  assign n12686 = x42 | n573 ;
  assign n12687 = n1760 & n12686 ;
  assign n12688 = n12687 ^ n10817 ^ 1'b0 ;
  assign n12689 = x78 & n12688 ;
  assign n12690 = n8578 | n11242 ;
  assign n12695 = n3865 ^ n2858 ^ 1'b0 ;
  assign n12696 = ~n3430 & n12695 ;
  assign n12697 = ~n3610 & n12696 ;
  assign n12698 = n12697 ^ n5079 ^ 1'b0 ;
  assign n12691 = ~n5530 & n7345 ;
  assign n12692 = n9463 & ~n12691 ;
  assign n12693 = n8699 | n12692 ;
  assign n12694 = n12693 ^ n12512 ^ 1'b0 ;
  assign n12699 = n12698 ^ n12694 ^ 1'b0 ;
  assign n12700 = n880 & ~n12699 ;
  assign n12701 = n5286 | n12458 ;
  assign n12702 = x223 | n12701 ;
  assign n12703 = n8691 ^ n1149 ^ 1'b0 ;
  assign n12704 = ~n2208 & n2511 ;
  assign n12705 = n7280 & n7689 ;
  assign n12706 = ~n1879 & n9913 ;
  assign n12707 = n12706 ^ n5059 ^ 1'b0 ;
  assign n12708 = n1308 | n4327 ;
  assign n12709 = n12708 ^ n9604 ^ 1'b0 ;
  assign n12710 = n12709 ^ n5253 ^ n2493 ;
  assign n12711 = ~x144 & n12695 ;
  assign n12712 = n12711 ^ n12049 ^ 1'b0 ;
  assign n12713 = n5057 & ~n12712 ;
  assign n12714 = n4313 | n12713 ;
  assign n12715 = n1128 | n6749 ;
  assign n12716 = n12715 ^ n540 ^ 1'b0 ;
  assign n12717 = n1199 & n2153 ;
  assign n12718 = ~n12716 & n12717 ;
  assign n12719 = n8152 & ~n12718 ;
  assign n12720 = ~n12714 & n12719 ;
  assign n12721 = n5675 ^ n3413 ^ 1'b0 ;
  assign n12722 = n12721 ^ n11093 ^ 1'b0 ;
  assign n12723 = n5293 | n12722 ;
  assign n12724 = n6490 & ~n9525 ;
  assign n12725 = n1684 & n12724 ;
  assign n12726 = x179 & n361 ;
  assign n12727 = ~n1630 & n12726 ;
  assign n12728 = n1195 & n12727 ;
  assign n12729 = n3399 & n3542 ;
  assign n12730 = n12728 | n12729 ;
  assign n12731 = n12730 ^ n3434 ^ 1'b0 ;
  assign n12732 = n11045 | n12731 ;
  assign n12733 = ~n3862 & n8433 ;
  assign n12734 = n1360 & n6281 ;
  assign n12735 = n10309 | n12734 ;
  assign n12736 = n5788 ^ n4793 ^ n1316 ;
  assign n12737 = n10636 | n12208 ;
  assign n12738 = n3824 ^ n2397 ^ 1'b0 ;
  assign n12739 = ~n8129 & n12738 ;
  assign n12740 = ~n3499 & n10288 ;
  assign n12741 = n12740 ^ x124 ^ 1'b0 ;
  assign n12742 = n661 | n1557 ;
  assign n12743 = n7291 | n12742 ;
  assign n12744 = n1268 & ~n2861 ;
  assign n12745 = n642 | n12744 ;
  assign n12746 = n12745 ^ n7766 ^ 1'b0 ;
  assign n12747 = n12743 & ~n12746 ;
  assign n12748 = ~n12305 & n12747 ;
  assign n12749 = n6791 & n7471 ;
  assign n12752 = x73 & n700 ;
  assign n12753 = n625 & n12752 ;
  assign n12754 = n12753 ^ n6978 ^ 1'b0 ;
  assign n12755 = ( n3476 & n6471 ) | ( n3476 & n12754 ) | ( n6471 & n12754 ) ;
  assign n12750 = n566 & ~n7822 ;
  assign n12751 = n9246 & n12750 ;
  assign n12756 = n12755 ^ n12751 ^ 1'b0 ;
  assign n12757 = n4972 ^ x98 ^ 1'b0 ;
  assign n12758 = n2082 | n12757 ;
  assign n12759 = n625 | n12758 ;
  assign n12760 = n3499 & ~n12759 ;
  assign n12765 = n1402 & ~n7014 ;
  assign n12761 = n3219 | n6571 ;
  assign n12762 = n452 | n12761 ;
  assign n12763 = ~n1366 & n6639 ;
  assign n12764 = n12762 & ~n12763 ;
  assign n12766 = n12765 ^ n12764 ^ 1'b0 ;
  assign n12767 = n6012 & n11443 ;
  assign n12768 = n1896 & n12767 ;
  assign n12769 = ( n2809 & ~n4783 ) | ( n2809 & n6621 ) | ( ~n4783 & n6621 ) ;
  assign n12770 = n9893 & ~n12769 ;
  assign n12771 = n6531 ^ n3498 ^ 1'b0 ;
  assign n12772 = n7928 & n12771 ;
  assign n12773 = n3198 | n3895 ;
  assign n12774 = ~n796 & n3988 ;
  assign n12775 = n12774 ^ n7002 ^ 1'b0 ;
  assign n12776 = n643 & ~n6523 ;
  assign n12777 = ~n9986 & n12776 ;
  assign n12778 = n12777 ^ n5189 ^ 1'b0 ;
  assign n12779 = n8443 & n12778 ;
  assign n12780 = ~n3414 & n12779 ;
  assign n12781 = n7434 ^ n4779 ^ 1'b0 ;
  assign n12782 = n1052 & ~n1133 ;
  assign n12783 = ~n11479 & n12782 ;
  assign n12784 = ~n1459 & n4380 ;
  assign n12785 = n8073 ^ n4173 ^ 1'b0 ;
  assign n12786 = n5847 ^ n3357 ^ 1'b0 ;
  assign n12787 = n12785 & ~n12786 ;
  assign n12788 = n7484 & n8036 ;
  assign n12789 = x226 & n8602 ;
  assign n12790 = ~x81 & n1241 ;
  assign n12791 = n12790 ^ x88 ^ 1'b0 ;
  assign n12792 = ~n5893 & n11961 ;
  assign n12793 = ~n949 & n3067 ;
  assign n12794 = n1046 & n12793 ;
  assign n12795 = ~n3914 & n12794 ;
  assign n12796 = n1605 | n12795 ;
  assign n12797 = n1764 | n12796 ;
  assign n12798 = n11856 & n12797 ;
  assign n12799 = n4888 ^ n886 ^ 1'b0 ;
  assign n12800 = ~n3473 & n3998 ;
  assign n12801 = n3097 & ~n4899 ;
  assign n12802 = n10711 ^ n7440 ^ 1'b0 ;
  assign n12803 = n12801 & n12802 ;
  assign n12804 = n12803 ^ n1093 ^ 1'b0 ;
  assign n12805 = n9254 ^ n4047 ^ 1'b0 ;
  assign n12806 = n5002 & n12172 ;
  assign n12807 = ~x95 & n12806 ;
  assign n12808 = n552 & ~n2382 ;
  assign n12809 = n12807 & n12808 ;
  assign n12810 = n12809 ^ n508 ^ 1'b0 ;
  assign n12811 = n1143 | n12810 ;
  assign n12812 = x154 & n4016 ;
  assign n12813 = ~n1605 & n12812 ;
  assign n12814 = n6108 & n12813 ;
  assign n12815 = n12811 & n12814 ;
  assign n12816 = n8733 ^ n2818 ^ 1'b0 ;
  assign n12817 = n7118 | n12816 ;
  assign n12818 = n12817 ^ n12317 ^ 1'b0 ;
  assign n12819 = ~n502 & n1760 ;
  assign n12820 = n12270 & ~n12819 ;
  assign n12821 = n3583 & ~n3922 ;
  assign n12823 = ~n535 & n2586 ;
  assign n12824 = ~x241 & n12823 ;
  assign n12822 = n2179 & ~n5015 ;
  assign n12825 = n12824 ^ n12822 ^ 1'b0 ;
  assign n12826 = n12825 ^ n7407 ^ 1'b0 ;
  assign n12827 = ~n2141 & n12826 ;
  assign n12828 = n8658 ^ n6028 ^ 1'b0 ;
  assign n12829 = ~n4037 & n12828 ;
  assign n12830 = n7847 & n12829 ;
  assign n12831 = n12830 ^ n3345 ^ 1'b0 ;
  assign n12832 = n2177 & n6668 ;
  assign n12833 = ~n10936 & n12832 ;
  assign n12834 = x200 & n4688 ;
  assign n12835 = n12834 ^ n4107 ^ 1'b0 ;
  assign n12836 = n12835 ^ n7135 ^ 1'b0 ;
  assign n12837 = n12833 | n12836 ;
  assign n12838 = n5146 & ~n8108 ;
  assign n12839 = ~n827 & n12838 ;
  assign n12840 = n2412 ^ n1864 ^ 1'b0 ;
  assign n12841 = ~n3115 & n12840 ;
  assign n12842 = x50 & ~n4995 ;
  assign n12843 = n12842 ^ n2330 ^ 1'b0 ;
  assign n12844 = n12843 ^ n4140 ^ 1'b0 ;
  assign n12845 = ~n12841 & n12844 ;
  assign n12846 = n3628 | n7971 ;
  assign n12847 = n12846 ^ n7720 ^ 1'b0 ;
  assign n12848 = ~n8290 & n12847 ;
  assign n12849 = n10647 ^ n7853 ^ 1'b0 ;
  assign n12850 = n2566 & n12849 ;
  assign n12851 = n5717 ^ n2022 ^ 1'b0 ;
  assign n12852 = ~n4063 & n12851 ;
  assign n12853 = n3974 ^ n2782 ^ 1'b0 ;
  assign n12854 = x94 & n7138 ;
  assign n12855 = n12854 ^ x27 ^ 1'b0 ;
  assign n12856 = ~n12853 & n12855 ;
  assign n12857 = n10751 & n12856 ;
  assign n12858 = n8480 ^ n4449 ^ 1'b0 ;
  assign n12859 = n9817 & ~n12858 ;
  assign n12860 = n3983 & ~n6560 ;
  assign n12861 = n825 & ~n12860 ;
  assign n12862 = n4178 ^ n401 ^ 1'b0 ;
  assign n12863 = n8874 | n12862 ;
  assign n12864 = n3948 ^ n3692 ^ 1'b0 ;
  assign n12865 = n7031 & n12864 ;
  assign n12866 = ~n2066 & n2361 ;
  assign n12867 = ~n6539 & n12866 ;
  assign n12868 = n6990 & ~n12867 ;
  assign n12869 = n4340 ^ n2728 ^ 1'b0 ;
  assign n12870 = n8118 & n12869 ;
  assign n12871 = n4350 | n12870 ;
  assign n12872 = n12871 ^ n2591 ^ 1'b0 ;
  assign n12873 = n10579 | n11612 ;
  assign n12874 = n5493 | n12873 ;
  assign n12875 = n11612 ^ n5914 ^ 1'b0 ;
  assign n12876 = x232 & ~n12875 ;
  assign n12877 = n6461 & ~n12876 ;
  assign n12878 = n7706 & ~n11150 ;
  assign n12879 = n2626 & ~n3302 ;
  assign n12880 = n5411 & n11718 ;
  assign n12881 = n4601 & n9428 ;
  assign n12882 = n12881 ^ n3105 ^ 1'b0 ;
  assign n12883 = n12880 & ~n12882 ;
  assign n12884 = n12879 & n12883 ;
  assign n12885 = n7671 ^ n2875 ^ 1'b0 ;
  assign n12886 = n3452 ^ x87 ^ 1'b0 ;
  assign n12887 = n4467 & n12886 ;
  assign n12888 = n3175 & n12887 ;
  assign n12889 = n6484 | n12888 ;
  assign n12890 = n12889 ^ n6236 ^ 1'b0 ;
  assign n12891 = n11010 & ~n12890 ;
  assign n12892 = n4012 ^ n3989 ^ n2129 ;
  assign n12893 = ( n3345 & ~n5694 ) | ( n3345 & n6540 ) | ( ~n5694 & n6540 ) ;
  assign n12894 = n5222 ^ n1159 ^ 1'b0 ;
  assign n12895 = ~n12893 & n12894 ;
  assign n12896 = n12895 ^ n10341 ^ 1'b0 ;
  assign n12897 = n957 & n1773 ;
  assign n12898 = ~n12543 & n12897 ;
  assign n12899 = n1651 & ~n9651 ;
  assign n12900 = ~n3171 & n12899 ;
  assign n12901 = ~n638 & n1740 ;
  assign n12902 = n6287 & ~n12901 ;
  assign n12903 = n7276 & n12902 ;
  assign n12904 = n4596 & n12147 ;
  assign n12905 = n12904 ^ x182 ^ 1'b0 ;
  assign n12906 = x76 | n3740 ;
  assign n12907 = n7411 & ~n8553 ;
  assign n12908 = n12907 ^ n11738 ^ 1'b0 ;
  assign n12909 = n535 & n1571 ;
  assign n12910 = n3064 ^ n512 ^ 1'b0 ;
  assign n12911 = ~n12909 & n12910 ;
  assign n12912 = n4814 ^ n876 ^ 1'b0 ;
  assign n12913 = n12912 ^ n8333 ^ 1'b0 ;
  assign n12914 = n298 & ~n12913 ;
  assign n12915 = n4897 ^ n4021 ^ 1'b0 ;
  assign n12916 = n5191 & n9948 ;
  assign n12917 = n4256 | n12916 ;
  assign n12918 = x157 | n2910 ;
  assign n12919 = n12918 ^ n11895 ^ 1'b0 ;
  assign n12920 = ~n1429 & n5261 ;
  assign n12921 = n3265 & ~n12920 ;
  assign n12922 = n12919 & ~n12921 ;
  assign n12923 = ( n4378 & ~n6895 ) | ( n4378 & n11488 ) | ( ~n6895 & n11488 ) ;
  assign n12924 = n7642 | n11814 ;
  assign n12925 = n6807 ^ n1324 ^ 1'b0 ;
  assign n12926 = n524 & n12925 ;
  assign n12927 = n12926 ^ n9173 ^ 1'b0 ;
  assign n12928 = n2887 & n12927 ;
  assign n12929 = n7828 | n12928 ;
  assign n12930 = n1723 & ~n12929 ;
  assign n12931 = n12930 ^ n4516 ^ 1'b0 ;
  assign n12932 = n7009 & n8797 ;
  assign n12933 = ~n10089 & n12932 ;
  assign n12934 = n3688 ^ n663 ^ 1'b0 ;
  assign n12940 = n936 | n3629 ;
  assign n12935 = n4565 ^ n3989 ^ 1'b0 ;
  assign n12936 = ~n456 & n12935 ;
  assign n12937 = n2392 & n10181 ;
  assign n12938 = ~n12936 & n12937 ;
  assign n12939 = n7127 & ~n12938 ;
  assign n12941 = n12940 ^ n12939 ^ 1'b0 ;
  assign n12943 = n1923 ^ n259 ^ x93 ;
  assign n12944 = n1368 & ~n12943 ;
  assign n12945 = n12944 ^ x47 ^ 1'b0 ;
  assign n12946 = x5 | n11330 ;
  assign n12947 = n12945 | n12946 ;
  assign n12948 = n3879 | n12947 ;
  assign n12942 = n7257 | n11657 ;
  assign n12949 = n12948 ^ n12942 ^ 1'b0 ;
  assign n12950 = ~n1383 & n11353 ;
  assign n12951 = n1285 & ~n7107 ;
  assign n12952 = n3878 & ~n12951 ;
  assign n12953 = n2394 & ~n11518 ;
  assign n12954 = n11518 & n12953 ;
  assign n12955 = n12703 ^ n5125 ^ 1'b0 ;
  assign n12956 = n5907 | n6969 ;
  assign n12957 = ( ~n2274 & n5574 ) | ( ~n2274 & n10330 ) | ( n5574 & n10330 ) ;
  assign n12958 = n12002 ^ n5025 ^ 1'b0 ;
  assign n12959 = n1700 & ~n12958 ;
  assign n12960 = n4180 ^ n1183 ^ 1'b0 ;
  assign n12961 = n2261 & ~n12960 ;
  assign n12962 = n12961 ^ n9693 ^ n1091 ;
  assign n12963 = n12962 ^ n8560 ^ n4304 ;
  assign n12964 = ~n840 & n10990 ;
  assign n12965 = n12964 ^ n1499 ^ 1'b0 ;
  assign n12966 = ~n12963 & n12965 ;
  assign n12967 = n5422 & ~n12966 ;
  assign n12968 = n967 & ~n5958 ;
  assign n12969 = ~n12420 & n12968 ;
  assign n12970 = n1492 ^ n750 ^ 1'b0 ;
  assign n12971 = n9721 & n12970 ;
  assign n12972 = n1797 & n12971 ;
  assign n12973 = ( n1825 & n2855 ) | ( n1825 & n12972 ) | ( n2855 & n12972 ) ;
  assign n12974 = n833 & ~n1572 ;
  assign n12975 = ~n532 & n4181 ;
  assign n12976 = n5200 ^ n2529 ^ 1'b0 ;
  assign n12977 = ~n3532 & n12976 ;
  assign n12978 = n12977 ^ n9084 ^ 1'b0 ;
  assign n12979 = n12975 & n12978 ;
  assign n12980 = n2411 & n5890 ;
  assign n12981 = n9438 ^ n3798 ^ 1'b0 ;
  assign n12982 = n528 & ~n5862 ;
  assign n12983 = n12495 | n12982 ;
  assign n12984 = n12137 ^ n337 ^ 1'b0 ;
  assign n12985 = n5125 | n12984 ;
  assign n12986 = n3308 & ~n10080 ;
  assign n12987 = n3140 & n10389 ;
  assign n12988 = n3153 & n12987 ;
  assign n12989 = n12988 ^ n10433 ^ 1'b0 ;
  assign n12990 = n2336 | n2366 ;
  assign n12991 = ~n1642 & n5898 ;
  assign n12992 = n12991 ^ n1740 ^ 1'b0 ;
  assign n12993 = n7179 | n12992 ;
  assign n12994 = n10721 & ~n12993 ;
  assign n12995 = n12990 & n12994 ;
  assign n12997 = n8412 ^ n3112 ^ 1'b0 ;
  assign n12996 = n4616 & n9795 ;
  assign n12998 = n12997 ^ n12996 ^ 1'b0 ;
  assign n12999 = n7601 | n8811 ;
  assign n13000 = n12999 ^ n8752 ^ 1'b0 ;
  assign n13001 = ~n808 & n2392 ;
  assign n13002 = n13001 ^ n8242 ^ 1'b0 ;
  assign n13003 = n10179 & n13002 ;
  assign n13004 = n11059 ^ n9820 ^ 1'b0 ;
  assign n13005 = ~n5373 & n13004 ;
  assign n13006 = ~n6061 & n7451 ;
  assign n13007 = ~n7451 & n13006 ;
  assign n13008 = n1028 & n2737 ;
  assign n13009 = n13007 & n13008 ;
  assign n13010 = n2190 | n13009 ;
  assign n13011 = n2161 ^ n486 ^ 1'b0 ;
  assign n13012 = n1173 & n13011 ;
  assign n13013 = n3558 & ~n10097 ;
  assign n13014 = ~n3558 & n13013 ;
  assign n13015 = n13012 & ~n13014 ;
  assign n13016 = ~n13012 & n13015 ;
  assign n13017 = n7115 | n13016 ;
  assign n13018 = n7115 & ~n13017 ;
  assign n13019 = n13010 & ~n13018 ;
  assign n13020 = n8150 ^ n6375 ^ 1'b0 ;
  assign n13021 = ~n7253 & n8428 ;
  assign n13022 = n10296 & n13021 ;
  assign n13023 = n1930 & n4779 ;
  assign n13024 = n1689 | n13023 ;
  assign n13025 = n13024 ^ n4189 ^ 1'b0 ;
  assign n13027 = n8679 ^ n803 ^ 1'b0 ;
  assign n13028 = n3936 ^ n378 ^ 1'b0 ;
  assign n13029 = n4222 & n13028 ;
  assign n13030 = x31 & ~n13029 ;
  assign n13031 = n12185 & ~n13030 ;
  assign n13032 = ~n13027 & n13031 ;
  assign n13026 = n4777 ^ n3249 ^ 1'b0 ;
  assign n13033 = n13032 ^ n13026 ^ 1'b0 ;
  assign n13034 = x176 ^ x20 ^ 1'b0 ;
  assign n13035 = n13034 ^ n12030 ^ 1'b0 ;
  assign n13036 = n11469 & n13035 ;
  assign n13037 = n1310 & n1666 ;
  assign n13038 = ~n4948 & n13037 ;
  assign n13039 = n1616 & ~n13038 ;
  assign n13040 = ~n3678 & n13039 ;
  assign n13041 = n7142 & ~n13040 ;
  assign n13042 = n552 & n13041 ;
  assign n13045 = n3768 ^ n2374 ^ 1'b0 ;
  assign n13046 = n13045 ^ n7006 ^ 1'b0 ;
  assign n13043 = n3442 ^ n2633 ^ 1'b0 ;
  assign n13044 = n6079 | n13043 ;
  assign n13047 = n13046 ^ n13044 ^ 1'b0 ;
  assign n13048 = n9431 ^ n3125 ^ 1'b0 ;
  assign n13049 = n1544 & ~n3578 ;
  assign n13050 = n12389 ^ n4794 ^ 1'b0 ;
  assign n13051 = n4539 & ~n13050 ;
  assign n13052 = n13051 ^ n5946 ^ n2193 ;
  assign n13053 = n13052 ^ n4480 ^ 1'b0 ;
  assign n13054 = ~x33 & n6964 ;
  assign n13055 = n4124 ^ n1217 ^ 1'b0 ;
  assign n13056 = n13054 & n13055 ;
  assign n13057 = n4469 & ~n13056 ;
  assign n13061 = n1949 ^ n323 ^ 1'b0 ;
  assign n13062 = n4874 & n13061 ;
  assign n13058 = n774 ^ n257 ^ 1'b0 ;
  assign n13059 = n6178 & ~n13058 ;
  assign n13060 = ~n7045 & n13059 ;
  assign n13063 = n13062 ^ n13060 ^ 1'b0 ;
  assign n13064 = n13063 ^ n7415 ^ 1'b0 ;
  assign n13065 = n1901 ^ n1320 ^ 1'b0 ;
  assign n13066 = n2431 & ~n13065 ;
  assign n13067 = n13066 ^ n423 ^ 1'b0 ;
  assign n13068 = n6322 ^ n2868 ^ 1'b0 ;
  assign n13069 = ~n13067 & n13068 ;
  assign n13070 = n772 | n10080 ;
  assign n13071 = n10237 ^ n6427 ^ 1'b0 ;
  assign n13072 = n8755 | n13071 ;
  assign n13073 = n13072 ^ n3611 ^ 1'b0 ;
  assign n13074 = n6940 ^ n5487 ^ 1'b0 ;
  assign n13075 = n13073 | n13074 ;
  assign n13077 = ~n488 & n2207 ;
  assign n13076 = n776 ^ n275 ^ x75 ;
  assign n13078 = n13077 ^ n13076 ^ 1'b0 ;
  assign n13079 = n2026 | n9170 ;
  assign n13080 = x241 | n13079 ;
  assign n13081 = n3891 | n7223 ;
  assign n13083 = n3671 ^ n1783 ^ 1'b0 ;
  assign n13084 = ~n573 & n13083 ;
  assign n13082 = n10821 ^ n3592 ^ 1'b0 ;
  assign n13085 = n13084 ^ n13082 ^ 1'b0 ;
  assign n13086 = n3143 & ~n13085 ;
  assign n13087 = n6823 ^ n3055 ^ 1'b0 ;
  assign n13088 = n11524 ^ n10716 ^ n4657 ;
  assign n13089 = n8821 ^ n5047 ^ 1'b0 ;
  assign n13090 = ~n4096 & n7272 ;
  assign n13091 = ~n1360 & n13090 ;
  assign n13092 = n7872 ^ n7864 ^ 1'b0 ;
  assign n13093 = n9981 ^ n6401 ^ n1880 ;
  assign n13094 = n3090 | n5818 ;
  assign n13095 = n2185 & ~n13094 ;
  assign n13096 = n10613 ^ n1732 ^ 1'b0 ;
  assign n13097 = x236 ^ x88 ^ 1'b0 ;
  assign n13098 = n2188 & n13097 ;
  assign n13099 = n9563 & ~n13098 ;
  assign n13100 = n13099 ^ n5311 ^ 1'b0 ;
  assign n13102 = x190 | n283 ;
  assign n13101 = n2588 & n3130 ;
  assign n13103 = n13102 ^ n13101 ^ 1'b0 ;
  assign n13104 = n4265 ^ n2437 ^ 1'b0 ;
  assign n13105 = n6668 & ~n7869 ;
  assign n13106 = ~n13104 & n13105 ;
  assign n13107 = n13106 ^ n12077 ^ 1'b0 ;
  assign n13108 = n13103 | n13107 ;
  assign n13109 = n552 & ~n13108 ;
  assign n13110 = n5642 ^ n3289 ^ x46 ;
  assign n13111 = ~n6300 & n7113 ;
  assign n13112 = n5928 | n7951 ;
  assign n13113 = n13112 ^ n2423 ^ 1'b0 ;
  assign n13114 = n2014 | n2179 ;
  assign n13115 = n13113 | n13114 ;
  assign n13116 = ~n8094 & n13115 ;
  assign n13117 = n13116 ^ n11218 ^ 1'b0 ;
  assign n13118 = n10731 & n13117 ;
  assign n13120 = x156 & n7561 ;
  assign n13121 = n13120 ^ n4970 ^ 1'b0 ;
  assign n13122 = n5625 | n13121 ;
  assign n13123 = n13122 ^ n11648 ^ 1'b0 ;
  assign n13119 = n12121 & n12695 ;
  assign n13124 = n13123 ^ n13119 ^ 1'b0 ;
  assign n13125 = x112 | n593 ;
  assign n13130 = n570 & ~n4271 ;
  assign n13131 = n13130 ^ n967 ^ 1'b0 ;
  assign n13132 = ~n1304 & n2057 ;
  assign n13133 = ~n3844 & n13132 ;
  assign n13134 = ~n901 & n1793 ;
  assign n13135 = n4101 | n5891 ;
  assign n13136 = n13134 & n13135 ;
  assign n13137 = n13133 & n13136 ;
  assign n13138 = n13131 | n13137 ;
  assign n13139 = n13138 ^ n3946 ^ 1'b0 ;
  assign n13126 = ~n1527 & n3929 ;
  assign n13127 = ~n8808 & n13126 ;
  assign n13128 = ~n798 & n8915 ;
  assign n13129 = n13127 & n13128 ;
  assign n13140 = n13139 ^ n13129 ^ n3046 ;
  assign n13141 = n6410 | n12196 ;
  assign n13142 = n13141 ^ n12924 ^ 1'b0 ;
  assign n13143 = n6117 ^ n4356 ^ 1'b0 ;
  assign n13144 = n13143 ^ n3187 ^ 1'b0 ;
  assign n13145 = n3186 & n7246 ;
  assign n13146 = n6041 & ~n7384 ;
  assign n13147 = n2914 & n13146 ;
  assign n13148 = n13147 ^ n11101 ^ 1'b0 ;
  assign n13149 = n13145 & n13148 ;
  assign n13150 = ~n9266 & n13149 ;
  assign n13151 = n13150 ^ n11183 ^ 1'b0 ;
  assign n13152 = n9035 ^ n7494 ^ 1'b0 ;
  assign n13153 = n1395 & n1494 ;
  assign n13154 = x101 | n13153 ;
  assign n13155 = n13154 ^ n10106 ^ 1'b0 ;
  assign n13159 = n5493 & ~n8687 ;
  assign n13156 = ~x189 & n2760 ;
  assign n13157 = n4177 & n13156 ;
  assign n13158 = n3522 & n13157 ;
  assign n13160 = n13159 ^ n13158 ^ 1'b0 ;
  assign n13161 = n4736 | n7144 ;
  assign n13162 = n6396 | n13161 ;
  assign n13163 = n13162 ^ n5376 ^ 1'b0 ;
  assign n13164 = ( x42 & ~n2765 ) | ( x42 & n3171 ) | ( ~n2765 & n3171 ) ;
  assign n13165 = n3082 & n13164 ;
  assign n13166 = ~n2345 & n13165 ;
  assign n13167 = n5189 ^ n1094 ^ 1'b0 ;
  assign n13168 = n1262 & ~n13167 ;
  assign n13169 = n10446 & n13168 ;
  assign n13170 = n13166 | n13169 ;
  assign n13171 = n13170 ^ n6401 ^ 1'b0 ;
  assign n13172 = ( n5213 & ~n10217 ) | ( n5213 & n13076 ) | ( ~n10217 & n13076 ) ;
  assign n13173 = n9191 ^ n2844 ^ 1'b0 ;
  assign n13174 = ~n8436 & n13173 ;
  assign n13175 = n13174 ^ n3620 ^ 1'b0 ;
  assign n13176 = n3661 ^ n1601 ^ 1'b0 ;
  assign n13177 = n7628 | n13176 ;
  assign n13178 = n9219 | n10122 ;
  assign n13179 = n2590 & n5154 ;
  assign n13180 = n7019 ^ n3308 ^ 1'b0 ;
  assign n13181 = ~n3747 & n6747 ;
  assign n13182 = ~x26 & n13181 ;
  assign n13183 = n6218 ^ n323 ^ 1'b0 ;
  assign n13184 = n13029 & ~n13183 ;
  assign n13186 = ( n3452 & n5682 ) | ( n3452 & n6065 ) | ( n5682 & n6065 ) ;
  assign n13187 = ( n1240 & ~n2828 ) | ( n1240 & n13186 ) | ( ~n2828 & n13186 ) ;
  assign n13188 = n5253 | n13187 ;
  assign n13189 = n10213 | n13188 ;
  assign n13185 = n11961 & n12119 ;
  assign n13190 = n13189 ^ n13185 ^ 1'b0 ;
  assign n13191 = n1415 & n1668 ;
  assign n13192 = ~n1266 & n13191 ;
  assign n13193 = ~n1772 & n13192 ;
  assign n13194 = n13193 ^ n4922 ^ 1'b0 ;
  assign n13195 = n5081 & n13194 ;
  assign n13196 = n3758 ^ n3280 ^ 1'b0 ;
  assign n13197 = n4652 & ~n13196 ;
  assign n13198 = ~n9183 & n13197 ;
  assign n13199 = n7448 & n13198 ;
  assign n13200 = n5370 | n13199 ;
  assign n13201 = n6788 | n13200 ;
  assign n13202 = ~x3 & n7366 ;
  assign n13203 = n9162 & n13202 ;
  assign n13204 = n1602 ^ n959 ^ x123 ;
  assign n13205 = n13204 ^ n1405 ^ 1'b0 ;
  assign n13206 = n5717 ^ n2250 ^ 1'b0 ;
  assign n13207 = ~n2951 & n13206 ;
  assign n13208 = n13207 ^ n4736 ^ 1'b0 ;
  assign n13209 = n6763 | n13208 ;
  assign n13210 = n8443 ^ n5627 ^ 1'b0 ;
  assign n13212 = x174 & ~n2352 ;
  assign n13213 = n13212 ^ n7232 ^ 1'b0 ;
  assign n13211 = n6241 & ~n10187 ;
  assign n13214 = n13213 ^ n13211 ^ 1'b0 ;
  assign n13215 = n12405 ^ n3403 ^ 1'b0 ;
  assign n13216 = n13215 ^ n820 ^ 1'b0 ;
  assign n13217 = n13214 & ~n13216 ;
  assign n13218 = x63 & ~n13217 ;
  assign n13219 = n3567 | n8637 ;
  assign n13220 = n7259 | n13219 ;
  assign n13221 = n7643 ^ n2350 ^ 1'b0 ;
  assign n13222 = n13220 & n13221 ;
  assign n13223 = n2476 & n7715 ;
  assign n13224 = n4389 ^ n2606 ^ 1'b0 ;
  assign n13225 = n1620 | n13224 ;
  assign n13226 = n3286 | n13225 ;
  assign n13227 = n2029 ^ n1266 ^ 1'b0 ;
  assign n13228 = ( n3250 & n9537 ) | ( n3250 & n13227 ) | ( n9537 & n13227 ) ;
  assign n13229 = n8233 ^ n6297 ^ 1'b0 ;
  assign n13230 = ~n5485 & n13229 ;
  assign n13231 = n11565 & n13230 ;
  assign n13232 = n5379 & n5468 ;
  assign n13233 = n13232 ^ n4228 ^ 1'b0 ;
  assign n13234 = n13231 & n13233 ;
  assign n13236 = n6944 ^ n2404 ^ 1'b0 ;
  assign n13237 = n372 & n13236 ;
  assign n13235 = n8031 | n11264 ;
  assign n13238 = n13237 ^ n13235 ^ 1'b0 ;
  assign n13239 = n9007 & n13238 ;
  assign n13240 = ~n8881 & n9951 ;
  assign n13241 = n13240 ^ n941 ^ 1'b0 ;
  assign n13242 = n273 & n6548 ;
  assign n13243 = n13242 ^ x224 ^ 1'b0 ;
  assign n13244 = n7011 ^ n4992 ^ 1'b0 ;
  assign n13245 = n2061 | n13244 ;
  assign n13246 = n7802 & ~n13245 ;
  assign n13247 = n13246 ^ n259 ^ 1'b0 ;
  assign n13248 = n3187 & n5368 ;
  assign n13249 = n13247 & ~n13248 ;
  assign n13250 = n13249 ^ n2953 ^ 1'b0 ;
  assign n13253 = n4796 & n11431 ;
  assign n13251 = n461 & n8820 ;
  assign n13252 = ~n5407 & n13251 ;
  assign n13254 = n13253 ^ n13252 ^ 1'b0 ;
  assign n13255 = n7408 | n13254 ;
  assign n13256 = n6320 ^ n4048 ^ 1'b0 ;
  assign n13257 = n13256 ^ n490 ^ 1'b0 ;
  assign n13258 = n13255 | n13257 ;
  assign n13259 = n3476 & ~n10908 ;
  assign n13260 = n13259 ^ n4024 ^ 1'b0 ;
  assign n13261 = n2652 ^ x37 ^ 1'b0 ;
  assign n13262 = n11910 ^ n5929 ^ 1'b0 ;
  assign n13263 = n4157 | n11804 ;
  assign n13264 = n13263 ^ n4611 ^ 1'b0 ;
  assign n13265 = n9001 & n10811 ;
  assign n13266 = n4539 & ~n13265 ;
  assign n13267 = n903 ^ x0 ^ 1'b0 ;
  assign n13268 = n13267 ^ x153 ^ 1'b0 ;
  assign n13269 = n1510 | n1678 ;
  assign n13270 = n13269 ^ n3721 ^ 1'b0 ;
  assign n13271 = n10777 ^ n2569 ^ 1'b0 ;
  assign n13274 = n9077 ^ n2982 ^ 1'b0 ;
  assign n13275 = n5086 & n13274 ;
  assign n13276 = n5134 ^ n1951 ^ 1'b0 ;
  assign n13277 = n13275 & n13276 ;
  assign n13272 = ~x98 & n10107 ;
  assign n13273 = n13272 ^ n2486 ^ 1'b0 ;
  assign n13278 = n13277 ^ n13273 ^ 1'b0 ;
  assign n13279 = n6080 | n13278 ;
  assign n13280 = n1697 & n13279 ;
  assign n13281 = n6229 ^ n5093 ^ n3589 ;
  assign n13282 = n8155 & ~n13281 ;
  assign n13283 = n13282 ^ n3882 ^ 1'b0 ;
  assign n13284 = n7301 & ~n8918 ;
  assign n13285 = n9796 & n13284 ;
  assign n13286 = n3447 & ~n13285 ;
  assign n13287 = n12758 | n13286 ;
  assign n13288 = n8435 & ~n13287 ;
  assign n13289 = n3764 ^ n1077 ^ 1'b0 ;
  assign n13290 = x2 & ~n13289 ;
  assign n13291 = n13290 ^ n2148 ^ 1'b0 ;
  assign n13292 = n13291 ^ n7076 ^ 1'b0 ;
  assign n13293 = n6662 | n13292 ;
  assign n13294 = n13293 ^ n7973 ^ 1'b0 ;
  assign n13295 = n8716 & ~n8890 ;
  assign n13296 = n9142 & n10087 ;
  assign n13300 = n1866 & n2143 ;
  assign n13301 = n13300 ^ n1223 ^ 1'b0 ;
  assign n13297 = n4351 ^ n3226 ^ 1'b0 ;
  assign n13298 = n8756 & ~n13297 ;
  assign n13299 = n6557 & n13298 ;
  assign n13302 = n13301 ^ n13299 ^ 1'b0 ;
  assign n13303 = n4928 & ~n10590 ;
  assign n13304 = n5312 | n13303 ;
  assign n13305 = x110 | n13304 ;
  assign n13306 = ( n1941 & n3536 ) | ( n1941 & n7792 ) | ( n3536 & n7792 ) ;
  assign n13307 = n4771 & n11816 ;
  assign n13308 = ~n3451 & n13307 ;
  assign n13309 = n7154 ^ n1634 ^ 1'b0 ;
  assign n13310 = n13308 & ~n13309 ;
  assign n13311 = n6412 ^ n1959 ^ 1'b0 ;
  assign n13312 = n3590 | n4142 ;
  assign n13313 = n2191 & ~n13312 ;
  assign n13314 = n2039 & n13313 ;
  assign n13315 = n675 & ~n2256 ;
  assign n13316 = n3485 & n7337 ;
  assign n13317 = n7982 & n13316 ;
  assign n13318 = n2357 & ~n13317 ;
  assign n13319 = n13318 ^ n3052 ^ 1'b0 ;
  assign n13320 = n3941 & n13319 ;
  assign n13321 = ~n10714 & n13320 ;
  assign n13322 = n864 ^ n553 ^ 1'b0 ;
  assign n13323 = n13322 ^ n12337 ^ 1'b0 ;
  assign n13324 = n9387 ^ n8929 ^ 1'b0 ;
  assign n13325 = x251 | n10893 ;
  assign n13326 = n1402 | n4013 ;
  assign n13327 = n1411 ^ x144 ^ 1'b0 ;
  assign n13328 = n1071 & n6974 ;
  assign n13329 = ~n2681 & n13328 ;
  assign n13330 = n3112 & ~n3499 ;
  assign n13331 = n5968 & n13330 ;
  assign n13332 = n1511 ^ x130 ^ 1'b0 ;
  assign n13333 = ~n4340 & n13332 ;
  assign n13334 = ~n3832 & n13333 ;
  assign n13335 = n13334 ^ n6712 ^ 1'b0 ;
  assign n13336 = n5324 | n13335 ;
  assign n13337 = n13335 & ~n13336 ;
  assign n13338 = x220 & ~n13337 ;
  assign n13339 = ~n4068 & n5581 ;
  assign n13340 = n2652 & ~n13339 ;
  assign n13341 = ~n13338 & n13340 ;
  assign n13342 = n2076 | n4118 ;
  assign n13343 = n6595 & ~n13342 ;
  assign n13344 = n7928 ^ x253 ^ 1'b0 ;
  assign n13345 = n13343 | n13344 ;
  assign n13346 = n13345 ^ n2885 ^ 1'b0 ;
  assign n13347 = n1675 & ~n12247 ;
  assign n13348 = ~x112 & n13347 ;
  assign n13349 = n456 & n6804 ;
  assign n13350 = n13349 ^ n7373 ^ 1'b0 ;
  assign n13351 = n3789 ^ n2837 ^ 1'b0 ;
  assign n13352 = n1415 & n13351 ;
  assign n13353 = n3982 ^ n313 ^ 1'b0 ;
  assign n13354 = n13352 & ~n13353 ;
  assign n13355 = ~n3563 & n13354 ;
  assign n13356 = ~n5676 & n11645 ;
  assign n13357 = n2324 & n3803 ;
  assign n13358 = n13357 ^ n5849 ^ 1'b0 ;
  assign n13359 = ~n1320 & n11100 ;
  assign n13362 = n8730 ^ n366 ^ 1'b0 ;
  assign n13363 = n3209 & ~n5170 ;
  assign n13364 = ~n13362 & n13363 ;
  assign n13365 = n6480 & n13364 ;
  assign n13360 = n1226 ^ n851 ^ 1'b0 ;
  assign n13361 = n602 & n13360 ;
  assign n13366 = n13365 ^ n13361 ^ 1'b0 ;
  assign n13367 = n13366 ^ n7494 ^ 1'b0 ;
  assign n13368 = n13359 & ~n13367 ;
  assign n13369 = n8246 | n10414 ;
  assign n13370 = n8324 ^ n3180 ^ 1'b0 ;
  assign n13371 = ~n6523 & n11122 ;
  assign n13372 = n13371 ^ n8295 ^ 1'b0 ;
  assign n13373 = n452 ^ x122 ^ 1'b0 ;
  assign n13374 = n4834 & n13373 ;
  assign n13375 = n13374 ^ x151 ^ 1'b0 ;
  assign n13376 = n13375 ^ n698 ^ 1'b0 ;
  assign n13377 = ~n13372 & n13376 ;
  assign n13378 = n9946 & n13377 ;
  assign n13379 = n13378 ^ n5907 ^ 1'b0 ;
  assign n13380 = n3878 ^ n2955 ^ 1'b0 ;
  assign n13381 = n5097 ^ n2936 ^ 1'b0 ;
  assign n13382 = n13381 ^ n9626 ^ n1822 ;
  assign n13383 = n13382 ^ n5443 ^ 1'b0 ;
  assign n13384 = n7993 | n12064 ;
  assign n13385 = n5481 & ~n13384 ;
  assign n13386 = ~n1951 & n8660 ;
  assign n13387 = ~n923 & n13386 ;
  assign n13388 = n3039 & ~n5250 ;
  assign n13389 = n13388 ^ n3756 ^ 1'b0 ;
  assign n13390 = n1402 & n7076 ;
  assign n13391 = n1693 & n13390 ;
  assign n13392 = n8624 ^ n8567 ^ 1'b0 ;
  assign n13393 = n313 | n13392 ;
  assign n13394 = n13393 ^ n6095 ^ 1'b0 ;
  assign n13395 = n3180 & n5837 ;
  assign n13396 = ~n818 & n13395 ;
  assign n13397 = n10551 ^ n2148 ^ n988 ;
  assign n13398 = n2537 ^ n1792 ^ 1'b0 ;
  assign n13399 = n6047 ^ n4579 ^ 1'b0 ;
  assign n13400 = n13398 & ~n13399 ;
  assign n13401 = n13400 ^ n1678 ^ 1'b0 ;
  assign n13402 = ~n3404 & n6344 ;
  assign n13403 = ~n4677 & n13402 ;
  assign n13404 = n5703 & ~n13403 ;
  assign n13405 = ~n13401 & n13404 ;
  assign n13408 = n4432 & n8397 ;
  assign n13409 = n13408 ^ n4491 ^ 1'b0 ;
  assign n13406 = n1841 ^ n395 ^ 1'b0 ;
  assign n13407 = n2452 & ~n13406 ;
  assign n13410 = n13409 ^ n13407 ^ 1'b0 ;
  assign n13411 = ~n3321 & n4151 ;
  assign n13412 = ~n3620 & n10367 ;
  assign n13413 = n13412 ^ n4224 ^ 1'b0 ;
  assign n13414 = n300 & ~n1298 ;
  assign n13415 = n2554 & ~n13414 ;
  assign n13416 = n2955 & n13415 ;
  assign n13417 = n9855 ^ n6195 ^ 1'b0 ;
  assign n13418 = n1685 & ~n13417 ;
  assign n13419 = n446 & n3807 ;
  assign n13420 = n6884 & n13419 ;
  assign n13421 = n13420 ^ n13152 ^ 1'b0 ;
  assign n13422 = n7163 & n13421 ;
  assign n13423 = n4024 & ~n7768 ;
  assign n13424 = ~n3093 & n13423 ;
  assign n13425 = n1029 & ~n7845 ;
  assign n13426 = n13425 ^ x179 ^ 1'b0 ;
  assign n13427 = n13426 ^ n8793 ^ 1'b0 ;
  assign n13428 = n7212 & n13427 ;
  assign n13429 = n6273 & n13428 ;
  assign n13430 = n13424 & n13429 ;
  assign n13431 = ( n2218 & n2252 ) | ( n2218 & n3447 ) | ( n2252 & n3447 ) ;
  assign n13432 = ~n2689 & n13431 ;
  assign n13433 = n518 & n13432 ;
  assign n13434 = n8367 & ~n11964 ;
  assign n13435 = n2954 | n8474 ;
  assign n13436 = ~n9918 & n13435 ;
  assign n13437 = ~n1819 & n13436 ;
  assign n13438 = n3365 & ~n5005 ;
  assign n13440 = n894 | n7146 ;
  assign n13441 = n13440 ^ n1178 ^ 1'b0 ;
  assign n13439 = n2973 ^ n1703 ^ 1'b0 ;
  assign n13442 = n13441 ^ n13439 ^ 1'b0 ;
  assign n13443 = n13438 & n13442 ;
  assign n13444 = n3782 & n4537 ;
  assign n13445 = ~x222 & n13444 ;
  assign n13446 = x218 & n13445 ;
  assign n13447 = n1361 | n1511 ;
  assign n13448 = n3021 ^ n1285 ^ 1'b0 ;
  assign n13449 = n13447 & ~n13448 ;
  assign n13450 = ~n3520 & n8716 ;
  assign n13451 = ~n13449 & n13450 ;
  assign n13452 = n10682 ^ n3140 ^ 1'b0 ;
  assign n13453 = n1243 | n1920 ;
  assign n13454 = n7898 ^ n1873 ^ 1'b0 ;
  assign n13455 = n5445 & n13454 ;
  assign n13456 = n5350 & n13455 ;
  assign n13457 = n5121 | n8246 ;
  assign n13458 = n13457 ^ n8760 ^ 1'b0 ;
  assign n13459 = n13456 & n13458 ;
  assign n13460 = n13459 ^ n9121 ^ n824 ;
  assign n13465 = n1888 & ~n4828 ;
  assign n13466 = ~n1888 & n13465 ;
  assign n13461 = n876 & ~n3993 ;
  assign n13462 = ~n876 & n13461 ;
  assign n13463 = n10296 & ~n13462 ;
  assign n13464 = n2857 & n13463 ;
  assign n13467 = n13466 ^ n13464 ^ 1'b0 ;
  assign n13468 = n11147 ^ n6905 ^ 1'b0 ;
  assign n13469 = n13468 ^ n7280 ^ 1'b0 ;
  assign n13470 = n3982 & n13469 ;
  assign n13471 = n13470 ^ n7847 ^ 1'b0 ;
  assign n13472 = ~n11713 & n13471 ;
  assign n13473 = n8803 | n12585 ;
  assign n13474 = n8825 ^ n1610 ^ 1'b0 ;
  assign n13475 = n12841 & n13474 ;
  assign n13476 = n10845 | n13475 ;
  assign n13477 = n414 & ~n3343 ;
  assign n13478 = n13477 ^ n2962 ^ 1'b0 ;
  assign n13479 = n11152 & ~n13478 ;
  assign n13480 = n4808 | n5151 ;
  assign n13481 = n9466 & ~n13480 ;
  assign n13482 = ~n3258 & n4562 ;
  assign n13483 = n13482 ^ n1883 ^ 1'b0 ;
  assign n13484 = n10844 | n13483 ;
  assign n13485 = n1266 & ~n13484 ;
  assign n13486 = x101 | n2373 ;
  assign n13487 = n6218 | n7187 ;
  assign n13488 = n4456 & n6262 ;
  assign n13489 = n4575 & n13488 ;
  assign n13490 = x198 & ~n1694 ;
  assign n13491 = n13489 & n13490 ;
  assign n13492 = n8437 | n13491 ;
  assign n13493 = n1646 & n6054 ;
  assign n13494 = n9181 & n11336 ;
  assign n13495 = n13494 ^ n1337 ^ 1'b0 ;
  assign n13496 = n3922 ^ n1360 ^ 1'b0 ;
  assign n13497 = ~n2281 & n13496 ;
  assign n13498 = n13497 ^ n7858 ^ 1'b0 ;
  assign n13499 = ~n3252 & n13498 ;
  assign n13500 = n2561 & n3060 ;
  assign n13501 = n8660 ^ n7275 ^ 1'b0 ;
  assign n13502 = n13191 ^ n6781 ^ n2718 ;
  assign n13503 = n13502 ^ x17 ^ 1'b0 ;
  assign n13504 = ~n8290 & n13503 ;
  assign n13505 = n13504 ^ n3583 ^ 1'b0 ;
  assign n13506 = n13505 ^ n9826 ^ 1'b0 ;
  assign n13507 = ~n4848 & n6674 ;
  assign n13508 = ~n12792 & n13507 ;
  assign n13509 = n934 & ~n8123 ;
  assign n13510 = ~n4751 & n13509 ;
  assign n13511 = ~n2079 & n13510 ;
  assign n13512 = n1736 & ~n6147 ;
  assign n13513 = ~n4671 & n13512 ;
  assign n13514 = n1600 & ~n13513 ;
  assign n13515 = ~n5660 & n13514 ;
  assign n13516 = n3265 & n6271 ;
  assign n13517 = n13516 ^ n5861 ^ 1'b0 ;
  assign n13519 = n4959 ^ n2465 ^ 1'b0 ;
  assign n13518 = n5781 & n7007 ;
  assign n13520 = n13519 ^ n13518 ^ 1'b0 ;
  assign n13521 = n6944 & ~n8207 ;
  assign n13522 = n13520 & n13521 ;
  assign n13523 = ~n13517 & n13522 ;
  assign n13526 = n2274 & ~n8774 ;
  assign n13527 = ~n2124 & n13526 ;
  assign n13528 = x21 & ~n13527 ;
  assign n13529 = n13527 & n13528 ;
  assign n13524 = n854 & ~n1295 ;
  assign n13525 = ~n12898 & n13524 ;
  assign n13530 = n13529 ^ n13525 ^ 1'b0 ;
  assign n13531 = n11120 ^ n378 ^ 1'b0 ;
  assign n13532 = n3057 & n13531 ;
  assign n13533 = n3390 ^ n726 ^ 1'b0 ;
  assign n13534 = ~n3880 & n13533 ;
  assign n13535 = n13534 ^ n7049 ^ 1'b0 ;
  assign n13536 = n552 | n6663 ;
  assign n13537 = n13536 ^ n752 ^ 1'b0 ;
  assign n13538 = n13537 ^ n452 ^ 1'b0 ;
  assign n13539 = n3956 & ~n5368 ;
  assign n13540 = n13539 ^ n4699 ^ 1'b0 ;
  assign n13541 = n2615 | n2941 ;
  assign n13542 = n13541 ^ n11233 ^ 1'b0 ;
  assign n13543 = n13542 ^ n12140 ^ 1'b0 ;
  assign n13544 = n9109 ^ n8507 ^ 1'b0 ;
  assign n13545 = n4497 ^ n3808 ^ 1'b0 ;
  assign n13546 = n13545 ^ n1831 ^ 1'b0 ;
  assign n13547 = n13237 & n13546 ;
  assign n13548 = n13547 ^ n12868 ^ 1'b0 ;
  assign n13549 = n13043 ^ n5810 ^ 1'b0 ;
  assign n13550 = n7582 | n13549 ;
  assign n13551 = n2303 & ~n13550 ;
  assign n13552 = n1035 & n7779 ;
  assign n13553 = n12467 & n13552 ;
  assign n13554 = n6640 & ~n9455 ;
  assign n13555 = n12912 ^ n8363 ^ n7391 ;
  assign n13556 = ~n1324 & n13555 ;
  assign n13557 = n13554 & n13556 ;
  assign n13558 = n13553 | n13557 ;
  assign n13559 = n13551 & ~n13558 ;
  assign n13560 = n1120 & ~n8843 ;
  assign n13561 = n7174 | n8356 ;
  assign n13562 = n12149 ^ n5240 ^ 1'b0 ;
  assign n13563 = n5759 | n7785 ;
  assign n13564 = n13563 ^ n3365 ^ 1'b0 ;
  assign n13565 = n13564 ^ n5804 ^ 1'b0 ;
  assign n13566 = n10151 | n13127 ;
  assign n13567 = n1698 & ~n13566 ;
  assign n13568 = n3266 ^ n978 ^ 1'b0 ;
  assign n13569 = n5066 ^ n4412 ^ 1'b0 ;
  assign n13570 = ~n4927 & n13569 ;
  assign n13571 = ~n5578 & n13570 ;
  assign n13572 = ~n13568 & n13571 ;
  assign n13573 = n7705 | n13572 ;
  assign n13574 = n13567 & ~n13573 ;
  assign n13575 = n7386 ^ n5982 ^ 1'b0 ;
  assign n13576 = n10407 & ~n13575 ;
  assign n13577 = n5120 & ~n9654 ;
  assign n13578 = n13577 ^ n8816 ^ 1'b0 ;
  assign n13579 = n1117 | n3371 ;
  assign n13580 = n13579 ^ n13352 ^ 1'b0 ;
  assign n13587 = ~n322 & n6972 ;
  assign n13588 = n13587 ^ n9256 ^ 1'b0 ;
  assign n13589 = ( n4745 & ~n7627 ) | ( n4745 & n13588 ) | ( ~n7627 & n13588 ) ;
  assign n13582 = n9706 ^ n667 ^ 1'b0 ;
  assign n13583 = ~n6032 & n13582 ;
  assign n13584 = n10178 ^ n1201 ^ 1'b0 ;
  assign n13585 = n13583 & ~n13584 ;
  assign n13581 = n1148 & n4816 ;
  assign n13586 = n13585 ^ n13581 ^ 1'b0 ;
  assign n13590 = n13589 ^ n13586 ^ 1'b0 ;
  assign n13591 = n7398 ^ n5012 ^ 1'b0 ;
  assign n13592 = ~n8179 & n13591 ;
  assign n13593 = n824 ^ n428 ^ 1'b0 ;
  assign n13594 = n13592 & n13593 ;
  assign n13595 = n13594 ^ n8540 ^ 1'b0 ;
  assign n13596 = x147 & ~n1169 ;
  assign n13597 = n4636 & n13596 ;
  assign n13598 = n2500 ^ n2314 ^ 1'b0 ;
  assign n13599 = n13598 ^ n5261 ^ 1'b0 ;
  assign n13600 = n5099 & ~n13599 ;
  assign n13601 = n13600 ^ n283 ^ 1'b0 ;
  assign n13602 = ~n1299 & n2223 ;
  assign n13603 = n13598 & ~n13602 ;
  assign n13604 = n12314 ^ n6905 ^ 1'b0 ;
  assign n13605 = n13603 | n13604 ;
  assign n13606 = n13398 ^ n2753 ^ 1'b0 ;
  assign n13607 = x87 & n13606 ;
  assign n13608 = n13605 | n13607 ;
  assign n13609 = n9387 & ~n13608 ;
  assign n13610 = n11050 ^ n1738 ^ 1'b0 ;
  assign n13611 = n9406 | n10104 ;
  assign n13612 = n13611 ^ n13077 ^ 1'b0 ;
  assign n13613 = n9066 | n9682 ;
  assign n13614 = n1773 | n4065 ;
  assign n13615 = n6975 & n7744 ;
  assign n13616 = n13615 ^ n4889 ^ 1'b0 ;
  assign n13617 = n2107 ^ x234 ^ 1'b0 ;
  assign n13618 = n4949 & n13617 ;
  assign n13619 = n13618 ^ n1475 ^ 1'b0 ;
  assign n13620 = n6606 | n13619 ;
  assign n13621 = n13620 ^ n4376 ^ 1'b0 ;
  assign n13622 = n1082 | n1988 ;
  assign n13623 = n2117 & ~n13622 ;
  assign n13624 = x101 & ~n13623 ;
  assign n13625 = ~n13621 & n13624 ;
  assign n13626 = n2477 | n9276 ;
  assign n13627 = ~n7406 & n13626 ;
  assign n13628 = n3866 ^ n1066 ^ 1'b0 ;
  assign n13629 = n4901 | n13628 ;
  assign n13630 = n10495 & n10880 ;
  assign n13631 = n8374 ^ n7291 ^ 1'b0 ;
  assign n13632 = n13630 & n13631 ;
  assign n13633 = n13632 ^ n11640 ^ 1'b0 ;
  assign n13634 = n6268 ^ n4513 ^ 1'b0 ;
  assign n13635 = n263 & n13634 ;
  assign n13636 = n13635 ^ n3983 ^ 1'b0 ;
  assign n13637 = n11055 & ~n13636 ;
  assign n13638 = n13637 ^ n6893 ^ 1'b0 ;
  assign n13639 = n3274 | n11571 ;
  assign n13640 = n13156 & ~n13639 ;
  assign n13641 = n1424 & ~n8378 ;
  assign n13642 = n13640 | n13641 ;
  assign n13643 = n6461 ^ n6220 ^ 1'b0 ;
  assign n13644 = n12196 | n13643 ;
  assign n13645 = n8551 ^ n2370 ^ 1'b0 ;
  assign n13646 = ~n3436 & n5808 ;
  assign n13647 = ~n13645 & n13646 ;
  assign n13650 = n570 & n1511 ;
  assign n13651 = n13650 ^ n5569 ^ 1'b0 ;
  assign n13648 = n4170 | n6079 ;
  assign n13649 = n13648 ^ n481 ^ 1'b0 ;
  assign n13652 = n13651 ^ n13649 ^ 1'b0 ;
  assign n13653 = n13647 | n13652 ;
  assign n13654 = n1453 ^ n1258 ^ 1'b0 ;
  assign n13655 = n5074 & ~n6813 ;
  assign n13656 = n13655 ^ n2475 ^ 1'b0 ;
  assign n13657 = n3726 | n13656 ;
  assign n13658 = n7502 | n13657 ;
  assign n13659 = n13658 ^ n9803 ^ 1'b0 ;
  assign n13660 = n8565 ^ n4293 ^ 1'b0 ;
  assign n13661 = n1066 | n13660 ;
  assign n13662 = ~n8297 & n11120 ;
  assign n13663 = n13662 ^ n2250 ^ 1'b0 ;
  assign n13664 = n7775 & n8058 ;
  assign n13665 = n12065 & ~n13664 ;
  assign n13666 = n3252 | n12167 ;
  assign n13667 = n7527 & ~n13666 ;
  assign n13668 = n10316 & ~n10430 ;
  assign n13669 = n13668 ^ n2697 ^ 1'b0 ;
  assign n13670 = n9116 & ~n13669 ;
  assign n13671 = ~n1089 & n13670 ;
  assign n13672 = n2652 ^ n1525 ^ 1'b0 ;
  assign n13673 = n1464 & n13672 ;
  assign n13674 = n5014 & n13673 ;
  assign n13675 = n1354 & n13674 ;
  assign n13676 = ~n2125 & n13675 ;
  assign n13677 = ~n7395 & n11058 ;
  assign n13678 = ~n919 & n4400 ;
  assign n13679 = n1366 & n13678 ;
  assign n13680 = n937 | n13679 ;
  assign n13681 = n11621 | n13680 ;
  assign n13682 = n3323 | n6400 ;
  assign n13683 = n3323 & ~n13682 ;
  assign n13684 = n6954 & n13683 ;
  assign n13685 = n7900 & ~n13684 ;
  assign n13686 = ~n7900 & n13685 ;
  assign n13687 = n7051 & ~n8270 ;
  assign n13688 = n8270 & n13687 ;
  assign n13689 = n13686 | n13688 ;
  assign n13690 = n13686 & ~n13689 ;
  assign n13691 = n3032 ^ n1580 ^ 1'b0 ;
  assign n13692 = n6421 ^ x76 ^ 1'b0 ;
  assign n13693 = n13691 & ~n13692 ;
  assign n13694 = n11082 ^ n7079 ^ 1'b0 ;
  assign n13695 = n4291 & ~n5426 ;
  assign n13696 = n5373 & n13695 ;
  assign n13697 = n3879 | n13696 ;
  assign n13698 = n9153 & ~n13697 ;
  assign n13699 = n6900 | n13698 ;
  assign n13700 = n13699 ^ n1415 ^ 1'b0 ;
  assign n13701 = n2824 ^ n2586 ^ 1'b0 ;
  assign n13702 = n11982 & n13701 ;
  assign n13703 = ~n7836 & n13702 ;
  assign n13704 = n2052 ^ x146 ^ 1'b0 ;
  assign n13705 = n13704 ^ n1102 ^ 1'b0 ;
  assign n13706 = n1312 | n3896 ;
  assign n13707 = n13706 ^ n2208 ^ 1'b0 ;
  assign n13708 = n13707 ^ n2187 ^ 1'b0 ;
  assign n13709 = n9809 & n13708 ;
  assign n13710 = n12470 & n13709 ;
  assign n13711 = n5059 ^ x155 ^ 1'b0 ;
  assign n13712 = n13710 | n13711 ;
  assign n13713 = n2838 & n4954 ;
  assign n13714 = ~n1525 & n13713 ;
  assign n13715 = n1368 & ~n13714 ;
  assign n13723 = n5399 & ~n8373 ;
  assign n13716 = n6744 ^ n6516 ^ 1'b0 ;
  assign n13717 = n3171 & n13716 ;
  assign n13718 = n4385 & n13717 ;
  assign n13719 = n13718 ^ x249 ^ 1'b0 ;
  assign n13720 = n657 | n13719 ;
  assign n13721 = n5126 & ~n13720 ;
  assign n13722 = n13026 | n13721 ;
  assign n13724 = n13723 ^ n13722 ^ 1'b0 ;
  assign n13725 = n12813 ^ n2252 ^ 1'b0 ;
  assign n13726 = n805 | n2668 ;
  assign n13727 = n13726 ^ n7350 ^ 1'b0 ;
  assign n13728 = ~n1049 & n13727 ;
  assign n13729 = n13728 ^ n8713 ^ 1'b0 ;
  assign n13731 = n12064 ^ n2854 ^ 1'b0 ;
  assign n13732 = n13731 ^ n7624 ^ n5819 ;
  assign n13730 = ~n705 & n9711 ;
  assign n13733 = n13732 ^ n13730 ^ 1'b0 ;
  assign n13734 = n4905 ^ n648 ^ 1'b0 ;
  assign n13735 = ~n5305 & n13734 ;
  assign n13736 = x143 & ~n921 ;
  assign n13737 = n13736 ^ n1920 ^ 1'b0 ;
  assign n13738 = n12177 ^ n4935 ^ 1'b0 ;
  assign n13741 = n2089 & ~n3477 ;
  assign n13739 = n2782 & n9834 ;
  assign n13740 = n13739 ^ n8218 ^ 1'b0 ;
  assign n13742 = n13741 ^ n13740 ^ 1'b0 ;
  assign n13743 = n3074 & ~n10511 ;
  assign n13744 = n296 & n1819 ;
  assign n13745 = ~n7737 & n13744 ;
  assign n13746 = n8923 & n13745 ;
  assign n13747 = n2237 | n2340 ;
  assign n13748 = n2278 ^ n1613 ^ 1'b0 ;
  assign n13749 = n13748 ^ n8020 ^ 1'b0 ;
  assign n13750 = n4865 | n5564 ;
  assign n13751 = n2038 | n3198 ;
  assign n13752 = n2725 & ~n13751 ;
  assign n13753 = ( ~n472 & n1964 ) | ( ~n472 & n2877 ) | ( n1964 & n2877 ) ;
  assign n13760 = n4236 & n7020 ;
  assign n13761 = n13760 ^ n3847 ^ 1'b0 ;
  assign n13756 = ~n6550 & n7622 ;
  assign n13754 = x110 & ~n3132 ;
  assign n13755 = n13754 ^ n5754 ^ 1'b0 ;
  assign n13757 = n13756 ^ n13755 ^ 1'b0 ;
  assign n13758 = n9967 & n13757 ;
  assign n13759 = n13758 ^ n3300 ^ 1'b0 ;
  assign n13762 = n13761 ^ n13759 ^ 1'b0 ;
  assign n13763 = n13753 & ~n13762 ;
  assign n13764 = n8801 ^ n7876 ^ 1'b0 ;
  assign n13765 = n387 | n7155 ;
  assign n13766 = n13765 ^ n7361 ^ 1'b0 ;
  assign n13767 = ~n5567 & n13766 ;
  assign n13768 = n2951 & ~n3119 ;
  assign n13769 = n8908 ^ n8516 ^ 1'b0 ;
  assign n13770 = ~n13768 & n13769 ;
  assign n13771 = n10469 ^ n9410 ^ 1'b0 ;
  assign n13772 = n13771 ^ n13248 ^ 1'b0 ;
  assign n13773 = n10672 & n13772 ;
  assign n13774 = ~n7748 & n8513 ;
  assign n13775 = ~n8425 & n13774 ;
  assign n13783 = x214 & ~n8077 ;
  assign n13777 = n2207 ^ n1698 ^ 1'b0 ;
  assign n13778 = n4048 & n13777 ;
  assign n13779 = n397 ^ x37 ^ 1'b0 ;
  assign n13780 = n397 & ~n13779 ;
  assign n13781 = n13780 ^ n5742 ^ 1'b0 ;
  assign n13782 = n13778 & ~n13781 ;
  assign n13784 = n13783 ^ n13782 ^ 1'b0 ;
  assign n13776 = ~n546 & n579 ;
  assign n13785 = n13784 ^ n13776 ^ n3512 ;
  assign n13786 = n6479 ^ n2765 ^ 1'b0 ;
  assign n13787 = n6218 & n13786 ;
  assign n13788 = n13787 ^ n5447 ^ 1'b0 ;
  assign n13789 = n920 | n12716 ;
  assign n13790 = n3050 | n13789 ;
  assign n13791 = n13790 ^ n807 ^ 1'b0 ;
  assign n13793 = n4584 ^ n3539 ^ 1'b0 ;
  assign n13792 = x75 & n5332 ;
  assign n13794 = n13793 ^ n13792 ^ 1'b0 ;
  assign n13795 = n10759 | n13794 ;
  assign n13796 = n13795 ^ n11653 ^ 1'b0 ;
  assign n13797 = n628 | n3845 ;
  assign n13798 = n10136 & ~n13797 ;
  assign n13799 = n12167 | n13798 ;
  assign n13800 = n13268 | n13799 ;
  assign n13801 = ~n4695 & n8572 ;
  assign n13802 = n5920 ^ n5173 ^ 1'b0 ;
  assign n13803 = n12397 ^ n2558 ^ 1'b0 ;
  assign n13804 = ~n13403 & n13803 ;
  assign n13805 = n3397 & n11519 ;
  assign n13806 = n8161 ^ n5558 ^ 1'b0 ;
  assign n13807 = n7652 & n13806 ;
  assign n13808 = n6396 | n13807 ;
  assign n13809 = n13808 ^ n11508 ^ 1'b0 ;
  assign n13810 = n859 & ~n13809 ;
  assign n13811 = n7448 ^ n4199 ^ 1'b0 ;
  assign n13812 = ~n516 & n529 ;
  assign n13813 = n4831 & ~n13812 ;
  assign n13814 = n13811 | n13813 ;
  assign n13815 = n6058 & ~n7115 ;
  assign n13816 = n13815 ^ n12559 ^ 1'b0 ;
  assign n13817 = n11960 ^ n5129 ^ 1'b0 ;
  assign n13818 = ~n9896 & n13447 ;
  assign n13819 = n10936 ^ n2546 ^ 1'b0 ;
  assign n13820 = n10485 ^ n1746 ^ 1'b0 ;
  assign n13821 = n13819 & n13820 ;
  assign n13822 = n13401 ^ n5343 ^ n1385 ;
  assign n13823 = n12443 & n13822 ;
  assign n13824 = n7100 ^ n5978 ^ 1'b0 ;
  assign n13825 = n13700 & ~n13824 ;
  assign n13826 = n12337 ^ n10744 ^ 1'b0 ;
  assign n13827 = n1405 & n9741 ;
  assign n13828 = n9356 | n12691 ;
  assign n13829 = n1883 & ~n13828 ;
  assign n13830 = n13829 ^ n6288 ^ 1'b0 ;
  assign n13831 = n4727 | n4957 ;
  assign n13832 = n13831 ^ n4889 ^ 1'b0 ;
  assign n13833 = n13832 ^ n2515 ^ 1'b0 ;
  assign n13834 = n3462 | n4620 ;
  assign n13835 = n13833 & ~n13834 ;
  assign n13836 = n8504 ^ n2539 ^ 1'b0 ;
  assign n13837 = ~n1657 & n7039 ;
  assign n13838 = n7290 | n13837 ;
  assign n13839 = ( n6273 & n7726 ) | ( n6273 & n13838 ) | ( n7726 & n13838 ) ;
  assign n13840 = n3361 | n10623 ;
  assign n13841 = n994 & ~n8201 ;
  assign n13842 = n3045 & n13841 ;
  assign n13843 = n3597 ^ n642 ^ 1'b0 ;
  assign n13844 = ~x59 & n13843 ;
  assign n13845 = n1337 & ~n13844 ;
  assign n13846 = n5168 | n13245 ;
  assign n13847 = x216 & ~n1693 ;
  assign n13848 = n4425 & ~n6128 ;
  assign n13849 = n13848 ^ x160 ^ 1'b0 ;
  assign n13850 = n6760 & ~n13849 ;
  assign n13851 = n7703 & n13850 ;
  assign n13852 = n13847 & n13851 ;
  assign n13853 = n9399 & n13507 ;
  assign n13854 = n13852 & n13853 ;
  assign n13855 = ~n13489 & n13854 ;
  assign n13856 = n1549 ^ n392 ^ 1'b0 ;
  assign n13857 = n3645 & ~n7287 ;
  assign n13858 = n7741 ^ n4586 ^ 1'b0 ;
  assign n13859 = x168 & n8709 ;
  assign n13860 = n3176 | n11704 ;
  assign n13861 = n6100 & n8406 ;
  assign n13862 = n1096 & ~n5279 ;
  assign n13863 = n13862 ^ n7197 ^ 1'b0 ;
  assign n13864 = n7371 & ~n8412 ;
  assign n13865 = ~n13863 & n13864 ;
  assign n13866 = ~n3175 & n9149 ;
  assign n13867 = n9475 & n13866 ;
  assign n13868 = n11916 ^ n4791 ^ n2338 ;
  assign n13869 = n13868 ^ n6205 ^ 1'b0 ;
  assign n13870 = ~n13867 & n13869 ;
  assign n13871 = n6339 | n6966 ;
  assign n13872 = ~n434 & n1822 ;
  assign n13873 = ~n13871 & n13872 ;
  assign n13874 = n4358 | n13873 ;
  assign n13875 = n13874 ^ n1344 ^ 1'b0 ;
  assign n13876 = ~n4116 & n13875 ;
  assign n13877 = n7518 | n9069 ;
  assign n13878 = n9484 | n13542 ;
  assign n13879 = n13877 & n13878 ;
  assign n13880 = ~n1233 & n10310 ;
  assign n13881 = n13880 ^ n5940 ^ 1'b0 ;
  assign n13882 = n11788 ^ n6118 ^ 1'b0 ;
  assign n13891 = n1703 | n11394 ;
  assign n13892 = n6498 & ~n13891 ;
  assign n13887 = n2926 ^ n2497 ^ 1'b0 ;
  assign n13888 = n2180 | n4393 ;
  assign n13889 = n13888 ^ n10763 ^ 1'b0 ;
  assign n13890 = n13887 & ~n13889 ;
  assign n13883 = n5272 | n11567 ;
  assign n13884 = n11330 & ~n13883 ;
  assign n13885 = ~n7448 & n8219 ;
  assign n13886 = n13884 & n13885 ;
  assign n13893 = n13892 ^ n13890 ^ n13886 ;
  assign n13894 = n1419 & n5974 ;
  assign n13895 = n13894 ^ n4751 ^ 1'b0 ;
  assign n13896 = n13895 ^ n13830 ^ 1'b0 ;
  assign n13897 = n7202 | n12531 ;
  assign n13898 = n3297 | n13897 ;
  assign n13899 = n3045 ^ n921 ^ 1'b0 ;
  assign n13900 = n11625 ^ n1488 ^ 1'b0 ;
  assign n13901 = n2232 | n13900 ;
  assign n13902 = n13899 & ~n13901 ;
  assign n13903 = ~n1343 & n4721 ;
  assign n13904 = ~n10012 & n13903 ;
  assign n13905 = n12429 ^ n8300 ^ 1'b0 ;
  assign n13906 = n4009 | n13905 ;
  assign n13907 = n1658 & ~n13906 ;
  assign n13908 = n13904 | n13907 ;
  assign n13909 = n1506 | n13908 ;
  assign n13910 = ~n6473 & n12861 ;
  assign n13911 = n13910 ^ n1353 ^ 1'b0 ;
  assign n13912 = ~n5255 & n6281 ;
  assign n13913 = n4211 ^ n3413 ^ 1'b0 ;
  assign n13914 = ( ~n4903 & n8165 ) | ( ~n4903 & n8556 ) | ( n8165 & n8556 ) ;
  assign n13915 = n10972 ^ x232 ^ 1'b0 ;
  assign n13916 = ~n1356 & n13915 ;
  assign n13917 = ~n4753 & n13916 ;
  assign n13918 = n13917 ^ n1628 ^ 1'b0 ;
  assign n13919 = n13918 ^ x151 ^ 1'b0 ;
  assign n13920 = ~n10171 & n12296 ;
  assign n13921 = ~n11458 & n13920 ;
  assign n13922 = ~n1658 & n4500 ;
  assign n13923 = n13922 ^ n2496 ^ 1'b0 ;
  assign n13924 = n7215 & ~n7694 ;
  assign n13925 = ~n6974 & n9066 ;
  assign n13926 = n11442 ^ n1360 ^ 1'b0 ;
  assign n13929 = n4871 & ~n6106 ;
  assign n13927 = ~n3318 & n4806 ;
  assign n13928 = n13927 ^ x86 ^ 1'b0 ;
  assign n13930 = n13929 ^ n13928 ^ 1'b0 ;
  assign n13931 = n4006 | n13930 ;
  assign n13932 = x41 & ~n3095 ;
  assign n13933 = n13932 ^ n10086 ^ 1'b0 ;
  assign n13934 = n8187 ^ n6091 ^ 1'b0 ;
  assign n13935 = ~n3939 & n13934 ;
  assign n13936 = n13935 ^ n7874 ^ 1'b0 ;
  assign n13937 = n6809 & n11911 ;
  assign n13938 = ~n4326 & n13937 ;
  assign n13939 = n5681 & ~n9212 ;
  assign n13940 = n5445 ^ n1684 ^ 1'b0 ;
  assign n13941 = n13940 ^ n2998 ^ n1633 ;
  assign n13942 = ~n505 & n7471 ;
  assign n13943 = n13942 ^ n2402 ^ 1'b0 ;
  assign n13944 = ~n9550 & n13943 ;
  assign n13945 = n13944 ^ n3177 ^ 1'b0 ;
  assign n13946 = n2764 & ~n6127 ;
  assign n13947 = ~n3269 & n5481 ;
  assign n13948 = n13947 ^ n10580 ^ 1'b0 ;
  assign n13949 = n4920 & n13948 ;
  assign n13950 = ~n13946 & n13949 ;
  assign n13951 = n8211 | n8553 ;
  assign n13952 = n1105 & ~n10845 ;
  assign n13953 = n10674 & ~n11176 ;
  assign n13954 = ~n7339 & n9150 ;
  assign n13955 = ~n7280 & n13954 ;
  assign n13956 = n9930 & n13955 ;
  assign n13957 = n800 & n13956 ;
  assign n13958 = n13957 ^ n4716 ^ 1'b0 ;
  assign n13959 = n3175 ^ n2796 ^ 1'b0 ;
  assign n13960 = n4865 ^ n4075 ^ 1'b0 ;
  assign n13961 = n5495 & ~n13960 ;
  assign n13962 = n13959 & ~n13961 ;
  assign n13963 = n5060 & n9276 ;
  assign n13964 = n3957 & ~n4579 ;
  assign n13965 = n13964 ^ x66 ^ 1'b0 ;
  assign n13966 = n13965 ^ n5110 ^ 1'b0 ;
  assign n13967 = n1148 & n13966 ;
  assign n13968 = ~x59 & n8018 ;
  assign n13969 = n11932 | n13968 ;
  assign n13970 = n2939 | n13969 ;
  assign n13972 = ( x160 & n552 ) | ( x160 & ~n7692 ) | ( n552 & ~n7692 ) ;
  assign n13971 = n9240 & n11377 ;
  assign n13973 = n13972 ^ n13971 ^ 1'b0 ;
  assign n13974 = n5531 ^ n5338 ^ 1'b0 ;
  assign n13975 = n4671 & ~n13974 ;
  assign n13976 = n5082 & n13975 ;
  assign n13977 = n5988 | n6647 ;
  assign n13978 = n7448 & ~n13977 ;
  assign n13979 = n633 & ~n6698 ;
  assign n13980 = ~n2503 & n2633 ;
  assign n13981 = n3982 | n6790 ;
  assign n13983 = n4769 & n11640 ;
  assign n13982 = x59 & n6587 ;
  assign n13984 = n13983 ^ n13982 ^ 1'b0 ;
  assign n13985 = n13981 & n13984 ;
  assign n13987 = n8154 ^ n7540 ^ 1'b0 ;
  assign n13988 = ( n633 & ~n4923 ) | ( n633 & n13987 ) | ( ~n4923 & n13987 ) ;
  assign n13986 = n1010 & n12505 ;
  assign n13989 = n13988 ^ n13986 ^ 1'b0 ;
  assign n13990 = n12560 | n13989 ;
  assign n13991 = n6083 & ~n11796 ;
  assign n13992 = n4006 & n13991 ;
  assign n13993 = n9008 ^ n6110 ^ 1'b0 ;
  assign n13997 = n2145 | n6762 ;
  assign n13998 = n13997 ^ n2762 ^ 1'b0 ;
  assign n13994 = x185 & ~n7957 ;
  assign n13995 = n13994 ^ n7216 ^ 1'b0 ;
  assign n13996 = n5471 & n13995 ;
  assign n13999 = n13998 ^ n13996 ^ 1'b0 ;
  assign n14000 = n13993 & n13999 ;
  assign n14001 = n994 & ~n3166 ;
  assign n14002 = n2867 & ~n14001 ;
  assign n14003 = n14002 ^ n1494 ^ 1'b0 ;
  assign n14004 = n14000 & ~n14003 ;
  assign n14007 = n10541 ^ n6149 ^ n1635 ;
  assign n14005 = ~n859 & n6647 ;
  assign n14006 = ~n7347 & n14005 ;
  assign n14008 = n14007 ^ n14006 ^ 1'b0 ;
  assign n14009 = n3118 & n8570 ;
  assign n14010 = n14009 ^ x21 ^ 1'b0 ;
  assign n14011 = n6401 & ~n14010 ;
  assign n14012 = n6065 & n9539 ;
  assign n14013 = n14012 ^ n4152 ^ 1'b0 ;
  assign n14014 = n14013 ^ n1840 ^ 1'b0 ;
  assign n14015 = n7559 | n14014 ;
  assign n14016 = n13409 ^ n1159 ^ 1'b0 ;
  assign n14017 = n2150 & n14016 ;
  assign n14022 = n2394 & ~n4053 ;
  assign n14023 = ~n9339 & n14022 ;
  assign n14018 = n3721 & ~n4209 ;
  assign n14019 = ~n2579 & n14018 ;
  assign n14020 = n14019 ^ n625 ^ 1'b0 ;
  assign n14021 = ~n1221 & n14020 ;
  assign n14024 = n14023 ^ n14021 ^ 1'b0 ;
  assign n14025 = n14024 ^ n8738 ^ 1'b0 ;
  assign n14026 = x75 & n13514 ;
  assign n14027 = ~n9639 & n14026 ;
  assign n14029 = ~n1930 & n10153 ;
  assign n14028 = ~n12032 & n12503 ;
  assign n14030 = n14029 ^ n14028 ^ 1'b0 ;
  assign n14031 = n14027 & ~n14030 ;
  assign n14032 = n4178 & n5185 ;
  assign n14033 = ~n12296 & n14032 ;
  assign n14034 = n4657 & ~n5508 ;
  assign n14035 = ~n9681 & n14034 ;
  assign n14036 = n6842 & n14035 ;
  assign n14037 = n10460 & ~n11516 ;
  assign n14038 = ~n8875 & n14037 ;
  assign n14039 = ~n2510 & n12414 ;
  assign n14040 = n14039 ^ n6560 ^ 1'b0 ;
  assign n14041 = ~n3073 & n13145 ;
  assign n14042 = ~n1324 & n9065 ;
  assign n14043 = n2003 & n14042 ;
  assign n14044 = n4160 ^ n2274 ^ 1'b0 ;
  assign n14045 = n7383 | n14044 ;
  assign n14046 = n14045 ^ n1713 ^ 1'b0 ;
  assign n14047 = n8941 | n14046 ;
  assign n14048 = n3272 & n5968 ;
  assign n14049 = n14048 ^ n6469 ^ 1'b0 ;
  assign n14050 = n12138 ^ n8228 ^ 1'b0 ;
  assign n14051 = n14049 & ~n14050 ;
  assign n14052 = n1635 & n8693 ;
  assign n14053 = ~n1622 & n14052 ;
  assign n14054 = n12818 | n14053 ;
  assign n14055 = n13453 & ~n14054 ;
  assign n14056 = n2633 ^ n1738 ^ 1'b0 ;
  assign n14057 = n11034 & n14056 ;
  assign n14058 = n14057 ^ n6012 ^ 1'b0 ;
  assign n14059 = n1326 | n5189 ;
  assign n14060 = n3485 | n14059 ;
  assign n14061 = n14060 ^ n8179 ^ 1'b0 ;
  assign n14062 = n1740 & n6009 ;
  assign n14063 = n14062 ^ n3027 ^ 1'b0 ;
  assign n14064 = n267 & n3702 ;
  assign n14065 = n11678 & n14064 ;
  assign n14071 = n6416 ^ n6279 ^ n5052 ;
  assign n14070 = n2302 | n4118 ;
  assign n14072 = n14071 ^ n14070 ^ 1'b0 ;
  assign n14066 = ( n1234 & n2496 ) | ( n1234 & n3100 ) | ( n2496 & n3100 ) ;
  assign n14067 = n2578 | n14066 ;
  assign n14068 = n14067 ^ n2027 ^ 1'b0 ;
  assign n14069 = n14068 ^ n8043 ^ 1'b0 ;
  assign n14073 = n14072 ^ n14069 ^ n3073 ;
  assign n14074 = ( ~x218 & n4986 ) | ( ~x218 & n14073 ) | ( n4986 & n14073 ) ;
  assign n14075 = n11001 & n13307 ;
  assign n14076 = n14075 ^ n7208 ^ 1'b0 ;
  assign n14077 = n14076 ^ n10210 ^ 1'b0 ;
  assign n14080 = ( n2866 & n9168 ) | ( n2866 & ~n13721 ) | ( n9168 & ~n13721 ) ;
  assign n14078 = n6606 & ~n8200 ;
  assign n14079 = n1683 | n14078 ;
  assign n14081 = n14080 ^ n14079 ^ 1'b0 ;
  assign n14082 = n4811 | n5851 ;
  assign n14083 = ~n9373 & n14082 ;
  assign n14084 = n14083 ^ n7892 ^ 1'b0 ;
  assign n14087 = ~n463 & n1429 ;
  assign n14088 = n10811 ^ n7569 ^ 1'b0 ;
  assign n14089 = ~n14087 & n14088 ;
  assign n14085 = n5617 & n5925 ;
  assign n14086 = n4734 | n14085 ;
  assign n14090 = n14089 ^ n14086 ^ 1'b0 ;
  assign n14091 = ~n2891 & n12792 ;
  assign n14092 = n4502 ^ n1690 ^ 1'b0 ;
  assign n14093 = n2973 & ~n14092 ;
  assign n14094 = ~n7814 & n14093 ;
  assign n14095 = x31 & n14094 ;
  assign n14096 = n11945 ^ n3577 ^ 1'b0 ;
  assign n14097 = ~n10070 & n14096 ;
  assign n14098 = ~n3040 & n14097 ;
  assign n14099 = n14095 & n14098 ;
  assign n14100 = n9201 ^ n2454 ^ 1'b0 ;
  assign n14101 = ~n4940 & n14100 ;
  assign n14102 = n2909 & n3901 ;
  assign n14103 = n1070 & n14102 ;
  assign n14104 = ~n2786 & n6747 ;
  assign n14105 = n14104 ^ n562 ^ 1'b0 ;
  assign n14106 = n2239 ^ n1909 ^ 1'b0 ;
  assign n14107 = n7064 | n14106 ;
  assign n14108 = n14106 & ~n14107 ;
  assign n14109 = n8079 & ~n14108 ;
  assign n14110 = n5607 & n14109 ;
  assign n14111 = n644 & n2755 ;
  assign n14112 = n6657 & n14111 ;
  assign n14113 = ~n2568 & n10152 ;
  assign n14114 = n4831 | n14113 ;
  assign n14116 = n1414 | n1757 ;
  assign n14115 = ~n8358 & n12239 ;
  assign n14117 = n14116 ^ n14115 ^ 1'b0 ;
  assign n14118 = ~n317 & n12535 ;
  assign n14119 = ~n13194 & n14118 ;
  assign n14120 = ~n703 & n6716 ;
  assign n14121 = n14120 ^ n415 ^ 1'b0 ;
  assign n14122 = n5908 ^ n1957 ^ 1'b0 ;
  assign n14123 = n2796 & ~n4301 ;
  assign n14124 = ( n1632 & n12667 ) | ( n1632 & n14123 ) | ( n12667 & n14123 ) ;
  assign n14125 = ~n3463 & n14124 ;
  assign n14126 = n4532 | n6979 ;
  assign n14127 = x188 | n14126 ;
  assign n14128 = n14127 ^ n7308 ^ 1'b0 ;
  assign n14129 = n11695 ^ n2725 ^ 1'b0 ;
  assign n14130 = n8392 & n14129 ;
  assign n14131 = n9836 | n10166 ;
  assign n14132 = n5326 & ~n13761 ;
  assign n14133 = n2485 & ~n4720 ;
  assign n14134 = n12813 ^ n12768 ^ 1'b0 ;
  assign n14135 = n14133 & ~n14134 ;
  assign n14136 = n8764 ^ n1160 ^ 1'b0 ;
  assign n14137 = n7174 & ~n14136 ;
  assign n14139 = n9100 ^ n5877 ^ 1'b0 ;
  assign n14138 = ~x81 & n3800 ;
  assign n14140 = n14139 ^ n14138 ^ 1'b0 ;
  assign n14152 = n488 | n1709 ;
  assign n14153 = n1709 & ~n14152 ;
  assign n14143 = n265 & n710 ;
  assign n14144 = ~n710 & n14143 ;
  assign n14145 = n836 & n853 ;
  assign n14146 = n14144 & n14145 ;
  assign n14147 = n2818 & ~n14146 ;
  assign n14148 = n14146 & n14147 ;
  assign n14149 = n8722 & ~n14148 ;
  assign n14150 = n14148 & n14149 ;
  assign n14141 = n2357 & n7436 ;
  assign n14142 = ~n7436 & n14141 ;
  assign n14151 = n14150 ^ n14142 ^ 1'b0 ;
  assign n14154 = n14153 ^ n14151 ^ 1'b0 ;
  assign n14155 = n1405 | n14154 ;
  assign n14156 = n666 & ~n10430 ;
  assign n14157 = n1369 & n14156 ;
  assign n14158 = ~n421 & n14157 ;
  assign n14159 = n2764 | n14158 ;
  assign n14160 = x185 & n14159 ;
  assign n14161 = n14160 ^ n894 ^ 1'b0 ;
  assign n14162 = n11661 ^ n5489 ^ 1'b0 ;
  assign n14163 = n6435 & n14162 ;
  assign n14164 = ~n3232 & n14163 ;
  assign n14165 = n5105 ^ n607 ^ 1'b0 ;
  assign n14166 = n5056 | n14165 ;
  assign n14167 = n4616 & ~n14166 ;
  assign n14168 = n4420 & n14167 ;
  assign n14169 = n4772 & ~n14168 ;
  assign n14170 = n14169 ^ n4671 ^ 1'b0 ;
  assign n14171 = ~n2335 & n7639 ;
  assign n14172 = n5188 & ~n14171 ;
  assign n14173 = n14172 ^ n3239 ^ 1'b0 ;
  assign n14175 = n666 & ~n981 ;
  assign n14174 = n1130 | n1308 ;
  assign n14176 = n14175 ^ n14174 ^ 1'b0 ;
  assign n14177 = ~n4473 & n14176 ;
  assign n14178 = n1623 & ~n3448 ;
  assign n14179 = n1205 | n14178 ;
  assign n14180 = n9855 | n14179 ;
  assign n14181 = n1409 & ~n8753 ;
  assign n14182 = n12443 & n14181 ;
  assign n14183 = n1191 & ~n2304 ;
  assign n14184 = n14183 ^ n8619 ^ 1'b0 ;
  assign n14185 = ~n4925 & n6951 ;
  assign n14186 = ~n1353 & n3537 ;
  assign n14187 = ~n5284 & n14186 ;
  assign n14188 = n14187 ^ n10714 ^ 1'b0 ;
  assign n14189 = n866 & n14188 ;
  assign n14190 = ~n4825 & n14189 ;
  assign n14191 = n5788 ^ n930 ^ 1'b0 ;
  assign n14192 = ~n7124 & n8833 ;
  assign n14193 = n500 | n10516 ;
  assign n14194 = n3328 ^ n1608 ^ 1'b0 ;
  assign n14195 = ~n14193 & n14194 ;
  assign n14196 = n14195 ^ n6884 ^ 1'b0 ;
  assign n14197 = n6790 | n11797 ;
  assign n14198 = n1474 & ~n4584 ;
  assign n14199 = n5222 & n5830 ;
  assign n14200 = n14198 & n14199 ;
  assign n14201 = n14197 & n14200 ;
  assign n14202 = n666 & n6070 ;
  assign n14203 = n7910 & n8528 ;
  assign n14204 = n11655 & n14203 ;
  assign n14205 = n1832 & n5629 ;
  assign n14207 = n9302 & n13400 ;
  assign n14208 = ~n9981 & n14207 ;
  assign n14206 = n7785 ^ n3676 ^ 1'b0 ;
  assign n14209 = n14208 ^ n14206 ^ 1'b0 ;
  assign n14210 = n14205 & n14209 ;
  assign n14211 = ~n14204 & n14210 ;
  assign n14212 = n12257 ^ n331 ^ 1'b0 ;
  assign n14213 = x82 & n14212 ;
  assign n14214 = n6882 & ~n9651 ;
  assign n14215 = n2359 & n11063 ;
  assign n14216 = x37 & n14215 ;
  assign n14217 = n6228 & ~n12393 ;
  assign n14218 = n14217 ^ n3334 ^ 1'b0 ;
  assign n14219 = n1293 & n2521 ;
  assign n14220 = ( n11589 & n12221 ) | ( n11589 & ~n14219 ) | ( n12221 & ~n14219 ) ;
  assign n14221 = n6997 & ~n12215 ;
  assign n14222 = n14124 ^ n6382 ^ 1'b0 ;
  assign n14223 = n754 & n14222 ;
  assign n14224 = n1221 & ~n2409 ;
  assign n14225 = n3469 & ~n8954 ;
  assign n14226 = n5869 & ~n7305 ;
  assign n14227 = n14226 ^ n3057 ^ 1'b0 ;
  assign n14228 = n14225 & ~n14227 ;
  assign n14229 = n10131 & ~n10330 ;
  assign n14230 = n11325 & n14229 ;
  assign n14231 = n4116 & ~n9557 ;
  assign n14232 = n7709 & n9761 ;
  assign n14233 = ~n7808 & n14232 ;
  assign n14234 = ~n14231 & n14233 ;
  assign n14235 = n4483 ^ n418 ^ 1'b0 ;
  assign n14236 = n2366 | n14235 ;
  assign n14237 = n14236 ^ n11302 ^ 1'b0 ;
  assign n14238 = n7880 & ~n14237 ;
  assign n14239 = n13750 ^ n11857 ^ n10706 ;
  assign n14240 = n7020 ^ n4384 ^ 1'b0 ;
  assign n14241 = ~n876 & n5060 ;
  assign n14242 = n14241 ^ n6421 ^ 1'b0 ;
  assign n14243 = n14240 & n14242 ;
  assign n14244 = ( n1050 & n11859 ) | ( n1050 & n13696 ) | ( n11859 & n13696 ) ;
  assign n14245 = n6298 | n7077 ;
  assign n14246 = n2505 & n5701 ;
  assign n14247 = ~n6381 & n14246 ;
  assign n14248 = n8237 ^ n2124 ^ 1'b0 ;
  assign n14249 = n1324 & n12202 ;
  assign n14250 = n5110 | n14249 ;
  assign n14251 = n1903 & n5192 ;
  assign n14252 = n14251 ^ n7846 ^ 1'b0 ;
  assign n14253 = n1544 | n4425 ;
  assign n14254 = n1544 & ~n14253 ;
  assign n14255 = x143 & ~n901 ;
  assign n14256 = ~x143 & n14255 ;
  assign n14257 = n1114 & ~n14256 ;
  assign n14258 = n14254 & n14257 ;
  assign n14259 = n14258 ^ n5828 ^ 1'b0 ;
  assign n14260 = n14252 & ~n14259 ;
  assign n14261 = n9178 & n9397 ;
  assign n14262 = ~n3153 & n7879 ;
  assign n14263 = n14262 ^ n1803 ^ 1'b0 ;
  assign n14264 = n4242 ^ n772 ^ 1'b0 ;
  assign n14265 = ~n4005 & n14264 ;
  assign n14266 = n2370 & ~n2863 ;
  assign n14267 = ~n2370 & n14266 ;
  assign n14268 = n1450 & n14267 ;
  assign n14269 = n8592 | n14268 ;
  assign n14270 = n2213 | n14269 ;
  assign n14271 = n14125 ^ n8554 ^ 1'b0 ;
  assign n14272 = n4310 & n14271 ;
  assign n14273 = x219 & n3768 ;
  assign n14274 = n14273 ^ n4151 ^ n3459 ;
  assign n14275 = ~n7023 & n12513 ;
  assign n14276 = n7922 ^ n7661 ^ n3402 ;
  assign n14277 = n10579 | n14276 ;
  assign n14278 = n14277 ^ n5959 ^ 1'b0 ;
  assign n14279 = n6167 & ~n14278 ;
  assign n14280 = ~n7828 & n14279 ;
  assign n14281 = n12525 & n14280 ;
  assign n14282 = n12767 ^ n10514 ^ 1'b0 ;
  assign n14283 = n2275 & n14282 ;
  assign n14284 = n2910 & ~n12154 ;
  assign n14285 = x23 & n14284 ;
  assign n14286 = n5047 & ~n14285 ;
  assign n14287 = ~n866 & n14286 ;
  assign n14288 = n12062 ^ n9026 ^ 1'b0 ;
  assign n14289 = n7006 | n8242 ;
  assign n14290 = n2276 & n4434 ;
  assign n14291 = n9639 & ~n12500 ;
  assign n14292 = ~n10296 & n14291 ;
  assign n14293 = n2254 ^ n376 ^ 1'b0 ;
  assign n14294 = ~n4454 & n14293 ;
  assign n14295 = n4910 | n14294 ;
  assign n14296 = n8740 ^ n6290 ^ 1'b0 ;
  assign n14297 = n994 & ~n9942 ;
  assign n14298 = n14297 ^ n3565 ^ 1'b0 ;
  assign n14299 = n14298 ^ n12797 ^ 1'b0 ;
  assign n14300 = n13265 ^ n5168 ^ 1'b0 ;
  assign n14301 = n2630 ^ n1952 ^ 1'b0 ;
  assign n14302 = n7320 ^ n6507 ^ 1'b0 ;
  assign n14303 = n3199 & n9797 ;
  assign n14304 = n8897 & n14303 ;
  assign n14305 = n3672 & ~n11034 ;
  assign n14306 = n4834 ^ n3662 ^ 1'b0 ;
  assign n14307 = ~n1524 & n7529 ;
  assign n14308 = n974 & n14307 ;
  assign n14309 = n14308 ^ x86 ^ 1'b0 ;
  assign n14310 = n3963 | n5963 ;
  assign n14311 = n14310 ^ n13603 ^ 1'b0 ;
  assign n14312 = ~n7171 & n13243 ;
  assign n14313 = n14312 ^ n11173 ^ 1'b0 ;
  assign n14314 = n1707 & ~n9362 ;
  assign n14315 = n14314 ^ n7556 ^ 1'b0 ;
  assign n14316 = ~n1651 & n2423 ;
  assign n14317 = n7337 & n14316 ;
  assign n14318 = n14315 & n14317 ;
  assign n14319 = n8256 ^ n1198 ^ 1'b0 ;
  assign n14320 = n6170 ^ n1981 ^ 1'b0 ;
  assign n14321 = ( n1540 & n2825 ) | ( n1540 & n9406 ) | ( n2825 & n9406 ) ;
  assign n14322 = n5024 ^ n2926 ^ 1'b0 ;
  assign n14323 = ~n4101 & n14322 ;
  assign n14324 = n4936 & n14323 ;
  assign n14325 = n14324 ^ n7880 ^ 1'b0 ;
  assign n14326 = n8773 & n14325 ;
  assign n14327 = n9629 & n14326 ;
  assign n14328 = n4103 ^ n2404 ^ 1'b0 ;
  assign n14329 = n3655 & n14328 ;
  assign n14330 = n2633 & ~n12020 ;
  assign n14331 = n14330 ^ n10292 ^ 1'b0 ;
  assign n14332 = n866 & ~n4576 ;
  assign n14333 = n13833 & n14332 ;
  assign n14335 = n6238 ^ n6028 ^ 1'b0 ;
  assign n14334 = n559 & n2909 ;
  assign n14336 = n14335 ^ n14334 ^ n2289 ;
  assign n14337 = ~n2476 & n12120 ;
  assign n14338 = n14337 ^ n8754 ^ 1'b0 ;
  assign n14339 = n4159 & ~n9437 ;
  assign n14341 = n6276 ^ n3655 ^ n1245 ;
  assign n14342 = n14341 ^ n4600 ^ 1'b0 ;
  assign n14343 = n2932 & n14342 ;
  assign n14340 = n2166 & ~n8474 ;
  assign n14344 = n14343 ^ n14340 ^ 1'b0 ;
  assign n14345 = n8976 & ~n14344 ;
  assign n14346 = n13199 & n14345 ;
  assign n14348 = n1006 | n1139 ;
  assign n14349 = n7293 & ~n14348 ;
  assign n14347 = n8902 | n9781 ;
  assign n14350 = n14349 ^ n14347 ^ 1'b0 ;
  assign n14351 = ~n10986 & n14350 ;
  assign n14352 = n4552 ^ n4526 ^ 1'b0 ;
  assign n14353 = n9173 ^ n3754 ^ 1'b0 ;
  assign n14354 = n14353 ^ n5067 ^ 1'b0 ;
  assign n14355 = n6684 ^ n4569 ^ 1'b0 ;
  assign n14358 = n6513 & ~n7202 ;
  assign n14356 = n7130 ^ x79 ^ 1'b0 ;
  assign n14357 = n4058 | n14356 ;
  assign n14359 = n14358 ^ n14357 ^ 1'b0 ;
  assign n14360 = ~n12429 & n14359 ;
  assign n14361 = n14360 ^ n11439 ^ n5296 ;
  assign n14362 = n3996 ^ n2858 ^ 1'b0 ;
  assign n14363 = n14362 ^ n4730 ^ 1'b0 ;
  assign n14364 = ( ~n747 & n6172 ) | ( ~n747 & n6372 ) | ( n6172 & n6372 ) ;
  assign n14365 = ( n1239 & n2298 ) | ( n1239 & n4291 ) | ( n2298 & n4291 ) ;
  assign n14366 = n12431 & ~n14365 ;
  assign n14367 = n14365 & n14366 ;
  assign n14368 = n14364 & n14367 ;
  assign n14369 = n11829 & n14368 ;
  assign n14370 = ~n11829 & n14369 ;
  assign n14371 = n11394 ^ n1451 ^ 1'b0 ;
  assign n14372 = n6369 ^ n2162 ^ 1'b0 ;
  assign n14373 = n6409 & n14372 ;
  assign n14374 = n4648 ^ n1720 ^ 1'b0 ;
  assign n14375 = n2476 ^ n394 ^ 1'b0 ;
  assign n14376 = n14353 ^ n2437 ^ 1'b0 ;
  assign n14377 = n1974 | n5278 ;
  assign n14384 = n10723 ^ n8241 ^ 1'b0 ;
  assign n14385 = n7936 | n14384 ;
  assign n14386 = n14385 ^ n13538 ^ 1'b0 ;
  assign n14378 = n7378 | n8184 ;
  assign n14379 = n519 & ~n1559 ;
  assign n14380 = n14379 ^ n8458 ^ 1'b0 ;
  assign n14381 = n2526 & ~n14380 ;
  assign n14382 = n14381 ^ n10118 ^ n8397 ;
  assign n14383 = ~n14378 & n14382 ;
  assign n14387 = n14386 ^ n14383 ^ 1'b0 ;
  assign n14388 = n7988 ^ n7164 ^ 1'b0 ;
  assign n14389 = ~n5667 & n14388 ;
  assign n14390 = n2562 ^ n1368 ^ 1'b0 ;
  assign n14391 = n8287 & n14390 ;
  assign n14392 = n7934 ^ n4345 ^ n1447 ;
  assign n14393 = n6496 & n14392 ;
  assign n14399 = ~n836 & n2443 ;
  assign n14398 = ~n3580 & n14323 ;
  assign n14400 = n14399 ^ n14398 ^ 1'b0 ;
  assign n14401 = n6189 & n14400 ;
  assign n14394 = n1444 & ~n4708 ;
  assign n14395 = n14394 ^ n12200 ^ 1'b0 ;
  assign n14396 = n6879 | n14395 ;
  assign n14397 = n14396 ^ n1217 ^ 1'b0 ;
  assign n14402 = n14401 ^ n14397 ^ 1'b0 ;
  assign n14403 = n14393 & n14402 ;
  assign n14404 = n8198 & n13933 ;
  assign n14405 = n5660 & ~n7835 ;
  assign n14406 = n2761 ^ n285 ^ 1'b0 ;
  assign n14407 = n1594 | n7520 ;
  assign n14408 = ~n5282 & n14407 ;
  assign n14409 = n12571 & n14408 ;
  assign n14410 = n2789 & n9078 ;
  assign n14411 = n4914 | n7933 ;
  assign n14412 = n5506 & ~n14411 ;
  assign n14413 = n14412 ^ n1559 ^ 1'b0 ;
  assign n14414 = ~n14410 & n14413 ;
  assign n14415 = n14414 ^ n956 ^ 1'b0 ;
  assign n14416 = n9708 ^ n9090 ^ 1'b0 ;
  assign n14417 = ~n3456 & n14416 ;
  assign n14418 = n3789 & n6809 ;
  assign n14419 = n14418 ^ n6500 ^ 1'b0 ;
  assign n14420 = n1772 | n8201 ;
  assign n14421 = n14419 | n14420 ;
  assign n14422 = n6248 | n14421 ;
  assign n14423 = n13418 ^ n5843 ^ 1'b0 ;
  assign n14424 = n3064 | n14423 ;
  assign n14425 = n4186 & ~n14424 ;
  assign n14426 = n4009 | n14425 ;
  assign n14427 = ~n2208 & n6886 ;
  assign n14428 = n5412 & n14427 ;
  assign n14429 = n14428 ^ n13905 ^ 1'b0 ;
  assign n14430 = n7491 & n14429 ;
  assign n14431 = ~n14426 & n14430 ;
  assign n14432 = n10935 ^ n6986 ^ 1'b0 ;
  assign n14433 = ~n3805 & n8553 ;
  assign n14434 = ~n9883 & n14433 ;
  assign n14435 = ~n368 & n2789 ;
  assign n14436 = ~n279 & n4720 ;
  assign n14437 = ~n6762 & n14436 ;
  assign n14438 = n7628 & n14437 ;
  assign n14439 = n2227 & n4999 ;
  assign n14440 = n2185 & n14439 ;
  assign n14441 = n4693 & ~n14440 ;
  assign n14442 = n14438 & n14441 ;
  assign n14443 = n8543 | n14442 ;
  assign n14444 = n1285 | n2954 ;
  assign n14445 = x176 & ~n14444 ;
  assign n14446 = n14445 ^ n13928 ^ 1'b0 ;
  assign n14447 = n3257 & n9916 ;
  assign n14448 = n6798 ^ n407 ^ 1'b0 ;
  assign n14449 = n2235 | n14448 ;
  assign n14450 = ~n10637 & n14449 ;
  assign n14451 = n14450 ^ n8877 ^ 1'b0 ;
  assign n14452 = ~n3810 & n7239 ;
  assign n14453 = n6443 & ~n8187 ;
  assign n14454 = ~n14452 & n14453 ;
  assign n14455 = n8173 & ~n14132 ;
  assign n14456 = n14455 ^ n5806 ^ 1'b0 ;
  assign n14457 = ~n628 & n7973 ;
  assign n14458 = n2047 & n14457 ;
  assign n14459 = n14458 ^ n681 ^ 1'b0 ;
  assign n14460 = n4276 | n6768 ;
  assign n14461 = n14460 ^ n6357 ^ 1'b0 ;
  assign n14462 = n9376 & ~n14461 ;
  assign n14463 = n14462 ^ n6693 ^ 1'b0 ;
  assign n14464 = n12364 ^ n6905 ^ 1'b0 ;
  assign n14465 = n7494 ^ n2495 ^ 1'b0 ;
  assign n14466 = n12260 ^ n1684 ^ 1'b0 ;
  assign n14467 = n2891 & ~n7826 ;
  assign n14468 = n4138 | n4142 ;
  assign n14469 = n14467 & ~n14468 ;
  assign n14470 = n14469 ^ n2820 ^ 1'b0 ;
  assign n14471 = n2210 & ~n14470 ;
  assign n14472 = ~n4855 & n14471 ;
  assign n14473 = ( n2314 & ~n14466 ) | ( n2314 & n14472 ) | ( ~n14466 & n14472 ) ;
  assign n14474 = n9222 ^ n864 ^ 1'b0 ;
  assign n14475 = n13878 ^ n8704 ^ 1'b0 ;
  assign n14476 = n14474 | n14475 ;
  assign n14477 = n6704 ^ x37 ^ 1'b0 ;
  assign n14478 = n7611 ^ x155 ^ 1'b0 ;
  assign n14479 = n3776 | n14478 ;
  assign n14480 = n14477 | n14479 ;
  assign n14481 = n14480 ^ n5050 ^ 1'b0 ;
  assign n14482 = n11530 & ~n14481 ;
  assign n14483 = n1923 | n2208 ;
  assign n14484 = n2397 & n9655 ;
  assign n14485 = n614 & n14484 ;
  assign n14486 = n6385 | n14348 ;
  assign n14487 = n6993 & ~n14486 ;
  assign n14488 = n14487 ^ n4179 ^ 1'b0 ;
  assign n14489 = ~n694 & n4564 ;
  assign n14490 = n1305 & n14489 ;
  assign n14491 = n14490 ^ n10198 ^ 1'b0 ;
  assign n14492 = x93 & ~n4018 ;
  assign n14493 = n4760 & n14492 ;
  assign n14494 = n12608 ^ n1914 ^ 1'b0 ;
  assign n14495 = n4899 & n14494 ;
  assign n14496 = n14495 ^ n8138 ^ 1'b0 ;
  assign n14497 = n2190 ^ n778 ^ 1'b0 ;
  assign n14498 = n6861 ^ n3114 ^ 1'b0 ;
  assign n14499 = n14498 ^ n1906 ^ 1'b0 ;
  assign n14500 = n4395 & n14499 ;
  assign n14501 = n14500 ^ n3980 ^ 1'b0 ;
  assign n14502 = n14501 ^ n6905 ^ n633 ;
  assign n14503 = n3491 ^ n2367 ^ 1'b0 ;
  assign n14504 = ~n3545 & n14503 ;
  assign n14505 = n4719 & n12494 ;
  assign n14506 = ~n6977 & n14505 ;
  assign n14507 = n14504 & n14506 ;
  assign n14508 = n5012 & ~n8957 ;
  assign n14509 = ~n5351 & n14508 ;
  assign n14510 = n12843 ^ n9971 ^ 1'b0 ;
  assign n14511 = ~n3803 & n14510 ;
  assign n14512 = n5830 & ~n6661 ;
  assign n14513 = ~n4065 & n14512 ;
  assign n14514 = n988 | n3003 ;
  assign n14515 = n14514 ^ n3454 ^ 1'b0 ;
  assign n14516 = ( ~n1426 & n14513 ) | ( ~n1426 & n14515 ) | ( n14513 & n14515 ) ;
  assign n14517 = n2848 & ~n14516 ;
  assign n14518 = ~x22 & n14517 ;
  assign n14519 = n13492 ^ n9418 ^ 1'b0 ;
  assign n14520 = n3331 & ~n7069 ;
  assign n14521 = ~n2809 & n8001 ;
  assign n14522 = n1787 | n14521 ;
  assign n14523 = ~n2097 & n2652 ;
  assign n14524 = n12754 ^ n2075 ^ n373 ;
  assign n14525 = ~n11541 & n14524 ;
  assign n14526 = n2895 & ~n14525 ;
  assign n14527 = n8129 ^ n5435 ^ 1'b0 ;
  assign n14528 = n4545 ^ n2600 ^ 1'b0 ;
  assign n14529 = ~n14527 & n14528 ;
  assign n14530 = ( n8594 & ~n11400 ) | ( n8594 & n12291 ) | ( ~n11400 & n12291 ) ;
  assign n14531 = n5845 & n9385 ;
  assign n14532 = n10464 | n13034 ;
  assign n14533 = n8442 & ~n11744 ;
  assign n14534 = n14533 ^ n4297 ^ 1'b0 ;
  assign n14535 = ~n3172 & n8923 ;
  assign n14536 = n10948 | n12990 ;
  assign n14537 = n1535 | n7335 ;
  assign n14538 = n3869 & ~n14537 ;
  assign n14539 = n14538 ^ n11774 ^ 1'b0 ;
  assign n14540 = x237 & ~n3565 ;
  assign n14541 = ~n7032 & n14540 ;
  assign n14542 = n5521 | n8532 ;
  assign n14543 = n14541 & ~n14542 ;
  assign n14544 = n1233 ^ n545 ^ 1'b0 ;
  assign n14545 = x100 | n14544 ;
  assign n14546 = n5714 | n7440 ;
  assign n14547 = ~n971 & n14546 ;
  assign n14548 = ~n6693 & n7880 ;
  assign n14549 = n14548 ^ n3793 ^ 1'b0 ;
  assign n14550 = ~n1124 & n6399 ;
  assign n14551 = n14550 ^ n8894 ^ n3224 ;
  assign n14552 = n9168 & ~n12775 ;
  assign n14553 = ~n14551 & n14552 ;
  assign n14554 = n10974 ^ n1549 ^ 1'b0 ;
  assign n14555 = ~n320 & n2968 ;
  assign n14556 = ~n1850 & n14555 ;
  assign n14557 = n6008 | n13507 ;
  assign n14558 = n4193 & ~n8035 ;
  assign n14559 = n13325 & n14558 ;
  assign n14560 = n10669 ^ n3432 ^ 1'b0 ;
  assign n14561 = n12911 ^ n887 ^ 1'b0 ;
  assign n14562 = n7306 | n14561 ;
  assign n14563 = n10689 ^ n4072 ^ 1'b0 ;
  assign n14564 = n4213 & n8613 ;
  assign n14565 = n4536 & n14564 ;
  assign n14566 = ~n2207 & n10607 ;
  assign n14567 = n14566 ^ n7200 ^ 1'b0 ;
  assign n14568 = n6696 & ~n7757 ;
  assign n14569 = n14568 ^ n2968 ^ 1'b0 ;
  assign n14570 = x95 & n14569 ;
  assign n14573 = n4161 ^ n3548 ^ 1'b0 ;
  assign n14571 = ~n1667 & n4741 ;
  assign n14572 = n14571 ^ x141 ^ 1'b0 ;
  assign n14574 = n14573 ^ n14572 ^ n3616 ;
  assign n14575 = x220 | n14574 ;
  assign n14576 = ( ~n1190 & n14570 ) | ( ~n1190 & n14575 ) | ( n14570 & n14575 ) ;
  assign n14577 = n6038 ^ n4767 ^ 1'b0 ;
  assign n14578 = n4412 & ~n14577 ;
  assign n14579 = x25 & ~n9038 ;
  assign n14580 = ~n14578 & n14579 ;
  assign n14581 = n1766 | n14580 ;
  assign n14582 = n7276 ^ n2469 ^ 1'b0 ;
  assign n14583 = n2418 & ~n14582 ;
  assign n14584 = n14583 ^ n3484 ^ 1'b0 ;
  assign n14585 = n14584 ^ n2368 ^ 1'b0 ;
  assign n14586 = n9493 & n14585 ;
  assign n14587 = ( n1450 & n4703 ) | ( n1450 & ~n14586 ) | ( n4703 & ~n14586 ) ;
  assign n14589 = ~n557 & n3533 ;
  assign n14590 = n14589 ^ n2704 ^ 1'b0 ;
  assign n14588 = n482 & n8706 ;
  assign n14591 = n14590 ^ n14588 ^ 1'b0 ;
  assign n14592 = n14591 ^ n1415 ^ 1'b0 ;
  assign n14593 = n9312 & ~n10637 ;
  assign n14594 = n1571 & n14013 ;
  assign n14595 = n672 & ~n7709 ;
  assign n14597 = n2328 & ~n3336 ;
  assign n14598 = n14597 ^ n3536 ^ 1'b0 ;
  assign n14596 = n1611 | n3022 ;
  assign n14599 = n14598 ^ n14596 ^ 1'b0 ;
  assign n14600 = n7884 | n14599 ;
  assign n14603 = n840 | n3963 ;
  assign n14604 = n14603 ^ n2700 ^ 1'b0 ;
  assign n14605 = n14604 ^ n4655 ^ 1'b0 ;
  assign n14601 = n11630 ^ n4304 ^ 1'b0 ;
  assign n14602 = n5844 & ~n14601 ;
  assign n14606 = n14605 ^ n14602 ^ 1'b0 ;
  assign n14607 = ~n1337 & n11206 ;
  assign n14608 = n14607 ^ n2283 ^ 1'b0 ;
  assign n14609 = n1124 | n14608 ;
  assign n14610 = n2431 & n7321 ;
  assign n14611 = n14610 ^ n5286 ^ 1'b0 ;
  assign n14612 = n12380 & n14611 ;
  assign n14613 = n2572 ^ n1596 ^ 1'b0 ;
  assign n14614 = n294 | n715 ;
  assign n14615 = n715 & ~n14614 ;
  assign n14616 = n2035 & ~n14615 ;
  assign n14617 = ~n2035 & n14616 ;
  assign n14618 = n778 & ~n14617 ;
  assign n14619 = n14617 & n14618 ;
  assign n14620 = n2218 & n8049 ;
  assign n14621 = n14619 & n14620 ;
  assign n14622 = ~n1474 & n3280 ;
  assign n14623 = ~n3280 & n14622 ;
  assign n14624 = n2037 | n14623 ;
  assign n14625 = n14623 & ~n14624 ;
  assign n14626 = n502 & ~n14625 ;
  assign n14627 = n14621 & n14626 ;
  assign n14628 = ~n7284 & n11514 ;
  assign n14629 = n6444 & n10316 ;
  assign n14630 = n2599 & n4414 ;
  assign n14631 = n1286 & ~n14630 ;
  assign n14632 = ~n14629 & n14631 ;
  assign n14633 = n1443 | n2787 ;
  assign n14634 = n14633 ^ x109 ^ 1'b0 ;
  assign n14635 = n12185 & ~n14634 ;
  assign n14636 = n6059 & ~n14635 ;
  assign n14637 = n14636 ^ n13918 ^ 1'b0 ;
  assign n14638 = n11988 ^ n8553 ^ 1'b0 ;
  assign n14639 = ~n13717 & n14638 ;
  assign n14640 = n14639 ^ n8089 ^ 1'b0 ;
  assign n14641 = n4745 & n14640 ;
  assign n14642 = n463 & n1826 ;
  assign n14643 = n14642 ^ n5650 ^ 1'b0 ;
  assign n14644 = n2733 | n9663 ;
  assign n14645 = n14643 | n14644 ;
  assign n14646 = n6162 ^ n4772 ^ 1'b0 ;
  assign n14647 = n1198 | n14646 ;
  assign n14648 = n14647 ^ n3337 ^ 1'b0 ;
  assign n14649 = n2954 | n10603 ;
  assign n14650 = n6173 & n6420 ;
  assign n14651 = n10500 ^ n5540 ^ 1'b0 ;
  assign n14652 = n7845 | n14651 ;
  assign n14653 = n4006 ^ n1537 ^ 1'b0 ;
  assign n14654 = ~n6900 & n14653 ;
  assign n14655 = ~n14652 & n14654 ;
  assign n14656 = ~n6228 & n14655 ;
  assign n14657 = ( n4172 & n5272 ) | ( n4172 & n14074 ) | ( n5272 & n14074 ) ;
  assign n14658 = n1801 & ~n3749 ;
  assign n14659 = ~n4475 & n14658 ;
  assign n14660 = n6769 ^ n3567 ^ 1'b0 ;
  assign n14661 = n13832 ^ n8657 ^ 1'b0 ;
  assign n14662 = n14660 & n14661 ;
  assign n14663 = n8656 & ~n9787 ;
  assign n14664 = n14663 ^ n9000 ^ 1'b0 ;
  assign n14665 = n9114 & ~n11226 ;
  assign n14666 = ~n1195 & n14665 ;
  assign n14667 = n14664 | n14666 ;
  assign n14668 = n736 | n2665 ;
  assign n14669 = n14668 ^ n7061 ^ n6539 ;
  assign n14670 = ( x84 & x180 ) | ( x84 & n10234 ) | ( x180 & n10234 ) ;
  assign n14671 = n5413 & n9764 ;
  assign n14672 = n14671 ^ n2503 ^ 1'b0 ;
  assign n14673 = n6988 ^ n1226 ^ 1'b0 ;
  assign n14674 = n4065 & n14673 ;
  assign n14675 = n14674 ^ n7715 ^ 1'b0 ;
  assign n14676 = ~n7040 & n14675 ;
  assign n14677 = x86 & n4753 ;
  assign n14678 = n8699 & n14677 ;
  assign n14681 = ~x186 & n13029 ;
  assign n14679 = n13780 & ~n14666 ;
  assign n14680 = n14679 ^ n1380 ^ 1'b0 ;
  assign n14682 = n14681 ^ n14680 ^ n3373 ;
  assign n14683 = n1243 | n9880 ;
  assign n14684 = n1518 ^ n1492 ^ 1'b0 ;
  assign n14685 = n365 & ~n14684 ;
  assign n14686 = n1643 ^ x11 ^ 1'b0 ;
  assign n14687 = n14685 & n14686 ;
  assign n14688 = ~n5370 & n14687 ;
  assign n14689 = n14688 ^ n4838 ^ 1'b0 ;
  assign n14690 = n14689 ^ n1360 ^ 1'b0 ;
  assign n14691 = n345 & ~n10465 ;
  assign n14692 = n3086 | n6464 ;
  assign n14693 = n14692 ^ n2714 ^ 1'b0 ;
  assign n14694 = n14693 ^ n6003 ^ 1'b0 ;
  assign n14695 = n14694 ^ n7528 ^ 1'b0 ;
  assign n14696 = n913 & n14695 ;
  assign n14697 = n4631 | n14696 ;
  assign n14698 = n14697 ^ n2302 ^ 1'b0 ;
  assign n14699 = n4295 & n6468 ;
  assign n14700 = n14699 ^ n14187 ^ 1'b0 ;
  assign n14701 = n1818 & n3390 ;
  assign n14702 = n14701 ^ n2082 ^ 1'b0 ;
  assign n14703 = n1468 & ~n14702 ;
  assign n14704 = n2899 & n14703 ;
  assign n14705 = n14704 ^ x148 ^ 1'b0 ;
  assign n14706 = ~n6834 & n10770 ;
  assign n14707 = ~n6627 & n14706 ;
  assign n14708 = ~n9796 & n14707 ;
  assign n14709 = n5955 & ~n13752 ;
  assign n14710 = n12863 & n14709 ;
  assign n14711 = n9260 & ~n10004 ;
  assign n14716 = ~n543 & n6287 ;
  assign n14717 = n2644 & n14716 ;
  assign n14713 = n3863 & n6256 ;
  assign n14714 = ~n1815 & n14713 ;
  assign n14712 = ~n1785 & n12803 ;
  assign n14715 = n14714 ^ n14712 ^ 1'b0 ;
  assign n14718 = n14717 ^ n14715 ^ 1'b0 ;
  assign n14719 = x219 & ~n327 ;
  assign n14720 = ~x219 & n14719 ;
  assign n14721 = ~n543 & n14720 ;
  assign n14722 = x59 ^ x30 ^ 1'b0 ;
  assign n14723 = n14721 & n14722 ;
  assign n14724 = n481 & ~n14723 ;
  assign n14725 = n4241 & n5468 ;
  assign n14726 = ~n5468 & n14725 ;
  assign n14727 = n1594 | n14726 ;
  assign n14728 = n1571 | n1691 ;
  assign n14729 = n1571 & ~n14728 ;
  assign n14730 = n877 | n14729 ;
  assign n14731 = n14729 & ~n14730 ;
  assign n14732 = n6735 & ~n14731 ;
  assign n14733 = n14731 & n14732 ;
  assign n14734 = n14727 | n14733 ;
  assign n14735 = n14727 & ~n14734 ;
  assign n14736 = n4611 | n14735 ;
  assign n14737 = n4611 & ~n14736 ;
  assign n14748 = ~n661 & n1252 ;
  assign n14749 = ~n1252 & n14748 ;
  assign n14750 = x136 & n14749 ;
  assign n14751 = n14750 ^ n651 ^ 1'b0 ;
  assign n14738 = x246 & ~n789 ;
  assign n14739 = n789 & n14738 ;
  assign n14740 = x123 & x194 ;
  assign n14741 = ~x194 & n14740 ;
  assign n14742 = n267 & n14741 ;
  assign n14743 = x232 & ~n14742 ;
  assign n14744 = ~n6706 & n14743 ;
  assign n14745 = n14739 & n14744 ;
  assign n14746 = n8614 | n8908 ;
  assign n14747 = n14745 & ~n14746 ;
  assign n14752 = n14751 ^ n14747 ^ 1'b0 ;
  assign n14753 = n14737 | n14752 ;
  assign n14754 = n14724 & ~n14753 ;
  assign n14755 = ~n2776 & n8153 ;
  assign n14756 = n11377 ^ n4215 ^ 1'b0 ;
  assign n14757 = n2825 | n11284 ;
  assign n14758 = n3581 & n14757 ;
  assign n14759 = n5021 | n9736 ;
  assign n14760 = n8689 & ~n14759 ;
  assign n14761 = ~n3750 & n12848 ;
  assign n14762 = n3750 & n14761 ;
  assign n14763 = n8507 | n10806 ;
  assign n14764 = n14763 ^ n6372 ^ 1'b0 ;
  assign n14771 = n8170 ^ n4143 ^ 1'b0 ;
  assign n14768 = n1941 ^ n1646 ^ 1'b0 ;
  assign n14765 = n8202 & ~n10346 ;
  assign n14766 = x98 & ~n14765 ;
  assign n14767 = n14766 ^ n3842 ^ 1'b0 ;
  assign n14769 = n14768 ^ n14767 ^ 1'b0 ;
  assign n14770 = n14769 ^ n5409 ^ 1'b0 ;
  assign n14772 = n14771 ^ n14770 ^ 1'b0 ;
  assign n14773 = n14764 & n14772 ;
  assign n14774 = n6934 ^ n4097 ^ 1'b0 ;
  assign n14775 = n5361 & ~n11999 ;
  assign n14776 = n6274 | n7259 ;
  assign n14777 = n14776 ^ n2877 ^ 1'b0 ;
  assign n14778 = ~n1896 & n10108 ;
  assign n14779 = n12440 ^ n4363 ^ 1'b0 ;
  assign n14780 = ~n6146 & n14779 ;
  assign n14781 = n14780 ^ n2798 ^ 1'b0 ;
  assign n14782 = ~n6134 & n14236 ;
  assign n14783 = n6036 ^ n2827 ^ 1'b0 ;
  assign n14784 = n11479 ^ n4968 ^ 1'b0 ;
  assign n14785 = n10957 ^ n8697 ^ 1'b0 ;
  assign n14786 = n14784 | n14785 ;
  assign n14787 = n2364 | n8644 ;
  assign n14788 = n905 & ~n14787 ;
  assign n14789 = ~n3770 & n13668 ;
  assign n14790 = n14789 ^ n10031 ^ 1'b0 ;
  assign n14791 = n9451 ^ n5961 ^ 1'b0 ;
  assign n14792 = n14790 & n14791 ;
  assign n14793 = ~n11042 & n11618 ;
  assign n14794 = ~n1760 & n14793 ;
  assign n14795 = n1383 & n14794 ;
  assign n14796 = ~n6276 & n14795 ;
  assign n14797 = n14796 ^ n7326 ^ 1'b0 ;
  assign n14798 = n3067 | n4466 ;
  assign n14799 = n14798 ^ n6997 ^ 1'b0 ;
  assign n14800 = x69 & ~n4715 ;
  assign n14801 = n14800 ^ n10398 ^ 1'b0 ;
  assign n14802 = n3760 | n14801 ;
  assign n14803 = n10564 ^ n1291 ^ 1'b0 ;
  assign n14805 = x186 & n1710 ;
  assign n14806 = n4656 & n14805 ;
  assign n14804 = ~n1799 & n10105 ;
  assign n14807 = n14806 ^ n14804 ^ 1'b0 ;
  assign n14808 = n14807 ^ n11187 ^ 1'b0 ;
  assign n14809 = n1536 & n1793 ;
  assign n14810 = n8378 ^ n5076 ^ 1'b0 ;
  assign n14811 = n5068 & ~n7026 ;
  assign n14812 = n14811 ^ n2521 ^ 1'b0 ;
  assign n14813 = n14812 ^ n7077 ^ 1'b0 ;
  assign n14814 = ~n3880 & n10617 ;
  assign n14815 = ~n14813 & n14814 ;
  assign n14816 = n9757 & n12355 ;
  assign n14817 = n14816 ^ n12977 ^ 1'b0 ;
  assign n14818 = n7255 ^ n5984 ^ 1'b0 ;
  assign n14819 = n14818 ^ n5194 ^ 1'b0 ;
  assign n14820 = n11105 ^ n1341 ^ 1'b0 ;
  assign n14821 = n12655 & n14820 ;
  assign n14822 = n2632 & ~n6786 ;
  assign n14823 = n4543 | n14822 ;
  assign n14824 = n11954 | n14823 ;
  assign n14825 = n14824 ^ n6271 ^ 1'b0 ;
  assign n14826 = n14825 ^ n8190 ^ n4128 ;
  assign n14827 = n7808 ^ n1594 ^ 1'b0 ;
  assign n14828 = n6281 | n14827 ;
  assign n14829 = n3601 & ~n9966 ;
  assign n14830 = n14829 ^ n5386 ^ 1'b0 ;
  assign n14831 = n4686 ^ n3191 ^ 1'b0 ;
  assign n14833 = n1807 & ~n2657 ;
  assign n14834 = ~n7637 & n14833 ;
  assign n14832 = ~n7359 & n7725 ;
  assign n14835 = n14834 ^ n14832 ^ 1'b0 ;
  assign n14836 = ~n14831 & n14835 ;
  assign n14837 = ~n14830 & n14836 ;
  assign n14838 = n11589 ^ n2581 ^ 1'b0 ;
  assign n14839 = n384 | n14838 ;
  assign n14845 = n2423 & n3641 ;
  assign n14840 = ~n2116 & n2848 ;
  assign n14841 = n14840 ^ n3776 ^ 1'b0 ;
  assign n14842 = ~n2776 & n4824 ;
  assign n14843 = n6499 | n14842 ;
  assign n14844 = n14841 | n14843 ;
  assign n14846 = n14845 ^ n14844 ^ 1'b0 ;
  assign n14847 = n1597 ^ x59 ^ 1'b0 ;
  assign n14851 = n2050 & n4181 ;
  assign n14852 = n14851 ^ n11479 ^ 1'b0 ;
  assign n14853 = n2261 & n14852 ;
  assign n14848 = ~x98 & n1531 ;
  assign n14849 = n3961 ^ n3180 ^ 1'b0 ;
  assign n14850 = n14848 & n14849 ;
  assign n14854 = n14853 ^ n14850 ^ 1'b0 ;
  assign n14855 = n6858 ^ n600 ^ 1'b0 ;
  assign n14856 = n3844 & n14855 ;
  assign n14857 = n11987 ^ n3634 ^ 1'b0 ;
  assign n14858 = n3713 & n14857 ;
  assign n14859 = n6587 ^ n2213 ^ 1'b0 ;
  assign n14860 = n12652 ^ n9797 ^ 1'b0 ;
  assign n14861 = n14859 | n14860 ;
  assign n14862 = ~n6274 & n12805 ;
  assign n14863 = n1461 & ~n6939 ;
  assign n14864 = n11037 ^ n10076 ^ 1'b0 ;
  assign n14865 = n13145 ^ x248 ^ 1'b0 ;
  assign n14866 = x77 & n14865 ;
  assign n14867 = ~n13143 & n13520 ;
  assign n14868 = ~n1447 & n13204 ;
  assign n14869 = ~n3300 & n14868 ;
  assign n14870 = n4959 & ~n14869 ;
  assign n14871 = n14870 ^ n6889 ^ 1'b0 ;
  assign n14872 = n1518 & ~n5481 ;
  assign n14873 = n14872 ^ n9563 ^ n2019 ;
  assign n14874 = n8294 ^ n3419 ^ 1'b0 ;
  assign n14875 = ~n13460 & n14874 ;
  assign n14876 = n1260 & ~n1923 ;
  assign n14877 = ~n7748 & n14876 ;
  assign n14878 = n14877 ^ n13870 ^ 1'b0 ;
  assign n14879 = n3920 | n4005 ;
  assign n14880 = ( n5026 & n7156 ) | ( n5026 & ~n14879 ) | ( n7156 & ~n14879 ) ;
  assign n14881 = n1919 | n5283 ;
  assign n14882 = n1704 ^ n1653 ^ 1'b0 ;
  assign n14883 = n14882 ^ n3910 ^ 1'b0 ;
  assign n14884 = n2152 | n6263 ;
  assign n14885 = n5163 & n7149 ;
  assign n14886 = n8443 & ~n11869 ;
  assign n14887 = ~n5269 & n14886 ;
  assign n14888 = n370 & n3053 ;
  assign n14890 = n3637 & ~n7155 ;
  assign n14891 = n14890 ^ n1841 ^ 1'b0 ;
  assign n14889 = n6428 ^ n3854 ^ 1'b0 ;
  assign n14892 = n14891 ^ n14889 ^ 1'b0 ;
  assign n14893 = ~n8377 & n12339 ;
  assign n14894 = n14893 ^ n2185 ^ 1'b0 ;
  assign n14895 = n1697 & ~n4395 ;
  assign n14896 = n3116 & ~n7058 ;
  assign n14897 = n14896 ^ n8187 ^ 1'b0 ;
  assign n14898 = n12974 ^ n9632 ^ 1'b0 ;
  assign n14899 = n9388 & ~n13108 ;
  assign n14900 = n14899 ^ n2731 ^ 1'b0 ;
  assign n14901 = n1339 | n1832 ;
  assign n14902 = n4664 ^ n4076 ^ 1'b0 ;
  assign n14903 = ~n6434 & n14902 ;
  assign n14904 = n2731 | n6432 ;
  assign n14905 = n14903 | n14904 ;
  assign n14906 = n11584 ^ n428 ^ 1'b0 ;
  assign n14907 = n597 | n14906 ;
  assign n14908 = n14082 | n14907 ;
  assign n14909 = n14557 & ~n14908 ;
  assign n14910 = ~n9186 & n14909 ;
  assign n14911 = n2331 & ~n11578 ;
  assign n14912 = n5999 & ~n7015 ;
  assign n14913 = n3740 & n14912 ;
  assign n14914 = n4536 & n13029 ;
  assign n14915 = n6002 & n14914 ;
  assign n14916 = n2755 & n7949 ;
  assign n14917 = n14916 ^ n7894 ^ 1'b0 ;
  assign n14918 = ~n8628 & n14917 ;
  assign n14919 = n10762 ^ n5163 ^ 1'b0 ;
  assign n14920 = n14919 ^ n5891 ^ 1'b0 ;
  assign n14921 = n14918 | n14920 ;
  assign n14922 = n7766 ^ n6461 ^ n1286 ;
  assign n14923 = n7613 & n14922 ;
  assign n14924 = n7674 & n10140 ;
  assign n14925 = ~n10005 & n12531 ;
  assign n14926 = n3670 & n7490 ;
  assign n14927 = n14926 ^ n9932 ^ 1'b0 ;
  assign n14928 = n492 & ~n3575 ;
  assign n14929 = x1 & n14928 ;
  assign n14930 = n14924 & ~n14929 ;
  assign n14931 = n5298 ^ n4631 ^ 1'b0 ;
  assign n14932 = n6735 | n14931 ;
  assign n14933 = n5031 & ~n14932 ;
  assign n14934 = n2106 | n7032 ;
  assign n14935 = n14934 ^ n7590 ^ 1'b0 ;
  assign n14936 = n6413 ^ n2946 ^ 1'b0 ;
  assign n14937 = n1396 & n14936 ;
  assign n14938 = ( x15 & n3248 ) | ( x15 & ~n8485 ) | ( n3248 & ~n8485 ) ;
  assign n14939 = ~n7768 & n14938 ;
  assign n14940 = ~n14937 & n14939 ;
  assign n14941 = ~n1488 & n14940 ;
  assign n14942 = n6727 | n12002 ;
  assign n14943 = n14942 ^ n1077 ^ 1'b0 ;
  assign n14944 = n7276 | n12691 ;
  assign n14945 = n2493 & ~n14944 ;
  assign n14946 = n9055 | n14945 ;
  assign n14947 = n7032 | n14946 ;
  assign n14948 = n1031 & ~n3346 ;
  assign n14949 = n313 & ~n14948 ;
  assign n14950 = n14949 ^ n12008 ^ n6247 ;
  assign n14951 = n1651 & n8878 ;
  assign n14952 = n9410 | n14951 ;
  assign n14953 = x129 | n4156 ;
  assign n14955 = n3182 | n11695 ;
  assign n14954 = n607 & ~n1059 ;
  assign n14956 = n14955 ^ n14954 ^ 1'b0 ;
  assign n14957 = ~n1169 & n4129 ;
  assign n14958 = n14957 ^ n1757 ^ n1212 ;
  assign n14959 = n14958 ^ n10555 ^ n4749 ;
  assign n14960 = n14956 & n14959 ;
  assign n14961 = n1564 | n13347 ;
  assign n14962 = ~n7170 & n14961 ;
  assign n14963 = n14962 ^ n5399 ^ 1'b0 ;
  assign n14964 = n1145 | n2609 ;
  assign n14965 = n14964 ^ n2228 ^ 1'b0 ;
  assign n14966 = n13793 ^ n9955 ^ 1'b0 ;
  assign n14967 = ~n14965 & n14966 ;
  assign n14968 = n8827 & n14967 ;
  assign n14969 = n1795 | n3678 ;
  assign n14971 = n3461 & n7115 ;
  assign n14970 = n5835 & ~n7493 ;
  assign n14972 = n14971 ^ n14970 ^ 1'b0 ;
  assign n14973 = n14818 ^ n3214 ^ 1'b0 ;
  assign n14974 = n5837 & ~n14973 ;
  assign n14975 = n2155 & n14545 ;
  assign n14976 = n13344 & n14975 ;
  assign n14977 = n14976 ^ n2737 ^ 1'b0 ;
  assign n14978 = n1715 & n10892 ;
  assign n14979 = n3123 & n8992 ;
  assign n14980 = ~n11431 & n14979 ;
  assign n14984 = n7833 ^ n6479 ^ 1'b0 ;
  assign n14985 = n8056 & n14984 ;
  assign n14986 = ~n7257 & n14985 ;
  assign n14981 = n1131 & n1459 ;
  assign n14982 = n14981 ^ n1178 ^ 1'b0 ;
  assign n14983 = n14157 | n14982 ;
  assign n14987 = n14986 ^ n14983 ^ 1'b0 ;
  assign n14990 = n4003 | n6605 ;
  assign n14991 = n14990 ^ n2415 ^ 1'b0 ;
  assign n14992 = n14991 ^ n4644 ^ n3111 ;
  assign n14993 = ~n8900 & n14992 ;
  assign n14988 = ~n3423 & n6997 ;
  assign n14989 = n7266 | n14988 ;
  assign n14994 = n14993 ^ n14989 ^ n4464 ;
  assign n14995 = n1799 & n4493 ;
  assign n14996 = n9193 ^ n3477 ^ 1'b0 ;
  assign n14997 = n14995 | n14996 ;
  assign n14998 = n3549 ^ x42 ^ 1'b0 ;
  assign n14999 = n14998 ^ n1358 ^ 1'b0 ;
  assign n15000 = n7668 & ~n13929 ;
  assign n15001 = n8253 ^ x127 ^ 1'b0 ;
  assign n15002 = n7136 | n15001 ;
  assign n15003 = n956 | n15002 ;
  assign n15004 = n8960 ^ n5613 ^ 1'b0 ;
  assign n15005 = n15003 | n15004 ;
  assign n15006 = n4021 | n6117 ;
  assign n15007 = n1939 & ~n15006 ;
  assign n15008 = n9717 ^ n9643 ^ 1'b0 ;
  assign n15009 = n12839 ^ n9368 ^ 1'b0 ;
  assign n15010 = n5091 ^ x191 ^ 1'b0 ;
  assign n15011 = n11063 & ~n15010 ;
  assign n15012 = n776 & n4331 ;
  assign n15013 = n840 & n15012 ;
  assign n15014 = n15013 ^ n11628 ^ n720 ;
  assign n15015 = n7456 ^ n644 ^ 1'b0 ;
  assign n15016 = n15014 | n15015 ;
  assign n15017 = n11356 ^ n5448 ^ 1'b0 ;
  assign n15018 = n3901 & n15017 ;
  assign n15019 = n573 | n15018 ;
  assign n15020 = n13397 ^ n5756 ^ 1'b0 ;
  assign n15021 = n15019 | n15020 ;
  assign n15022 = n3531 ^ n3076 ^ 1'b0 ;
  assign n15026 = x38 & x198 ;
  assign n15027 = n15026 ^ n2497 ^ 1'b0 ;
  assign n15023 = n2507 & n8408 ;
  assign n15024 = n15023 ^ n5091 ^ 1'b0 ;
  assign n15025 = n11469 & n15024 ;
  assign n15028 = n15027 ^ n15025 ^ n14433 ;
  assign n15029 = ~n2322 & n15028 ;
  assign n15030 = ~n15022 & n15029 ;
  assign n15031 = n666 & ~n2517 ;
  assign n15032 = n2632 & n11124 ;
  assign n15033 = ~n6797 & n15032 ;
  assign n15034 = x50 & n15033 ;
  assign n15035 = n15034 ^ n6801 ^ 1'b0 ;
  assign n15036 = n12288 ^ n8229 ^ 1'b0 ;
  assign n15037 = n6198 | n15036 ;
  assign n15038 = n8578 ^ x226 ^ 1'b0 ;
  assign n15039 = n420 & ~n15038 ;
  assign n15040 = n4537 & n15039 ;
  assign n15041 = n15040 ^ n12636 ^ 1'b0 ;
  assign n15042 = n13619 | n14355 ;
  assign n15043 = n9709 & ~n15042 ;
  assign n15044 = n11937 ^ n8887 ^ 1'b0 ;
  assign n15045 = n13504 & n15044 ;
  assign n15046 = ~n4246 & n15045 ;
  assign n15047 = n2887 & n6570 ;
  assign n15048 = n9421 & ~n12557 ;
  assign n15050 = n1641 ^ n821 ^ 1'b0 ;
  assign n15049 = ~n2497 & n13940 ;
  assign n15051 = n15050 ^ n15049 ^ 1'b0 ;
  assign n15052 = n14846 ^ n4555 ^ 1'b0 ;
  assign n15053 = ~n3575 & n15052 ;
  assign n15054 = ~n5534 & n9185 ;
  assign n15055 = x106 & n15054 ;
  assign n15056 = ~n2678 & n15055 ;
  assign n15057 = ~n11638 & n12176 ;
  assign n15058 = ~n6560 & n15057 ;
  assign n15059 = n2450 | n6128 ;
  assign n15060 = n5389 | n7461 ;
  assign n15061 = n2867 | n15060 ;
  assign n15062 = n7826 ^ x92 ^ 1'b0 ;
  assign n15063 = n15061 & ~n15062 ;
  assign n15064 = n15063 ^ n7833 ^ 1'b0 ;
  assign n15065 = n15059 | n15064 ;
  assign n15066 = n915 & ~n10855 ;
  assign n15067 = n15066 ^ n3064 ^ 1'b0 ;
  assign n15068 = n7734 & n15067 ;
  assign n15069 = n15068 ^ n2855 ^ 1'b0 ;
  assign n15070 = n10895 ^ n817 ^ 1'b0 ;
  assign n15071 = n15069 | n15070 ;
  assign n15072 = n7879 & ~n15071 ;
  assign n15073 = n15072 ^ n4276 ^ 1'b0 ;
  assign n15074 = n958 & ~n12615 ;
  assign n15075 = n15074 ^ n14076 ^ 1'b0 ;
  assign n15076 = n4230 ^ n2274 ^ 1'b0 ;
  assign n15077 = ~n6550 & n15076 ;
  assign n15078 = n5837 & n15077 ;
  assign n15079 = ~n7194 & n9226 ;
  assign n15080 = n15079 ^ n5848 ^ 1'b0 ;
  assign n15090 = ~n1678 & n5314 ;
  assign n15081 = n4356 & ~n9643 ;
  assign n15082 = n12385 ^ n1680 ^ 1'b0 ;
  assign n15083 = n5175 & ~n15082 ;
  assign n15084 = ~n15081 & n15083 ;
  assign n15085 = n5170 & n15084 ;
  assign n15086 = n9621 ^ n3434 ^ 1'b0 ;
  assign n15087 = ~n3662 & n15086 ;
  assign n15088 = n15085 & n15087 ;
  assign n15089 = n15088 ^ n2696 ^ 1'b0 ;
  assign n15091 = n15090 ^ n15089 ^ 1'b0 ;
  assign n15092 = n7298 | n8432 ;
  assign n15093 = ~n700 & n2664 ;
  assign n15094 = n15092 & n15093 ;
  assign n15095 = n1859 & ~n2503 ;
  assign n15096 = n8276 ^ n4377 ^ 1'b0 ;
  assign n15097 = n1307 | n9137 ;
  assign n15098 = n15097 ^ n2071 ^ 1'b0 ;
  assign n15099 = n590 & n1663 ;
  assign n15100 = n15099 ^ n3780 ^ 1'b0 ;
  assign n15101 = n6821 ^ n2435 ^ 1'b0 ;
  assign n15102 = n15100 | n15101 ;
  assign n15103 = n15102 ^ n6014 ^ 1'b0 ;
  assign n15104 = n14178 ^ n1935 ^ 1'b0 ;
  assign n15105 = ~x218 & n5407 ;
  assign n15106 = n7323 & n15105 ;
  assign n15107 = n11933 ^ n2997 ^ 1'b0 ;
  assign n15108 = ~n15106 & n15107 ;
  assign n15109 = ~n7148 & n8976 ;
  assign n15110 = ~x14 & n15109 ;
  assign n15112 = ~n4808 & n7179 ;
  assign n15113 = n4808 & n15112 ;
  assign n15111 = x101 & n8192 ;
  assign n15114 = n15113 ^ n15111 ^ 1'b0 ;
  assign n15115 = ~n1683 & n6178 ;
  assign n15116 = n1683 & n15115 ;
  assign n15117 = ~x3 & n15116 ;
  assign n15118 = ~n3039 & n15117 ;
  assign n15119 = ~n15114 & n15118 ;
  assign n15120 = n6372 & ~n13380 ;
  assign n15121 = ~n2395 & n15120 ;
  assign n15122 = n12592 ^ n1900 ^ 1'b0 ;
  assign n15123 = ( n9389 & n10038 ) | ( n9389 & ~n10344 ) | ( n10038 & ~n10344 ) ;
  assign n15124 = n9090 ^ x116 ^ 1'b0 ;
  assign n15125 = n4491 | n15124 ;
  assign n15126 = n15123 | n15125 ;
  assign n15127 = n8840 ^ n6590 ^ x161 ;
  assign n15128 = n6143 & n15127 ;
  assign n15129 = n8821 ^ n3475 ^ 1'b0 ;
  assign n15130 = n5493 & n15129 ;
  assign n15131 = n4828 ^ x62 ^ 1'b0 ;
  assign n15132 = ~n2743 & n15131 ;
  assign n15133 = n15132 ^ n10553 ^ 1'b0 ;
  assign n15134 = n1038 & n9040 ;
  assign n15135 = n15134 ^ n3264 ^ 1'b0 ;
  assign n15136 = n2761 | n3280 ;
  assign n15137 = n5237 | n15136 ;
  assign n15138 = n3217 & ~n7479 ;
  assign n15139 = ~n15137 & n15138 ;
  assign n15140 = n8514 ^ n880 ^ 1'b0 ;
  assign n15141 = n3013 | n15140 ;
  assign n15142 = n4261 | n15141 ;
  assign n15143 = ~n4314 & n5911 ;
  assign n15144 = n1431 & ~n2462 ;
  assign n15145 = n15144 ^ n13628 ^ 1'b0 ;
  assign n15146 = ~n4373 & n12128 ;
  assign n15147 = n15145 & ~n15146 ;
  assign n15148 = ~n15143 & n15147 ;
  assign n15149 = n500 & n2998 ;
  assign n15150 = ~n3221 & n15149 ;
  assign n15151 = n15150 ^ n3145 ^ 1'b0 ;
  assign n15152 = ~n4101 & n15151 ;
  assign n15153 = ~n4720 & n15152 ;
  assign n15154 = n4789 & n9445 ;
  assign n15155 = n15153 & n15154 ;
  assign n15156 = n12420 & ~n15155 ;
  assign n15157 = ~n8888 & n15156 ;
  assign n15158 = ~n9759 & n10498 ;
  assign n15159 = n14895 & n15158 ;
  assign n15161 = n662 | n4006 ;
  assign n15160 = n3604 & ~n11469 ;
  assign n15162 = n15161 ^ n15160 ^ 1'b0 ;
  assign n15163 = n1646 & ~n15162 ;
  assign n15164 = n2613 ^ n341 ^ 1'b0 ;
  assign n15165 = n15164 ^ n11173 ^ 1'b0 ;
  assign n15166 = n722 & ~n3518 ;
  assign n15167 = n15166 ^ n3905 ^ 1'b0 ;
  assign n15168 = n12514 | n14842 ;
  assign n15169 = n12574 ^ n5288 ^ 1'b0 ;
  assign n15170 = n465 & n13192 ;
  assign n15171 = ~n2164 & n15170 ;
  assign n15172 = n3462 ^ n1170 ^ 1'b0 ;
  assign n15173 = n8094 ^ n3468 ^ x176 ;
  assign n15174 = ~n6574 & n15173 ;
  assign n15175 = n9219 & n15174 ;
  assign n15176 = n8365 ^ x101 ^ 1'b0 ;
  assign n15177 = ~n15175 & n15176 ;
  assign n15178 = n3431 ^ n1588 ^ 1'b0 ;
  assign n15179 = n15178 ^ n9740 ^ 1'b0 ;
  assign n15180 = n10298 | n15179 ;
  assign n15181 = ~n5485 & n10665 ;
  assign n15182 = ~n3865 & n8997 ;
  assign n15183 = n14053 ^ n896 ^ 1'b0 ;
  assign n15184 = n7321 ^ n3331 ^ 1'b0 ;
  assign n15185 = n3015 | n15184 ;
  assign n15186 = n1670 & n15185 ;
  assign n15187 = n15183 & n15186 ;
  assign n15191 = ~n9184 & n13381 ;
  assign n15188 = n4039 & ~n6421 ;
  assign n15189 = ~x247 & n15188 ;
  assign n15190 = n12207 | n15189 ;
  assign n15192 = n15191 ^ n15190 ^ 1'b0 ;
  assign n15193 = n853 | n2661 ;
  assign n15194 = n15193 ^ n13201 ^ 1'b0 ;
  assign n15195 = n10682 & ~n11747 ;
  assign n15196 = n374 & n15195 ;
  assign n15197 = n1488 & n3234 ;
  assign n15198 = x218 & n1523 ;
  assign n15199 = ~n2600 & n15198 ;
  assign n15200 = n12536 ^ n9778 ^ 1'b0 ;
  assign n15201 = n12014 & ~n15200 ;
  assign n15202 = ~n698 & n1643 ;
  assign n15203 = n2185 & n15202 ;
  assign n15204 = n15203 ^ n10175 ^ n1626 ;
  assign n15205 = n6599 | n9860 ;
  assign n15206 = n15204 & ~n15205 ;
  assign n15207 = n14957 ^ n5255 ^ 1'b0 ;
  assign n15208 = n5385 & ~n15207 ;
  assign n15209 = n13738 ^ n11380 ^ 1'b0 ;
  assign n15210 = n8336 & ~n15209 ;
  assign n15211 = n3308 ^ n2861 ^ 1'b0 ;
  assign n15212 = n3756 & n15211 ;
  assign n15213 = ~n8462 & n15212 ;
  assign n15214 = n3678 & n15213 ;
  assign n15215 = n9084 & n15214 ;
  assign n15216 = n15215 ^ n3836 ^ 1'b0 ;
  assign n15217 = n15216 ^ n11109 ^ n892 ;
  assign n15218 = ~n14003 & n14858 ;
  assign n15219 = ~n3247 & n15218 ;
  assign n15220 = n1393 & ~n7860 ;
  assign n15221 = ~n3533 & n15220 ;
  assign n15222 = n11124 & ~n15221 ;
  assign n15223 = n15222 ^ n3830 ^ 1'b0 ;
  assign n15224 = ( n4594 & n5989 ) | ( n4594 & ~n15193 ) | ( n5989 & ~n15193 ) ;
  assign n15225 = n15224 ^ n13344 ^ n10629 ;
  assign n15226 = n4540 ^ x53 ^ 1'b0 ;
  assign n15227 = n15225 | n15226 ;
  assign n15228 = n1436 & n8600 ;
  assign n15229 = n1188 | n1907 ;
  assign n15230 = n15229 ^ n7206 ^ 1'b0 ;
  assign n15231 = n4730 | n15230 ;
  assign n15232 = n1905 & n7555 ;
  assign n15233 = ~n7869 & n15232 ;
  assign n15234 = n2562 & ~n6331 ;
  assign n15235 = ~n15233 & n15234 ;
  assign n15236 = n9728 & n11034 ;
  assign n15237 = n2081 & ~n2437 ;
  assign n15238 = n11196 ^ n7268 ^ 1'b0 ;
  assign n15239 = n8280 & n15238 ;
  assign n15240 = n5600 & ~n11544 ;
  assign n15241 = n13447 ^ n1531 ^ 1'b0 ;
  assign n15242 = n7914 ^ n2431 ^ 1'b0 ;
  assign n15243 = n15242 ^ n4113 ^ 1'b0 ;
  assign n15244 = n4558 ^ n1195 ^ 1'b0 ;
  assign n15245 = n642 & ~n15244 ;
  assign n15246 = ~n13899 & n15245 ;
  assign n15247 = n4872 ^ n4868 ^ 1'b0 ;
  assign n15248 = n10564 & n15247 ;
  assign n15249 = n15248 ^ n9381 ^ 1'b0 ;
  assign n15250 = ~n6764 & n7185 ;
  assign n15252 = ~n10691 & n12190 ;
  assign n15251 = n1839 | n9560 ;
  assign n15253 = n15252 ^ n15251 ^ 1'b0 ;
  assign n15254 = n15253 ^ n2370 ^ 1'b0 ;
  assign n15255 = n722 | n3681 ;
  assign n15256 = n7720 | n15255 ;
  assign n15257 = ~n5293 & n10300 ;
  assign n15258 = n15257 ^ n1025 ^ 1'b0 ;
  assign n15259 = n15258 ^ n4643 ^ 1'b0 ;
  assign n15260 = n9745 & ~n15259 ;
  assign n15261 = n2246 ^ n620 ^ 1'b0 ;
  assign n15262 = n15261 ^ n432 ^ 1'b0 ;
  assign n15263 = x85 & ~n15262 ;
  assign n15264 = n6674 | n15263 ;
  assign n15265 = ~n15101 & n15264 ;
  assign n15266 = n15265 ^ n9341 ^ 1'b0 ;
  assign n15267 = n4545 | n15266 ;
  assign n15268 = n2044 & ~n15267 ;
  assign n15269 = ~n15260 & n15268 ;
  assign n15270 = x118 & n666 ;
  assign n15271 = ~x118 & n15270 ;
  assign n15272 = x226 | n785 ;
  assign n15273 = n785 & ~n15272 ;
  assign n15274 = x239 & ~n15273 ;
  assign n15275 = n15271 & n15274 ;
  assign n15276 = n376 | n15275 ;
  assign n15277 = n15275 & ~n15276 ;
  assign n15278 = ~n2872 & n15277 ;
  assign n15279 = n7934 ^ n3153 ^ 1'b0 ;
  assign n15280 = n5507 & ~n15279 ;
  assign n15281 = n5316 & n15280 ;
  assign n15282 = ~n15280 & n15281 ;
  assign n15283 = n15278 | n15282 ;
  assign n15284 = n1780 | n15283 ;
  assign n15285 = n3786 ^ n3718 ^ 1'b0 ;
  assign n15286 = n15285 ^ n10608 ^ n3800 ;
  assign n15287 = n5378 ^ n1177 ^ 1'b0 ;
  assign n15288 = n8320 ^ n1841 ^ 1'b0 ;
  assign n15289 = n1700 & n15288 ;
  assign n15290 = n1301 & n15289 ;
  assign n15291 = ~n15287 & n15290 ;
  assign n15292 = n12949 & n15291 ;
  assign n15293 = n15286 & ~n15292 ;
  assign n15294 = n15293 ^ n2175 ^ 1'b0 ;
  assign n15295 = n14022 ^ n281 ^ 1'b0 ;
  assign n15296 = n15295 ^ n14705 ^ 1'b0 ;
  assign n15297 = n6407 & n15296 ;
  assign n15298 = x212 | n2076 ;
  assign n15299 = n10387 & n15298 ;
  assign n15300 = n15299 ^ n1694 ^ 1'b0 ;
  assign n15301 = n3710 & ~n6981 ;
  assign n15302 = ~n7615 & n15301 ;
  assign n15305 = n6657 ^ n6646 ^ 1'b0 ;
  assign n15306 = n15305 ^ n9944 ^ 1'b0 ;
  assign n15303 = n14984 ^ n5139 ^ 1'b0 ;
  assign n15304 = ~n9819 & n15303 ;
  assign n15307 = n15306 ^ n15304 ^ 1'b0 ;
  assign n15308 = n3878 ^ n387 ^ 1'b0 ;
  assign n15309 = n5343 & ~n15308 ;
  assign n15310 = n15309 ^ n11271 ^ 1'b0 ;
  assign n15311 = ~n2024 & n4957 ;
  assign n15312 = n4273 & ~n15311 ;
  assign n15313 = x229 & n4881 ;
  assign n15314 = n15313 ^ n2185 ^ 1'b0 ;
  assign n15315 = n1541 & ~n15314 ;
  assign n15316 = n15312 | n15315 ;
  assign n15317 = n2572 & ~n3551 ;
  assign n15318 = n15317 ^ n9185 ^ n6610 ;
  assign n15319 = n5739 | n13821 ;
  assign n15320 = n14861 & n15319 ;
  assign n15325 = ~n1435 & n2860 ;
  assign n15326 = n15325 ^ n5915 ^ 1'b0 ;
  assign n15321 = n6017 & ~n10275 ;
  assign n15322 = n8184 & n15321 ;
  assign n15323 = n15322 ^ n2872 ^ 1'b0 ;
  assign n15324 = n853 & n15323 ;
  assign n15327 = n15326 ^ n15324 ^ 1'b0 ;
  assign n15328 = n2786 & n13401 ;
  assign n15329 = n2730 & ~n9781 ;
  assign n15330 = n2037 | n4806 ;
  assign n15331 = n257 & n1514 ;
  assign n15332 = n9687 ^ n2845 ^ 1'b0 ;
  assign n15333 = ~n10004 & n10672 ;
  assign n15334 = ~n3862 & n15333 ;
  assign n15335 = n4416 | n15334 ;
  assign n15336 = n5615 & ~n8035 ;
  assign n15337 = n2330 & n5551 ;
  assign n15338 = n12791 & ~n15337 ;
  assign n15339 = n15338 ^ n5983 ^ 1'b0 ;
  assign n15340 = n6494 ^ n4741 ^ 1'b0 ;
  assign n15341 = n13664 & n15340 ;
  assign n15342 = ~n557 & n15341 ;
  assign n15343 = n15342 ^ n4980 ^ 1'b0 ;
  assign n15344 = n5498 & n11532 ;
  assign n15345 = ~n4556 & n12502 ;
  assign n15346 = ~n15344 & n15345 ;
  assign n15347 = n4300 | n14658 ;
  assign n15348 = n3441 | n15347 ;
  assign n15349 = n12118 & n12926 ;
  assign n15350 = n405 & n15349 ;
  assign n15351 = ~n3065 & n5175 ;
  assign n15352 = ~n4246 & n15351 ;
  assign n15353 = ~n7563 & n15352 ;
  assign n15354 = n15353 ^ n11102 ^ 1'b0 ;
  assign n15355 = ~n7791 & n15354 ;
  assign n15356 = ~n12729 & n14560 ;
  assign n15357 = n15356 ^ n10178 ^ 1'b0 ;
  assign n15358 = n6186 & ~n13549 ;
  assign n15359 = ~n4265 & n15358 ;
  assign n15360 = n5872 & ~n15359 ;
  assign n15361 = n15360 ^ n14666 ^ 1'b0 ;
  assign n15362 = n13426 ^ n4703 ^ 1'b0 ;
  assign n15363 = n2356 & n4298 ;
  assign n15364 = ~n15362 & n15363 ;
  assign n15365 = ~n8371 & n15364 ;
  assign n15366 = n14103 ^ n13182 ^ 1'b0 ;
  assign n15367 = n1951 & ~n4162 ;
  assign n15368 = n7108 & n15367 ;
  assign n15369 = ~n3459 & n15368 ;
  assign n15370 = n15369 ^ n8970 ^ 1'b0 ;
  assign n15371 = n4784 & ~n13029 ;
  assign n15372 = n6391 | n15371 ;
  assign n15373 = x21 & n7117 ;
  assign n15374 = n5665 & n9366 ;
  assign n15375 = n2620 & ~n11645 ;
  assign n15376 = n15374 & n15375 ;
  assign n15379 = n14538 ^ n13205 ^ 1'b0 ;
  assign n15377 = x182 | n1791 ;
  assign n15378 = n14362 & n15377 ;
  assign n15380 = n15379 ^ n15378 ^ 1'b0 ;
  assign n15381 = n5622 ^ n2098 ^ 1'b0 ;
  assign n15382 = ~n12138 & n15381 ;
  assign n15384 = n1062 ^ x31 ^ 1'b0 ;
  assign n15383 = n2898 & n14275 ;
  assign n15385 = n15384 ^ n15383 ^ 1'b0 ;
  assign n15386 = n3065 | n5964 ;
  assign n15387 = n3850 ^ n2901 ^ 1'b0 ;
  assign n15388 = n6626 ^ n3516 ^ 1'b0 ;
  assign n15389 = n15388 ^ n1475 ^ 1'b0 ;
  assign n15390 = n8279 & n13576 ;
  assign n15391 = n15390 ^ n1002 ^ 1'b0 ;
  assign n15392 = n2161 & ~n14707 ;
  assign n15396 = ~n2796 & n10997 ;
  assign n15394 = ~n397 & n2428 ;
  assign n15395 = ~n6250 & n15394 ;
  assign n15393 = n2345 ^ n1525 ^ 1'b0 ;
  assign n15397 = n15396 ^ n15395 ^ n15393 ;
  assign n15398 = n6106 ^ n3040 ^ 1'b0 ;
  assign n15399 = ( ~n3123 & n4824 ) | ( ~n3123 & n15398 ) | ( n4824 & n15398 ) ;
  assign n15400 = n5712 & ~n12765 ;
  assign n15401 = n11775 ^ n5911 ^ n2764 ;
  assign n15402 = ~n1017 & n10567 ;
  assign n15403 = ~n15401 & n15402 ;
  assign n15404 = n12720 ^ n11210 ^ 1'b0 ;
  assign n15405 = n8933 ^ n1896 ^ 1'b0 ;
  assign n15406 = n4784 & n15405 ;
  assign n15407 = n15406 ^ n14957 ^ 1'b0 ;
  assign n15408 = n15407 ^ n9483 ^ 1'b0 ;
  assign n15409 = n6455 ^ n1693 ^ 1'b0 ;
  assign n15410 = n15409 ^ n7483 ^ 1'b0 ;
  assign n15411 = n13431 & ~n15410 ;
  assign n15412 = n6945 ^ n6536 ^ 1'b0 ;
  assign n15413 = n15411 & n15412 ;
  assign n15414 = ~n1682 & n13066 ;
  assign n15415 = n15414 ^ n12314 ^ 1'b0 ;
  assign n15416 = n6258 | n15415 ;
  assign n15417 = n5157 & ~n9463 ;
  assign n15418 = n3239 & ~n3995 ;
  assign n15419 = n15418 ^ n2519 ^ 1'b0 ;
  assign n15420 = ~n600 & n9771 ;
  assign n15421 = n15420 ^ n10495 ^ 1'b0 ;
  assign n15422 = n1361 & ~n4396 ;
  assign n15423 = ~n4556 & n14068 ;
  assign n15424 = ~n11375 & n15423 ;
  assign n15425 = ~n2078 & n15424 ;
  assign n15426 = n7107 | n9867 ;
  assign n15427 = n15426 ^ n2957 ^ 1'b0 ;
  assign n15428 = n3465 ^ n2350 ^ 1'b0 ;
  assign n15429 = n13899 | n15428 ;
  assign n15430 = n15427 & ~n15429 ;
  assign n15431 = n1556 & ~n8543 ;
  assign n15432 = n15431 ^ x207 ^ 1'b0 ;
  assign n15433 = n11931 ^ n6816 ^ 1'b0 ;
  assign n15434 = n8079 ^ n6021 ^ 1'b0 ;
  assign n15435 = n4750 | n15434 ;
  assign n15436 = ~n2846 & n14106 ;
  assign n15437 = ~n1505 & n15280 ;
  assign n15438 = n15437 ^ n4549 ^ 1'b0 ;
  assign n15439 = ~n3832 & n10498 ;
  assign n15440 = n15439 ^ n1820 ^ 1'b0 ;
  assign n15441 = n15440 ^ n1605 ^ 1'b0 ;
  assign n15443 = n6154 | n9212 ;
  assign n15444 = n6605 & ~n15443 ;
  assign n15442 = n1368 & ~n5750 ;
  assign n15445 = n15444 ^ n15442 ^ 1'b0 ;
  assign n15447 = n1360 ^ x59 ^ 1'b0 ;
  assign n15446 = n4821 & n6617 ;
  assign n15448 = n15447 ^ n15446 ^ 1'b0 ;
  assign n15449 = n5023 & ~n15448 ;
  assign n15450 = n444 & n9196 ;
  assign n15451 = ~n1191 & n15450 ;
  assign n15452 = n2194 & n14589 ;
  assign n15453 = n15452 ^ n12625 ^ 1'b0 ;
  assign n15454 = n1272 | n15453 ;
  assign n15455 = n6760 ^ n320 ^ 1'b0 ;
  assign n15456 = n7320 & ~n15455 ;
  assign n15457 = x212 & n2582 ;
  assign n15458 = n15456 & n15457 ;
  assign n15459 = n2892 | n15458 ;
  assign n15460 = n3837 | n15459 ;
  assign n15461 = n3353 | n7383 ;
  assign n15462 = n15461 ^ n7929 ^ 1'b0 ;
  assign n15463 = n15462 ^ n1302 ^ 1'b0 ;
  assign n15464 = n15463 ^ n642 ^ 1'b0 ;
  assign n15465 = n14077 | n15464 ;
  assign n15466 = n3235 | n15465 ;
  assign n15467 = n3611 & n4851 ;
  assign n15468 = n15467 ^ n7557 ^ 1'b0 ;
  assign n15469 = n12848 ^ n1339 ^ 1'b0 ;
  assign n15470 = n14458 ^ x161 ^ 1'b0 ;
  assign n15471 = n8722 ^ n747 ^ 1'b0 ;
  assign n15472 = n15471 ^ n11689 ^ 1'b0 ;
  assign n15473 = ~n11308 & n13049 ;
  assign n15474 = n9886 & n15473 ;
  assign n15475 = ~n363 & n5882 ;
  assign n15476 = ~n2866 & n15475 ;
  assign n15477 = ~n2241 & n15476 ;
  assign n15478 = n1421 & n1762 ;
  assign n15479 = n15478 ^ n3270 ^ 1'b0 ;
  assign n15480 = n11207 ^ x84 ^ 1'b0 ;
  assign n15481 = n5215 & n7757 ;
  assign n15482 = n1847 & n2558 ;
  assign n15483 = ~n3803 & n15482 ;
  assign n15484 = n2106 & n5203 ;
  assign n15485 = ~n3366 & n15484 ;
  assign n15486 = ( n2063 & n9523 ) | ( n2063 & n15485 ) | ( n9523 & n15485 ) ;
  assign n15487 = n15486 ^ n538 ^ 1'b0 ;
  assign n15488 = ~n9199 & n15487 ;
  assign n15489 = n15488 ^ n927 ^ 1'b0 ;
  assign n15490 = n7161 | n15489 ;
  assign n15491 = n15483 & ~n15490 ;
  assign n15492 = ~n4739 & n12174 ;
  assign n15493 = ~n860 & n15492 ;
  assign n15494 = n2776 | n4223 ;
  assign n15495 = n1397 | n15494 ;
  assign n15496 = n1767 & n8968 ;
  assign n15497 = ~n15495 & n15496 ;
  assign n15498 = x67 & ~n3071 ;
  assign n15499 = n6062 ^ n1535 ^ 1'b0 ;
  assign n15500 = n15499 ^ n8516 ^ 1'b0 ;
  assign n15501 = n15498 | n15500 ;
  assign n15502 = n5392 & ~n5796 ;
  assign n15503 = n15502 ^ n13638 ^ 1'b0 ;
  assign n15504 = n7177 & ~n9354 ;
  assign n15505 = n15504 ^ n11336 ^ 1'b0 ;
  assign n15513 = n1337 ^ n415 ^ 1'b0 ;
  assign n15509 = ~n1877 & n11291 ;
  assign n15506 = n8529 ^ n6214 ^ 1'b0 ;
  assign n15507 = n445 | n15506 ;
  assign n15508 = n6739 | n15507 ;
  assign n15510 = n15509 ^ n15508 ^ 1'b0 ;
  assign n15511 = n5300 | n15510 ;
  assign n15512 = n14942 | n15511 ;
  assign n15514 = n15513 ^ n15512 ^ 1'b0 ;
  assign n15515 = ~n6834 & n7628 ;
  assign n15516 = n5047 ^ n1273 ^ 1'b0 ;
  assign n15517 = n13286 ^ n766 ^ 1'b0 ;
  assign n15518 = n6283 | n15517 ;
  assign n15519 = n15518 ^ n571 ^ 1'b0 ;
  assign n15520 = n5879 & n10886 ;
  assign n15521 = n15520 ^ n14828 ^ 1'b0 ;
  assign n15522 = n1272 ^ n809 ^ 1'b0 ;
  assign n15523 = n2022 | n4600 ;
  assign n15524 = n11135 | n15523 ;
  assign n15525 = n15057 ^ n14177 ^ n11363 ;
  assign n15526 = n6646 | n10513 ;
  assign n15527 = n15526 ^ n9737 ^ 1'b0 ;
  assign n15528 = n13312 ^ n4189 ^ 1'b0 ;
  assign n15529 = n8167 | n15528 ;
  assign n15530 = n15212 ^ x86 ^ 1'b0 ;
  assign n15531 = n5263 ^ n2279 ^ 1'b0 ;
  assign n15532 = n12118 ^ n720 ^ 1'b0 ;
  assign n15533 = n10997 | n15532 ;
  assign n15534 = n635 | n15533 ;
  assign n15535 = n15534 ^ n12756 ^ 1'b0 ;
  assign n15536 = n10495 ^ n3397 ^ 1'b0 ;
  assign n15537 = ~n5818 & n15536 ;
  assign n15538 = ~n1511 & n2562 ;
  assign n15539 = n15538 ^ n2830 ^ 1'b0 ;
  assign n15540 = n15537 & n15539 ;
  assign n15541 = n15540 ^ n5106 ^ 1'b0 ;
  assign n15542 = n15535 & ~n15541 ;
  assign n15543 = ~n1139 & n8672 ;
  assign n15544 = n5418 ^ n840 ^ 1'b0 ;
  assign n15545 = ~n2833 & n15544 ;
  assign n15546 = n15545 ^ n9765 ^ 1'b0 ;
  assign n15547 = n15546 ^ n9379 ^ 1'b0 ;
  assign n15548 = n12941 ^ n7043 ^ 1'b0 ;
  assign n15549 = n14031 ^ n4074 ^ 1'b0 ;
  assign n15550 = n15258 | n15549 ;
  assign n15551 = n2215 | n7274 ;
  assign n15552 = n2129 | n15551 ;
  assign n15553 = ~n4586 & n6372 ;
  assign n15554 = n15553 ^ x125 ^ 1'b0 ;
  assign n15555 = n13441 ^ n1410 ^ 1'b0 ;
  assign n15556 = n3868 | n15555 ;
  assign n15557 = n4549 & n4788 ;
  assign n15558 = ~n4296 & n15557 ;
  assign n15559 = x202 & ~n15558 ;
  assign n15560 = n6895 & n15559 ;
  assign n15561 = n4190 | n13978 ;
  assign n15562 = n864 | n6811 ;
  assign n15563 = n1591 & ~n15562 ;
  assign n15564 = n8484 | n8609 ;
  assign n15565 = x182 & n2720 ;
  assign n15566 = n2632 & ~n3578 ;
  assign n15567 = n6847 & ~n15566 ;
  assign n15568 = n3417 & n15567 ;
  assign n15569 = ~n872 & n15568 ;
  assign n15570 = n5079 & n9576 ;
  assign n15571 = ~x24 & n15570 ;
  assign n15572 = n15571 ^ n15340 ^ 1'b0 ;
  assign n15573 = ~n4363 & n8382 ;
  assign n15574 = n6295 & n15573 ;
  assign n15575 = n6888 ^ n4538 ^ 1'b0 ;
  assign n15576 = n3914 & n15575 ;
  assign n15577 = n3591 ^ x185 ^ 1'b0 ;
  assign n15578 = ~n2191 & n15577 ;
  assign n15579 = n14589 | n15578 ;
  assign n15580 = n3105 & ~n6217 ;
  assign n15581 = ~n3591 & n4728 ;
  assign n15582 = n7105 & ~n14534 ;
  assign n15583 = n10344 & ~n12809 ;
  assign n15584 = n7077 & ~n13447 ;
  assign n15585 = n15584 ^ n10418 ^ 1'b0 ;
  assign n15588 = n5909 ^ n1864 ^ 1'b0 ;
  assign n15589 = n5598 & n15588 ;
  assign n15590 = ~n1955 & n15589 ;
  assign n15591 = n6238 & n15590 ;
  assign n15586 = n4478 & n4668 ;
  assign n15587 = ~n4946 & n15586 ;
  assign n15592 = n15591 ^ n15587 ^ 1'b0 ;
  assign n15593 = n4903 & n15592 ;
  assign n15594 = n15593 ^ n11197 ^ 1'b0 ;
  assign n15595 = n2186 | n15594 ;
  assign n15596 = n15595 ^ n11694 ^ 1'b0 ;
  assign n15597 = n1436 & n15596 ;
  assign n15598 = ~n5626 & n14572 ;
  assign n15599 = n2904 & n15598 ;
  assign n15600 = ~n6431 & n15599 ;
  assign n15601 = ( ~n8458 & n9982 ) | ( ~n8458 & n15600 ) | ( n9982 & n15600 ) ;
  assign n15602 = n10270 ^ n10158 ^ 1'b0 ;
  assign n15603 = n14670 ^ n6258 ^ 1'b0 ;
  assign n15604 = n8553 ^ n4334 ^ 1'b0 ;
  assign n15605 = n2087 | n15484 ;
  assign n15606 = n3489 | n15605 ;
  assign n15607 = n2476 | n15606 ;
  assign n15608 = n4569 ^ n949 ^ 1'b0 ;
  assign n15609 = n15607 & ~n15608 ;
  assign n15611 = n1000 | n1939 ;
  assign n15612 = ~n8725 & n15611 ;
  assign n15610 = ~n2318 & n2764 ;
  assign n15613 = n15612 ^ n15610 ^ 1'b0 ;
  assign n15616 = n6786 ^ n4124 ^ 1'b0 ;
  assign n15614 = n13668 ^ n7098 ^ 1'b0 ;
  assign n15615 = n11723 & n15614 ;
  assign n15617 = n15616 ^ n15615 ^ 1'b0 ;
  assign n15622 = n6028 ^ n4276 ^ 1'b0 ;
  assign n15623 = n9487 & ~n15622 ;
  assign n15624 = ~n8214 & n15623 ;
  assign n15625 = n15624 ^ n10908 ^ 1'b0 ;
  assign n15626 = ~n6396 & n15625 ;
  assign n15627 = n8212 & n15626 ;
  assign n15618 = ( n589 & n2006 ) | ( n589 & n3847 ) | ( n2006 & n3847 ) ;
  assign n15619 = n2661 | n15618 ;
  assign n15620 = n8169 & ~n15619 ;
  assign n15621 = n1356 | n15620 ;
  assign n15628 = n15627 ^ n15621 ^ 1'b0 ;
  assign n15629 = n2652 ^ n812 ^ n683 ;
  assign n15630 = x160 | n3624 ;
  assign n15631 = n15630 ^ n7671 ^ 1'b0 ;
  assign n15632 = ~n13953 & n15631 ;
  assign n15635 = x34 & n11451 ;
  assign n15636 = n13056 ^ n3532 ^ n1793 ;
  assign n15637 = n15635 & ~n15636 ;
  assign n15633 = n3325 & ~n7310 ;
  assign n15634 = n2818 & n15633 ;
  assign n15638 = n15637 ^ n15634 ^ 1'b0 ;
  assign n15639 = n838 & ~n4054 ;
  assign n15640 = n15639 ^ n4645 ^ 1'b0 ;
  assign n15641 = n1050 & ~n10495 ;
  assign n15642 = n15641 ^ n562 ^ 1'b0 ;
  assign n15643 = n15640 | n15642 ;
  assign n15644 = ~n4671 & n12055 ;
  assign n15645 = n15643 | n15644 ;
  assign n15646 = n7179 & ~n15645 ;
  assign n15647 = n2443 & ~n15646 ;
  assign n15648 = n4267 ^ x254 ^ 1'b0 ;
  assign n15649 = n7164 | n15648 ;
  assign n15650 = n15649 ^ n5493 ^ 1'b0 ;
  assign n15651 = n2102 ^ n748 ^ n361 ;
  assign n15652 = n7140 ^ n6411 ^ 1'b0 ;
  assign n15653 = n7326 & ~n15652 ;
  assign n15654 = n2989 & n6243 ;
  assign n15655 = x182 & ~n1202 ;
  assign n15656 = ~n15654 & n15655 ;
  assign n15657 = n3780 ^ x50 ^ x43 ;
  assign n15658 = n13261 ^ n2254 ^ 1'b0 ;
  assign n15659 = n4431 & n15658 ;
  assign n15660 = ~n6553 & n15659 ;
  assign n15661 = n9066 ^ n3774 ^ 1'b0 ;
  assign n15664 = ~n3093 & n5378 ;
  assign n15665 = n15664 ^ n7474 ^ 1'b0 ;
  assign n15662 = n540 & n6563 ;
  assign n15663 = n2470 & n15662 ;
  assign n15666 = n15665 ^ n15663 ^ 1'b0 ;
  assign n15667 = n15666 ^ n8364 ^ 1'b0 ;
  assign n15668 = n4874 & ~n8808 ;
  assign n15669 = n3714 & n10082 ;
  assign n15670 = n15669 ^ n9000 ^ 1'b0 ;
  assign n15671 = n8976 | n15670 ;
  assign n15672 = n3830 & n5101 ;
  assign n15673 = ~n2235 & n8765 ;
  assign n15674 = n15673 ^ n5717 ^ 1'b0 ;
  assign n15675 = n14551 & ~n15674 ;
  assign n15676 = n9387 & ~n15675 ;
  assign n15677 = n5372 & n15676 ;
  assign n15678 = n15677 ^ n3255 ^ n354 ;
  assign n15679 = n3710 & n14117 ;
  assign n15680 = n4598 & n15679 ;
  assign n15681 = n14919 ^ n9731 ^ 1'b0 ;
  assign n15682 = n8872 & ~n13599 ;
  assign n15683 = n4811 & ~n15682 ;
  assign n15684 = n15683 ^ n2402 ^ 1'b0 ;
  assign n15685 = n13538 ^ n1021 ^ 1'b0 ;
  assign n15686 = n9416 ^ n6729 ^ 1'b0 ;
  assign n15687 = n5750 & ~n14365 ;
  assign n15688 = n15687 ^ n2901 ^ 1'b0 ;
  assign n15689 = ~n15686 & n15688 ;
  assign n15690 = n6383 ^ n2944 ^ 1'b0 ;
  assign n15691 = n15690 ^ n5000 ^ 1'b0 ;
  assign n15692 = n7214 | n15691 ;
  assign n15693 = n6022 | n15692 ;
  assign n15694 = n7170 ^ n2824 ^ 1'b0 ;
  assign n15695 = n15694 ^ n4838 ^ 1'b0 ;
  assign n15696 = n6499 & ~n9654 ;
  assign n15698 = n9687 ^ x206 ^ 1'b0 ;
  assign n15699 = n15698 ^ n7526 ^ 1'b0 ;
  assign n15697 = ~n994 & n1618 ;
  assign n15700 = n15699 ^ n15697 ^ 1'b0 ;
  assign n15701 = ( ~n3348 & n5658 ) | ( ~n3348 & n15261 ) | ( n5658 & n15261 ) ;
  assign n15702 = ~n10969 & n14498 ;
  assign n15703 = n15702 ^ n1826 ^ 1'b0 ;
  assign n15704 = n3073 & ~n8354 ;
  assign n15705 = n15704 ^ n2272 ^ 1'b0 ;
  assign n15706 = n11343 ^ n6089 ^ 1'b0 ;
  assign n15707 = ~n10157 & n15706 ;
  assign n15712 = ~n7021 & n7578 ;
  assign n15708 = n1247 & ~n8298 ;
  assign n15709 = ~n6777 & n15708 ;
  assign n15710 = n780 | n15709 ;
  assign n15711 = n15710 ^ n6008 ^ 1'b0 ;
  assign n15713 = n15712 ^ n15711 ^ x57 ;
  assign n15714 = n15707 & n15713 ;
  assign n15715 = n3964 & ~n15714 ;
  assign n15716 = n11611 ^ n1914 ^ 1'b0 ;
  assign n15717 = n15716 ^ n9368 ^ 1'b0 ;
  assign n15718 = n12077 | n15678 ;
  assign n15719 = n3556 ^ n2702 ^ n964 ;
  assign n15720 = ~n5958 & n15719 ;
  assign n15721 = n1605 & n11172 ;
  assign n15722 = ~n1116 & n4701 ;
  assign n15723 = n15722 ^ n964 ^ 1'b0 ;
  assign n15724 = n7695 | n8286 ;
  assign n15725 = n14272 & ~n15724 ;
  assign n15726 = ~n415 & n15725 ;
  assign n15727 = n12553 ^ n1195 ^ 1'b0 ;
  assign n15728 = n4279 & n15727 ;
  assign n15729 = n15728 ^ n12298 ^ 1'b0 ;
  assign n15730 = n3331 | n8311 ;
  assign n15731 = n15730 ^ n10152 ^ 1'b0 ;
  assign n15732 = n1961 & ~n10201 ;
  assign n15733 = n15732 ^ n3817 ^ 1'b0 ;
  assign n15734 = n7449 & n15733 ;
  assign n15735 = n10059 ^ n6276 ^ 1'b0 ;
  assign n15736 = n2630 & ~n3182 ;
  assign n15737 = n859 & n4166 ;
  assign n15738 = ~n2944 & n3698 ;
  assign n15739 = n15738 ^ n1790 ^ 1'b0 ;
  assign n15740 = n10333 ^ n2242 ^ 1'b0 ;
  assign n15741 = n1591 | n15740 ;
  assign n15742 = n15739 & ~n15741 ;
  assign n15743 = n15742 ^ n3837 ^ 1'b0 ;
  assign n15744 = n2100 & ~n15743 ;
  assign n15747 = ~n1694 & n8006 ;
  assign n15748 = ~n3171 & n15747 ;
  assign n15745 = n10322 ^ n1112 ^ 1'b0 ;
  assign n15746 = n15745 ^ n11763 ^ n10089 ;
  assign n15749 = n15748 ^ n15746 ^ n3703 ;
  assign n15750 = n3507 & ~n4189 ;
  assign n15751 = n15750 ^ n497 ^ 1'b0 ;
  assign n15752 = x186 & n15751 ;
  assign n15753 = n11906 & ~n15752 ;
  assign n15754 = n14784 & n15753 ;
  assign n15755 = n10689 ^ n355 ^ 1'b0 ;
  assign n15756 = n5988 | n15755 ;
  assign n15757 = n5924 ^ n2061 ^ 1'b0 ;
  assign n15758 = n2310 & ~n5648 ;
  assign n15759 = ~n2310 & n15758 ;
  assign n15760 = n313 & ~n956 ;
  assign n15761 = n956 & n15760 ;
  assign n15762 = n754 & n15761 ;
  assign n15763 = n5336 | n15762 ;
  assign n15764 = n5336 & ~n15763 ;
  assign n15765 = n11654 & n15764 ;
  assign n15766 = n15759 | n15765 ;
  assign n15767 = n15759 & ~n15766 ;
  assign n15768 = n3083 ^ x229 ^ 1'b0 ;
  assign n15769 = n698 | n5256 ;
  assign n15770 = n15768 | n15769 ;
  assign n15771 = n2848 & n2881 ;
  assign n15772 = n15771 ^ n1576 ^ 1'b0 ;
  assign n15773 = n15772 ^ n15547 ^ 1'b0 ;
  assign n15774 = ( n2765 & n4429 ) | ( n2765 & n8706 ) | ( n4429 & n8706 ) ;
  assign n15775 = n4739 & ~n15774 ;
  assign n15776 = n8737 & n11439 ;
  assign n15777 = ~n1556 & n15776 ;
  assign n15778 = ~n3856 & n14675 ;
  assign n15779 = n15777 & n15778 ;
  assign n15780 = ( ~n3632 & n5529 ) | ( ~n3632 & n9503 ) | ( n5529 & n9503 ) ;
  assign n15781 = n14646 & ~n15780 ;
  assign n15782 = n3091 & ~n6295 ;
  assign n15783 = n15782 ^ n1740 ^ 1'b0 ;
  assign n15784 = n8082 & ~n10473 ;
  assign n15785 = ~n8179 & n11711 ;
  assign n15786 = n6771 & n15785 ;
  assign n15787 = n1701 | n7922 ;
  assign n15788 = n15787 ^ n6049 ^ 1'b0 ;
  assign n15789 = ~n15786 & n15788 ;
  assign n15790 = n2816 & n4398 ;
  assign n15791 = n2854 & n15790 ;
  assign n15792 = n15032 | n15791 ;
  assign n15793 = n10908 & ~n15792 ;
  assign n15794 = n3807 & n11647 ;
  assign n15795 = n4589 ^ n1370 ^ 1'b0 ;
  assign n15796 = n5036 & n15795 ;
  assign n15797 = n15796 ^ n15477 ^ n6552 ;
  assign n15798 = n12578 ^ n7297 ^ 1'b0 ;
  assign n15799 = n5370 | n15798 ;
  assign n15800 = n14127 ^ n9815 ^ 1'b0 ;
  assign n15801 = n361 & ~n2412 ;
  assign n15802 = n366 | n1681 ;
  assign n15803 = n15802 ^ n10797 ^ 1'b0 ;
  assign n15804 = n6207 | n15803 ;
  assign n15805 = n10433 ^ n8657 ^ 1'b0 ;
  assign n15806 = n3812 & n15805 ;
  assign n15807 = n15465 | n15806 ;
  assign n15808 = n5015 | n14759 ;
  assign n15809 = n14105 & ~n15808 ;
  assign n15810 = n7792 | n10465 ;
  assign n15811 = n887 | n6109 ;
  assign n15812 = n5356 | n15811 ;
  assign n15813 = ~n3965 & n15812 ;
  assign n15814 = n5418 ^ n978 ^ 1'b0 ;
  assign n15815 = n397 & ~n3703 ;
  assign n15816 = ~n3960 & n15815 ;
  assign n15817 = n15816 ^ n14030 ^ 1'b0 ;
  assign n15818 = n2082 & ~n10777 ;
  assign n15819 = n8760 & ~n14113 ;
  assign n15820 = n3590 | n7002 ;
  assign n15821 = n10763 | n14298 ;
  assign n15822 = n5162 & ~n15821 ;
  assign n15823 = ~n623 & n12714 ;
  assign n15824 = n12041 & n15823 ;
  assign n15825 = n8801 ^ n2752 ^ n1968 ;
  assign n15826 = n15825 ^ n8419 ^ 1'b0 ;
  assign n15827 = n15824 | n15826 ;
  assign n15828 = n7878 & n11511 ;
  assign n15829 = n15828 ^ n4260 ^ 1'b0 ;
  assign n15830 = n1608 & ~n4913 ;
  assign n15831 = n15830 ^ n2867 ^ 1'b0 ;
  assign n15832 = ~n1031 & n4147 ;
  assign n15833 = ~n1076 & n6944 ;
  assign n15834 = ~n6944 & n15833 ;
  assign n15835 = n7218 ^ n1905 ^ 1'b0 ;
  assign n15836 = n1682 & ~n7559 ;
  assign n15837 = ~n1682 & n15836 ;
  assign n15838 = n15835 & ~n15837 ;
  assign n15839 = n15834 & n15838 ;
  assign n15840 = n7980 | n15839 ;
  assign n15841 = n1302 & n2858 ;
  assign n15842 = n15841 ^ n5658 ^ n1632 ;
  assign n15843 = n11487 ^ n851 ^ 1'b0 ;
  assign n15844 = n15842 & n15843 ;
  assign n15845 = n1562 ^ n797 ^ 1'b0 ;
  assign n15846 = ~n5222 & n15845 ;
  assign n15847 = n15846 ^ n5266 ^ 1'b0 ;
  assign n15848 = n5235 & n6539 ;
  assign n15849 = n2852 & n15848 ;
  assign n15850 = n15849 ^ n11065 ^ 1'b0 ;
  assign n15851 = n10740 & ~n15850 ;
  assign n15852 = n12266 ^ n3083 ^ 1'b0 ;
  assign n15853 = n6685 & n13144 ;
  assign n15854 = n10276 | n10953 ;
  assign n15855 = n8212 ^ n2623 ^ 1'b0 ;
  assign n15856 = n14275 ^ n4993 ^ 1'b0 ;
  assign n15857 = n15856 ^ n6969 ^ 1'b0 ;
  assign n15858 = n7750 | n15857 ;
  assign n15859 = n1639 & ~n5382 ;
  assign n15860 = n1563 & ~n7775 ;
  assign n15861 = ~n3223 & n14241 ;
  assign n15863 = n12509 ^ n2519 ^ 1'b0 ;
  assign n15864 = n11457 & n15863 ;
  assign n15862 = n10551 | n13159 ;
  assign n15865 = n15864 ^ n15862 ^ 1'b0 ;
  assign n15866 = n5586 & ~n13595 ;
  assign n15868 = ~n311 & n2517 ;
  assign n15869 = n15868 ^ n2186 ^ 1'b0 ;
  assign n15867 = n4899 | n8129 ;
  assign n15870 = n15869 ^ n15867 ^ 1'b0 ;
  assign n15871 = n1537 & ~n15870 ;
  assign n15872 = n9174 | n15871 ;
  assign n15873 = n15872 ^ n809 ^ 1'b0 ;
  assign n15874 = n6383 & n15873 ;
  assign n15879 = n8348 ^ n5904 ^ 1'b0 ;
  assign n15880 = n717 & n15879 ;
  assign n15878 = n7265 | n10126 ;
  assign n15881 = n15880 ^ n15878 ^ n2629 ;
  assign n15875 = n778 & ~n6438 ;
  assign n15876 = ~n12359 & n15875 ;
  assign n15877 = n1442 | n15876 ;
  assign n15882 = n15881 ^ n15877 ^ n14591 ;
  assign n15887 = n6667 ^ n2629 ^ 1'b0 ;
  assign n15888 = n15887 ^ n4321 ^ 1'b0 ;
  assign n15889 = n8442 & n15888 ;
  assign n15883 = n3174 ^ n2470 ^ 1'b0 ;
  assign n15884 = n7358 & ~n15883 ;
  assign n15885 = n3830 & ~n7816 ;
  assign n15886 = ~n15884 & n15885 ;
  assign n15890 = n15889 ^ n15886 ^ 1'b0 ;
  assign n15891 = n7994 ^ n6241 ^ 1'b0 ;
  assign n15892 = n415 | n15891 ;
  assign n15893 = n1390 | n2861 ;
  assign n15894 = n15893 ^ n6578 ^ 1'b0 ;
  assign n15895 = n3789 & ~n15894 ;
  assign n15899 = ~n920 & n3985 ;
  assign n15900 = ~n286 & n15899 ;
  assign n15897 = n1269 | n3176 ;
  assign n15898 = n15897 ^ n2011 ^ 1'b0 ;
  assign n15896 = n3144 & n6696 ;
  assign n15901 = n15900 ^ n15898 ^ n15896 ;
  assign n15902 = n14036 ^ n2647 ^ 1'b0 ;
  assign n15903 = n9876 | n15902 ;
  assign n15904 = n13118 ^ n3858 ^ 1'b0 ;
  assign n15905 = n6974 ^ n5659 ^ 1'b0 ;
  assign n15906 = n11908 | n15905 ;
  assign n15907 = n8548 & n10284 ;
  assign n15908 = ~n5262 & n11438 ;
  assign n15909 = ( ~n1125 & n2230 ) | ( ~n1125 & n10138 ) | ( n2230 & n10138 ) ;
  assign n15910 = ~n10843 & n10991 ;
  assign n15911 = ( n4067 & n4840 ) | ( n4067 & n11191 ) | ( n4840 & n11191 ) ;
  assign n15919 = n7924 ^ n6861 ^ n2858 ;
  assign n15912 = n6173 ^ n5909 ^ 1'b0 ;
  assign n15913 = n5672 & n15912 ;
  assign n15914 = n573 | n3059 ;
  assign n15915 = n7431 | n15914 ;
  assign n15916 = ( ~n3729 & n15913 ) | ( ~n3729 & n15915 ) | ( n15913 & n15915 ) ;
  assign n15917 = n3957 & n8660 ;
  assign n15918 = ~n15916 & n15917 ;
  assign n15920 = n15919 ^ n15918 ^ 1'b0 ;
  assign n15921 = n15911 & ~n15920 ;
  assign n15922 = n15616 & n15921 ;
  assign n15923 = n2184 & n3163 ;
  assign n15924 = n15923 ^ n12360 ^ 1'b0 ;
  assign n15925 = n8768 ^ n4598 ^ 1'b0 ;
  assign n15926 = n7649 ^ n6095 ^ 1'b0 ;
  assign n15927 = n15736 & n15926 ;
  assign n15930 = n2402 | n4955 ;
  assign n15931 = n15930 ^ n1291 ^ 1'b0 ;
  assign n15928 = n11218 ^ n2400 ^ n641 ;
  assign n15929 = ~n5904 & n15928 ;
  assign n15932 = n15931 ^ n15929 ^ 1'b0 ;
  assign n15933 = n2127 | n9785 ;
  assign n15934 = n15933 ^ n6444 ^ 1'b0 ;
  assign n15935 = ~n2709 & n15934 ;
  assign n15936 = ~n814 & n11895 ;
  assign n15937 = n15936 ^ n6422 ^ 1'b0 ;
  assign n15938 = x100 & ~n15743 ;
  assign n15939 = n4526 & n14955 ;
  assign n15940 = n1512 & ~n12157 ;
  assign n15941 = n12157 & n15940 ;
  assign n15942 = n7202 ^ n6537 ^ n5207 ;
  assign n15943 = ( ~n13675 & n15941 ) | ( ~n13675 & n15942 ) | ( n15941 & n15942 ) ;
  assign n15948 = ~n605 & n1477 ;
  assign n15949 = n4558 & n15948 ;
  assign n15944 = n5481 ^ n1512 ^ 1'b0 ;
  assign n15945 = n9229 & ~n15944 ;
  assign n15946 = ~n2636 & n15945 ;
  assign n15947 = n15946 ^ n8092 ^ 1'b0 ;
  assign n15950 = n15949 ^ n15947 ^ 1'b0 ;
  assign n15951 = n11859 | n15950 ;
  assign n15952 = x22 | n2136 ;
  assign n15953 = x3 & n15952 ;
  assign n15954 = n1251 & n9341 ;
  assign n15955 = n15954 ^ n420 ^ 1'b0 ;
  assign n15956 = n6104 | n10331 ;
  assign n15959 = n1353 & n8900 ;
  assign n15957 = ~n5110 & n7631 ;
  assign n15958 = ~n7305 & n15957 ;
  assign n15960 = n15959 ^ n15958 ^ 1'b0 ;
  assign n15961 = n10844 ^ n2844 ^ 1'b0 ;
  assign n15962 = n7454 & n14925 ;
  assign n15963 = n15962 ^ n5567 ^ 1'b0 ;
  assign n15964 = n15961 & n15963 ;
  assign n15965 = n3454 & ~n11013 ;
  assign n15966 = n9256 ^ n5259 ^ 1'b0 ;
  assign n15967 = n4112 ^ n942 ^ 1'b0 ;
  assign n15968 = n7783 | n9993 ;
  assign n15969 = n15968 ^ n14940 ^ 1'b0 ;
  assign n15970 = n2983 | n3626 ;
  assign n15971 = n8212 | n15970 ;
  assign n15972 = n2681 & ~n9095 ;
  assign n15973 = n15972 ^ n14116 ^ 1'b0 ;
  assign n15974 = ( n2354 & n5129 ) | ( n2354 & n13938 ) | ( n5129 & n13938 ) ;
  assign n15975 = n8748 ^ n380 ^ 1'b0 ;
  assign n15977 = ( n4671 & ~n7281 ) | ( n4671 & n12221 ) | ( ~n7281 & n12221 ) ;
  assign n15976 = n1694 | n15384 ;
  assign n15978 = n15977 ^ n15976 ^ 1'b0 ;
  assign n15979 = n14667 ^ n2310 ^ 1'b0 ;
  assign n15980 = ~n4495 & n15979 ;
  assign n15981 = n3729 | n4189 ;
  assign n15982 = n3729 & ~n15981 ;
  assign n15983 = n6211 ^ n4558 ^ 1'b0 ;
  assign n15984 = n15983 ^ n3237 ^ 1'b0 ;
  assign n15985 = ~n15982 & n15984 ;
  assign n15986 = n3705 & ~n3759 ;
  assign n15987 = n8644 & n15986 ;
  assign n15988 = n5859 & ~n15987 ;
  assign n15989 = n14573 ^ n2866 ^ 1'b0 ;
  assign n15990 = n9787 ^ n9234 ^ 1'b0 ;
  assign n15991 = n15989 | n15990 ;
  assign n15992 = n12986 ^ n5231 ^ 1'b0 ;
  assign n15993 = n15992 ^ n15897 ^ n9177 ;
  assign n15994 = n9185 ^ n4828 ^ 1'b0 ;
  assign n15995 = n1010 & ~n15994 ;
  assign n15996 = x47 & n15995 ;
  assign n15997 = n15996 ^ x43 ^ 1'b0 ;
  assign n15998 = n561 & ~n12524 ;
  assign n15999 = n8965 ^ n5285 ^ 1'b0 ;
  assign n16000 = n13113 & n14672 ;
  assign n16001 = n5828 & ~n15440 ;
  assign n16002 = n9940 & n16001 ;
  assign n16003 = n16002 ^ n3740 ^ 1'b0 ;
  assign n16004 = n8827 ^ n2660 ^ n785 ;
  assign n16005 = n8773 ^ n6224 ^ 1'b0 ;
  assign n16006 = n2052 & ~n2700 ;
  assign n16007 = n16006 ^ n2997 ^ 1'b0 ;
  assign n16008 = n16007 ^ n7160 ^ 1'b0 ;
  assign n16009 = n16008 ^ n4578 ^ n2475 ;
  assign n16010 = ~n12216 & n16009 ;
  assign n16011 = n16010 ^ n13413 ^ 1'b0 ;
  assign n16012 = n6948 & ~n9863 ;
  assign n16013 = n13561 & ~n16012 ;
  assign n16014 = n16011 & n16013 ;
  assign n16015 = n8497 ^ n2008 ^ n1507 ;
  assign n16016 = n15935 ^ n12512 ^ 1'b0 ;
  assign n16017 = n926 & ~n9162 ;
  assign n16018 = ~n7713 & n16017 ;
  assign n16019 = n4972 ^ n928 ^ 1'b0 ;
  assign n16020 = n15225 ^ n7390 ^ 1'b0 ;
  assign n16021 = n8359 ^ n3458 ^ 1'b0 ;
  assign n16022 = ~n6595 & n16021 ;
  assign n16023 = ~n10096 & n16022 ;
  assign n16024 = n6585 & n16023 ;
  assign n16025 = n16024 ^ n6506 ^ 1'b0 ;
  assign n16026 = n4949 | n11776 ;
  assign n16027 = ~n512 & n8875 ;
  assign n16028 = n16027 ^ n5303 ^ 1'b0 ;
  assign n16029 = ~n2289 & n3026 ;
  assign n16030 = n4318 & n16029 ;
  assign n16031 = n16030 ^ n9225 ^ 1'b0 ;
  assign n16032 = n16028 & ~n16031 ;
  assign n16033 = ~n5325 & n11951 ;
  assign n16034 = n14589 ^ n3649 ^ 1'b0 ;
  assign n16035 = ~n1704 & n16034 ;
  assign n16036 = n7567 & n16035 ;
  assign n16037 = n3251 & n16036 ;
  assign n16038 = n9280 ^ n8656 ^ 1'b0 ;
  assign n16039 = n11322 ^ n8792 ^ n1920 ;
  assign n16040 = n9165 | n11421 ;
  assign n16041 = n8700 | n16040 ;
  assign n16042 = n7750 ^ n2352 ^ 1'b0 ;
  assign n16043 = ~n425 & n11871 ;
  assign n16044 = n15672 & ~n16043 ;
  assign n16045 = n16044 ^ n747 ^ 1'b0 ;
  assign n16046 = ~n3095 & n9723 ;
  assign n16047 = n3842 & ~n16046 ;
  assign n16048 = n16047 ^ n6944 ^ 1'b0 ;
  assign n16049 = ~n6461 & n7009 ;
  assign n16050 = n16049 ^ n8503 ^ 1'b0 ;
  assign n16051 = n12592 & ~n16050 ;
  assign n16052 = n16051 ^ n2983 ^ 1'b0 ;
  assign n16053 = n3496 & n7341 ;
  assign n16054 = n16053 ^ n979 ^ 1'b0 ;
  assign n16055 = n3884 ^ n3795 ^ 1'b0 ;
  assign n16056 = n6827 ^ n5880 ^ 1'b0 ;
  assign n16057 = n16055 | n16056 ;
  assign n16058 = n1139 & ~n6055 ;
  assign n16059 = n10813 & n16058 ;
  assign n16060 = n16057 & ~n16059 ;
  assign n16061 = n361 | n5443 ;
  assign n16062 = n6548 & ~n16061 ;
  assign n16063 = n2887 | n16062 ;
  assign n16064 = n16063 ^ n4576 ^ 1'b0 ;
  assign n16065 = n8811 & ~n16064 ;
  assign n16066 = n10112 ^ n3479 ^ 1'b0 ;
  assign n16067 = n2443 & n16066 ;
  assign n16068 = n2466 & n16067 ;
  assign n16069 = n6365 & n16068 ;
  assign n16070 = n12279 ^ n552 ^ 1'b0 ;
  assign n16071 = n16069 | n16070 ;
  assign n16072 = x141 & n1886 ;
  assign n16073 = n14166 ^ n11628 ^ 1'b0 ;
  assign n16074 = ( n1252 & ~n16072 ) | ( n1252 & n16073 ) | ( ~n16072 & n16073 ) ;
  assign n16075 = ~n16071 & n16074 ;
  assign n16076 = n5134 ^ n1646 ^ n1477 ;
  assign n16077 = n16076 ^ n10717 ^ 1'b0 ;
  assign n16078 = n2466 & n4652 ;
  assign n16079 = n2343 & n16078 ;
  assign n16081 = n2185 & ~n14565 ;
  assign n16082 = n16081 ^ n10416 ^ 1'b0 ;
  assign n16080 = n13836 & n14131 ;
  assign n16083 = n16082 ^ n16080 ^ 1'b0 ;
  assign n16084 = ~n5077 & n5823 ;
  assign n16085 = n1111 & n16084 ;
  assign n16086 = n16085 ^ n12310 ^ 1'b0 ;
  assign n16087 = n7479 | n9702 ;
  assign n16088 = n16087 ^ x201 ^ 1'b0 ;
  assign n16089 = n12948 & ~n16088 ;
  assign n16090 = n2855 & n3052 ;
  assign n16091 = n9408 ^ n5953 ^ 1'b0 ;
  assign n16092 = ~n16090 & n16091 ;
  assign n16095 = x206 & n4118 ;
  assign n16096 = n16095 ^ n10077 ^ 1'b0 ;
  assign n16093 = n434 & n7641 ;
  assign n16094 = ~n2256 & n16093 ;
  assign n16097 = n16096 ^ n16094 ^ 1'b0 ;
  assign n16098 = ~n2791 & n3571 ;
  assign n16099 = n8903 ^ n8392 ^ 1'b0 ;
  assign n16100 = n703 | n16099 ;
  assign n16101 = n16100 ^ n6478 ^ 1'b0 ;
  assign n16102 = ~n5054 & n16101 ;
  assign n16103 = n2063 | n4111 ;
  assign n16104 = n16103 ^ n9793 ^ 1'b0 ;
  assign n16105 = n16102 & n16104 ;
  assign n16106 = n2081 & n7739 ;
  assign n16107 = n16106 ^ n9090 ^ n4957 ;
  assign n16108 = n8017 & n15844 ;
  assign n16109 = ~n8968 & n16108 ;
  assign n16111 = n7998 ^ n2450 ^ n858 ;
  assign n16110 = x75 & ~n1423 ;
  assign n16112 = n16111 ^ n16110 ^ 1'b0 ;
  assign n16113 = n14304 ^ n12619 ^ 1'b0 ;
  assign n16114 = ~n16112 & n16113 ;
  assign n16115 = n3198 | n5625 ;
  assign n16116 = n16115 ^ n15498 ^ 1'b0 ;
  assign n16117 = ~n4367 & n9982 ;
  assign n16118 = n2035 & n12777 ;
  assign n16119 = n13468 & ~n16118 ;
  assign n16120 = n12669 ^ n4509 ^ 1'b0 ;
  assign n16121 = n13157 ^ n5775 ^ 1'b0 ;
  assign n16122 = n10858 & ~n16121 ;
  assign n16124 = n3874 | n4674 ;
  assign n16125 = n16124 ^ n8283 ^ 1'b0 ;
  assign n16126 = n372 & ~n4267 ;
  assign n16127 = ~n16125 & n16126 ;
  assign n16128 = n1533 | n16127 ;
  assign n16123 = ~n15171 & n16048 ;
  assign n16129 = n16128 ^ n16123 ^ 1'b0 ;
  assign n16130 = n12452 & n13738 ;
  assign n16131 = ~n2910 & n4586 ;
  assign n16132 = ( x18 & n14208 ) | ( x18 & n16131 ) | ( n14208 & n16131 ) ;
  assign n16133 = n5021 & n6207 ;
  assign n16134 = n16133 ^ n8223 ^ 1'b0 ;
  assign n16135 = ~n5144 & n16134 ;
  assign n16137 = n5047 ^ n3817 ^ 1'b0 ;
  assign n16138 = ~n7301 & n16137 ;
  assign n16136 = n1856 & n5793 ;
  assign n16139 = n16138 ^ n16136 ^ 1'b0 ;
  assign n16140 = n972 & n13062 ;
  assign n16141 = n3263 & n9688 ;
  assign n16142 = n16140 & n16141 ;
  assign n16143 = n4147 | n16142 ;
  assign n16144 = n16143 ^ n8123 ^ 1'b0 ;
  assign n16145 = n13907 ^ n4020 ^ 1'b0 ;
  assign n16146 = n11532 & n16145 ;
  assign n16147 = ~n2193 & n2652 ;
  assign n16148 = n1877 & n16147 ;
  assign n16150 = n4361 & ~n11937 ;
  assign n16149 = x176 & n12362 ;
  assign n16151 = n16150 ^ n16149 ^ 1'b0 ;
  assign n16152 = n4432 & ~n10334 ;
  assign n16153 = n16152 ^ n8631 ^ 1'b0 ;
  assign n16154 = ~n16151 & n16153 ;
  assign n16155 = n16154 ^ n897 ^ 1'b0 ;
  assign n16156 = ~n16148 & n16155 ;
  assign n16157 = n5898 & n11074 ;
  assign n16158 = n14924 ^ n766 ^ 1'b0 ;
  assign n16159 = n3479 ^ n352 ^ 1'b0 ;
  assign n16160 = n6891 & n16159 ;
  assign n16161 = x153 & ~n16160 ;
  assign n16162 = n11268 & n16161 ;
  assign n16163 = n16162 ^ n3628 ^ 1'b0 ;
  assign n16164 = n15539 ^ n9585 ^ 1'b0 ;
  assign n16165 = n5330 & ~n12346 ;
  assign n16166 = n16165 ^ n8127 ^ 1'b0 ;
  assign n16167 = n5311 ^ n2093 ^ 1'b0 ;
  assign n16168 = ~n11519 & n16167 ;
  assign n16169 = n13628 ^ n13173 ^ 1'b0 ;
  assign n16170 = ~n10229 & n10666 ;
  assign n16171 = n7164 ^ n2187 ^ 1'b0 ;
  assign n16172 = n7527 ^ n7181 ^ 1'b0 ;
  assign n16173 = x3 & ~n5440 ;
  assign n16174 = ~n5907 & n16173 ;
  assign n16175 = ~n2082 & n14876 ;
  assign n16176 = n16174 & n16175 ;
  assign n16177 = ~n6840 & n8888 ;
  assign n16178 = n2110 | n12519 ;
  assign n16179 = n12956 & ~n16178 ;
  assign n16180 = ~n7323 & n10316 ;
  assign n16181 = n16180 ^ n6167 ^ 1'b0 ;
  assign n16184 = n2065 & n8448 ;
  assign n16182 = n5512 | n12131 ;
  assign n16183 = n14089 & ~n16182 ;
  assign n16185 = n16184 ^ n16183 ^ 1'b0 ;
  assign n16186 = ~n4518 & n8481 ;
  assign n16187 = n14961 & n16186 ;
  assign n16188 = n16187 ^ n7738 ^ 1'b0 ;
  assign n16189 = n9959 ^ n2826 ^ 1'b0 ;
  assign n16190 = ( ~n4676 & n13759 ) | ( ~n4676 & n16189 ) | ( n13759 & n16189 ) ;
  assign n16191 = n4695 & ~n10523 ;
  assign n16192 = n5002 & n8444 ;
  assign n16193 = n4378 | n16192 ;
  assign n16194 = n8850 | n16193 ;
  assign n16195 = n16194 ^ n11057 ^ 1'b0 ;
  assign n16196 = n9477 ^ n894 ^ 1'b0 ;
  assign n16197 = n1832 & n16196 ;
  assign n16198 = n16197 ^ n8768 ^ 1'b0 ;
  assign n16199 = n16198 ^ n8008 ^ 1'b0 ;
  assign n16200 = ~n16195 & n16199 ;
  assign n16201 = ~n11012 & n16200 ;
  assign n16202 = n16191 & n16201 ;
  assign n16203 = n5155 ^ n4619 ^ 1'b0 ;
  assign n16204 = n3045 & ~n16203 ;
  assign n16205 = n4868 ^ n2526 ^ 1'b0 ;
  assign n16206 = n16204 & n16205 ;
  assign n16208 = n1080 | n1997 ;
  assign n16207 = ~x73 & n15039 ;
  assign n16209 = n16208 ^ n16207 ^ 1'b0 ;
  assign n16210 = n1775 & ~n14604 ;
  assign n16211 = ~n2469 & n16210 ;
  assign n16212 = n4075 | n16211 ;
  assign n16213 = n16212 ^ n7070 ^ 1'b0 ;
  assign n16214 = n5922 & n16213 ;
  assign n16215 = n7688 ^ n3229 ^ 1'b0 ;
  assign n16216 = n1237 & ~n16215 ;
  assign n16217 = n16216 ^ n11597 ^ 1'b0 ;
  assign n16218 = n15777 & n16217 ;
  assign n16219 = n1018 & n6420 ;
  assign n16220 = n11392 ^ n1617 ^ 1'b0 ;
  assign n16221 = x130 & ~n16220 ;
  assign n16222 = ~n1537 & n15507 ;
  assign n16223 = n16221 & n16222 ;
  assign n16224 = n16223 ^ n3431 ^ 1'b0 ;
  assign n16225 = n3774 & ~n16224 ;
  assign n16226 = ~n9483 & n16225 ;
  assign n16227 = n2304 & n13555 ;
  assign n16228 = n16227 ^ n3524 ^ 1'b0 ;
  assign n16229 = ~n3060 & n7580 ;
  assign n16230 = n3520 ^ n2582 ^ 1'b0 ;
  assign n16231 = n2804 | n16230 ;
  assign n16232 = n16231 ^ n12988 ^ 1'b0 ;
  assign n16233 = n8792 ^ n4483 ^ 1'b0 ;
  assign n16234 = n16233 ^ n2793 ^ 1'b0 ;
  assign n16235 = n11000 ^ n5293 ^ 1'b0 ;
  assign n16236 = n307 | n16235 ;
  assign n16237 = n3153 | n6963 ;
  assign n16238 = n1651 & ~n16237 ;
  assign n16239 = n3709 | n16238 ;
  assign n16240 = n16239 ^ n9156 ^ 1'b0 ;
  assign n16241 = n14554 ^ n13315 ^ n6357 ;
  assign n16242 = ~n5665 & n10798 ;
  assign n16243 = n10835 ^ n8175 ^ 1'b0 ;
  assign n16244 = ~n6553 & n16243 ;
  assign n16245 = ~n7149 & n16244 ;
  assign n16246 = n3292 | n8960 ;
  assign n16247 = x56 & n538 ;
  assign n16248 = ~x56 & n16247 ;
  assign n16249 = n6034 & n16248 ;
  assign n16250 = n16249 ^ n6147 ^ 1'b0 ;
  assign n16251 = n761 | n858 ;
  assign n16252 = n858 & ~n16251 ;
  assign n16253 = n1353 & ~n16252 ;
  assign n16254 = ~n1353 & n16253 ;
  assign n16255 = x189 & ~n16254 ;
  assign n16256 = ~x189 & n16255 ;
  assign n16257 = n972 | n1243 ;
  assign n16258 = n972 & ~n16257 ;
  assign n16259 = x250 & ~n16258 ;
  assign n16260 = n16258 & n16259 ;
  assign n16261 = n16256 | n16260 ;
  assign n16262 = n16256 & ~n16261 ;
  assign n16263 = ~n3521 & n5164 ;
  assign n16264 = n16263 ^ n4705 ^ 1'b0 ;
  assign n16265 = n16262 & n16264 ;
  assign n16266 = n2089 & ~n4580 ;
  assign n16267 = ~n2089 & n16266 ;
  assign n16268 = n6605 ^ n4268 ^ 1'b0 ;
  assign n16269 = n4293 & ~n16268 ;
  assign n16270 = ~n1474 & n16269 ;
  assign n16271 = n1474 & n16270 ;
  assign n16272 = n1847 & n16271 ;
  assign n16273 = x15 & ~n2470 ;
  assign n16274 = ~x15 & n16273 ;
  assign n16275 = n3778 | n3825 ;
  assign n16276 = n16274 & ~n16275 ;
  assign n16277 = ~n16272 & n16276 ;
  assign n16278 = n16277 ^ n4831 ^ 1'b0 ;
  assign n16279 = n16267 | n16278 ;
  assign n16280 = n16265 & ~n16279 ;
  assign n16281 = n16280 ^ n14077 ^ 1'b0 ;
  assign n16282 = ~n16250 & n16281 ;
  assign n16283 = n11274 ^ x254 ^ 1'b0 ;
  assign n16284 = n10633 & n16283 ;
  assign n16285 = n5278 ^ n1453 ^ 1'b0 ;
  assign n16286 = n1290 | n1857 ;
  assign n16287 = n16286 ^ n5990 ^ 1'b0 ;
  assign n16288 = n3567 & n16287 ;
  assign n16289 = n15316 | n16288 ;
  assign n16290 = ~n505 & n4242 ;
  assign n16291 = ~n4024 & n16290 ;
  assign n16292 = n12425 ^ n6203 ^ 1'b0 ;
  assign n16293 = n5048 & n16292 ;
  assign n16294 = n2658 & n3713 ;
  assign n16295 = ~n16293 & n16294 ;
  assign n16296 = n12804 & n14955 ;
  assign n16297 = ~n9565 & n16296 ;
  assign n16298 = n10733 & ~n16297 ;
  assign n16299 = ~n614 & n12241 ;
  assign n16300 = n16299 ^ n6343 ^ 1'b0 ;
  assign n16301 = ~n11187 & n12033 ;
  assign n16302 = n552 & ~n1062 ;
  assign n16303 = n16302 ^ n717 ^ 1'b0 ;
  assign n16304 = ~n4818 & n6399 ;
  assign n16305 = ~n744 & n16304 ;
  assign n16306 = n16305 ^ n10281 ^ 1'b0 ;
  assign n16307 = ~n16303 & n16306 ;
  assign n16308 = n2794 | n7112 ;
  assign n16309 = n16308 ^ n3604 ^ 1'b0 ;
  assign n16310 = ~n503 & n1991 ;
  assign n16311 = n2517 & n8438 ;
  assign n16312 = n16311 ^ n10216 ^ n5796 ;
  assign n16313 = n16053 | n16312 ;
  assign n16314 = n13679 ^ n9880 ^ 1'b0 ;
  assign n16315 = n485 & ~n5275 ;
  assign n16316 = n10116 & ~n16315 ;
  assign n16317 = n16316 ^ n3033 ^ 1'b0 ;
  assign n16318 = ~n13710 & n15967 ;
  assign n16319 = n12972 ^ n8293 ^ 1'b0 ;
  assign n16320 = n8438 & ~n16319 ;
  assign n16321 = n16320 ^ n468 ^ 1'b0 ;
  assign n16322 = n6978 ^ n5238 ^ 1'b0 ;
  assign n16323 = n679 | n9327 ;
  assign n16324 = n16322 & ~n16323 ;
  assign n16325 = n9543 ^ n2669 ^ 1'b0 ;
  assign n16326 = ~n2776 & n16325 ;
  assign n16327 = n1447 & n16326 ;
  assign n16328 = n16327 ^ n1521 ^ 1'b0 ;
  assign n16329 = n800 | n2731 ;
  assign n16330 = n3928 | n16329 ;
  assign n16331 = ~n12157 & n16330 ;
  assign n16332 = ~n8907 & n16331 ;
  assign n16333 = n5490 & ~n16332 ;
  assign n16334 = n3071 & ~n7835 ;
  assign n16335 = n16334 ^ n12392 ^ 1'b0 ;
  assign n16336 = n10107 ^ n7345 ^ 1'b0 ;
  assign n16337 = ~n6026 & n9276 ;
  assign n16338 = n6343 & ~n16337 ;
  assign n16339 = n16338 ^ n1046 ^ 1'b0 ;
  assign n16340 = n11619 ^ n7783 ^ n6780 ;
  assign n16341 = n6665 & ~n16340 ;
  assign n16342 = n16341 ^ n8451 ^ 1'b0 ;
  assign n16343 = n2283 & n4389 ;
  assign n16344 = n9000 | n15665 ;
  assign n16346 = ( ~n936 & n6209 ) | ( ~n936 & n8048 ) | ( n6209 & n8048 ) ;
  assign n16347 = n8045 & ~n16346 ;
  assign n16345 = ~n575 & n5192 ;
  assign n16348 = n16347 ^ n16345 ^ 1'b0 ;
  assign n16349 = n6154 | n16348 ;
  assign n16350 = n6368 | n11972 ;
  assign n16351 = n16350 ^ n4793 ^ 1'b0 ;
  assign n16352 = ~n5401 & n14496 ;
  assign n16353 = n10555 & n16352 ;
  assign n16354 = ~n6466 & n9942 ;
  assign n16355 = ~n1450 & n16354 ;
  assign n16356 = n9188 ^ n4753 ^ 1'b0 ;
  assign n16357 = ~n13245 & n16356 ;
  assign n16358 = n10725 & n16357 ;
  assign n16359 = n16358 ^ n4753 ^ 1'b0 ;
  assign n16360 = n6478 & n7400 ;
  assign n16361 = n2014 & n16360 ;
  assign n16362 = n3608 ^ n1822 ^ 1'b0 ;
  assign n16363 = n9659 & ~n12434 ;
  assign n16364 = n3242 & ~n11096 ;
  assign n16365 = n956 & ~n7347 ;
  assign n16367 = n11675 & ~n14436 ;
  assign n16366 = x128 & ~n1703 ;
  assign n16368 = n16367 ^ n16366 ^ 1'b0 ;
  assign n16369 = n988 | n1919 ;
  assign n16370 = n6562 & ~n16369 ;
  assign n16371 = n2455 & ~n16370 ;
  assign n16372 = n8574 | n16371 ;
  assign n16373 = n2293 | n16372 ;
  assign n16374 = n4668 ^ n4130 ^ 1'b0 ;
  assign n16375 = x206 & ~n16374 ;
  assign n16376 = ~n5217 & n5845 ;
  assign n16377 = n10396 & ~n16376 ;
  assign n16378 = n4350 | n16377 ;
  assign n16379 = n653 & ~n4223 ;
  assign n16382 = n4211 | n8485 ;
  assign n16383 = n7298 | n16382 ;
  assign n16384 = n16383 ^ n3667 ^ 1'b0 ;
  assign n16381 = n1080 & ~n10756 ;
  assign n16385 = n16384 ^ n16381 ^ 1'b0 ;
  assign n16380 = n8823 & ~n13657 ;
  assign n16386 = n16385 ^ n16380 ^ 1'b0 ;
  assign n16387 = n2044 & n3811 ;
  assign n16388 = n16387 ^ n10646 ^ 1'b0 ;
  assign n16389 = n15892 & ~n16388 ;
  assign n16390 = n456 | n2672 ;
  assign n16391 = n8883 & n16390 ;
  assign n16392 = n3895 & n16391 ;
  assign n16393 = n15421 & n16392 ;
  assign n16394 = n8130 ^ n2190 ^ 1'b0 ;
  assign n16395 = ~n6682 & n16394 ;
  assign n16396 = n6572 & n11122 ;
  assign n16397 = n16396 ^ n7687 ^ n5418 ;
  assign n16398 = ~n4329 & n8072 ;
  assign n16399 = ~n9404 & n16398 ;
  assign n16400 = n13256 & n16399 ;
  assign n16405 = n2682 ^ n2157 ^ 1'b0 ;
  assign n16406 = ~n5215 & n16405 ;
  assign n16401 = n11218 ^ n7856 ^ 1'b0 ;
  assign n16402 = n1564 & n16401 ;
  assign n16403 = n16402 ^ n5945 ^ 1'b0 ;
  assign n16404 = n14523 & ~n16403 ;
  assign n16407 = n16406 ^ n16404 ^ 1'b0 ;
  assign n16408 = n6378 | n10014 ;
  assign n16409 = x192 & ~n16408 ;
  assign n16410 = n10804 ^ n4350 ^ 1'b0 ;
  assign n16411 = n2961 ^ n937 ^ 1'b0 ;
  assign n16412 = n11335 & ~n16411 ;
  assign n16413 = n9703 ^ n8365 ^ 1'b0 ;
  assign n16414 = ~n11596 & n16413 ;
  assign n16415 = n14007 & n16414 ;
  assign n16416 = n9477 ^ n7237 ^ 1'b0 ;
  assign n16417 = n16416 ^ n10511 ^ n5864 ;
  assign n16418 = n11900 ^ n11206 ^ 1'b0 ;
  assign n16419 = n1990 & n16418 ;
  assign n16420 = n16419 ^ n4976 ^ 1'b0 ;
  assign n16421 = n16420 ^ n9560 ^ 1'b0 ;
  assign n16422 = x252 & ~n3842 ;
  assign n16423 = n16422 ^ n11177 ^ 1'b0 ;
  assign n16424 = n9989 | n16423 ;
  assign n16425 = n955 & ~n5874 ;
  assign n16426 = ~n11147 & n16425 ;
  assign n16427 = n16426 ^ n9406 ^ n3636 ;
  assign n16428 = x25 | n5635 ;
  assign n16429 = n16428 ^ n16329 ^ 1'b0 ;
  assign n16430 = ~n10395 & n16429 ;
  assign n16431 = n16430 ^ n9363 ^ 1'b0 ;
  assign n16432 = n12843 & ~n16431 ;
  assign n16433 = n10084 ^ n3870 ^ 1'b0 ;
  assign n16434 = n16432 & ~n16433 ;
  assign n16435 = n13794 ^ n5091 ^ 1'b0 ;
  assign n16436 = n13829 | n16435 ;
  assign n16437 = n13884 ^ n8507 ^ 1'b0 ;
  assign n16438 = n1814 | n1900 ;
  assign n16439 = n16438 ^ n9991 ^ 1'b0 ;
  assign n16440 = ~n1740 & n16439 ;
  assign n16441 = ( ~x141 & n1724 ) | ( ~x141 & n2663 ) | ( n1724 & n2663 ) ;
  assign n16442 = n7733 & ~n16441 ;
  assign n16443 = ~n1048 & n16442 ;
  assign n16445 = n774 & n3388 ;
  assign n16444 = n461 & ~n5290 ;
  assign n16446 = n16445 ^ n16444 ^ 1'b0 ;
  assign n16447 = n887 & ~n16099 ;
  assign n16448 = n3430 & n16447 ;
  assign n16449 = n3252 & ~n16448 ;
  assign n16450 = n5337 | n11856 ;
  assign n16451 = n16450 ^ n8663 ^ 1'b0 ;
  assign n16452 = n2018 & ~n16451 ;
  assign n16453 = n2210 | n7469 ;
  assign n16454 = n12777 & ~n16453 ;
  assign n16455 = n16454 ^ n747 ^ 1'b0 ;
  assign n16456 = n12071 & n16455 ;
  assign n16457 = n13576 ^ n1427 ^ 1'b0 ;
  assign n16458 = n7536 | n13924 ;
  assign n16459 = n16458 ^ n2185 ^ 1'b0 ;
  assign n16460 = x14 & ~n1156 ;
  assign n16461 = n3578 ^ n820 ^ 1'b0 ;
  assign n16462 = n16460 & n16461 ;
  assign n16463 = n1770 & ~n5490 ;
  assign n16464 = ~n2264 & n11708 ;
  assign n16465 = ~n1654 & n16464 ;
  assign n16466 = n13727 & n16465 ;
  assign n16467 = n3060 & ~n10404 ;
  assign n16468 = ~n10726 & n16467 ;
  assign n16469 = ~n9898 & n13325 ;
  assign n16470 = n5489 ^ n1176 ^ 1'b0 ;
  assign n16471 = n6322 & ~n14871 ;
  assign n16472 = n16471 ^ n2980 ^ 1'b0 ;
  assign n16473 = n10939 | n16472 ;
  assign n16474 = n16472 & ~n16473 ;
  assign n16475 = n16474 ^ n14087 ^ 1'b0 ;
  assign n16476 = n11066 & n16475 ;
  assign n16477 = n11252 & n16476 ;
  assign n16478 = n3893 | n5222 ;
  assign n16479 = ( ~n7341 & n7851 ) | ( ~n7341 & n16478 ) | ( n7851 & n16478 ) ;
  assign n16480 = n7362 ^ x157 ^ 1'b0 ;
  assign n16481 = n8072 & n16480 ;
  assign n16482 = n787 & n16481 ;
  assign n16483 = ~n6401 & n16482 ;
  assign n16484 = n10275 | n12763 ;
  assign n16485 = n16484 ^ n1378 ^ 1'b0 ;
  assign n16486 = n4538 ^ n448 ^ 1'b0 ;
  assign n16487 = n1291 & ~n12242 ;
  assign n16488 = n16487 ^ n13509 ^ 1'b0 ;
  assign n16489 = n3624 ^ n690 ^ 1'b0 ;
  assign n16490 = n2350 | n16489 ;
  assign n16491 = n9121 | n14376 ;
  assign n16492 = n16491 ^ n7414 ^ 1'b0 ;
  assign n16494 = n1328 & ~n13156 ;
  assign n16495 = n16494 ^ n2970 ^ 1'b0 ;
  assign n16496 = n16495 ^ n1472 ^ 1'b0 ;
  assign n16497 = n7604 & ~n16496 ;
  assign n16493 = n8312 ^ n6451 ^ 1'b0 ;
  assign n16498 = n16497 ^ n16493 ^ 1'b0 ;
  assign n16499 = n14955 ^ n4645 ^ 1'b0 ;
  assign n16500 = ~n7117 & n16499 ;
  assign n16501 = n4260 ^ n2120 ^ 1'b0 ;
  assign n16502 = n3979 | n16501 ;
  assign n16503 = n2611 | n16502 ;
  assign n16504 = n6052 & ~n16503 ;
  assign n16505 = n2590 | n16504 ;
  assign n16506 = n10314 ^ n7609 ^ 1'b0 ;
  assign n16507 = n5587 & n6025 ;
  assign n16508 = n16507 ^ n2395 ^ 1'b0 ;
  assign n16509 = n16506 & ~n16508 ;
  assign n16510 = n6571 & n16509 ;
  assign n16511 = n9944 | n16510 ;
  assign n16512 = n4169 | n16511 ;
  assign n16513 = n816 & n3807 ;
  assign n16514 = n11256 & n16513 ;
  assign n16515 = n1477 | n16514 ;
  assign n16516 = n2575 ^ n2426 ^ 1'b0 ;
  assign n16517 = n2647 & n5867 ;
  assign n16518 = n15959 ^ n6985 ^ 1'b0 ;
  assign n16519 = ~n928 & n2431 ;
  assign n16520 = n2185 & ~n3415 ;
  assign n16521 = n12016 ^ n2794 ^ 1'b0 ;
  assign n16522 = n662 & n16521 ;
  assign n16523 = n6080 & n16522 ;
  assign n16524 = ~n10890 & n16523 ;
  assign n16525 = ~n16520 & n16524 ;
  assign n16526 = n385 & ~n3445 ;
  assign n16527 = n3445 & n16526 ;
  assign n16528 = n16527 ^ n16150 ^ 1'b0 ;
  assign n16529 = ~n5034 & n9007 ;
  assign n16530 = ~n9007 & n16529 ;
  assign n16531 = x186 & ~n16530 ;
  assign n16532 = n5386 & n16531 ;
  assign n16533 = ~n16528 & n16532 ;
  assign n16534 = n2466 & ~n3436 ;
  assign n16535 = ~n2466 & n16534 ;
  assign n16541 = x235 & n561 ;
  assign n16542 = ~n561 & n16541 ;
  assign n16543 = n16542 ^ n401 ^ 1'b0 ;
  assign n16536 = n1723 | n2179 ;
  assign n16537 = n2179 & ~n16536 ;
  assign n16538 = n1514 & ~n16537 ;
  assign n16539 = ~n1514 & n16538 ;
  assign n16540 = n14545 & ~n16539 ;
  assign n16544 = n16543 ^ n16540 ^ 1'b0 ;
  assign n16545 = ~n16535 & n16544 ;
  assign n16546 = n14531 ^ n11798 ^ 1'b0 ;
  assign n16547 = n11394 | n16546 ;
  assign n16548 = n16547 ^ n15368 ^ 1'b0 ;
  assign n16549 = n502 & n2702 ;
  assign n16550 = n16549 ^ n4675 ^ 1'b0 ;
  assign n16551 = n16550 ^ n11683 ^ 1'b0 ;
  assign n16552 = ~n10509 & n16551 ;
  assign n16553 = n5126 ^ n3742 ^ 1'b0 ;
  assign n16554 = n9550 & ~n10561 ;
  assign n16555 = ~n4229 & n16554 ;
  assign n16556 = n14116 ^ n7720 ^ 1'b0 ;
  assign n16557 = n1126 | n14977 ;
  assign n16558 = n13267 ^ n12061 ^ n2164 ;
  assign n16559 = n10744 | n15018 ;
  assign n16560 = n16558 | n16559 ;
  assign n16561 = n10608 | n12559 ;
  assign n16562 = n5944 & n16561 ;
  assign n16563 = n11057 ^ n5943 ^ 1'b0 ;
  assign n16564 = n7367 ^ n5262 ^ 1'b0 ;
  assign n16565 = n3243 & ~n9252 ;
  assign n16566 = n5586 ^ n1922 ^ 1'b0 ;
  assign n16567 = ~n16565 & n16566 ;
  assign n16568 = ( n1837 & ~n9553 ) | ( n1837 & n9930 ) | ( ~n9553 & n9930 ) ;
  assign n16569 = n8493 & n16568 ;
  assign n16570 = n11647 ^ n8008 ^ 1'b0 ;
  assign n16571 = n12760 | n16570 ;
  assign n16572 = n5984 ^ n859 ^ 1'b0 ;
  assign n16573 = ( n937 & n7683 ) | ( n937 & ~n16572 ) | ( n7683 & ~n16572 ) ;
  assign n16574 = n16573 ^ n12756 ^ x20 ;
  assign n16575 = n2809 | n9099 ;
  assign n16576 = n16575 ^ n8518 ^ 1'b0 ;
  assign n16577 = n14354 ^ n5463 ^ 1'b0 ;
  assign n16578 = n6252 | n16577 ;
  assign n16579 = n4724 | n9932 ;
  assign n16580 = n2807 & n4380 ;
  assign n16581 = ( n4424 & n13802 ) | ( n4424 & ~n16580 ) | ( n13802 & ~n16580 ) ;
  assign n16582 = n9363 & n10922 ;
  assign n16583 = n3287 & ~n4980 ;
  assign n16584 = ~n16582 & n16583 ;
  assign n16585 = n2061 | n15013 ;
  assign n16586 = n7791 | n16585 ;
  assign n16587 = n5978 ^ n1165 ^ 1'b0 ;
  assign n16588 = n16586 & ~n16587 ;
  assign n16589 = n15011 ^ n5163 ^ 1'b0 ;
  assign n16590 = n5275 & n16589 ;
  assign n16591 = n6455 ^ n2856 ^ 1'b0 ;
  assign n16592 = n6945 & ~n16591 ;
  assign n16593 = ~n9177 & n16592 ;
  assign n16594 = n8722 & n16376 ;
  assign n16595 = n16594 ^ n3189 ^ 1'b0 ;
  assign n16596 = n9299 & n16595 ;
  assign n16597 = n16463 ^ n1597 ^ 1'b0 ;
  assign n16598 = n1569 ^ n919 ^ 1'b0 ;
  assign n16599 = n14287 | n16598 ;
  assign n16600 = n16599 ^ n6661 ^ 1'b0 ;
  assign n16601 = n5707 ^ n3979 ^ 1'b0 ;
  assign n16602 = n16601 ^ n9344 ^ 1'b0 ;
  assign n16603 = n4118 ^ n354 ^ 1'b0 ;
  assign n16604 = n1334 & ~n16603 ;
  assign n16605 = n11785 ^ n7680 ^ 1'b0 ;
  assign n16606 = x55 & ~n16605 ;
  assign n16607 = n5530 ^ n3393 ^ 1'b0 ;
  assign n16608 = n1341 & ~n6313 ;
  assign n16609 = n16607 | n16608 ;
  assign n16610 = n2161 & ~n16609 ;
  assign n16611 = n2085 | n8055 ;
  assign n16612 = x112 & ~n16611 ;
  assign n16613 = n12592 ^ n305 ^ 1'b0 ;
  assign n16614 = ~n16612 & n16613 ;
  assign n16615 = n16610 & n16614 ;
  assign n16616 = n6012 ^ n4421 ^ 1'b0 ;
  assign n16617 = n2395 & n3370 ;
  assign n16618 = n2826 ^ n2495 ^ 1'b0 ;
  assign n16619 = x43 & n16618 ;
  assign n16623 = n3622 ^ n1186 ^ 1'b0 ;
  assign n16624 = x157 & n16623 ;
  assign n16625 = ~n1149 & n16624 ;
  assign n16626 = n16625 ^ n1525 ^ 1'b0 ;
  assign n16627 = n4645 & n16626 ;
  assign n16628 = n11621 & n16627 ;
  assign n16620 = n5176 ^ n3248 ^ 1'b0 ;
  assign n16621 = n10310 & ~n16620 ;
  assign n16622 = n5493 & n16621 ;
  assign n16629 = n16628 ^ n16622 ^ 1'b0 ;
  assign n16630 = n3318 & ~n10795 ;
  assign n16631 = n16630 ^ n10188 ^ 1'b0 ;
  assign n16632 = n2630 & n16631 ;
  assign n16633 = n5817 | n14589 ;
  assign n16634 = n9554 & n11131 ;
  assign n16635 = n16634 ^ n3140 ^ 1'b0 ;
  assign n16636 = n5987 | n15909 ;
  assign n16637 = n6964 & n14948 ;
  assign n16638 = ~n824 & n1791 ;
  assign n16639 = n5360 & n16638 ;
  assign n16640 = n1688 & n16639 ;
  assign n16641 = n8948 ^ n1130 ^ 1'b0 ;
  assign n16642 = ~n3381 & n16641 ;
  assign n16643 = n16597 ^ n12444 ^ 1'b0 ;
  assign n16644 = n7634 | n16643 ;
  assign n16645 = n651 | n15649 ;
  assign n16646 = ( n888 & ~n1865 ) | ( n888 & n13273 ) | ( ~n1865 & n13273 ) ;
  assign n16647 = n3020 ^ x87 ^ 1'b0 ;
  assign n16648 = n16647 ^ n9020 ^ 1'b0 ;
  assign n16649 = n1618 | n3148 ;
  assign n16650 = ~n12345 & n16649 ;
  assign n16651 = ~n6020 & n16650 ;
  assign n16652 = ~n4801 & n4920 ;
  assign n16653 = n16652 ^ n12753 ^ 1'b0 ;
  assign n16654 = n3469 & ~n16653 ;
  assign n16655 = n9990 & n13115 ;
  assign n16656 = ~n16654 & n16655 ;
  assign n16657 = n1968 & n12440 ;
  assign n16658 = x182 & ~n1397 ;
  assign n16659 = ~n1236 & n16658 ;
  assign n16660 = n16659 ^ n10682 ^ 1'b0 ;
  assign n16661 = n2853 | n6790 ;
  assign n16662 = n6790 & ~n16661 ;
  assign n16663 = n969 & n16662 ;
  assign n16664 = n16663 ^ n3895 ^ 1'b0 ;
  assign n16665 = n16664 ^ n10155 ^ 1'b0 ;
  assign n16666 = ~n3986 & n16665 ;
  assign n16667 = n4116 & ~n6756 ;
  assign n16668 = n9778 & n16667 ;
  assign n16669 = ~n8280 & n16668 ;
  assign n16670 = n14798 ^ n12595 ^ 1'b0 ;
  assign n16671 = ~n16669 & n16670 ;
  assign n16672 = n12729 ^ n3143 ^ 1'b0 ;
  assign n16673 = n5530 & n15928 ;
  assign n16674 = n16673 ^ n3281 ^ 1'b0 ;
  assign n16675 = n3021 | n4982 ;
  assign n16676 = n16675 ^ n2959 ^ 1'b0 ;
  assign n16677 = n15537 ^ n3334 ^ 1'b0 ;
  assign n16678 = n8408 & n16677 ;
  assign n16679 = n16678 ^ n3558 ^ 1'b0 ;
  assign n16680 = ~n2009 & n16679 ;
  assign n16681 = n11105 ^ n2175 ^ 1'b0 ;
  assign n16682 = x76 & n16681 ;
  assign n16683 = n11370 & n16682 ;
  assign n16684 = n1724 | n4318 ;
  assign n16685 = ~n12735 & n16684 ;
  assign n16686 = n16685 ^ x166 ^ 1'b0 ;
  assign n16687 = n15739 ^ n2185 ^ 1'b0 ;
  assign n16688 = n6597 & ~n16687 ;
  assign n16689 = n4308 & n15841 ;
  assign n16690 = n4917 & ~n8954 ;
  assign n16691 = n16690 ^ n14524 ^ 1'b0 ;
  assign n16692 = n2989 & ~n16691 ;
  assign n16693 = n1336 & n14497 ;
  assign n16694 = ~n5192 & n16693 ;
  assign n16695 = n12389 ^ n2616 ^ 1'b0 ;
  assign n16696 = ~n1324 & n3718 ;
  assign n16697 = n16696 ^ n860 ^ 1'b0 ;
  assign n16698 = n13585 & n16697 ;
  assign n16699 = n9720 ^ n6816 ^ 1'b0 ;
  assign n16700 = n1661 & ~n6104 ;
  assign n16701 = n16700 ^ x6 ^ 1'b0 ;
  assign n16702 = n6953 | n8468 ;
  assign n16703 = n16702 ^ n4532 ^ 1'b0 ;
  assign n16704 = n8632 ^ n2148 ^ 1'b0 ;
  assign n16705 = n8545 & ~n16704 ;
  assign n16706 = n2543 & n4587 ;
  assign n16707 = ~n2626 & n16706 ;
  assign n16708 = n16707 ^ n14589 ^ 1'b0 ;
  assign n16709 = ~n485 & n16708 ;
  assign n16710 = n10123 & ~n16709 ;
  assign n16711 = n11587 & n16710 ;
  assign n16712 = n5812 ^ n3331 ^ 1'b0 ;
  assign n16713 = n2083 | n12525 ;
  assign n16714 = n7042 ^ n4122 ^ 1'b0 ;
  assign n16715 = n1765 & ~n16714 ;
  assign n16716 = ~n10674 & n16715 ;
  assign n16717 = n5090 & ~n7597 ;
  assign n16718 = n16717 ^ n14090 ^ n2868 ;
  assign n16719 = n16111 ^ n1638 ^ 1'b0 ;
  assign n16720 = ~n8332 & n16719 ;
  assign n16721 = n16720 ^ n3940 ^ 1'b0 ;
  assign n16722 = n8841 ^ n4934 ^ 1'b0 ;
  assign n16723 = n9477 ^ n4179 ^ 1'b0 ;
  assign n16724 = n16722 | n16723 ;
  assign n16725 = n2486 | n5564 ;
  assign n16726 = n4274 ^ n533 ^ 1'b0 ;
  assign n16727 = n8956 | n11368 ;
  assign n16728 = n13793 ^ n4903 ^ 1'b0 ;
  assign n16729 = n16728 ^ n519 ^ 1'b0 ;
  assign n16730 = n16729 ^ n4814 ^ 1'b0 ;
  assign n16731 = n5018 ^ x95 ^ 1'b0 ;
  assign n16732 = n4161 & n5950 ;
  assign n16733 = n16732 ^ n6798 ^ 1'b0 ;
  assign n16734 = n2588 & n16733 ;
  assign n16735 = ~n13059 & n14882 ;
  assign n16736 = ( n16731 & n16734 ) | ( n16731 & n16735 ) | ( n16734 & n16735 ) ;
  assign n16737 = n5571 | n12948 ;
  assign n16739 = n3181 & ~n4933 ;
  assign n16738 = n4678 ^ n1393 ^ 1'b0 ;
  assign n16740 = n16739 ^ n16738 ^ 1'b0 ;
  assign n16741 = n16740 ^ n9781 ^ 1'b0 ;
  assign n16742 = n6556 ^ n1845 ^ 1'b0 ;
  assign n16743 = n3931 ^ n2066 ^ 1'b0 ;
  assign n16744 = n4827 & n16743 ;
  assign n16745 = n11402 & n16744 ;
  assign n16746 = n4176 & n10041 ;
  assign n16747 = n6523 ^ n1285 ^ 1'b0 ;
  assign n16748 = n7542 & n15445 ;
  assign n16749 = ~n16747 & n16748 ;
  assign n16750 = n8803 ^ n8056 ^ 1'b0 ;
  assign n16751 = n2731 | n8693 ;
  assign n16752 = n12596 & ~n16751 ;
  assign n16753 = ~n16750 & n16752 ;
  assign n16754 = ~n9793 & n16753 ;
  assign n16755 = n1027 | n8074 ;
  assign n16756 = n16755 ^ n16085 ^ 1'b0 ;
  assign n16757 = n1880 | n7800 ;
  assign n16758 = n16756 & ~n16757 ;
  assign n16759 = ~n1058 & n10281 ;
  assign n16760 = n10528 ^ n8695 ^ 1'b0 ;
  assign n16761 = n2689 & n13791 ;
  assign n16762 = n16761 ^ n3606 ^ 1'b0 ;
  assign n16763 = x87 & ~n562 ;
  assign n16764 = n3024 & n16763 ;
  assign n16765 = n4160 & ~n9823 ;
  assign n16766 = n16765 ^ n8120 ^ 1'b0 ;
  assign n16767 = n16766 ^ n14635 ^ 1'b0 ;
  assign n16768 = ( n1214 & ~n6797 ) | ( n1214 & n13848 ) | ( ~n6797 & n13848 ) ;
  assign n16769 = ~n6062 & n13875 ;
  assign n16770 = ~n10650 & n16769 ;
  assign n16771 = n521 | n2668 ;
  assign n16772 = n16771 ^ n11751 ^ 1'b0 ;
  assign n16773 = n2172 ^ n452 ^ 1'b0 ;
  assign n16774 = n14071 | n16773 ;
  assign n16775 = n1657 | n16774 ;
  assign n16776 = n16772 & ~n16775 ;
  assign n16777 = n13108 ^ n4022 ^ 1'b0 ;
  assign n16778 = n6226 & n16777 ;
  assign n16779 = n16778 ^ n5681 ^ n3961 ;
  assign n16780 = n5844 & n16779 ;
  assign n16781 = ~n7697 & n10396 ;
  assign n16782 = n16781 ^ n1694 ^ 1'b0 ;
  assign n16783 = n10877 & n16782 ;
  assign n16784 = n11504 ^ n2190 ^ 1'b0 ;
  assign n16785 = n7175 ^ n6439 ^ 1'b0 ;
  assign n16786 = n9963 | n16785 ;
  assign n16787 = n16786 ^ n426 ^ 1'b0 ;
  assign n16788 = n6899 | n16787 ;
  assign n16789 = n2665 | n6986 ;
  assign n16790 = n6582 ^ n2350 ^ 1'b0 ;
  assign n16791 = n5529 & n16790 ;
  assign n16792 = n16791 ^ n13395 ^ 1'b0 ;
  assign n16793 = n12829 & ~n13428 ;
  assign n16794 = n16793 ^ n2820 ^ 1'b0 ;
  assign n16796 = n5379 & n14352 ;
  assign n16797 = ~n5293 & n16796 ;
  assign n16795 = n9153 & n12888 ;
  assign n16798 = n16797 ^ n16795 ^ 1'b0 ;
  assign n16799 = n16798 ^ n5099 ^ 1'b0 ;
  assign n16800 = n3083 & ~n10266 ;
  assign n16801 = n2389 & n16800 ;
  assign n16802 = n390 & ~n3472 ;
  assign n16803 = n9436 ^ n7251 ^ 1'b0 ;
  assign n16804 = n7808 & n16803 ;
  assign n16805 = ~n16802 & n16804 ;
  assign n16810 = ( ~n273 & n897 ) | ( ~n273 & n10488 ) | ( n897 & n10488 ) ;
  assign n16806 = n3591 & ~n8080 ;
  assign n16807 = ~n5307 & n16806 ;
  assign n16808 = x213 & ~n16807 ;
  assign n16809 = ~n1638 & n16808 ;
  assign n16811 = n16810 ^ n16809 ^ 1'b0 ;
  assign n16812 = n3040 & n6055 ;
  assign n16813 = ~n11150 & n16812 ;
  assign n16814 = n8849 & ~n16813 ;
  assign n16815 = n5819 | n7570 ;
  assign n16816 = n8403 ^ n3632 ^ 1'b0 ;
  assign n16817 = ~n3676 & n16816 ;
  assign n16818 = ~n16815 & n16817 ;
  assign n16819 = n16818 ^ n13499 ^ 1'b0 ;
  assign n16820 = n3943 & ~n8245 ;
  assign n16821 = n16820 ^ n16647 ^ 1'b0 ;
  assign n16822 = n2515 | n7062 ;
  assign n16823 = ( n15884 & n16288 ) | ( n15884 & ~n16822 ) | ( n16288 & ~n16822 ) ;
  assign n16824 = n16823 ^ n1004 ^ 1'b0 ;
  assign n16825 = n8087 ^ n3018 ^ 1'b0 ;
  assign n16826 = n15630 & ~n16825 ;
  assign n16827 = n9445 | n11596 ;
  assign n16828 = n625 ^ x245 ^ 1'b0 ;
  assign n16829 = n3024 | n16828 ;
  assign n16830 = n12151 | n16829 ;
  assign n16831 = n16830 ^ n12048 ^ 1'b0 ;
  assign n16832 = n4685 & ~n9690 ;
  assign n16833 = n12827 & n14356 ;
  assign n16834 = n10677 ^ n6200 ^ 1'b0 ;
  assign n16835 = ~n3081 & n16834 ;
  assign n16836 = n2841 | n3142 ;
  assign n16837 = ~n3727 & n14468 ;
  assign n16838 = n937 | n8548 ;
  assign n16839 = n16838 ^ n7007 ^ 1'b0 ;
  assign n16840 = n5050 | n11908 ;
  assign n16841 = n16840 ^ n10195 ^ 1'b0 ;
  assign n16842 = ~n1473 & n10081 ;
  assign n16843 = n9270 ^ n1012 ^ 1'b0 ;
  assign n16846 = x182 & ~n700 ;
  assign n16845 = n3917 | n8291 ;
  assign n16847 = n16846 ^ n16845 ^ 1'b0 ;
  assign n16844 = n2304 & ~n14376 ;
  assign n16848 = n16847 ^ n16844 ^ 1'b0 ;
  assign n16849 = ~n2429 & n16848 ;
  assign n16850 = ~n5667 & n13360 ;
  assign n16851 = n16850 ^ n1378 ^ 1'b0 ;
  assign n16852 = n5564 ^ n4399 ^ 1'b0 ;
  assign n16853 = n10678 & n16852 ;
  assign n16854 = n10192 ^ n774 ^ 1'b0 ;
  assign n16855 = n8514 | n16854 ;
  assign n16856 = n3982 & n16855 ;
  assign n16857 = n1914 & ~n16856 ;
  assign n16858 = n16857 ^ n10926 ^ 1'b0 ;
  assign n16859 = n3191 | n16858 ;
  assign n16860 = n3527 ^ x253 ^ 1'b0 ;
  assign n16861 = n3181 | n8068 ;
  assign n16862 = n1703 & n3171 ;
  assign n16863 = n4013 ^ n2157 ^ 1'b0 ;
  assign n16864 = n16863 ^ n13124 ^ 1'b0 ;
  assign n16865 = n11192 & ~n16864 ;
  assign n16866 = ~n6386 & n14130 ;
  assign n16867 = n16866 ^ n12304 ^ 1'b0 ;
  assign n16868 = ( n2691 & ~n2785 ) | ( n2691 & n3687 ) | ( ~n2785 & n3687 ) ;
  assign n16869 = ~n6543 & n15409 ;
  assign n16870 = n8424 & n16869 ;
  assign n16871 = n10136 | n16870 ;
  assign n16872 = n5413 | n16871 ;
  assign n16873 = n4510 & n5140 ;
  assign n16874 = n9292 & n16873 ;
  assign n16875 = x159 & ~n3521 ;
  assign n16876 = n16875 ^ n867 ^ 1'b0 ;
  assign n16877 = n6276 ^ n2753 ^ 1'b0 ;
  assign n16878 = n16876 & ~n16877 ;
  assign n16879 = x148 & n2112 ;
  assign n16880 = n9964 & n16879 ;
  assign n16881 = n8889 ^ n1622 ^ 1'b0 ;
  assign n16882 = n13701 & n16881 ;
  assign n16883 = n13832 ^ n361 ^ 1'b0 ;
  assign n16884 = n10221 & ~n16883 ;
  assign n16885 = n4999 | n6691 ;
  assign n16886 = n16833 ^ n14660 ^ 1'b0 ;
  assign n16887 = n14572 | n16886 ;
  assign n16888 = n5658 ^ n2486 ^ 1'b0 ;
  assign n16889 = n10505 & ~n16888 ;
  assign n16890 = n16889 ^ n1423 ^ 1'b0 ;
  assign n16891 = ~n8663 & n16890 ;
  assign n16892 = n16733 ^ n6359 ^ 1'b0 ;
  assign n16893 = n11585 | n12088 ;
  assign n16894 = ~n307 & n786 ;
  assign n16895 = ~n10922 & n16894 ;
  assign n16896 = n15298 & n16895 ;
  assign n16897 = n8217 & ~n15515 ;
  assign n16898 = n10697 ^ n3608 ^ 1'b0 ;
  assign n16899 = n1291 | n7832 ;
  assign n16900 = n1822 & ~n16899 ;
  assign n16901 = n3604 & n6156 ;
  assign n16902 = n16901 ^ n3045 ^ 1'b0 ;
  assign n16903 = n7924 ^ n1474 ^ 1'b0 ;
  assign n16904 = n2142 | n2228 ;
  assign n16905 = n16904 ^ n1814 ^ 1'b0 ;
  assign n16906 = ~n2403 & n16905 ;
  assign n16907 = n4489 & n16906 ;
  assign n16908 = n2770 | n16907 ;
  assign n16909 = n16908 ^ n10612 ^ 1'b0 ;
  assign n16910 = n4041 & n16909 ;
  assign n16915 = x115 | n696 ;
  assign n16916 = n696 & ~n16915 ;
  assign n16917 = n5896 & ~n16916 ;
  assign n16918 = ~n5896 & n16917 ;
  assign n16919 = n7814 | n16918 ;
  assign n16911 = n2322 & ~n2700 ;
  assign n16912 = n1400 & ~n16911 ;
  assign n16913 = ~n1400 & n16912 ;
  assign n16914 = n9576 & ~n16913 ;
  assign n16920 = n16919 ^ n16914 ^ 1'b0 ;
  assign n16921 = ~n7616 & n16330 ;
  assign n16922 = n16921 ^ n15513 ^ 1'b0 ;
  assign n16923 = n8457 & ~n16922 ;
  assign n16924 = n2274 & n2879 ;
  assign n16925 = ~n13741 & n16924 ;
  assign n16926 = n16925 ^ n14956 ^ 1'b0 ;
  assign n16927 = n12813 ^ n4824 ^ n2736 ;
  assign n16928 = n5323 ^ n1907 ^ 1'b0 ;
  assign n16929 = ~n16927 & n16928 ;
  assign n16930 = n10922 ^ n3370 ^ 1'b0 ;
  assign n16931 = n13220 ^ n3468 ^ 1'b0 ;
  assign n16932 = n4860 & ~n5964 ;
  assign n16933 = ~n4860 & n16932 ;
  assign n16934 = n9033 & n9810 ;
  assign n16935 = ~n9810 & n16934 ;
  assign n16936 = n16933 & ~n16935 ;
  assign n16937 = ~n16933 & n16936 ;
  assign n16938 = n16937 ^ n12779 ^ 1'b0 ;
  assign n16939 = n15436 ^ n9059 ^ 1'b0 ;
  assign n16940 = ~n5928 & n15624 ;
  assign n16941 = n15150 ^ n11695 ^ 1'b0 ;
  assign n16942 = n16941 ^ n12676 ^ n458 ;
  assign n16943 = n13671 ^ n2566 ^ 1'b0 ;
  assign n16944 = n1578 & n16943 ;
  assign n16945 = n7185 | n7575 ;
  assign n16946 = n16945 ^ n9217 ^ 1'b0 ;
  assign n16947 = n4122 | n15175 ;
  assign n16948 = ~n10177 & n12687 ;
  assign n16949 = n8403 ^ n2361 ^ n532 ;
  assign n16950 = n16642 & n16949 ;
  assign n16951 = n16950 ^ n6196 ^ 1'b0 ;
  assign n16952 = ~n9108 & n10280 ;
  assign n16953 = n16952 ^ n3703 ^ 1'b0 ;
  assign n16954 = n11158 ^ n2852 ^ 1'b0 ;
  assign n16955 = ~n14508 & n14677 ;
  assign n16956 = n4304 & n7533 ;
  assign n16957 = n16956 ^ n4661 ^ 1'b0 ;
  assign n16958 = n8589 ^ n1690 ^ 1'b0 ;
  assign n16959 = ~n1239 & n16958 ;
  assign n16960 = n4261 & n16959 ;
  assign n16961 = ~n16957 & n16960 ;
  assign n16962 = x182 & ~n14668 ;
  assign n16963 = n803 & n3112 ;
  assign n16964 = x84 | n1926 ;
  assign n16965 = n5744 | n12345 ;
  assign n16966 = n4954 & ~n9222 ;
  assign n16967 = n16966 ^ n5203 ^ 1'b0 ;
  assign n16968 = n5890 & ~n14336 ;
  assign n16969 = n3606 ^ n1557 ^ 1'b0 ;
  assign n16970 = ~n4204 & n16969 ;
  assign n16971 = ( n2194 & n6868 ) | ( n2194 & ~n16970 ) | ( n6868 & ~n16970 ) ;
  assign n16972 = ~n7926 & n14323 ;
  assign n16973 = ~x136 & n16972 ;
  assign n16974 = n12317 & ~n16973 ;
  assign n16975 = n15960 ^ n6281 ^ 1'b0 ;
  assign n16976 = n2275 & n16975 ;
  assign n16977 = n1732 & n14093 ;
  assign n16978 = ~n570 & n16977 ;
  assign n16979 = n1459 & n16978 ;
  assign n16980 = ~n1076 & n13617 ;
  assign n16981 = n718 & n16980 ;
  assign n16982 = n16981 ^ n13675 ^ 1'b0 ;
  assign n16983 = n16982 ^ n5225 ^ 1'b0 ;
  assign n16984 = n16979 | n16983 ;
  assign n16985 = ( x165 & ~n5176 ) | ( x165 & n15791 ) | ( ~n5176 & n15791 ) ;
  assign n16986 = x160 & n16576 ;
  assign n16988 = n7278 ^ n6292 ^ n966 ;
  assign n16987 = ~n1896 & n4322 ;
  assign n16989 = n16988 ^ n16987 ^ 1'b0 ;
  assign n16990 = n7310 & ~n16989 ;
  assign n16991 = n14799 ^ n3590 ^ 1'b0 ;
  assign n16992 = n8131 | n16991 ;
  assign n16993 = n7421 | n8551 ;
  assign n16994 = n5748 | n16993 ;
  assign n16995 = n8074 ^ n1691 ^ 1'b0 ;
  assign n16996 = n9380 & n16995 ;
  assign n16997 = n16417 ^ x84 ^ 1'b0 ;
  assign n16998 = n16996 & ~n16997 ;
  assign n16999 = n15485 ^ n10571 ^ 1'b0 ;
  assign n17000 = n7293 ^ n3011 ^ 1'b0 ;
  assign n17001 = n10525 & ~n14919 ;
  assign n17002 = n17001 ^ n11272 ^ 1'b0 ;
  assign n17009 = n9558 & ~n11103 ;
  assign n17003 = n8472 ^ n7733 ^ 1'b0 ;
  assign n17004 = n17003 ^ x130 ^ 1'b0 ;
  assign n17005 = n5627 ^ n4680 ^ 1'b0 ;
  assign n17006 = ~n6420 & n17005 ;
  assign n17007 = n17006 ^ n10545 ^ 1'b0 ;
  assign n17008 = n17004 & n17007 ;
  assign n17010 = n17009 ^ n17008 ^ 1'b0 ;
  assign n17011 = n10325 ^ n540 ^ 1'b0 ;
  assign n17012 = n12571 ^ n886 ^ 1'b0 ;
  assign n17013 = x195 & ~n13156 ;
  assign n17014 = n17013 ^ n4668 ^ 1'b0 ;
  assign n17015 = n12915 ^ n11702 ^ 1'b0 ;
  assign n17016 = x65 & ~n1863 ;
  assign n17017 = ~x65 & n17016 ;
  assign n17018 = n9071 ^ n956 ^ 1'b0 ;
  assign n17019 = n17017 | n17018 ;
  assign n17020 = ( n1295 & n8599 ) | ( n1295 & n17019 ) | ( n8599 & n17019 ) ;
  assign n17021 = n1221 | n5650 ;
  assign n17022 = n3052 & ~n17021 ;
  assign n17023 = n10668 | n17022 ;
  assign n17024 = n17023 ^ n4136 ^ 1'b0 ;
  assign n17025 = n2207 ^ n327 ^ 1'b0 ;
  assign n17026 = n17024 & n17025 ;
  assign n17027 = n2433 & ~n4138 ;
  assign n17028 = ~n16160 & n17027 ;
  assign n17029 = n1810 & ~n13830 ;
  assign n17030 = ~n3784 & n16389 ;
  assign n17031 = n331 | n2944 ;
  assign n17032 = n17031 ^ n12463 ^ 1'b0 ;
  assign n17033 = ~n3319 & n5994 ;
  assign n17034 = n17032 & n17033 ;
  assign n17035 = n15571 & ~n17034 ;
  assign n17036 = ~n12379 & n17035 ;
  assign n17037 = n15875 ^ n5968 ^ 1'b0 ;
  assign n17038 = n1890 | n8551 ;
  assign n17039 = n2537 & n17038 ;
  assign n17040 = x222 & ~n1658 ;
  assign n17041 = n17040 ^ n445 ^ 1'b0 ;
  assign n17042 = n508 & n5597 ;
  assign n17043 = ~n4293 & n17042 ;
  assign n17044 = ~n1473 & n2373 ;
  assign n17045 = n17043 & n17044 ;
  assign n17046 = n3362 & n17045 ;
  assign n17047 = n17046 ^ n2505 ^ 1'b0 ;
  assign n17048 = n7280 & n17047 ;
  assign n17049 = ~n5683 & n17048 ;
  assign n17050 = ~n13155 & n17049 ;
  assign n17051 = n1177 & n15866 ;
  assign n17052 = n17050 & n17051 ;
  assign n17053 = n7465 & ~n13178 ;
  assign n17054 = ( n2893 & n7483 ) | ( n2893 & n14774 ) | ( n7483 & n14774 ) ;
  assign n17055 = n7385 ^ n1738 ^ 1'b0 ;
  assign n17056 = ~n2301 & n17055 ;
  assign n17057 = n17056 ^ n14022 ^ 1'b0 ;
  assign n17058 = n1045 & n17057 ;
  assign n17059 = n7552 ^ n7549 ^ 1'b0 ;
  assign n17060 = n17059 ^ n1736 ^ 1'b0 ;
  assign n17061 = ~n3283 & n17060 ;
  assign n17062 = n5468 & n11255 ;
  assign n17063 = n2366 & n4323 ;
  assign n17064 = ~n16022 & n17063 ;
  assign n17065 = n7185 ^ n2887 ^ 1'b0 ;
  assign n17066 = n17065 ^ n11204 ^ 1'b0 ;
  assign n17067 = n11442 ^ n10158 ^ 1'b0 ;
  assign n17068 = n3630 | n7241 ;
  assign n17069 = n977 | n9381 ;
  assign n17070 = ~n6263 & n8297 ;
  assign n17071 = n8468 ^ n6146 ^ n1029 ;
  assign n17072 = x36 & ~n4181 ;
  assign n17073 = n9446 ^ n2814 ^ 1'b0 ;
  assign n17074 = n17072 & n17073 ;
  assign n17075 = n6742 & n11481 ;
  assign n17076 = n17075 ^ n10711 ^ 1'b0 ;
  assign n17077 = ~n3834 & n7288 ;
  assign n17078 = n16057 & n17077 ;
  assign n17079 = ~n10689 & n12370 ;
  assign n17080 = n17078 & n17079 ;
  assign n17081 = n5607 | n15664 ;
  assign n17082 = n3028 | n17081 ;
  assign n17083 = ~n3324 & n17082 ;
  assign n17084 = n6573 | n17083 ;
  assign n17085 = n13795 ^ n8718 ^ 1'b0 ;
  assign n17086 = n2657 | n10606 ;
  assign n17087 = n17086 ^ n2511 ^ 1'b0 ;
  assign n17088 = n14344 & ~n17087 ;
  assign n17089 = ~n12878 & n15707 ;
  assign n17090 = n17089 ^ n15705 ^ 1'b0 ;
  assign n17091 = n17090 ^ n15678 ^ 1'b0 ;
  assign n17092 = n343 & ~n17091 ;
  assign n17093 = ~n522 & n16848 ;
  assign n17094 = n5779 ^ n1693 ^ 1'b0 ;
  assign n17095 = n7901 & ~n8150 ;
  assign n17096 = n2936 | n17095 ;
  assign n17097 = n691 | n17096 ;
  assign n17098 = n14895 ^ n7148 ^ 1'b0 ;
  assign n17099 = n5027 & ~n16895 ;
  assign n17100 = ~n16463 & n17099 ;
  assign n17101 = n2310 | n9954 ;
  assign n17102 = n1111 & ~n6370 ;
  assign n17103 = n17101 & n17102 ;
  assign n17104 = n15605 ^ n8511 ^ 1'b0 ;
  assign n17105 = n1336 & ~n5399 ;
  assign n17106 = n17105 ^ n11654 ^ 1'b0 ;
  assign n17107 = n9015 | n17106 ;
  assign n17108 = n12531 ^ n5105 ^ 1'b0 ;
  assign n17109 = n8422 ^ n7996 ^ 1'b0 ;
  assign n17110 = ~n8004 & n17109 ;
  assign n17111 = ~n4488 & n12410 ;
  assign n17112 = n3304 & ~n15483 ;
  assign n17113 = n5023 & n8324 ;
  assign n17114 = ~n1070 & n17113 ;
  assign n17115 = n17112 | n17114 ;
  assign n17116 = n14778 & n17115 ;
  assign n17117 = n2845 & n5168 ;
  assign n17118 = n10988 ^ n9925 ^ 1'b0 ;
  assign n17119 = n17117 & ~n17118 ;
  assign n17120 = ~n401 & n3230 ;
  assign n17121 = n401 & n17120 ;
  assign n17122 = n9323 & ~n17121 ;
  assign n17123 = ~n9323 & n17122 ;
  assign n17124 = ( n10146 & ~n11477 ) | ( n10146 & n15235 ) | ( ~n11477 & n15235 ) ;
  assign n17125 = n4270 & n6106 ;
  assign n17126 = n17125 ^ n2230 ^ 1'b0 ;
  assign n17127 = n17126 ^ n2809 ^ 1'b0 ;
  assign n17128 = n4524 & ~n17127 ;
  assign n17129 = n6999 & n11431 ;
  assign n17130 = n17129 ^ n4932 ^ 1'b0 ;
  assign n17131 = n17128 & n17130 ;
  assign n17132 = n17131 ^ n3531 ^ 1'b0 ;
  assign n17133 = n4579 ^ n959 ^ 1'b0 ;
  assign n17134 = ~n12777 & n17133 ;
  assign n17135 = n2006 & n17134 ;
  assign n17136 = ~n12293 & n16463 ;
  assign n17137 = n16150 ^ n9771 ^ 1'b0 ;
  assign n17138 = n6782 ^ n4925 ^ 1'b0 ;
  assign n17139 = n8580 & n17138 ;
  assign n17140 = n17139 ^ n6180 ^ 1'b0 ;
  assign n17141 = n17140 ^ n9210 ^ 1'b0 ;
  assign n17142 = n9651 ^ n6060 ^ 1'b0 ;
  assign n17143 = n6954 & n17142 ;
  assign n17144 = ~n4655 & n17143 ;
  assign n17145 = ~n13056 & n17144 ;
  assign n17146 = n7031 ^ x66 ^ 1'b0 ;
  assign n17147 = n14000 ^ n6442 ^ n440 ;
  assign n17148 = n15256 ^ n663 ^ 1'b0 ;
  assign n17149 = n2374 & n8386 ;
  assign n17150 = n17149 ^ n3239 ^ 1'b0 ;
  assign n17151 = n17150 ^ n8616 ^ 1'b0 ;
  assign n17152 = n8806 | n17151 ;
  assign n17153 = n4767 & n16157 ;
  assign n17154 = n2602 & n8570 ;
  assign n17155 = n9247 | n10440 ;
  assign n17156 = ( ~n1535 & n1657 ) | ( ~n1535 & n17155 ) | ( n1657 & n17155 ) ;
  assign n17157 = ~n8514 & n17156 ;
  assign n17158 = ~n15712 & n17157 ;
  assign n17159 = ~n5678 & n14116 ;
  assign n17160 = n13586 | n15872 ;
  assign n17161 = n17160 ^ n8084 ^ 1'b0 ;
  assign n17162 = n17159 & ~n17161 ;
  assign n17163 = n8967 ^ n8808 ^ 1'b0 ;
  assign n17164 = n2747 | n8572 ;
  assign n17165 = n17164 ^ n3891 ^ 1'b0 ;
  assign n17166 = ~n6391 & n17165 ;
  assign n17167 = n553 & ~n2861 ;
  assign n17168 = n2476 & ~n9909 ;
  assign n17169 = ( n5842 & ~n17167 ) | ( n5842 & n17168 ) | ( ~n17167 & n17168 ) ;
  assign n17170 = n14033 | n14995 ;
  assign n17171 = n17170 ^ n3536 ^ 1'b0 ;
  assign n17172 = ~n3243 & n6192 ;
  assign n17175 = n1877 & ~n15640 ;
  assign n17176 = ~x216 & n17175 ;
  assign n17173 = n2467 & n13585 ;
  assign n17174 = ~n2074 & n17173 ;
  assign n17177 = n17176 ^ n17174 ^ 1'b0 ;
  assign n17178 = n638 & ~n3784 ;
  assign n17179 = n17178 ^ n2470 ^ 1'b0 ;
  assign n17180 = n8169 | n17179 ;
  assign n17181 = n7769 & n17180 ;
  assign n17182 = n8448 ^ n6094 ^ n5151 ;
  assign n17184 = ( n2660 & n4310 ) | ( n2660 & n7512 ) | ( n4310 & n7512 ) ;
  assign n17183 = n1869 | n12473 ;
  assign n17185 = n17184 ^ n17183 ^ 1'b0 ;
  assign n17186 = n387 & ~n12302 ;
  assign n17187 = n12586 | n16060 ;
  assign n17188 = n5552 & ~n17187 ;
  assign n17189 = ( n7966 & n8919 ) | ( n7966 & ~n10108 ) | ( n8919 & ~n10108 ) ;
  assign n17190 = n8511 ^ n2366 ^ 1'b0 ;
  assign n17191 = ~n11783 & n12645 ;
  assign n17192 = n17191 ^ n13778 ^ 1'b0 ;
  assign n17194 = n1775 & ~n10328 ;
  assign n17195 = n5203 & n17194 ;
  assign n17193 = n8239 ^ n2274 ^ 1'b0 ;
  assign n17196 = n17195 ^ n17193 ^ 1'b0 ;
  assign n17197 = ~n9220 & n13588 ;
  assign n17198 = n8108 | n17197 ;
  assign n17206 = n3089 ^ n529 ^ 1'b0 ;
  assign n17207 = n607 & n17206 ;
  assign n17199 = x80 & ~n7688 ;
  assign n17200 = n936 & n17199 ;
  assign n17201 = n12709 & n17200 ;
  assign n17203 = n305 & n13780 ;
  assign n17202 = n4089 | n6315 ;
  assign n17204 = n17203 ^ n17202 ^ 1'b0 ;
  assign n17205 = ~n17201 & n17204 ;
  assign n17208 = n17207 ^ n17205 ^ 1'b0 ;
  assign n17210 = n3939 | n7244 ;
  assign n17211 = n6700 | n17210 ;
  assign n17209 = n8875 ^ x73 ^ 1'b0 ;
  assign n17212 = n17211 ^ n17209 ^ 1'b0 ;
  assign n17213 = n6962 ^ x70 ^ 1'b0 ;
  assign n17214 = n613 & ~n17213 ;
  assign n17215 = n7012 ^ n3756 ^ 1'b0 ;
  assign n17216 = n2973 & n5830 ;
  assign n17217 = ~n17215 & n17216 ;
  assign n17218 = n7002 ^ n4047 ^ 1'b0 ;
  assign n17219 = ~n1950 & n2633 ;
  assign n17220 = n3167 | n17219 ;
  assign n17221 = n17218 | n17220 ;
  assign n17222 = n3040 ^ n1066 ^ 1'b0 ;
  assign n17223 = n5259 | n9122 ;
  assign n17224 = n6686 & n6802 ;
  assign n17225 = ~n14448 & n17224 ;
  assign n17226 = ~n677 & n17225 ;
  assign n17227 = ~n12592 & n17226 ;
  assign n17228 = n11246 ^ n9817 ^ 1'b0 ;
  assign n17229 = n3883 | n5317 ;
  assign n17230 = ~n2735 & n17229 ;
  assign n17231 = n7515 ^ n2283 ^ 1'b0 ;
  assign n17232 = n968 | n17231 ;
  assign n17233 = n5503 & ~n11920 ;
  assign n17234 = n17233 ^ n1164 ^ 1'b0 ;
  assign n17235 = n17234 ^ n3648 ^ 1'b0 ;
  assign n17238 = ~n1573 & n10322 ;
  assign n17236 = n4454 | n10833 ;
  assign n17237 = ( ~n4302 & n6730 ) | ( ~n4302 & n17236 ) | ( n6730 & n17236 ) ;
  assign n17239 = n17238 ^ n17237 ^ 1'b0 ;
  assign n17240 = n17235 & n17239 ;
  assign n17241 = n17240 ^ n10042 ^ 1'b0 ;
  assign n17242 = n9041 & ~n17241 ;
  assign n17243 = ~n965 & n11075 ;
  assign n17244 = n17243 ^ n7385 ^ 1'b0 ;
  assign n17245 = n7461 & ~n10363 ;
  assign n17246 = n17245 ^ n16460 ^ 1'b0 ;
  assign n17247 = ~x76 & n13791 ;
  assign n17248 = n6798 & ~n11638 ;
  assign n17249 = n17248 ^ n5442 ^ 1'b0 ;
  assign n17250 = x11 & n17249 ;
  assign n17251 = ~n2470 & n17250 ;
  assign n17252 = n5635 & n5804 ;
  assign n17253 = n5712 & n13290 ;
  assign n17254 = ~n904 & n17253 ;
  assign n17255 = n17254 ^ x226 ^ 1'b0 ;
  assign n17256 = ~n370 & n8558 ;
  assign n17257 = n17256 ^ n13827 ^ 1'b0 ;
  assign n17258 = ( n2835 & n8055 ) | ( n2835 & n14818 ) | ( n8055 & n14818 ) ;
  assign n17259 = ~n5373 & n5692 ;
  assign n17260 = ~n6253 & n17259 ;
  assign n17261 = n4831 & ~n17260 ;
  assign n17262 = n17258 & n17261 ;
  assign n17264 = n1341 ^ n562 ^ 1'b0 ;
  assign n17263 = n9834 & ~n11685 ;
  assign n17265 = n17264 ^ n17263 ^ 1'b0 ;
  assign n17266 = ~n4934 & n5039 ;
  assign n17267 = n998 & ~n7901 ;
  assign n17268 = n17267 ^ n1221 ^ 1'b0 ;
  assign n17269 = n17266 & ~n17268 ;
  assign n17270 = n519 & ~n9292 ;
  assign n17271 = ~n1820 & n4238 ;
  assign n17272 = n5095 & n17271 ;
  assign n17273 = ~n5207 & n7695 ;
  assign n17274 = ~n8529 & n16160 ;
  assign n17275 = ~n12342 & n15647 ;
  assign n17276 = n17274 & n17275 ;
  assign n17277 = ~n4821 & n9836 ;
  assign n17278 = n9415 ^ n7220 ^ 1'b0 ;
  assign n17279 = ~n3649 & n9972 ;
  assign n17280 = n17279 ^ n4261 ^ 1'b0 ;
  assign n17281 = n5273 & ~n17280 ;
  assign n17282 = ~n17278 & n17281 ;
  assign n17283 = ~n1660 & n4118 ;
  assign n17284 = ~n5937 & n17283 ;
  assign n17285 = n17284 ^ n6826 ^ n5955 ;
  assign n17286 = ~n11722 & n17285 ;
  assign n17287 = n14842 & n15651 ;
  assign n17288 = n4695 | n16872 ;
  assign n17289 = n538 & ~n1553 ;
  assign n17290 = n5916 ^ n5638 ^ 1'b0 ;
  assign n17291 = n17290 ^ n10629 ^ 1'b0 ;
  assign n17292 = n17289 & n17291 ;
  assign n17293 = n8122 ^ n1414 ^ 1'b0 ;
  assign n17294 = ~n6784 & n9236 ;
  assign n17295 = n3216 & n7079 ;
  assign n17296 = n1181 & n11135 ;
  assign n17297 = ~x161 & n3424 ;
  assign n17298 = n10211 & n16876 ;
  assign n17301 = n2237 ^ n388 ^ 1'b0 ;
  assign n17300 = n2263 & ~n3331 ;
  assign n17302 = n17301 ^ n17300 ^ 1'b0 ;
  assign n17299 = ~n3181 & n4329 ;
  assign n17303 = n17302 ^ n17299 ^ 1'b0 ;
  assign n17304 = n354 & ~n2371 ;
  assign n17305 = n6954 ^ n1976 ^ 1'b0 ;
  assign n17306 = n2642 & n17305 ;
  assign n17307 = n519 | n15325 ;
  assign n17308 = n9626 & ~n17307 ;
  assign n17309 = n12753 ^ n10049 ^ n5273 ;
  assign n17310 = n17309 ^ n9752 ^ 1'b0 ;
  assign n17311 = ~n643 & n9982 ;
  assign n17312 = ~n1766 & n3437 ;
  assign n17313 = n8055 | n17312 ;
  assign n17314 = n17311 & ~n17313 ;
  assign n17315 = ~n7172 & n14302 ;
  assign n17316 = n17315 ^ n4336 ^ 1'b0 ;
  assign n17317 = n15260 ^ n9396 ^ 1'b0 ;
  assign n17318 = n5487 & n17317 ;
  assign n17319 = ~n788 & n4939 ;
  assign n17320 = n15983 & n17319 ;
  assign n17321 = n2071 & n6759 ;
  assign n17322 = n17321 ^ n9166 ^ 1'b0 ;
  assign n17323 = n1762 & n17322 ;
  assign n17324 = n17323 ^ n8010 ^ 1'b0 ;
  assign n17325 = n1779 & n17324 ;
  assign n17326 = n8770 & ~n13220 ;
  assign n17327 = ~n15315 & n17326 ;
  assign n17328 = n12041 | n17327 ;
  assign n17329 = n8628 & ~n17328 ;
  assign n17330 = n17329 ^ n14314 ^ 1'b0 ;
  assign n17331 = n14523 & n17330 ;
  assign n17334 = x12 & ~n8236 ;
  assign n17335 = n17334 ^ n1521 ^ 1'b0 ;
  assign n17332 = n4012 & ~n7836 ;
  assign n17333 = n10342 | n17332 ;
  assign n17336 = n17335 ^ n17333 ^ 1'b0 ;
  assign n17337 = n6681 ^ n2750 ^ 1'b0 ;
  assign n17338 = n15630 & ~n17337 ;
  assign n17339 = n17338 ^ n12035 ^ 1'b0 ;
  assign n17340 = n6602 & ~n17339 ;
  assign n17341 = ( n4671 & n9561 ) | ( n4671 & ~n17340 ) | ( n9561 & ~n17340 ) ;
  assign n17342 = ( n8563 & n17336 ) | ( n8563 & ~n17341 ) | ( n17336 & ~n17341 ) ;
  assign n17343 = n15990 & ~n17342 ;
  assign n17344 = n17343 ^ n3221 ^ 1'b0 ;
  assign n17345 = n8969 & ~n10059 ;
  assign n17346 = n1368 & n3780 ;
  assign n17347 = n15261 ^ n3790 ^ 1'b0 ;
  assign n17348 = n11899 | n17347 ;
  assign n17350 = n8529 | n8653 ;
  assign n17351 = ~n4043 & n11302 ;
  assign n17352 = n17350 & n17351 ;
  assign n17349 = n2185 & ~n5110 ;
  assign n17353 = n17352 ^ n17349 ^ 1'b0 ;
  assign n17354 = n3001 & ~n17353 ;
  assign n17355 = n6676 ^ n3687 ^ 1'b0 ;
  assign n17356 = n6225 & ~n16493 ;
  assign n17357 = ~n17143 & n17356 ;
  assign n17358 = n10968 ^ n1514 ^ 1'b0 ;
  assign n17359 = n8653 | n17358 ;
  assign n17360 = n17359 ^ n498 ^ 1'b0 ;
  assign n17361 = n2366 | n9693 ;
  assign n17362 = n16246 | n17361 ;
  assign n17363 = n10528 ^ n8695 ^ n1021 ;
  assign n17364 = n1678 & n7899 ;
  assign n17365 = n5639 | n15886 ;
  assign n17366 = n6158 & ~n17365 ;
  assign n17367 = n6967 ^ n4031 ^ 1'b0 ;
  assign n17368 = n15533 | n17367 ;
  assign n17369 = n17368 ^ x216 ^ 1'b0 ;
  assign n17370 = ( n6617 & n12781 ) | ( n6617 & ~n16973 ) | ( n12781 & ~n16973 ) ;
  assign n17371 = n12478 ^ n1264 ^ 1'b0 ;
  assign n17372 = n3729 & n17371 ;
  assign n17373 = n3756 & ~n4777 ;
  assign n17374 = n12943 ^ n4772 ^ 1'b0 ;
  assign n17375 = ~n1999 & n12342 ;
  assign n17376 = n17374 & n17375 ;
  assign n17377 = n17373 & n17376 ;
  assign n17378 = n6322 ^ n3143 ^ 1'b0 ;
  assign n17379 = ( ~n5851 & n10284 ) | ( ~n5851 & n17378 ) | ( n10284 & n17378 ) ;
  assign n17380 = n17379 ^ n5192 ^ 1'b0 ;
  assign n17381 = ~n12468 & n13088 ;
  assign n17382 = ~n13570 & n17381 ;
  assign n17383 = n11222 ^ n7179 ^ 1'b0 ;
  assign n17384 = n3469 ^ n2861 ^ 1'b0 ;
  assign n17385 = n6300 ^ n3210 ^ 1'b0 ;
  assign n17386 = ~n8654 & n17385 ;
  assign n17387 = n3721 | n17386 ;
  assign n17388 = n17387 ^ n8695 ^ 1'b0 ;
  assign n17389 = x43 & ~n17388 ;
  assign n17390 = ~n17384 & n17389 ;
  assign n17391 = n9696 ^ n5604 ^ 1'b0 ;
  assign n17392 = n5597 & n9597 ;
  assign n17393 = ~n10258 & n17392 ;
  assign n17394 = ~n2403 & n14093 ;
  assign n17395 = n17394 ^ n3980 ^ 1'b0 ;
  assign n17396 = n581 & n6355 ;
  assign n17397 = ~n6355 & n17396 ;
  assign n17398 = ~n397 & n1814 ;
  assign n17399 = n17397 & n17398 ;
  assign n17400 = n17395 | n17399 ;
  assign n17401 = n17395 & ~n17400 ;
  assign n17403 = x50 & ~n1910 ;
  assign n17404 = n1910 & n17403 ;
  assign n17405 = x172 & ~n17404 ;
  assign n17406 = ~x172 & n17405 ;
  assign n17402 = n9123 | n15764 ;
  assign n17407 = n17406 ^ n17402 ^ 1'b0 ;
  assign n17408 = n17401 | n17407 ;
  assign n17409 = n5061 | n6725 ;
  assign n17410 = n10332 & ~n17409 ;
  assign n17411 = n8127 ^ n1599 ^ 1'b0 ;
  assign n17412 = ( n6109 & ~n17410 ) | ( n6109 & n17411 ) | ( ~n17410 & n17411 ) ;
  assign n17413 = n17412 ^ n14452 ^ n5269 ;
  assign n17414 = n3805 | n17346 ;
  assign n17415 = n10935 ^ n1775 ^ 1'b0 ;
  assign n17416 = n16768 ^ n7905 ^ 1'b0 ;
  assign n17417 = n4470 & ~n17416 ;
  assign n17418 = n1391 & n17417 ;
  assign n17419 = n3390 ^ n781 ^ 1'b0 ;
  assign n17420 = n5748 ^ n842 ^ 1'b0 ;
  assign n17421 = n17419 & n17420 ;
  assign n17422 = n12159 ^ n6350 ^ 1'b0 ;
  assign n17423 = n8843 & ~n14066 ;
  assign n17424 = n14815 ^ n7692 ^ 1'b0 ;
  assign n17425 = n14356 ^ n1438 ^ 1'b0 ;
  assign n17426 = n16163 ^ n5081 ^ 1'b0 ;
  assign n17428 = ~n753 & n1318 ;
  assign n17429 = n753 & n17428 ;
  assign n17430 = x3 | n17429 ;
  assign n17427 = n2856 | n4373 ;
  assign n17431 = n17430 ^ n17427 ^ 1'b0 ;
  assign n17432 = n11120 ^ n2629 ^ 1'b0 ;
  assign n17433 = n17431 | n17432 ;
  assign n17434 = n1459 | n17433 ;
  assign n17437 = ~n4520 & n11093 ;
  assign n17438 = n4520 & n17437 ;
  assign n17439 = n7519 | n17438 ;
  assign n17440 = n7519 & ~n17439 ;
  assign n17435 = ~n2256 & n16657 ;
  assign n17436 = n2256 & n17435 ;
  assign n17441 = n17440 ^ n17436 ^ 1'b0 ;
  assign n17442 = ~n1903 & n17441 ;
  assign n17443 = ~n387 & n10198 ;
  assign n17444 = n16652 ^ n1621 ^ 1'b0 ;
  assign n17445 = n5728 | n11308 ;
  assign n17446 = n4523 | n10186 ;
  assign n17447 = n7252 & ~n17446 ;
  assign n17448 = ~n17445 & n17447 ;
  assign n17449 = n5998 | n8957 ;
  assign n17450 = n6408 ^ n2689 ^ 1'b0 ;
  assign n17451 = n3362 & n17450 ;
  assign n17452 = n1495 & n17451 ;
  assign n17453 = n1061 & n17452 ;
  assign n17454 = n17453 ^ n844 ^ 1'b0 ;
  assign n17455 = n17449 | n17454 ;
  assign n17456 = n17455 ^ n12951 ^ 1'b0 ;
  assign n17457 = n7775 | n17456 ;
  assign n17458 = n730 & n5199 ;
  assign n17459 = n1240 | n8814 ;
  assign n17460 = n3316 | n17459 ;
  assign n17462 = n6065 ^ n2599 ^ 1'b0 ;
  assign n17463 = n1544 & ~n17462 ;
  assign n17464 = n17463 ^ n17284 ^ 1'b0 ;
  assign n17461 = n16855 ^ n15995 ^ 1'b0 ;
  assign n17465 = n17464 ^ n17461 ^ 1'b0 ;
  assign n17466 = ~n1727 & n4408 ;
  assign n17467 = n4619 ^ n2423 ^ 1'b0 ;
  assign n17468 = n5030 & n17467 ;
  assign n17469 = n17466 & n17468 ;
  assign n17470 = n3177 & n14710 ;
  assign n17471 = n8067 ^ n5070 ^ 1'b0 ;
  assign n17472 = n17471 ^ n4625 ^ 1'b0 ;
  assign n17473 = n7529 & n17472 ;
  assign n17474 = n3526 & ~n6857 ;
  assign n17475 = n7469 & n17474 ;
  assign n17476 = n10056 & ~n17475 ;
  assign n17477 = n13537 & n17476 ;
  assign n17478 = n1707 & n10418 ;
  assign n17479 = n4553 & ~n15091 ;
  assign n17480 = n17479 ^ n6049 ^ 1'b0 ;
  assign n17481 = n17477 ^ n4545 ^ 1'b0 ;
  assign n17482 = ~n8041 & n17481 ;
  assign n17483 = n1693 | n2854 ;
  assign n17484 = n16034 ^ n13549 ^ 1'b0 ;
  assign n17485 = n1037 ^ n988 ^ 1'b0 ;
  assign n17486 = n2203 & ~n17485 ;
  assign n17487 = ~n16770 & n17486 ;
  assign n17488 = ( n1049 & n8422 ) | ( n1049 & ~n11356 ) | ( n8422 & ~n11356 ) ;
  assign n17489 = n10567 & ~n17488 ;
  assign n17490 = n6402 | n7841 ;
  assign n17491 = n3132 | n13539 ;
  assign n17492 = n4661 & ~n17491 ;
  assign n17494 = ~n3888 & n3905 ;
  assign n17495 = ~n8685 & n17494 ;
  assign n17493 = ~n2138 & n4433 ;
  assign n17496 = n17495 ^ n17493 ^ 1'b0 ;
  assign n17497 = ( n566 & n17492 ) | ( n566 & n17496 ) | ( n17492 & n17496 ) ;
  assign n17498 = n17497 ^ n9386 ^ 1'b0 ;
  assign n17499 = ~n17490 & n17498 ;
  assign n17500 = n12216 ^ n6568 ^ 1'b0 ;
  assign n17501 = n8907 & n17500 ;
  assign n17502 = n11927 ^ n6553 ^ 1'b0 ;
  assign n17503 = n7465 ^ n385 ^ 1'b0 ;
  assign n17504 = n7971 ^ n363 ^ 1'b0 ;
  assign n17505 = n3690 ^ n691 ^ 1'b0 ;
  assign n17506 = n7109 ^ n4166 ^ 1'b0 ;
  assign n17507 = n17506 ^ n14493 ^ 1'b0 ;
  assign n17508 = n5748 | n13576 ;
  assign n17509 = n11900 ^ n1801 ^ 1'b0 ;
  assign n17510 = ~n4982 & n17509 ;
  assign n17511 = n887 & ~n6884 ;
  assign n17512 = n728 & ~n17511 ;
  assign n17513 = n849 | n1980 ;
  assign n17514 = n17512 & ~n17513 ;
  assign n17515 = n10346 ^ n8367 ^ 1'b0 ;
  assign n17516 = n14677 ^ n5646 ^ 1'b0 ;
  assign n17518 = n6442 ^ x84 ^ 1'b0 ;
  assign n17519 = n4079 & ~n8180 ;
  assign n17520 = n17518 & ~n17519 ;
  assign n17517 = ~n1698 & n3817 ;
  assign n17521 = n17520 ^ n17517 ^ 1'b0 ;
  assign n17522 = x211 & ~n327 ;
  assign n17523 = ~n1337 & n17522 ;
  assign n17524 = n6716 ^ n5020 ^ 1'b0 ;
  assign n17525 = ~n11656 & n17524 ;
  assign n17526 = n4824 & n17525 ;
  assign n17527 = n5510 ^ n3980 ^ 1'b0 ;
  assign n17528 = n16200 & ~n17527 ;
  assign n17529 = n5390 & n17528 ;
  assign n17530 = ( n1850 & ~n8727 ) | ( n1850 & n10087 ) | ( ~n8727 & n10087 ) ;
  assign n17531 = n6371 | n12331 ;
  assign n17532 = n17531 ^ n6788 ^ 1'b0 ;
  assign n17534 = n11288 ^ n9534 ^ n1393 ;
  assign n17535 = n14338 & n17534 ;
  assign n17533 = n2254 | n11771 ;
  assign n17536 = n17535 ^ n17533 ^ 1'b0 ;
  assign n17539 = n12087 ^ n4126 ^ 1'b0 ;
  assign n17537 = n10865 ^ n6372 ^ 1'b0 ;
  assign n17538 = ~n5444 & n17537 ;
  assign n17540 = n17539 ^ n17538 ^ 1'b0 ;
  assign n17541 = n10615 & n17540 ;
  assign n17542 = n10157 & n17541 ;
  assign n17543 = n14027 | n17542 ;
  assign n17544 = n17543 ^ x219 ^ 1'b0 ;
  assign n17545 = n4560 & ~n9941 ;
  assign n17546 = n2115 | n17545 ;
  assign n17547 = n17546 ^ n13933 ^ 1'b0 ;
  assign n17549 = n2319 ^ n1919 ^ n820 ;
  assign n17548 = n2853 & ~n6766 ;
  assign n17550 = n17549 ^ n17548 ^ 1'b0 ;
  assign n17551 = n502 ^ x150 ^ 1'b0 ;
  assign n17552 = n17551 ^ n8617 ^ n2416 ;
  assign n17553 = n17552 ^ n10357 ^ 1'b0 ;
  assign n17554 = n2701 & n17553 ;
  assign n17555 = n13319 ^ x212 ^ 1'b0 ;
  assign n17556 = ~n10004 & n17555 ;
  assign n17557 = n5758 ^ n5023 ^ 1'b0 ;
  assign n17558 = n8001 | n10552 ;
  assign n17559 = n14205 | n17558 ;
  assign n17560 = n4644 & n12930 ;
  assign n17561 = n17560 ^ n11991 ^ 1'b0 ;
  assign n17562 = n6939 & n17561 ;
  assign n17563 = ~n930 & n17562 ;
  assign n17564 = n17563 ^ n5384 ^ 1'b0 ;
  assign n17565 = ~n2062 & n3499 ;
  assign n17566 = n8068 ^ n3221 ^ 1'b0 ;
  assign n17567 = n17566 ^ n2926 ^ 1'b0 ;
  assign n17568 = n15312 ^ n6708 ^ 1'b0 ;
  assign n17569 = n13059 ^ n5135 ^ 1'b0 ;
  assign n17570 = n630 & n1738 ;
  assign n17571 = n8758 ^ n1523 ^ 1'b0 ;
  assign n17572 = ~n17570 & n17571 ;
  assign n17573 = n14438 ^ n1195 ^ 1'b0 ;
  assign n17574 = n17573 ^ n3249 ^ 1'b0 ;
  assign n17575 = n2018 | n17574 ;
  assign n17576 = n1596 & ~n16799 ;
  assign n17577 = ~n1596 & n17576 ;
  assign n17578 = ~n7232 & n7734 ;
  assign n17579 = n923 & ~n1240 ;
  assign n17580 = n3511 & n4296 ;
  assign n17581 = n13481 | n16295 ;
  assign n17582 = n17580 | n17581 ;
  assign n17583 = n4928 & ~n14790 ;
  assign n17584 = n14992 & ~n17583 ;
  assign n17585 = n9111 ^ n1337 ^ 1'b0 ;
  assign n17586 = ~n1746 & n17585 ;
  assign n17589 = n2581 | n8284 ;
  assign n17590 = n4959 | n17589 ;
  assign n17591 = n3533 & n17590 ;
  assign n17587 = n675 & ~n7693 ;
  assign n17588 = n8268 & n17587 ;
  assign n17592 = n17591 ^ n17588 ^ 1'b0 ;
  assign n17593 = n17586 & ~n17592 ;
  assign n17594 = ~n7210 & n10396 ;
  assign n17595 = ~n8703 & n17594 ;
  assign n17596 = n17593 & n17595 ;
  assign n17597 = n6473 & n9764 ;
  assign n17598 = n1742 & ~n11673 ;
  assign n17599 = ~n5852 & n17598 ;
  assign n17600 = n7278 & ~n17599 ;
  assign n17601 = n17600 ^ n1501 ^ 1'b0 ;
  assign n17602 = n17597 & n17601 ;
  assign n17603 = ~n7297 & n8928 ;
  assign n17604 = n17603 ^ n14818 ^ 1'b0 ;
  assign n17605 = n9643 ^ n2970 ^ 1'b0 ;
  assign n17606 = n17605 ^ n1925 ^ 1'b0 ;
  assign n17607 = ~n1068 & n17606 ;
  assign n17608 = ~n7956 & n17607 ;
  assign n17609 = n13403 & n17608 ;
  assign n17610 = n17609 ^ n3729 ^ 1'b0 ;
  assign n17611 = n17604 & n17610 ;
  assign n17612 = n5752 | n11866 ;
  assign n17613 = n9789 & ~n17612 ;
  assign n17614 = ~x232 & n1426 ;
  assign n17615 = n14781 & n17614 ;
  assign n17616 = n13871 ^ n7263 ^ 1'b0 ;
  assign n17617 = n2507 & n5159 ;
  assign n17618 = n17616 & n17617 ;
  assign n17619 = n4913 | n17618 ;
  assign n17620 = n17619 ^ n6794 ^ 1'b0 ;
  assign n17621 = n2846 & n12033 ;
  assign n17623 = n9389 | n12990 ;
  assign n17624 = n9444 | n17623 ;
  assign n17622 = n2887 & ~n3223 ;
  assign n17625 = n17624 ^ n17622 ^ 1'b0 ;
  assign n17626 = ( ~n3799 & n7391 ) | ( ~n3799 & n17625 ) | ( n7391 & n17625 ) ;
  assign n17627 = n6259 & n10364 ;
  assign n17631 = ~n2704 & n15537 ;
  assign n17628 = n8153 ^ n305 ^ 1'b0 ;
  assign n17629 = n9184 & n12801 ;
  assign n17630 = n17628 | n17629 ;
  assign n17632 = n17631 ^ n17630 ^ 1'b0 ;
  assign n17633 = n2933 & ~n3740 ;
  assign n17642 = n11557 ^ n1701 ^ 1'b0 ;
  assign n17635 = n1263 & ~n4109 ;
  assign n17636 = n4109 & n17635 ;
  assign n17637 = ~n8538 & n11029 ;
  assign n17638 = ~n17636 & n17637 ;
  assign n17639 = ~n974 & n17638 ;
  assign n17640 = ~n17638 & n17639 ;
  assign n17641 = n4698 | n17640 ;
  assign n17643 = n17642 ^ n17641 ^ 1'b0 ;
  assign n17634 = ~n1334 & n1738 ;
  assign n17644 = n17643 ^ n17634 ^ 1'b0 ;
  assign n17645 = ~n981 & n1105 ;
  assign n17646 = ~n1105 & n17645 ;
  assign n17647 = n1318 & n17646 ;
  assign n17648 = x93 | n17647 ;
  assign n17649 = x93 & ~n17648 ;
  assign n17650 = n4009 | n17649 ;
  assign n17651 = n17650 ^ n692 ^ 1'b0 ;
  assign n17652 = n1679 & ~n15743 ;
  assign n17653 = n16652 & n17652 ;
  assign n17654 = n16071 & n17653 ;
  assign n17657 = x85 & ~n4104 ;
  assign n17658 = n4104 & n17657 ;
  assign n17655 = x54 & ~n1709 ;
  assign n17656 = ~x54 & n17655 ;
  assign n17659 = n17658 ^ n17656 ^ 1'b0 ;
  assign n17660 = ~n1886 & n17018 ;
  assign n17661 = n17521 | n17660 ;
  assign n17662 = n17659 & ~n17661 ;
  assign n17663 = n3187 & n10746 ;
  assign n17664 = ~n2995 & n7725 ;
  assign n17665 = n17664 ^ n4840 ^ 1'b0 ;
  assign n17666 = n16855 ^ n4256 ^ 1'b0 ;
  assign n17667 = n17665 & n17666 ;
  assign n17668 = n10433 ^ n6721 ^ 1'b0 ;
  assign n17669 = ~n5324 & n17668 ;
  assign n17670 = n12052 ^ n7628 ^ 1'b0 ;
  assign n17671 = n1228 & ~n4556 ;
  assign n17672 = ~n2169 & n17671 ;
  assign n17673 = x59 | n1499 ;
  assign n17679 = ~n1071 & n15913 ;
  assign n17680 = n17679 ^ n5998 ^ 1'b0 ;
  assign n17676 = n4824 | n10090 ;
  assign n17677 = n17676 ^ n3862 ^ 1'b0 ;
  assign n17675 = n7483 | n13551 ;
  assign n17678 = n17677 ^ n17675 ^ 1'b0 ;
  assign n17674 = n4598 | n14695 ;
  assign n17681 = n17680 ^ n17678 ^ n17674 ;
  assign n17682 = n8850 ^ n1660 ^ 1'b0 ;
  assign n17683 = ~n8112 & n17682 ;
  assign n17684 = n16811 ^ n13275 ^ 1'b0 ;
  assign n17685 = n4140 | n6357 ;
  assign n17689 = x26 & ~n1879 ;
  assign n17686 = n10976 & n15164 ;
  assign n17687 = ~n3768 & n17686 ;
  assign n17688 = n10089 | n17687 ;
  assign n17690 = n17689 ^ n17688 ^ 1'b0 ;
  assign n17691 = ~n17685 & n17690 ;
  assign n17692 = n8436 ^ n1648 ^ 1'b0 ;
  assign n17693 = n2320 & ~n17692 ;
  assign n17694 = ~n14839 & n17014 ;
  assign n17695 = ~n2445 & n11682 ;
  assign n17696 = n13329 ^ n7998 ^ 1'b0 ;
  assign n17697 = n2034 & n4367 ;
  assign n17698 = ~n3562 & n17697 ;
  assign n17699 = n17238 ^ n12170 ^ 1'b0 ;
  assign n17700 = n8795 ^ n8002 ^ n1886 ;
  assign n17701 = n532 & ~n2733 ;
  assign n17702 = ~n532 & n17701 ;
  assign n17703 = n903 | n17702 ;
  assign n17704 = n9043 | n10135 ;
  assign n17705 = n17703 & ~n17704 ;
  assign n17706 = ~n950 & n6174 ;
  assign n17707 = n313 & n4836 ;
  assign n17708 = n17707 ^ n3694 ^ 1'b0 ;
  assign n17709 = n17708 ^ n6328 ^ 1'b0 ;
  assign n17710 = n17706 | n17709 ;
  assign n17711 = n17710 ^ n9926 ^ 1'b0 ;
  assign n17712 = x43 & ~n8616 ;
  assign n17713 = n17712 ^ n5317 ^ 1'b0 ;
  assign n17714 = n11899 ^ n7262 ^ 1'b0 ;
  assign n17715 = x118 & ~n6073 ;
  assign n17716 = ~n3226 & n17715 ;
  assign n17717 = ~n11256 & n17716 ;
  assign n17718 = ( n2389 & n4238 ) | ( n2389 & ~n17717 ) | ( n4238 & ~n17717 ) ;
  assign n17719 = n16970 ^ n4300 ^ 1'b0 ;
  assign n17720 = n5808 & n17719 ;
  assign n17721 = n5973 & n17720 ;
  assign n17722 = n2516 | n6564 ;
  assign n17723 = n17721 | n17722 ;
  assign n17724 = ~n7488 & n14214 ;
  assign n17725 = n4481 & n5496 ;
  assign n17726 = n17725 ^ n4166 ^ 1'b0 ;
  assign n17727 = ~n4796 & n17726 ;
  assign n17728 = x68 & n17727 ;
  assign n17729 = n17728 ^ n465 ^ 1'b0 ;
  assign n17730 = n10487 ^ n10229 ^ 1'b0 ;
  assign n17731 = ~n17729 & n17730 ;
  assign n17732 = n3675 & n9543 ;
  assign n17733 = n3476 ^ n1620 ^ 1'b0 ;
  assign n17734 = n17732 | n17733 ;
  assign n17735 = n1616 ^ n722 ^ 1'b0 ;
  assign n17736 = n1085 & ~n17735 ;
  assign n17737 = ~n320 & n532 ;
  assign n17738 = n17737 ^ n1283 ^ 1'b0 ;
  assign n17739 = n17738 ^ n8653 ^ 1'b0 ;
  assign n17740 = n2517 & n5100 ;
  assign n17741 = n5620 ^ n929 ^ 1'b0 ;
  assign n17742 = n853 & ~n2259 ;
  assign n17743 = n17742 ^ n3534 ^ 1'b0 ;
  assign n17744 = n9258 & n17743 ;
  assign n17745 = n11140 & n17744 ;
  assign n17746 = n17745 ^ n2632 ^ 1'b0 ;
  assign n17747 = n1926 ^ n1836 ^ 1'b0 ;
  assign n17748 = n12404 ^ n2839 ^ 1'b0 ;
  assign n17749 = n4500 | n12835 ;
  assign n17750 = n1629 & n8261 ;
  assign n17751 = n4608 & n17750 ;
  assign n17752 = n1385 & n8735 ;
  assign n17753 = n10767 & n17752 ;
  assign n17757 = n1239 ^ n442 ^ 1'b0 ;
  assign n17754 = n5505 ^ n1045 ^ 1'b0 ;
  assign n17755 = n17451 | n17754 ;
  assign n17756 = n6722 | n17755 ;
  assign n17758 = n17757 ^ n17756 ^ 1'b0 ;
  assign n17759 = ~n5328 & n17628 ;
  assign n17760 = n8195 ^ n7683 ^ 1'b0 ;
  assign n17761 = n11197 | n17760 ;
  assign n17762 = n17761 ^ n5492 ^ 1'b0 ;
  assign n17763 = n5418 & ~n13905 ;
  assign n17764 = n4737 & ~n10671 ;
  assign n17765 = n17764 ^ n5505 ^ 1'b0 ;
  assign n17766 = ~n5861 & n17765 ;
  assign n17767 = n17766 ^ n7518 ^ n3871 ;
  assign n17768 = n12371 ^ n6412 ^ 1'b0 ;
  assign n17769 = n7168 & n17768 ;
  assign n17770 = n12596 & ~n17769 ;
  assign n17771 = n3524 & ~n16797 ;
  assign n17772 = n17771 ^ n1597 ^ 1'b0 ;
  assign n17773 = n3387 ^ n829 ^ 1'b0 ;
  assign n17774 = ( n7908 & n8223 ) | ( n7908 & n17773 ) | ( n8223 & n17773 ) ;
  assign n17775 = n14982 ^ x220 ^ 1'b0 ;
  assign n17776 = n6490 & ~n17775 ;
  assign n17777 = n3899 | n17776 ;
  assign n17778 = n17361 ^ n13110 ^ 1'b0 ;
  assign n17779 = n6616 | n12720 ;
  assign n17780 = n17779 ^ n16071 ^ 1'b0 ;
  assign n17781 = n862 | n17780 ;
  assign n17782 = n2072 | n4914 ;
  assign n17783 = n2482 & ~n17782 ;
  assign n17784 = n3556 & ~n17783 ;
  assign n17785 = n17784 ^ n6056 ^ 1'b0 ;
  assign n17786 = n4675 & n8485 ;
  assign n17787 = n8281 ^ n2099 ^ 1'b0 ;
  assign n17788 = ~n17786 & n17787 ;
  assign n17789 = n1282 & n17788 ;
  assign n17790 = ~n1499 & n14461 ;
  assign n17791 = n15975 ^ n7225 ^ 1'b0 ;
  assign n17792 = ~n7473 & n8338 ;
  assign n17793 = n8089 & ~n9254 ;
  assign n17794 = n17793 ^ n9033 ^ 1'b0 ;
  assign n17795 = ~n3528 & n16596 ;
  assign n17796 = n1505 & n17795 ;
  assign n17797 = n8004 & ~n9468 ;
  assign n17798 = n307 & ~n12423 ;
  assign n17799 = ~n1527 & n8974 ;
  assign n17800 = ~n1981 & n17799 ;
  assign n17801 = n7287 & ~n10559 ;
  assign n17802 = ~n1518 & n17801 ;
  assign n17803 = ~n15884 & n17802 ;
  assign n17804 = n7404 ^ n1249 ^ 1'b0 ;
  assign n17805 = ~n4395 & n17804 ;
  assign n17806 = x130 | n14246 ;
  assign n17807 = n10370 ^ n1190 ^ 1'b0 ;
  assign n17808 = n2072 | n17807 ;
  assign n17809 = n17806 | n17808 ;
  assign n17810 = ~n3197 & n6338 ;
  assign n17811 = n17810 ^ n8399 ^ 1'b0 ;
  assign n17812 = n6945 ^ n553 ^ 1'b0 ;
  assign n17813 = n955 & ~n17812 ;
  assign n17814 = n17813 ^ n1573 ^ 1'b0 ;
  assign n17815 = n8915 & ~n17814 ;
  assign n17816 = ~n14466 & n17815 ;
  assign n17817 = ( ~n7309 & n11705 ) | ( ~n7309 & n17816 ) | ( n11705 & n17816 ) ;
  assign n17818 = n17811 | n17817 ;
  assign n17819 = n5877 | n17818 ;
  assign n17820 = n4286 ^ n2315 ^ n1178 ;
  assign n17821 = n14382 ^ n5076 ^ 1'b0 ;
  assign n17822 = n16069 ^ n3237 ^ 1'b0 ;
  assign n17823 = n6617 ^ n950 ^ 1'b0 ;
  assign n17824 = n17822 & n17823 ;
  assign n17826 = n5343 ^ n4862 ^ n2116 ;
  assign n17825 = n15317 ^ n10885 ^ 1'b0 ;
  assign n17827 = n17826 ^ n17825 ^ 1'b0 ;
  assign n17828 = n17824 & ~n17827 ;
  assign n17829 = n2489 | n6665 ;
  assign n17830 = n5021 & ~n17829 ;
  assign n17831 = n15711 ^ n12614 ^ 1'b0 ;
  assign n17832 = n17831 ^ n2164 ^ 1'b0 ;
  assign n17833 = ~n11516 & n17832 ;
  assign n17834 = n15021 | n17833 ;
  assign n17835 = n557 & ~n4063 ;
  assign n17836 = n17835 ^ n5088 ^ 1'b0 ;
  assign n17837 = n17836 ^ n2469 ^ 1'b0 ;
  assign n17838 = n8947 ^ n7654 ^ 1'b0 ;
  assign n17839 = ~n1596 & n17838 ;
  assign n17840 = n17837 & n17839 ;
  assign n17841 = n14696 | n16902 ;
  assign n17842 = ~n11727 & n17841 ;
  assign n17843 = ~n442 & n4258 ;
  assign n17844 = n15719 & n17843 ;
  assign n17845 = n2891 & ~n6826 ;
  assign n17846 = ~n2291 & n6020 ;
  assign n17847 = n6986 | n17846 ;
  assign n17848 = n17847 ^ n14419 ^ 1'b0 ;
  assign n17849 = ~n5103 & n17848 ;
  assign n17851 = n14967 ^ n11172 ^ 1'b0 ;
  assign n17852 = n4331 & n17851 ;
  assign n17853 = n17852 ^ n4352 ^ 1'b0 ;
  assign n17850 = n5203 | n5440 ;
  assign n17854 = n17853 ^ n17850 ^ 1'b0 ;
  assign n17855 = n2949 | n15455 ;
  assign n17856 = n691 & ~n17855 ;
  assign n17857 = n8283 & ~n17856 ;
  assign n17858 = ~n2148 & n17857 ;
  assign n17859 = n2172 | n15322 ;
  assign n17860 = n2315 | n7851 ;
  assign n17861 = n8043 & ~n17860 ;
  assign n17862 = ~n17859 & n17861 ;
  assign n17863 = n7542 ^ n2791 ^ 1'b0 ;
  assign n17864 = n17560 & ~n17863 ;
  assign n17865 = n605 | n3870 ;
  assign n17866 = n2274 | n17865 ;
  assign n17867 = n17866 ^ n5926 ^ 1'b0 ;
  assign n17868 = n17867 ^ n2750 ^ 1'b0 ;
  assign n17869 = ( ~x226 & n7986 ) | ( ~x226 & n13717 ) | ( n7986 & n13717 ) ;
  assign n17870 = n17869 ^ n15316 ^ 1'b0 ;
  assign n17871 = n5613 ^ n3331 ^ n1684 ;
  assign n17872 = n14628 & n15745 ;
  assign n17873 = n1070 & n13551 ;
  assign n17874 = ~n3239 & n14418 ;
  assign n17875 = x191 & ~n3114 ;
  assign n17876 = n17874 & n17875 ;
  assign n17877 = n5225 & ~n11284 ;
  assign n17878 = n17876 | n17877 ;
  assign n17879 = n1159 | n17878 ;
  assign n17880 = x176 | n17219 ;
  assign n17881 = n17880 ^ n896 ^ 1'b0 ;
  assign n17882 = n5634 | n17881 ;
  assign n17883 = n3015 & n13630 ;
  assign n17884 = ~n1126 & n17883 ;
  assign n17885 = ~n13270 & n17884 ;
  assign n17886 = n16594 ^ n9717 ^ n7236 ;
  assign n17887 = n9661 ^ n6519 ^ 1'b0 ;
  assign n17888 = ~n1395 & n15673 ;
  assign n17889 = n6905 & n17888 ;
  assign n17890 = n2639 & ~n3595 ;
  assign n17891 = ~n2687 & n17890 ;
  assign n17892 = n3687 & ~n3875 ;
  assign n17893 = ~n8572 & n17892 ;
  assign n17894 = ( ~n2305 & n17891 ) | ( ~n2305 & n17893 ) | ( n17891 & n17893 ) ;
  assign n17895 = ~x124 & n3791 ;
  assign n17896 = n2893 ^ n2406 ^ x12 ;
  assign n17897 = ~x34 & n15340 ;
  assign n17898 = ~n1952 & n17897 ;
  assign n17899 = n11383 & n17898 ;
  assign n17900 = n16002 & n17806 ;
  assign n17901 = n2185 & n14504 ;
  assign n17902 = ~n3801 & n17901 ;
  assign n17903 = n17902 ^ n426 ^ 1'b0 ;
  assign n17904 = n8258 & ~n10955 ;
  assign n17905 = ~n666 & n17904 ;
  assign n17906 = n17905 ^ n6531 ^ 1'b0 ;
  assign n17907 = n8280 ^ n7108 ^ n2037 ;
  assign n17908 = n7696 ^ n1819 ^ 1'b0 ;
  assign n17909 = n3890 | n5396 ;
  assign n17910 = n5341 | n17909 ;
  assign n17911 = ( ~n13325 & n17908 ) | ( ~n13325 & n17910 ) | ( n17908 & n17910 ) ;
  assign n17912 = n4730 ^ x234 ^ 1'b0 ;
  assign n17913 = n12190 & n17061 ;
  assign n17914 = ~n2806 & n17913 ;
  assign n17915 = ~n9153 & n11680 ;
  assign n17916 = n305 | n16557 ;
  assign n17917 = ~x225 & n7419 ;
  assign n17918 = n7684 ^ n6993 ^ 1'b0 ;
  assign n17919 = n17917 & ~n17918 ;
  assign n17920 = n4071 | n11900 ;
  assign n17921 = n17920 ^ n2685 ^ 1'b0 ;
  assign n17922 = n6045 & ~n11486 ;
  assign n17923 = n11469 & n17922 ;
  assign n17924 = ~n6039 & n8524 ;
  assign n17925 = ~n4787 & n14426 ;
  assign n17926 = n876 & n9769 ;
  assign n17927 = n6330 & n11689 ;
  assign n17928 = n17927 ^ n2704 ^ 1'b0 ;
  assign n17929 = n13814 & ~n17928 ;
  assign n17930 = n17929 ^ n4491 ^ 1'b0 ;
  assign n17931 = n2839 | n8087 ;
  assign n17932 = n17931 ^ n7922 ^ 1'b0 ;
  assign n17933 = n10064 | n17932 ;
  assign n17934 = ~n4271 & n11419 ;
  assign n17935 = ~n4388 & n17934 ;
  assign n17936 = n5043 ^ n2852 ^ 1'b0 ;
  assign n17937 = n17936 ^ n4437 ^ 1'b0 ;
  assign n17938 = n2078 & n5707 ;
  assign n17939 = ~n7014 & n17938 ;
  assign n17940 = n4412 & n6493 ;
  assign n17941 = ~n2309 & n17940 ;
  assign n17942 = n6792 ^ n6205 ^ 1'b0 ;
  assign n17943 = ~n946 & n2354 ;
  assign n17944 = n4162 & ~n17943 ;
  assign n17945 = n10584 & ~n17944 ;
  assign n17946 = n17945 ^ n3240 ^ 1'b0 ;
  assign n17947 = n1404 | n5382 ;
  assign n17948 = n4313 & ~n17947 ;
  assign n17949 = n2232 & n17948 ;
  assign n17950 = n9052 | n14292 ;
  assign n17951 = n14114 ^ n7868 ^ 1'b0 ;
  assign n17952 = ~n6834 & n17951 ;
  assign n17953 = n3481 & n12071 ;
  assign n17954 = n14027 & n17953 ;
  assign n17955 = n8909 & ~n15611 ;
  assign n17956 = n5607 ^ n887 ^ 1'b0 ;
  assign n17957 = n840 & ~n17956 ;
  assign n17958 = n4395 & ~n15636 ;
  assign n17959 = n5984 | n13628 ;
  assign n17960 = n9629 | n17959 ;
  assign n17961 = n5711 | n11645 ;
  assign n17962 = n17961 ^ n2861 ^ 1'b0 ;
  assign n17963 = n13295 ^ n552 ^ 1'b0 ;
  assign n17964 = ~n17962 & n17963 ;
  assign n17965 = n17127 | n17209 ;
  assign n17966 = n8101 | n10385 ;
  assign n17967 = n17966 ^ n6084 ^ 1'b0 ;
  assign n17968 = n4185 & ~n17876 ;
  assign n17969 = n13679 & n17968 ;
  assign n17970 = n17969 ^ n4899 ^ 1'b0 ;
  assign n17971 = ~n5964 & n6328 ;
  assign n17975 = n880 & ~n6551 ;
  assign n17972 = n552 | n2021 ;
  assign n17973 = n17972 ^ n833 ^ 1'b0 ;
  assign n17974 = n4099 | n17973 ;
  assign n17976 = n17975 ^ n17974 ^ 1'b0 ;
  assign n17977 = n17976 ^ n11350 ^ 1'b0 ;
  assign n17978 = ~n17971 & n17977 ;
  assign n17979 = x28 | n14168 ;
  assign n17980 = n17979 ^ n3652 ^ n3348 ;
  assign n17981 = ~n736 & n17980 ;
  assign n17982 = n8408 ^ n5069 ^ 1'b0 ;
  assign n17983 = n3854 ^ n2964 ^ 1'b0 ;
  assign n17984 = n4691 & n17983 ;
  assign n17985 = ~n17982 & n17984 ;
  assign n17986 = n2336 & n15312 ;
  assign n17987 = ~n2336 & n17986 ;
  assign n17988 = n7477 | n17987 ;
  assign n17989 = n5509 ^ n4418 ^ 1'b0 ;
  assign n17990 = ~n17988 & n17989 ;
  assign n17991 = ~n3747 & n5193 ;
  assign n17992 = n10886 ^ n6023 ^ 1'b0 ;
  assign n17993 = x174 & n17992 ;
  assign n17994 = n10759 ^ n3052 ^ 1'b0 ;
  assign n17995 = n13783 & n17994 ;
  assign n17997 = ~n1006 & n5140 ;
  assign n17998 = n1006 & n17997 ;
  assign n17999 = ~n4257 & n17998 ;
  assign n18000 = ~n7210 & n17999 ;
  assign n18001 = n7210 & n18000 ;
  assign n17996 = n12568 & ~n14195 ;
  assign n18002 = n18001 ^ n17996 ^ 1'b0 ;
  assign n18003 = ~n2173 & n18002 ;
  assign n18004 = n18003 ^ x78 ^ 1'b0 ;
  assign n18005 = ~n13108 & n16619 ;
  assign n18006 = ~n5489 & n16627 ;
  assign n18007 = n4307 ^ n2080 ^ 1'b0 ;
  assign n18008 = ~n972 & n1668 ;
  assign n18009 = ~n1668 & n18008 ;
  assign n18010 = ~n994 & n18009 ;
  assign n18011 = n16919 | n18010 ;
  assign n18012 = n16919 & ~n18011 ;
  assign n18013 = n8390 & ~n16774 ;
  assign n18014 = n766 | n7194 ;
  assign n18015 = x1 & ~n18014 ;
  assign n18016 = n18015 ^ n10182 ^ 1'b0 ;
  assign n18020 = n1282 | n2836 ;
  assign n18021 = n1282 & ~n18020 ;
  assign n18017 = n786 & ~n2534 ;
  assign n18018 = n2534 & n18017 ;
  assign n18019 = n2035 & ~n18018 ;
  assign n18022 = n18021 ^ n18019 ^ 1'b0 ;
  assign n18023 = ~n1638 & n18022 ;
  assign n18024 = ~n9576 & n18023 ;
  assign n18025 = n10915 | n11856 ;
  assign n18026 = n18025 ^ n6931 ^ 1'b0 ;
  assign n18029 = n5417 & n7585 ;
  assign n18027 = n6208 & ~n8132 ;
  assign n18028 = n12736 & n18027 ;
  assign n18030 = n18029 ^ n18028 ^ 1'b0 ;
  assign n18031 = n2099 | n6907 ;
  assign n18032 = n8563 & ~n18031 ;
  assign n18033 = ~n8563 & n18032 ;
  assign n18034 = n2012 | n16776 ;
  assign n18035 = n6509 ^ n6073 ^ n3115 ;
  assign n18036 = ~n6842 & n18035 ;
  assign n18037 = n6297 ^ n4172 ^ 1'b0 ;
  assign n18038 = n3834 | n18037 ;
  assign n18039 = n18038 ^ n9589 ^ 1'b0 ;
  assign n18040 = n2909 | n8377 ;
  assign n18041 = n18040 ^ n1135 ^ 1'b0 ;
  assign n18042 = n6288 & n7559 ;
  assign n18043 = n18042 ^ n13003 ^ 1'b0 ;
  assign n18044 = n1723 | n8765 ;
  assign n18045 = n18044 ^ n2505 ^ 1'b0 ;
  assign n18046 = n1656 | n18045 ;
  assign n18047 = n1928 | n18046 ;
  assign n18048 = n3948 & n18047 ;
  assign n18049 = n3172 ^ n2314 ^ 1'b0 ;
  assign n18050 = n18049 ^ n10237 ^ 1'b0 ;
  assign n18051 = n956 & n13356 ;
  assign n18052 = n1658 & ~n6098 ;
  assign n18053 = n11495 & n18052 ;
  assign n18054 = n8430 | n18053 ;
  assign n18055 = n1345 | n18054 ;
  assign n18056 = ~n8631 & n9083 ;
  assign n18057 = n18056 ^ n6425 ^ 1'b0 ;
  assign n18058 = n14335 ^ n566 ^ 1'b0 ;
  assign n18059 = n7133 ^ n4526 ^ 1'b0 ;
  assign n18060 = n18059 ^ n7042 ^ 1'b0 ;
  assign n18061 = ~n18058 & n18060 ;
  assign n18062 = x124 & ~n1514 ;
  assign n18063 = n18062 ^ n13386 ^ 1'b0 ;
  assign n18064 = ( ~n9397 & n18061 ) | ( ~n9397 & n18063 ) | ( n18061 & n18063 ) ;
  assign n18065 = n444 & ~n15674 ;
  assign n18066 = n488 & n18065 ;
  assign n18067 = n8127 & ~n18066 ;
  assign n18068 = n3956 | n7493 ;
  assign n18069 = ( n4215 & n5942 ) | ( n4215 & ~n18068 ) | ( n5942 & ~n18068 ) ;
  assign n18070 = n18069 ^ n1068 ^ 1'b0 ;
  assign n18073 = ~n981 & n7431 ;
  assign n18074 = ~n4328 & n18073 ;
  assign n18071 = n3871 | n7507 ;
  assign n18072 = n18071 ^ n3666 ^ 1'b0 ;
  assign n18075 = n18074 ^ n18072 ^ 1'b0 ;
  assign n18076 = ~n13549 & n13931 ;
  assign n18077 = n14694 ^ n10217 ^ 1'b0 ;
  assign n18078 = ~n3005 & n18077 ;
  assign n18079 = n1703 & ~n18078 ;
  assign n18080 = ~n2331 & n6696 ;
  assign n18081 = n2210 | n3561 ;
  assign n18082 = n18081 ^ n5384 ^ 1'b0 ;
  assign n18083 = n3720 & n4375 ;
  assign n18084 = n18083 ^ n1861 ^ 1'b0 ;
  assign n18085 = n13981 & ~n18084 ;
  assign n18086 = n6180 & n18085 ;
  assign n18087 = n1487 & ~n18086 ;
  assign n18088 = n18087 ^ n2970 ^ 1'b0 ;
  assign n18089 = n18088 ^ n14815 ^ n2018 ;
  assign n18094 = ~n1656 & n13435 ;
  assign n18095 = n781 & n18094 ;
  assign n18090 = ~n5229 & n8773 ;
  assign n18091 = ~n1651 & n10642 ;
  assign n18092 = n18091 ^ n14022 ^ 1'b0 ;
  assign n18093 = n18090 & n18092 ;
  assign n18096 = n18095 ^ n18093 ^ 1'b0 ;
  assign n18097 = n9734 & ~n9986 ;
  assign n18098 = n18097 ^ n685 ^ 1'b0 ;
  assign n18099 = ~n9290 & n13547 ;
  assign n18100 = n4724 | n14930 ;
  assign n18101 = n18100 ^ n2411 ^ 1'b0 ;
  assign n18102 = n3045 | n3935 ;
  assign n18103 = n2311 ^ n2022 ^ 1'b0 ;
  assign n18104 = n18103 ^ n696 ^ 1'b0 ;
  assign n18105 = ~n9327 & n10689 ;
  assign n18106 = ~n918 & n16803 ;
  assign n18107 = n8667 | n11385 ;
  assign n18112 = ~n877 & n3920 ;
  assign n18108 = n3493 & n15626 ;
  assign n18109 = n18108 ^ n5709 ^ 1'b0 ;
  assign n18110 = n417 & ~n18109 ;
  assign n18111 = n18110 ^ n2421 ^ 1'b0 ;
  assign n18113 = n18112 ^ n18111 ^ n5521 ;
  assign n18114 = n3745 & ~n5971 ;
  assign n18115 = ~n1599 & n9769 ;
  assign n18116 = n18115 ^ n6432 ^ 1'b0 ;
  assign n18117 = n12785 & n18116 ;
  assign n18118 = n18117 ^ n12154 ^ n5955 ;
  assign n18119 = ~n331 & n392 ;
  assign n18120 = n7808 ^ n1698 ^ 1'b0 ;
  assign n18121 = n18119 & n18120 ;
  assign n18122 = n3059 ^ n343 ^ 1'b0 ;
  assign n18123 = n12256 & n17562 ;
  assign n18125 = ~n2011 & n3405 ;
  assign n18124 = n7789 | n13789 ;
  assign n18126 = n18125 ^ n18124 ^ 1'b0 ;
  assign n18127 = n17566 ^ x27 ^ 1'b0 ;
  assign n18128 = n18126 | n18127 ;
  assign n18129 = ~n2009 & n7039 ;
  assign n18130 = ~n1691 & n18129 ;
  assign n18131 = n6173 ^ n2320 ^ 1'b0 ;
  assign n18132 = n7241 ^ n663 ^ 1'b0 ;
  assign n18133 = ~n6102 & n15071 ;
  assign n18134 = n16002 ^ n3444 ^ 1'b0 ;
  assign n18135 = n1481 & n13802 ;
  assign n18136 = n18135 ^ n3659 ^ 1'b0 ;
  assign n18137 = ( n9786 & n18134 ) | ( n9786 & n18136 ) | ( n18134 & n18136 ) ;
  assign n18138 = n18137 ^ n11385 ^ 1'b0 ;
  assign n18139 = n15210 & n17900 ;
  assign n18140 = ~n11752 & n18139 ;
  assign n18141 = ~n896 & n1028 ;
  assign n18142 = n18141 ^ n18103 ^ 1'b0 ;
  assign n18143 = n1735 & n18142 ;
  assign n18144 = n3426 & ~n12012 ;
  assign n18145 = n18144 ^ n11607 ^ 1'b0 ;
  assign n18146 = n8584 ^ n1330 ^ 1'b0 ;
  assign n18147 = n2314 & ~n18146 ;
  assign n18148 = x100 | n12260 ;
  assign n18149 = ~n6527 & n18148 ;
  assign n18150 = n18149 ^ n498 ^ 1'b0 ;
  assign n18151 = ~n4336 & n15441 ;
  assign n18152 = n7486 & n18151 ;
  assign n18153 = ( ~n3575 & n6605 ) | ( ~n3575 & n8553 ) | ( n6605 & n8553 ) ;
  assign n18154 = n5929 | n11241 ;
  assign n18155 = n14099 ^ n13661 ^ 1'b0 ;
  assign n18157 = n2117 | n17046 ;
  assign n18158 = n12242 ^ n3437 ^ 1'b0 ;
  assign n18159 = n18157 & ~n18158 ;
  assign n18156 = n864 | n9122 ;
  assign n18160 = n18159 ^ n18156 ^ 1'b0 ;
  assign n18161 = n18160 ^ n5235 ^ n4576 ;
  assign n18162 = n9153 | n16489 ;
  assign n18163 = n4523 ^ n1139 ^ 1'b0 ;
  assign n18164 = n1336 & ~n18163 ;
  assign n18165 = n2342 & n12793 ;
  assign n18166 = ~n8547 & n18165 ;
  assign n18167 = n18166 ^ n4452 ^ 1'b0 ;
  assign n18168 = n7709 & ~n9545 ;
  assign n18169 = n6523 & n18168 ;
  assign n18170 = n18169 ^ n3461 ^ 1'b0 ;
  assign n18171 = ~n18167 & n18170 ;
  assign n18172 = n1657 & ~n5262 ;
  assign n18173 = n7367 & ~n18172 ;
  assign n18174 = n2276 & ~n18173 ;
  assign n18175 = n18174 ^ n774 ^ 1'b0 ;
  assign n18176 = n2640 ^ x160 ^ 1'b0 ;
  assign n18177 = n2185 ^ n708 ^ 1'b0 ;
  assign n18178 = ~n16717 & n18177 ;
  assign n18179 = n9029 & n18178 ;
  assign n18180 = n5312 & ~n8415 ;
  assign n18181 = n9029 ^ n5765 ^ 1'b0 ;
  assign n18182 = n12145 | n18181 ;
  assign n18183 = n5665 ^ x147 ^ 1'b0 ;
  assign n18184 = n8855 | n13110 ;
  assign n18185 = n12512 & ~n18184 ;
  assign n18186 = n4579 ^ n2814 ^ 1'b0 ;
  assign n18187 = n8211 ^ n5286 ^ 1'b0 ;
  assign n18188 = x176 & ~n3931 ;
  assign n18189 = n18188 ^ x92 ^ 1'b0 ;
  assign n18190 = n18187 | n18189 ;
  assign n18191 = n6213 ^ n2691 ^ 1'b0 ;
  assign n18196 = n8011 & n15233 ;
  assign n18192 = n7627 ^ n4158 ^ 1'b0 ;
  assign n18193 = n14238 ^ n9067 ^ 1'b0 ;
  assign n18194 = n14381 | n18193 ;
  assign n18195 = n18192 | n18194 ;
  assign n18197 = n18196 ^ n18195 ^ 1'b0 ;
  assign n18198 = ~n18191 & n18197 ;
  assign n18201 = n2246 & ~n5845 ;
  assign n18199 = n9208 & n16820 ;
  assign n18200 = n11520 & n18199 ;
  assign n18202 = n18201 ^ n18200 ^ n17928 ;
  assign n18203 = n17551 ^ n7340 ^ 1'b0 ;
  assign n18204 = n6991 | n18203 ;
  assign n18205 = n5519 ^ x219 ^ 1'b0 ;
  assign n18206 = n16744 & ~n18205 ;
  assign n18207 = n18206 ^ n2858 ^ 1'b0 ;
  assign n18208 = n18204 | n18207 ;
  assign n18209 = n2168 ^ n729 ^ 1'b0 ;
  assign n18210 = n17225 ^ n2855 ^ 1'b0 ;
  assign n18211 = n12563 & n18210 ;
  assign n18212 = ~n18209 & n18211 ;
  assign n18213 = ~n3308 & n5670 ;
  assign n18214 = n4104 ^ n2230 ^ 1'b0 ;
  assign n18215 = n3227 & n18214 ;
  assign n18216 = n18215 ^ n1128 ^ 1'b0 ;
  assign n18217 = n18213 & ~n18216 ;
  assign n18218 = n5907 & n13919 ;
  assign n18219 = ~n16390 & n18218 ;
  assign n18220 = ~n1569 & n4836 ;
  assign n18221 = n18220 ^ n6083 ^ 1'b0 ;
  assign n18222 = n1847 & ~n18221 ;
  assign n18223 = n5072 | n12069 ;
  assign n18224 = n18223 ^ n12460 ^ 1'b0 ;
  assign n18225 = n325 | n2065 ;
  assign n18226 = n18225 ^ n1195 ^ 1'b0 ;
  assign n18227 = n18226 ^ n4077 ^ 1'b0 ;
  assign n18228 = n8768 & n18227 ;
  assign n18229 = n860 & n9323 ;
  assign n18230 = n2011 & n8430 ;
  assign n18231 = n18229 & n18230 ;
  assign n18233 = n10758 & n16396 ;
  assign n18234 = n18233 ^ n17973 ^ n2343 ;
  assign n18232 = n5950 & n7162 ;
  assign n18235 = n18234 ^ n18232 ^ 1'b0 ;
  assign n18236 = n8632 | n14800 ;
  assign n18237 = n18236 ^ n16884 ^ 1'b0 ;
  assign n18238 = n16867 ^ n13956 ^ 1'b0 ;
  assign n18239 = n1094 & n18238 ;
  assign n18240 = n7288 ^ n5176 ^ 1'b0 ;
  assign n18241 = n3102 & ~n6337 ;
  assign n18242 = n18241 ^ n14381 ^ 1'b0 ;
  assign n18243 = n3551 & ~n18242 ;
  assign n18244 = n8499 & n18243 ;
  assign n18245 = n6684 ^ n5433 ^ 1'b0 ;
  assign n18246 = n5838 & n10530 ;
  assign n18247 = ~n2776 & n3210 ;
  assign n18248 = n3466 ^ n1709 ^ 1'b0 ;
  assign n18249 = n1451 | n18248 ;
  assign n18250 = x248 & ~n10425 ;
  assign n18251 = ~n5653 & n18250 ;
  assign n18253 = n3982 ^ n1974 ^ 1'b0 ;
  assign n18252 = n1451 & n18103 ;
  assign n18254 = n18253 ^ n18252 ^ 1'b0 ;
  assign n18255 = n10407 & n10692 ;
  assign n18256 = n7830 & ~n9863 ;
  assign n18257 = n4497 & ~n11226 ;
  assign n18258 = ~n9548 & n18257 ;
  assign n18259 = ~n5023 & n10942 ;
  assign n18260 = ~n5027 & n18259 ;
  assign n18261 = n2632 | n12163 ;
  assign n18262 = n18260 & ~n18261 ;
  assign n18263 = n10112 ^ n7020 ^ n4611 ;
  assign n18264 = n18263 ^ n728 ^ 1'b0 ;
  assign n18265 = ~n4938 & n10869 ;
  assign n18266 = n1610 & ~n14755 ;
  assign n18273 = n1831 & ~n15646 ;
  assign n18267 = n872 & n4295 ;
  assign n18268 = n18267 ^ x27 ^ 1'b0 ;
  assign n18269 = x235 & n2896 ;
  assign n18270 = n18268 & n18269 ;
  assign n18271 = n1604 & ~n18270 ;
  assign n18272 = n9978 & n18271 ;
  assign n18274 = n18273 ^ n18272 ^ 1'b0 ;
  assign n18275 = n5591 & n7446 ;
  assign n18276 = ~n1828 & n2443 ;
  assign n18277 = n6832 & n18276 ;
  assign n18278 = n18277 ^ n5442 ^ 1'b0 ;
  assign n18279 = n13470 ^ n3541 ^ 1'b0 ;
  assign n18280 = n12930 ^ n4094 ^ 1'b0 ;
  assign n18281 = n9326 ^ n7266 ^ 1'b0 ;
  assign n18282 = n14524 ^ n273 ^ 1'b0 ;
  assign n18283 = n16154 & ~n18282 ;
  assign n18284 = n2557 & ~n5136 ;
  assign n18285 = ( n4500 & ~n13077 ) | ( n4500 & n13572 ) | ( ~n13077 & n13572 ) ;
  assign n18286 = n16580 ^ n9932 ^ 1'b0 ;
  assign n18287 = n18286 ^ n1661 ^ 1'b0 ;
  assign n18288 = ~n5571 & n18287 ;
  assign n18289 = n5875 ^ n552 ^ 1'b0 ;
  assign n18290 = n1512 & n14299 ;
  assign n18291 = ~n510 & n18290 ;
  assign n18292 = n15853 ^ n14581 ^ 1'b0 ;
  assign n18293 = n1073 & ~n16175 ;
  assign n18294 = n14940 ^ n412 ^ 1'b0 ;
  assign n18295 = n8376 ^ n2371 ^ 1'b0 ;
  assign n18298 = n2640 & ~n10488 ;
  assign n18299 = n18298 ^ n3970 ^ 1'b0 ;
  assign n18296 = n11171 ^ n1415 ^ 1'b0 ;
  assign n18297 = n9835 | n18296 ;
  assign n18300 = n18299 ^ n18297 ^ 1'b0 ;
  assign n18306 = n15598 ^ n10437 ^ 1'b0 ;
  assign n18307 = n4799 & ~n18306 ;
  assign n18308 = ~n7902 & n11474 ;
  assign n18309 = ~n18307 & n18308 ;
  assign n18310 = n18309 ^ n15532 ^ 1'b0 ;
  assign n18301 = n14187 ^ n11231 ^ 1'b0 ;
  assign n18302 = n397 | n18301 ;
  assign n18303 = n8457 & ~n18302 ;
  assign n18304 = ~n10144 & n18303 ;
  assign n18305 = n5799 & ~n18304 ;
  assign n18311 = n18310 ^ n18305 ^ n1974 ;
  assign n18312 = n7133 & n17486 ;
  assign n18313 = n3333 | n5250 ;
  assign n18314 = n17971 | n18313 ;
  assign n18315 = n18314 ^ n16734 ^ n11171 ;
  assign n18316 = n14000 ^ n2466 ^ 1'b0 ;
  assign n18317 = n8645 & n18316 ;
  assign n18318 = n3331 ^ x67 ^ 1'b0 ;
  assign n18319 = n3217 | n18318 ;
  assign n18323 = n1146 | n2546 ;
  assign n18324 = n782 | n18323 ;
  assign n18320 = n9515 ^ n2706 ^ 1'b0 ;
  assign n18321 = n6023 & n18320 ;
  assign n18322 = n18321 ^ n8703 ^ 1'b0 ;
  assign n18325 = n18324 ^ n18322 ^ 1'b0 ;
  assign n18326 = n15546 & ~n18325 ;
  assign n18327 = ( ~x253 & n4749 ) | ( ~x253 & n11607 ) | ( n4749 & n11607 ) ;
  assign n18328 = n8083 & ~n15605 ;
  assign n18329 = n18328 ^ n11729 ^ 1'b0 ;
  assign n18330 = ~n7384 & n18329 ;
  assign n18331 = n14497 | n17506 ;
  assign n18332 = x61 & x169 ;
  assign n18333 = n18268 & n18332 ;
  assign n18334 = ~n3016 & n18333 ;
  assign n18335 = n5338 | n13723 ;
  assign n18336 = n18335 ^ n10430 ^ 1'b0 ;
  assign n18337 = n10323 ^ x82 ^ 1'b0 ;
  assign n18338 = x89 & ~n2046 ;
  assign n18339 = n10440 ^ n5659 ^ 1'b0 ;
  assign n18340 = ~n18338 & n18339 ;
  assign n18341 = n12128 ^ n6772 ^ 1'b0 ;
  assign n18342 = n18341 ^ n3195 ^ 1'b0 ;
  assign n18343 = ~n4115 & n7646 ;
  assign n18344 = n18343 ^ n3725 ^ 1'b0 ;
  assign n18345 = ~n2846 & n2977 ;
  assign n18346 = n18345 ^ n3213 ^ 1'b0 ;
  assign n18347 = n6493 & n7634 ;
  assign n18348 = ~n4080 & n18347 ;
  assign n18349 = n877 | n8754 ;
  assign n18350 = n7712 | n18349 ;
  assign n18351 = n18350 ^ n6308 ^ 1'b0 ;
  assign n18352 = n6087 ^ n354 ^ 1'b0 ;
  assign n18353 = n7845 | n18352 ;
  assign n18355 = n5575 | n10189 ;
  assign n18354 = n16843 & n17887 ;
  assign n18356 = n18355 ^ n18354 ^ 1'b0 ;
  assign n18357 = n1402 & n13651 ;
  assign n18358 = n2972 & n18357 ;
  assign n18359 = n18358 ^ n12926 ^ 1'b0 ;
  assign n18360 = n1360 & ~n15203 ;
  assign n18361 = n12922 & ~n17814 ;
  assign n18362 = ~n18360 & n18361 ;
  assign n18363 = ~n2993 & n3842 ;
  assign n18364 = n1673 & n18363 ;
  assign n18365 = n3917 | n18364 ;
  assign n18366 = n18365 ^ n6842 ^ 1'b0 ;
  assign n18367 = n18362 & ~n18366 ;
  assign n18368 = ~n18362 & n18367 ;
  assign n18369 = ~n8944 & n15224 ;
  assign n18370 = n18369 ^ n3819 ^ 1'b0 ;
  assign n18371 = n2720 & n18370 ;
  assign n18372 = ~n1451 & n15130 ;
  assign n18373 = ~n15130 & n18372 ;
  assign n18374 = n11397 & ~n18373 ;
  assign n18375 = n18373 & n18374 ;
  assign n18376 = n16903 & ~n18364 ;
  assign n18377 = n9737 & n18376 ;
  assign n18378 = x24 & ~n3473 ;
  assign n18379 = n18378 ^ n15537 ^ 1'b0 ;
  assign n18380 = n9076 ^ n4376 ^ 1'b0 ;
  assign n18381 = n18380 ^ n2507 ^ n1299 ;
  assign n18382 = n5914 ^ n4815 ^ 1'b0 ;
  assign n18383 = n18381 & ~n18382 ;
  assign n18384 = ~n3741 & n7419 ;
  assign n18385 = n1537 | n2687 ;
  assign n18386 = n18384 & ~n18385 ;
  assign n18387 = ( ~n1453 & n2629 ) | ( ~n1453 & n9440 ) | ( n2629 & n9440 ) ;
  assign n18388 = n18387 ^ n15532 ^ n4919 ;
  assign n18389 = n5564 & ~n7907 ;
  assign n18390 = ~n6049 & n12057 ;
  assign n18392 = n1944 ^ n1529 ^ 1'b0 ;
  assign n18391 = n1882 | n2307 ;
  assign n18393 = n18392 ^ n18391 ^ 1'b0 ;
  assign n18394 = n2519 | n18393 ;
  assign n18395 = n1252 & ~n9617 ;
  assign n18396 = n18395 ^ n2822 ^ 1'b0 ;
  assign n18397 = n2827 | n9484 ;
  assign n18398 = n13252 ^ n1831 ^ 1'b0 ;
  assign n18399 = n7166 & ~n18398 ;
  assign n18400 = n18399 ^ n8947 ^ 1'b0 ;
  assign n18401 = n5746 & ~n9019 ;
  assign n18402 = n7516 ^ n482 ^ 1'b0 ;
  assign n18403 = n1247 & n4799 ;
  assign n18404 = n17363 & n18403 ;
  assign n18405 = n14158 ^ n13988 ^ n3676 ;
  assign n18407 = ~n1050 & n11402 ;
  assign n18406 = n3140 & n3727 ;
  assign n18408 = n18407 ^ n18406 ^ 1'b0 ;
  assign n18409 = n15887 & n18408 ;
  assign n18411 = n1186 & n14693 ;
  assign n18412 = ~n12803 & n18411 ;
  assign n18410 = n18165 ^ n6370 ^ 1'b0 ;
  assign n18413 = n18412 ^ n18410 ^ 1'b0 ;
  assign n18414 = n3524 ^ n3180 ^ 1'b0 ;
  assign n18415 = n887 | n18414 ;
  assign n18416 = n1337 ^ n992 ^ 1'b0 ;
  assign n18417 = n2107 & ~n18416 ;
  assign n18418 = n1049 & n18417 ;
  assign n18419 = n6582 | n9475 ;
  assign n18420 = ~n3247 & n9926 ;
  assign n18422 = n7190 ^ n1965 ^ 1'b0 ;
  assign n18421 = n6071 & n9996 ;
  assign n18423 = n18422 ^ n18421 ^ 1'b0 ;
  assign n18424 = n8242 | n18423 ;
  assign n18425 = ~n9177 & n18424 ;
  assign n18426 = n2918 & ~n5311 ;
  assign n18427 = n18426 ^ n5005 ^ 1'b0 ;
  assign n18428 = ~n10663 & n12658 ;
  assign n18429 = n18428 ^ n12351 ^ 1'b0 ;
  assign n18430 = n18427 & ~n18429 ;
  assign n18431 = n10120 & ~n18430 ;
  assign n18432 = n3212 & n10334 ;
  assign n18433 = x155 & ~n18432 ;
  assign n18434 = n9823 | n10221 ;
  assign n18435 = n8386 ^ n2457 ^ 1'b0 ;
  assign n18436 = n8386 & ~n18435 ;
  assign n18437 = ~n8655 & n18436 ;
  assign n18438 = n15898 | n18437 ;
  assign n18439 = n4145 ^ n3150 ^ 1'b0 ;
  assign n18440 = n4120 & n5217 ;
  assign n18441 = n4351 & ~n10166 ;
  assign n18442 = n3618 & ~n18441 ;
  assign n18443 = n11857 & ~n12569 ;
  assign n18444 = n2697 & n7450 ;
  assign n18447 = n9915 ^ n6974 ^ n3308 ;
  assign n18448 = n18447 ^ n13778 ^ n4671 ;
  assign n18445 = n793 & n7868 ;
  assign n18446 = n14897 & n18445 ;
  assign n18449 = n18448 ^ n18446 ^ 1'b0 ;
  assign n18450 = n7773 & ~n17542 ;
  assign n18451 = n18450 ^ n16911 ^ 1'b0 ;
  assign n18452 = n1366 | n6803 ;
  assign n18453 = n18451 & ~n18452 ;
  assign n18454 = n6672 ^ n5288 ^ 1'b0 ;
  assign n18455 = ~n3127 & n14492 ;
  assign n18456 = n14244 ^ n11004 ^ 1'b0 ;
  assign n18457 = n5420 | n15675 ;
  assign n18458 = n12178 | n18457 ;
  assign n18459 = ~n2103 & n6266 ;
  assign n18460 = n18459 ^ n974 ^ 1'b0 ;
  assign n18461 = n3038 & ~n18460 ;
  assign n18462 = n18461 ^ n6171 ^ 1'b0 ;
  assign n18463 = n11424 & n14276 ;
  assign n18464 = ~n2978 & n18463 ;
  assign n18465 = n18464 ^ n975 ^ 1'b0 ;
  assign n18466 = n3580 & ~n10005 ;
  assign n18467 = n5107 & ~n18466 ;
  assign n18468 = n551 | n4076 ;
  assign n18469 = ~n2929 & n18468 ;
  assign n18470 = n18469 ^ n12016 ^ 1'b0 ;
  assign n18471 = n1087 | n5591 ;
  assign n18472 = n12021 ^ n5031 ^ 1'b0 ;
  assign n18473 = ~n10374 & n18472 ;
  assign n18474 = n18471 ^ n8246 ^ 1'b0 ;
  assign n18475 = n6434 | n9781 ;
  assign n18476 = n18475 ^ n14066 ^ 1'b0 ;
  assign n18477 = n6570 ^ n1261 ^ 1'b0 ;
  assign n18478 = n3022 & n7108 ;
  assign n18479 = n18477 & n18478 ;
  assign n18480 = n18479 ^ n7362 ^ 1'b0 ;
  assign n18481 = ~n5400 & n18480 ;
  assign n18482 = n13952 & ~n15822 ;
  assign n18483 = n5848 ^ x25 ^ 1'b0 ;
  assign n18484 = n2116 | n18483 ;
  assign n18485 = n9352 ^ n7280 ^ 1'b0 ;
  assign n18486 = ~n7144 & n9018 ;
  assign n18487 = n8388 | n11271 ;
  assign n18488 = n18487 ^ n3181 ^ 1'b0 ;
  assign n18489 = n1402 & n18488 ;
  assign n18490 = n7595 & ~n8415 ;
  assign n18491 = n18490 ^ n3076 ^ 1'b0 ;
  assign n18492 = n6273 ^ n3451 ^ 1'b0 ;
  assign n18493 = n2466 & n4199 ;
  assign n18494 = n18493 ^ n12230 ^ 1'b0 ;
  assign n18495 = n1139 ^ x172 ^ 1'b0 ;
  assign n18496 = n18494 | n18495 ;
  assign n18497 = n3371 | n18496 ;
  assign n18498 = n18497 ^ n11241 ^ 1'b0 ;
  assign n18499 = n8012 & ~n8092 ;
  assign n18500 = n8092 & n18499 ;
  assign n18502 = n9477 ^ n7992 ^ n5879 ;
  assign n18501 = n1105 & ~n4002 ;
  assign n18503 = n18502 ^ n18501 ^ 1'b0 ;
  assign n18504 = n5442 | n18503 ;
  assign n18505 = n4138 ^ n3841 ^ 1'b0 ;
  assign n18506 = n18505 ^ n1974 ^ 1'b0 ;
  assign n18507 = n1062 & n12680 ;
  assign n18508 = n1223 | n8748 ;
  assign n18509 = n13030 ^ n7430 ^ 1'b0 ;
  assign n18510 = n18508 | n18509 ;
  assign n18511 = n18507 & ~n18510 ;
  assign n18512 = ~x115 & n18511 ;
  assign n18513 = x23 & n2910 ;
  assign n18514 = n2860 | n8254 ;
  assign n18515 = n18514 ^ n16883 ^ 1'b0 ;
  assign n18516 = n10678 & n10716 ;
  assign n18517 = n18516 ^ n1622 ^ 1'b0 ;
  assign n18518 = n9004 ^ n2330 ^ 1'b0 ;
  assign n18519 = n5577 | n18518 ;
  assign n18520 = n18519 ^ n14442 ^ 1'b0 ;
  assign n18521 = n7914 ^ n4879 ^ 1'b0 ;
  assign n18522 = n9530 | n15509 ;
  assign n18523 = n651 & ~n18522 ;
  assign n18524 = n12957 & ~n18107 ;
  assign n18525 = x86 & ~n5399 ;
  assign n18526 = n15309 & n18525 ;
  assign n18527 = ~n13051 & n18526 ;
  assign n18528 = n9339 | n18527 ;
  assign n18529 = n5938 & ~n18528 ;
  assign n18530 = n3186 & n5887 ;
  assign n18531 = n4629 | n4972 ;
  assign n18533 = n1740 & n13507 ;
  assign n18534 = n10931 & n18533 ;
  assign n18532 = n988 | n18212 ;
  assign n18535 = n18534 ^ n18532 ^ 1'b0 ;
  assign n18536 = n12351 ^ n10049 ^ 1'b0 ;
  assign n18537 = n7603 & ~n18536 ;
  assign n18538 = x140 & ~n3323 ;
  assign n18539 = ~n841 & n18538 ;
  assign n18540 = n18539 ^ n6193 ^ 1'b0 ;
  assign n18541 = n5027 & ~n18540 ;
  assign n18542 = n3965 & n13727 ;
  assign n18543 = n7516 & n18542 ;
  assign n18544 = ~n1126 & n14972 ;
  assign n18545 = n13366 & n18544 ;
  assign n18546 = n1337 & n8303 ;
  assign n18547 = n18546 ^ n17958 ^ 1'b0 ;
  assign n18548 = n1732 & ~n3540 ;
  assign n18549 = n18548 ^ n926 ^ 1'b0 ;
  assign n18550 = n3359 & ~n18549 ;
  assign n18551 = n18550 ^ n1588 ^ 1'b0 ;
  assign n18552 = n18547 & ~n18551 ;
  assign n18553 = n5643 ^ n1701 ^ 1'b0 ;
  assign n18554 = n17563 ^ n15033 ^ 1'b0 ;
  assign n18555 = n9236 & n11395 ;
  assign n18557 = ~n16778 & n18302 ;
  assign n18556 = x213 & n836 ;
  assign n18558 = n18557 ^ n18556 ^ 1'b0 ;
  assign n18559 = n13062 ^ n1379 ^ 1'b0 ;
  assign n18560 = n10092 ^ n4701 ^ 1'b0 ;
  assign n18561 = n18559 | n18560 ;
  assign n18562 = ~n2555 & n13365 ;
  assign n18563 = n18562 ^ n8485 ^ 1'b0 ;
  assign n18564 = n4949 & n8051 ;
  assign n18565 = n7959 & n18564 ;
  assign n18566 = n18565 ^ n17301 ^ 1'b0 ;
  assign n18567 = x169 & n1112 ;
  assign n18568 = n18567 ^ n3377 ^ 1'b0 ;
  assign n18569 = ~n3518 & n3966 ;
  assign n18570 = ~n4510 & n18569 ;
  assign n18571 = n18568 & ~n18570 ;
  assign n18572 = n2159 & n2977 ;
  assign n18573 = n17618 ^ n11999 ^ 1'b0 ;
  assign n18574 = n13271 ^ n6322 ^ 1'b0 ;
  assign n18575 = n3358 & ~n4313 ;
  assign n18576 = n18575 ^ n1727 ^ 1'b0 ;
  assign n18577 = n2097 ^ n1742 ^ 1'b0 ;
  assign n18578 = n13727 & n18577 ;
  assign n18579 = ~n18119 & n18578 ;
  assign n18580 = ~n18576 & n18579 ;
  assign n18581 = n9781 ^ x27 ^ 1'b0 ;
  assign n18582 = n18581 ^ n12084 ^ n2577 ;
  assign n18583 = n11888 ^ n3331 ^ 1'b0 ;
  assign n18584 = n4290 & ~n18583 ;
  assign n18585 = n5195 ^ n327 ^ 1'b0 ;
  assign n18586 = ~n456 & n1859 ;
  assign n18587 = n3741 & ~n18586 ;
  assign n18588 = n18587 ^ n998 ^ 1'b0 ;
  assign n18589 = n17926 & n18588 ;
  assign n18590 = n10935 ^ n9027 ^ 1'b0 ;
  assign n18591 = n2655 | n14757 ;
  assign n18592 = n8492 ^ n4126 ^ 1'b0 ;
  assign n18593 = n18591 & n18592 ;
  assign n18594 = ~n18590 & n18593 ;
  assign n18595 = n18594 ^ x219 ^ 1'b0 ;
  assign n18596 = n6477 & ~n8796 ;
  assign n18597 = n8796 & n18596 ;
  assign n18598 = n16503 ^ n692 ^ 1'b0 ;
  assign n18599 = n5316 & n12279 ;
  assign n18600 = n1546 & n4512 ;
  assign n18601 = n18600 ^ n11751 ^ 1'b0 ;
  assign n18602 = x106 & ~n18601 ;
  assign n18603 = n18602 ^ n2590 ^ 1'b0 ;
  assign n18604 = n2720 ^ x244 ^ 1'b0 ;
  assign n18605 = n10175 ^ n8767 ^ n4370 ;
  assign n18606 = n8245 ^ n7355 ^ 1'b0 ;
  assign n18607 = n18605 & n18606 ;
  assign n18608 = ~n3462 & n18289 ;
  assign n18609 = ( n7151 & n7509 ) | ( n7151 & ~n18608 ) | ( n7509 & ~n18608 ) ;
  assign n18610 = n18609 ^ n9966 ^ 1'b0 ;
  assign n18611 = n15898 | n18610 ;
  assign n18612 = n11148 ^ n4485 ^ 1'b0 ;
  assign n18613 = n1247 & n18612 ;
  assign n18614 = n2275 & n15911 ;
  assign n18615 = ~n18613 & n18614 ;
  assign n18616 = n3676 ^ n2841 ^ 1'b0 ;
  assign n18617 = n754 & n18616 ;
  assign n18618 = n3953 & ~n6938 ;
  assign n18619 = n9592 & n18618 ;
  assign n18620 = ( ~n1062 & n18617 ) | ( ~n1062 & n18619 ) | ( n18617 & n18619 ) ;
  assign n18622 = n17005 ^ n4350 ^ 1'b0 ;
  assign n18621 = x211 & n15515 ;
  assign n18623 = n18622 ^ n18621 ^ 1'b0 ;
  assign n18624 = ~n476 & n4039 ;
  assign n18625 = n18624 ^ n6412 ^ n1232 ;
  assign n18626 = n10144 & n18625 ;
  assign n18627 = ~n3054 & n7212 ;
  assign n18628 = x106 & ~n4267 ;
  assign n18629 = ~n18627 & n18628 ;
  assign n18630 = n18629 ^ n7144 ^ 1'b0 ;
  assign n18632 = n2606 & n6315 ;
  assign n18633 = n18632 ^ n5645 ^ n5107 ;
  assign n18631 = ~x226 & n16640 ;
  assign n18634 = n18633 ^ n18631 ^ 1'b0 ;
  assign n18635 = n5665 & ~n16228 ;
  assign n18636 = n13890 & n18635 ;
  assign n18637 = n2968 ^ x141 ^ 1'b0 ;
  assign n18638 = n6642 & n18637 ;
  assign n18640 = n7361 ^ n5292 ^ 1'b0 ;
  assign n18639 = n12798 & ~n14682 ;
  assign n18641 = n18640 ^ n18639 ^ 1'b0 ;
  assign n18642 = ~n9464 & n9902 ;
  assign n18643 = ~n10555 & n18642 ;
  assign n18644 = n18643 ^ n4564 ^ 1'b0 ;
  assign n18645 = n18644 ^ n14563 ^ 1'b0 ;
  assign n18646 = n8967 & n18645 ;
  assign n18647 = n1009 | n14410 ;
  assign n18648 = n3059 & ~n18647 ;
  assign n18649 = n16186 ^ x251 ^ 1'b0 ;
  assign n18650 = n793 & n3235 ;
  assign n18651 = ~n2006 & n18650 ;
  assign n18655 = n728 & n4949 ;
  assign n18656 = n17629 ^ n8724 ^ 1'b0 ;
  assign n18657 = n18655 & n18656 ;
  assign n18658 = n3505 & n18657 ;
  assign n18659 = n1447 | n18658 ;
  assign n18660 = n18659 ^ n1221 ^ 1'b0 ;
  assign n18652 = x224 & ~n703 ;
  assign n18653 = n4361 & n18652 ;
  assign n18654 = n18653 ^ n2589 ^ 1'b0 ;
  assign n18661 = n18660 ^ n18654 ^ 1'b0 ;
  assign n18662 = ~n8602 & n16463 ;
  assign n18663 = ~n3033 & n18662 ;
  assign n18664 = n12860 ^ n1529 ^ 1'b0 ;
  assign n18665 = x125 | n1663 ;
  assign n18666 = n15003 ^ n10942 ^ 1'b0 ;
  assign n18667 = n5095 | n9277 ;
  assign n18668 = n18667 ^ n2061 ^ 1'b0 ;
  assign n18669 = n8600 ^ n6036 ^ 1'b0 ;
  assign n18670 = n13439 & n18669 ;
  assign n18671 = ( n8438 & n18668 ) | ( n8438 & ~n18670 ) | ( n18668 & ~n18670 ) ;
  assign n18672 = ~x163 & n7039 ;
  assign n18673 = ~n2855 & n4393 ;
  assign n18675 = n5114 ^ n305 ^ 1'b0 ;
  assign n18676 = n1214 & ~n18675 ;
  assign n18677 = n18676 ^ n13603 ^ n4086 ;
  assign n18674 = n4731 | n7036 ;
  assign n18678 = n18677 ^ n18674 ^ 1'b0 ;
  assign n18679 = n18678 ^ n10432 ^ n1404 ;
  assign n18680 = n9597 ^ n800 ^ 1'b0 ;
  assign n18681 = n3342 & n8673 ;
  assign n18682 = n18680 & n18681 ;
  assign n18683 = n18530 ^ n14560 ^ 1'b0 ;
  assign n18684 = ~n1145 & n18683 ;
  assign n18685 = n5271 | n18600 ;
  assign n18686 = n13845 ^ n3703 ^ 1'b0 ;
  assign n18687 = n6149 ^ n5253 ^ x202 ;
  assign n18688 = n5519 & ~n14794 ;
  assign n18689 = n17386 | n18236 ;
  assign n18690 = n4650 & n6271 ;
  assign n18691 = n2513 & ~n10815 ;
  assign n18692 = n1697 | n12708 ;
  assign n18693 = ~n5399 & n18692 ;
  assign n18694 = n8195 | n10473 ;
  assign n18695 = n3552 | n8730 ;
  assign n18696 = n18695 ^ n17550 ^ 1'b0 ;
  assign n18697 = x208 | n9802 ;
  assign n18698 = n18697 ^ n1623 ^ 1'b0 ;
  assign n18699 = n611 & ~n8474 ;
  assign n18700 = ~n8685 & n18699 ;
  assign n18701 = n18700 ^ n3181 ^ 1'b0 ;
  assign n18702 = ~n10692 & n18701 ;
  assign n18703 = n8921 ^ n4724 ^ 1'b0 ;
  assign n18704 = ~n17282 & n18703 ;
  assign n18705 = n16109 ^ n8256 ^ 1'b0 ;
  assign n18706 = n354 & ~n7894 ;
  assign n18707 = n12236 ^ n5835 ^ 1'b0 ;
  assign n18708 = n1880 & ~n8359 ;
  assign n18709 = n18708 ^ x24 ^ 1'b0 ;
  assign n18710 = x254 | n6363 ;
  assign n18711 = n18709 & ~n18710 ;
  assign n18713 = ~n10321 & n15054 ;
  assign n18714 = n13020 & n18713 ;
  assign n18712 = n8256 | n10838 ;
  assign n18715 = n18714 ^ n18712 ^ 1'b0 ;
  assign n18716 = n2526 | n8693 ;
  assign n18717 = n10653 | n18716 ;
  assign n18718 = ~n3235 & n7637 ;
  assign n18719 = n18718 ^ n15537 ^ 1'b0 ;
  assign n18720 = n18719 ^ n2762 ^ 1'b0 ;
  assign n18721 = n17110 & ~n18720 ;
  assign n18722 = n5314 & ~n7858 ;
  assign n18723 = ~n3414 & n18722 ;
  assign n18724 = n3020 & ~n18723 ;
  assign n18725 = ~n3980 & n18724 ;
  assign n18726 = n3377 & ~n18725 ;
  assign n18727 = n18726 ^ n12030 ^ 1'b0 ;
  assign n18728 = n17572 & n18727 ;
  assign n18729 = n18728 ^ n4743 ^ 1'b0 ;
  assign n18733 = n1974 ^ n638 ^ 1'b0 ;
  assign n18734 = x103 & ~n18733 ;
  assign n18735 = n6403 & n18734 ;
  assign n18736 = n8189 & n18735 ;
  assign n18730 = n1544 & n4327 ;
  assign n18731 = n4459 ^ n700 ^ 1'b0 ;
  assign n18732 = n18730 | n18731 ;
  assign n18737 = n18736 ^ n18732 ^ 1'b0 ;
  assign n18738 = n7103 & ~n9126 ;
  assign n18739 = n8465 & n18738 ;
  assign n18740 = n4532 & n8645 ;
  assign n18741 = n6541 & n8340 ;
  assign n18742 = n18741 ^ n11469 ^ 1'b0 ;
  assign n18743 = n9035 ^ n5064 ^ 1'b0 ;
  assign n18744 = ~n11578 & n18743 ;
  assign n18745 = n11131 & n12293 ;
  assign n18746 = ~n11285 & n18745 ;
  assign n18747 = n4412 & n11218 ;
  assign n18748 = ~n1556 & n18747 ;
  assign n18749 = ~n18746 & n18748 ;
  assign n18750 = n16546 ^ n5008 ^ n1423 ;
  assign n18751 = n3333 & ~n3676 ;
  assign n18752 = n5341 ^ n3458 ^ 1'b0 ;
  assign n18753 = n11014 | n18752 ;
  assign n18754 = n7708 & n18753 ;
  assign n18755 = ~n14908 & n18754 ;
  assign n18756 = n18755 ^ n11658 ^ 1'b0 ;
  assign n18757 = n7471 & ~n18756 ;
  assign n18758 = n18315 ^ n897 ^ 1'b0 ;
  assign n18759 = ~n12157 & n18758 ;
  assign n18760 = ~n828 & n924 ;
  assign n18761 = n3995 & n18760 ;
  assign n18762 = n12721 & n18761 ;
  assign n18763 = n13821 & ~n18762 ;
  assign n18764 = n18763 ^ n18633 ^ 1'b0 ;
  assign n18765 = n3910 | n17807 ;
  assign n18766 = n18765 ^ n913 ^ 1'b0 ;
  assign n18767 = ~n2029 & n18766 ;
  assign n18768 = n2426 ^ n360 ^ 1'b0 ;
  assign n18769 = ~n734 & n18768 ;
  assign n18770 = n18769 ^ n4813 ^ 1'b0 ;
  assign n18771 = ~n16362 & n18770 ;
  assign n18772 = ~n5844 & n16229 ;
  assign n18773 = n18191 ^ n875 ^ 1'b0 ;
  assign n18774 = n7350 & n18773 ;
  assign n18775 = ~n3390 & n18774 ;
  assign n18776 = ~n4204 & n18775 ;
  assign n18777 = n18776 ^ n17463 ^ 1'b0 ;
  assign n18778 = n3052 & ~n18777 ;
  assign n18779 = n3469 ^ x193 ^ 1'b0 ;
  assign n18780 = ~n540 & n12503 ;
  assign n18781 = n15245 ^ n15032 ^ 1'b0 ;
  assign n18782 = n11187 ^ n6550 ^ 1'b0 ;
  assign n18783 = n18782 ^ n11888 ^ 1'b0 ;
  assign n18784 = n18783 ^ n9761 ^ n3340 ;
  assign n18785 = n9555 & ~n18333 ;
  assign n18786 = n18785 ^ x209 ^ 1'b0 ;
  assign n18787 = n2310 & ~n6558 ;
  assign n18788 = ( ~n4804 & n15286 ) | ( ~n4804 & n16855 ) | ( n15286 & n16855 ) ;
  assign n18789 = n2896 ^ n1346 ^ 1'b0 ;
  assign n18790 = n6740 & n18789 ;
  assign n18791 = n1826 & n18790 ;
  assign n18792 = ~n1826 & n18791 ;
  assign n18793 = n10445 & n12789 ;
  assign n18794 = n18792 & n18793 ;
  assign n18795 = n1847 ^ n493 ^ 1'b0 ;
  assign n18796 = n3678 & ~n12997 ;
  assign n18797 = n13538 & n18796 ;
  assign n18798 = n5838 & n18797 ;
  assign n18799 = ~n18795 & n18798 ;
  assign n18800 = ~n2740 & n7820 ;
  assign n18801 = ~n8677 & n10501 ;
  assign n18802 = n18801 ^ n13101 ^ 1'b0 ;
  assign n18803 = n5047 & ~n10516 ;
  assign n18804 = ~n11281 & n18803 ;
  assign n18805 = n4026 ^ n1395 ^ 1'b0 ;
  assign n18806 = ~n4189 & n18805 ;
  assign n18807 = n5361 ^ n2124 ^ 1'b0 ;
  assign n18808 = n10580 ^ n3263 ^ 1'b0 ;
  assign n18809 = ~n2632 & n18808 ;
  assign n18810 = n8830 & n18809 ;
  assign n18811 = n1302 | n2009 ;
  assign n18812 = n955 & n971 ;
  assign n18813 = n15600 ^ n12760 ^ 1'b0 ;
  assign n18814 = ~n18812 & n18813 ;
  assign n18815 = n10684 | n11348 ;
  assign n18816 = n18815 ^ n13242 ^ 1'b0 ;
  assign n18817 = ~n3365 & n8843 ;
  assign n18818 = n18817 ^ n8560 ^ 1'b0 ;
  assign n18819 = n16326 & n18422 ;
  assign n18820 = n18819 ^ n10833 ^ n10342 ;
  assign n18821 = n2910 & ~n6097 ;
  assign n18822 = n18821 ^ n6243 ^ 1'b0 ;
  assign n18823 = n18820 & ~n18822 ;
  assign n18824 = n4536 & n18823 ;
  assign n18825 = n18824 ^ n7951 ^ 1'b0 ;
  assign n18826 = ~n12039 & n18825 ;
  assign n18827 = n992 | n9420 ;
  assign n18828 = n6780 | n18827 ;
  assign n18829 = ( n12324 & n15511 ) | ( n12324 & ~n18828 ) | ( n15511 & ~n18828 ) ;
  assign n18830 = n11338 & n18829 ;
  assign n18831 = n2636 & ~n4813 ;
  assign n18832 = n11083 ^ n456 ^ 1'b0 ;
  assign n18833 = n964 & n5045 ;
  assign n18834 = ~n7397 & n16967 ;
  assign n18835 = n2425 ^ n2414 ^ 1'b0 ;
  assign n18836 = n12735 ^ n11573 ^ 1'b0 ;
  assign n18837 = ~n10918 & n13475 ;
  assign n18838 = n18837 ^ n9183 ^ 1'b0 ;
  assign n18839 = ~x157 & n14436 ;
  assign n18840 = n18839 ^ n4859 ^ 1'b0 ;
  assign n18841 = n14658 ^ n8064 ^ 1'b0 ;
  assign n18842 = n18841 ^ n14538 ^ n8242 ;
  assign n18843 = ~n774 & n2728 ;
  assign n18844 = ~n2728 & n18843 ;
  assign n18845 = x74 & n18844 ;
  assign n18846 = n6048 ^ n2577 ^ 1'b0 ;
  assign n18847 = n18846 ^ n5730 ^ 1'b0 ;
  assign n18848 = n18845 & n18847 ;
  assign n18853 = n7888 | n9439 ;
  assign n18854 = n15664 & ~n18853 ;
  assign n18855 = n6602 & ~n18854 ;
  assign n18856 = n13302 & n18855 ;
  assign n18849 = n3226 ^ n884 ^ 1'b0 ;
  assign n18850 = n1743 | n4676 ;
  assign n18851 = n8387 & ~n18850 ;
  assign n18852 = n18849 | n18851 ;
  assign n18857 = n18856 ^ n18852 ^ 1'b0 ;
  assign n18858 = n13513 ^ x185 ^ 1'b0 ;
  assign n18859 = n18857 & n18858 ;
  assign n18860 = n15723 ^ n2259 ^ 1'b0 ;
  assign n18861 = n15875 & n18860 ;
  assign n18862 = n5287 & n18861 ;
  assign n18863 = n4970 | n6555 ;
  assign n18864 = n14066 ^ n11632 ^ 1'b0 ;
  assign n18865 = n15965 ^ n13241 ^ 1'b0 ;
  assign n18866 = ~n9539 & n13438 ;
  assign n18867 = n7888 & n18866 ;
  assign n18868 = ~n17475 & n18867 ;
  assign n18869 = ~n2158 & n7777 ;
  assign n18870 = n17665 ^ n12734 ^ 1'b0 ;
  assign n18871 = n4241 & ~n7710 ;
  assign n18872 = n12366 & n18871 ;
  assign n18873 = n18872 ^ n3749 ^ 1'b0 ;
  assign n18874 = n18870 & n18873 ;
  assign n18875 = n3430 ^ n444 ^ 1'b0 ;
  assign n18876 = n3760 & n18875 ;
  assign n18877 = n1732 & ~n2237 ;
  assign n18878 = n1120 & n14166 ;
  assign n18879 = ~n1447 & n1788 ;
  assign n18880 = n11157 ^ x94 ^ 1'b0 ;
  assign n18881 = ~n3973 & n16923 ;
  assign n18882 = n1512 & ~n9736 ;
  assign n18883 = n8896 | n18882 ;
  assign n18884 = x160 & ~n6527 ;
  assign n18885 = ~n10659 & n18884 ;
  assign n18887 = n3426 ^ n290 ^ 1'b0 ;
  assign n18888 = n2503 | n18887 ;
  assign n18886 = n6769 & n13029 ;
  assign n18889 = n18888 ^ n18886 ^ 1'b0 ;
  assign n18890 = n11107 & n18889 ;
  assign n18891 = ~n1694 & n18890 ;
  assign n18892 = n8921 ^ n5031 ^ 1'b0 ;
  assign n18893 = n700 | n16584 ;
  assign n18894 = n4219 ^ x67 ^ 1'b0 ;
  assign n18895 = n744 & n18894 ;
  assign n18896 = n18895 ^ n1775 ^ 1'b0 ;
  assign n18897 = n1521 & ~n18896 ;
  assign n18898 = ~n14866 & n18897 ;
  assign n18899 = n6744 ^ n3593 ^ 1'b0 ;
  assign n18900 = n12671 ^ n3996 ^ 1'b0 ;
  assign n18901 = n18900 ^ n18333 ^ 1'b0 ;
  assign n18902 = n337 & n13776 ;
  assign n18903 = n1988 & n18902 ;
  assign n18904 = n3819 & ~n18903 ;
  assign n18905 = n4204 ^ n1815 ^ 1'b0 ;
  assign n18906 = n18905 ^ n519 ^ 1'b0 ;
  assign n18907 = n14602 ^ n7208 ^ n6681 ;
  assign n18908 = n18906 & ~n18907 ;
  assign n18909 = n7039 ^ n5433 ^ 1'b0 ;
  assign n18910 = n9376 & ~n18909 ;
  assign n18911 = n18910 ^ n926 ^ 1'b0 ;
  assign n18912 = n2046 & ~n7695 ;
  assign n18913 = n14279 ^ n639 ^ 1'b0 ;
  assign n18914 = n17501 ^ n7657 ^ 1'b0 ;
  assign n18915 = n12682 ^ n4940 ^ 1'b0 ;
  assign n18916 = ~n12022 & n18915 ;
  assign n18917 = n322 & n15705 ;
  assign n18918 = n18916 & ~n18917 ;
  assign n18919 = n7716 & n18918 ;
  assign n18920 = n2241 & ~n3314 ;
  assign n18921 = n18920 ^ n16815 ^ 1'b0 ;
  assign n18922 = ~n2486 & n18921 ;
  assign n18923 = n9454 ^ n492 ^ 1'b0 ;
  assign n18924 = n8710 & n18923 ;
  assign n18925 = ~n10102 & n17560 ;
  assign n18926 = n781 | n18136 ;
  assign n18927 = n8698 ^ n3431 ^ 1'b0 ;
  assign n18928 = n6255 | n18927 ;
  assign n18929 = x221 & ~n1117 ;
  assign n18930 = n18928 & n18929 ;
  assign n18931 = n4587 | n14477 ;
  assign n18932 = ~n17711 & n18931 ;
  assign n18933 = n13220 ^ n3943 ^ 1'b0 ;
  assign n18936 = n2356 ^ n1510 ^ 1'b0 ;
  assign n18937 = n3366 & ~n18936 ;
  assign n18938 = ~n10744 & n18937 ;
  assign n18939 = ~n11192 & n18938 ;
  assign n18934 = n1321 & ~n4493 ;
  assign n18935 = n18934 ^ n7174 ^ 1'b0 ;
  assign n18940 = n18939 ^ n18935 ^ n6146 ;
  assign n18941 = n3678 ^ n445 ^ 1'b0 ;
  assign n18942 = n9994 & ~n18941 ;
  assign n18943 = n4464 ^ n3960 ^ 1'b0 ;
  assign n18944 = n6000 & n18943 ;
  assign n18945 = n3095 & ~n14470 ;
  assign n18946 = n15445 & ~n18945 ;
  assign n18947 = ~n18944 & n18946 ;
  assign n18948 = n1936 | n14632 ;
  assign n18949 = x39 | n18948 ;
  assign n18950 = n8628 ^ n6741 ^ 1'b0 ;
  assign n18951 = n15335 | n18950 ;
  assign n18952 = n5256 & n15309 ;
  assign n18953 = n8052 | n18952 ;
  assign n18954 = n577 & ~n5207 ;
  assign n18955 = n6525 & ~n18954 ;
  assign n18956 = n18955 ^ n3158 ^ 1'b0 ;
  assign n18957 = n10423 & n14695 ;
  assign n18958 = n18956 & n18957 ;
  assign n18959 = ~n10917 & n17266 ;
  assign n18960 = n1356 & n18959 ;
  assign n18961 = n18960 ^ n12230 ^ 1'b0 ;
  assign n18962 = n17587 ^ n5703 ^ 1'b0 ;
  assign n18963 = n9832 ^ n411 ^ 1'b0 ;
  assign n18964 = n4889 & ~n18963 ;
  assign n18965 = n9895 & n18964 ;
  assign n18966 = n18965 ^ n5507 ^ 1'b0 ;
  assign n18967 = n13195 | n18966 ;
  assign n18968 = n18967 ^ n12919 ^ 1'b0 ;
  assign n18969 = n18962 | n18968 ;
  assign n18970 = n2804 | n18969 ;
  assign n18971 = n18970 ^ x240 ^ 1'b0 ;
  assign n18972 = n12920 ^ n1310 ^ 1'b0 ;
  assign n18973 = n18972 ^ n4622 ^ 1'b0 ;
  assign n18974 = n1837 | n18973 ;
  assign n18975 = n2078 | n18974 ;
  assign n18976 = n18975 ^ n9269 ^ 1'b0 ;
  assign n18977 = n2404 & n3999 ;
  assign n18978 = n8373 & n12232 ;
  assign n18979 = n725 | n8326 ;
  assign n18980 = n18172 ^ n7039 ^ 1'b0 ;
  assign n18981 = ~n18979 & n18980 ;
  assign n18982 = n17788 ^ n1089 ^ 1'b0 ;
  assign n18983 = n8821 & n18982 ;
  assign n18984 = n1221 & n4882 ;
  assign n18985 = n8424 | n10024 ;
  assign n18986 = n18984 & ~n18985 ;
  assign n18987 = n3324 | n18986 ;
  assign n18988 = n13307 | n18987 ;
  assign n18989 = ~n8412 & n10353 ;
  assign n18990 = n3671 & n18989 ;
  assign n18991 = n1116 | n18990 ;
  assign n18992 = n14252 | n18991 ;
  assign n18993 = n2691 | n3951 ;
  assign n18994 = n18993 ^ n2149 ^ 1'b0 ;
  assign n18995 = n18992 | n18994 ;
  assign n18997 = n7049 | n8908 ;
  assign n18998 = n18997 ^ n13598 ^ 1'b0 ;
  assign n18996 = n5154 & n15937 ;
  assign n18999 = n18998 ^ n18996 ^ 1'b0 ;
  assign n19000 = n4868 ^ n4497 ^ 1'b0 ;
  assign n19001 = n3328 & ~n14686 ;
  assign n19002 = ~n15960 & n16974 ;
  assign n19003 = n19001 & n19002 ;
  assign n19004 = n8572 ^ n8348 ^ 1'b0 ;
  assign n19005 = ~n1443 & n19004 ;
  assign n19006 = n5575 & n19005 ;
  assign n19007 = n4416 ^ n3915 ^ x3 ;
  assign n19008 = n19007 ^ n3403 ^ 1'b0 ;
  assign n19009 = n5242 & ~n19008 ;
  assign n19010 = n1616 & ~n11207 ;
  assign n19011 = n19010 ^ n11611 ^ 1'b0 ;
  assign n19012 = ~n9152 & n19011 ;
  assign n19013 = n11895 ^ n2074 ^ 1'b0 ;
  assign n19014 = n5686 & ~n19013 ;
  assign n19015 = n9930 & n19014 ;
  assign n19016 = ~n14058 & n14135 ;
  assign n19017 = n13932 ^ n1280 ^ n327 ;
  assign n19018 = n19017 ^ n15425 ^ n14311 ;
  assign n19022 = n11662 ^ n2846 ^ n832 ;
  assign n19019 = n967 & n6854 ;
  assign n19020 = n19019 ^ n7296 ^ 1'b0 ;
  assign n19021 = n5714 & ~n19020 ;
  assign n19023 = n19022 ^ n19021 ^ 1'b0 ;
  assign n19024 = n2277 & n19023 ;
  assign n19025 = n3872 & n8139 ;
  assign n19026 = n1523 & ~n18622 ;
  assign n19027 = ~n7448 & n16340 ;
  assign n19028 = ~n2523 & n19027 ;
  assign n19029 = n19028 ^ n9786 ^ 1'b0 ;
  assign n19030 = n3632 | n19029 ;
  assign n19031 = n18690 ^ x144 ^ 1'b0 ;
  assign n19032 = ~n10349 & n19031 ;
  assign n19033 = ~n1606 & n13661 ;
  assign n19034 = ~n3953 & n17072 ;
  assign n19035 = n19034 ^ x100 ^ 1'b0 ;
  assign n19036 = n7349 ^ n3269 ^ 1'b0 ;
  assign n19037 = n9260 & n19036 ;
  assign n19038 = n19037 ^ n6637 ^ 1'b0 ;
  assign n19040 = n6423 | n6822 ;
  assign n19039 = ~n4318 & n11191 ;
  assign n19041 = n19040 ^ n19039 ^ 1'b0 ;
  assign n19042 = ~n3825 & n10408 ;
  assign n19043 = n19042 ^ n7520 ^ 1'b0 ;
  assign n19044 = n18433 ^ n9454 ^ 1'b0 ;
  assign n19045 = n1358 & n7395 ;
  assign n19046 = ~n3295 & n19045 ;
  assign n19047 = n7634 | n19046 ;
  assign n19048 = n12616 | n19047 ;
  assign n19049 = n8806 ^ n5450 ^ n456 ;
  assign n19050 = ( n930 & ~n7720 ) | ( n930 & n10729 ) | ( ~n7720 & n10729 ) ;
  assign n19051 = n19050 ^ n9043 ^ 1'b0 ;
  assign n19052 = n19049 & ~n19051 ;
  assign n19053 = n19052 ^ n16860 ^ 1'b0 ;
  assign n19054 = n11653 ^ n1988 ^ n825 ;
  assign n19055 = n14060 & ~n19054 ;
  assign n19056 = n5850 & n7539 ;
  assign n19057 = ( n2441 & ~n2806 ) | ( n2441 & n13315 ) | ( ~n2806 & n13315 ) ;
  assign n19058 = n4888 ^ n1336 ^ 1'b0 ;
  assign n19059 = n11323 ^ n1912 ^ 1'b0 ;
  assign n19060 = n8919 & n19059 ;
  assign n19061 = n10056 ^ n6401 ^ 1'b0 ;
  assign n19062 = n12878 & ~n18105 ;
  assign n19063 = n6574 ^ n4302 ^ n3908 ;
  assign n19064 = n8160 ^ n2006 ^ 1'b0 ;
  assign n19065 = ~n2776 & n19064 ;
  assign n19066 = n19065 ^ n3983 ^ 1'b0 ;
  assign n19067 = n12071 & n19066 ;
  assign n19068 = ~n3043 & n4291 ;
  assign n19069 = n19068 ^ n2511 ^ 1'b0 ;
  assign n19070 = n8565 | n19069 ;
  assign n19071 = n13675 | n18608 ;
  assign n19072 = n19070 & ~n19071 ;
  assign n19073 = n10505 & ~n15511 ;
  assign n19074 = n19073 ^ n17395 ^ n13833 ;
  assign n19078 = n11543 ^ n9174 ^ 1'b0 ;
  assign n19075 = n7291 ^ n979 ^ 1'b0 ;
  assign n19076 = n8837 ^ n7934 ^ 1'b0 ;
  assign n19077 = n19075 & ~n19076 ;
  assign n19079 = n19078 ^ n19077 ^ 1'b0 ;
  assign n19080 = ~n12616 & n13269 ;
  assign n19081 = n19080 ^ n3518 ^ 1'b0 ;
  assign n19082 = n1930 & ~n15959 ;
  assign n19083 = n9576 & ~n16372 ;
  assign n19084 = ~n2408 & n8294 ;
  assign n19085 = n385 & ~n6517 ;
  assign n19086 = n5050 ^ n2962 ^ 1'b0 ;
  assign n19087 = n19086 ^ n6200 ^ 1'b0 ;
  assign n19088 = n19085 & n19087 ;
  assign n19089 = n19088 ^ n6845 ^ 1'b0 ;
  assign n19090 = n7343 | n19089 ;
  assign n19091 = ( ~n8354 & n19084 ) | ( ~n8354 & n19090 ) | ( n19084 & n19090 ) ;
  assign n19092 = n1784 | n19091 ;
  assign n19093 = ~n1181 & n1773 ;
  assign n19094 = n5223 & n19093 ;
  assign n19095 = n19094 ^ n2392 ^ 1'b0 ;
  assign n19096 = n18327 ^ n10671 ^ 1'b0 ;
  assign n19097 = n6207 & n19096 ;
  assign n19098 = x12 & ~n4940 ;
  assign n19099 = ~n6192 & n19098 ;
  assign n19100 = n4222 ^ n1402 ^ 1'b0 ;
  assign n19101 = ( n1018 & n2319 ) | ( n1018 & ~n19100 ) | ( n2319 & ~n19100 ) ;
  assign n19102 = n14302 ^ n9002 ^ 1'b0 ;
  assign n19103 = ~n1337 & n17770 ;
  assign n19104 = n19103 ^ n18890 ^ 1'b0 ;
  assign n19105 = n19001 ^ n3440 ^ 1'b0 ;
  assign n19106 = n12803 & n19105 ;
  assign n19107 = n8849 ^ x241 ^ 1'b0 ;
  assign n19108 = ~n3187 & n6225 ;
  assign n19109 = n4294 & n19108 ;
  assign n19110 = ~n8374 & n14456 ;
  assign n19111 = n19110 ^ n901 ^ 1'b0 ;
  assign n19112 = n19109 | n19111 ;
  assign n19113 = ~n10774 & n15900 ;
  assign n19114 = n9276 ^ n6950 ^ 1'b0 ;
  assign n19115 = n7994 & ~n19114 ;
  assign n19116 = n19115 ^ n17470 ^ 1'b0 ;
  assign n19117 = n19113 & n19116 ;
  assign n19118 = n10715 ^ n3465 ^ 1'b0 ;
  assign n19119 = n12579 & ~n19118 ;
  assign n19120 = n14159 & n14773 ;
  assign n19121 = n19120 ^ n3643 ^ 1'b0 ;
  assign n19124 = n10042 ^ n4810 ^ 1'b0 ;
  assign n19125 = n19124 ^ n10325 ^ 1'b0 ;
  assign n19122 = n3329 & ~n5982 ;
  assign n19123 = n6360 & n19122 ;
  assign n19126 = n19125 ^ n19123 ^ 1'b0 ;
  assign n19127 = n4655 | n4749 ;
  assign n19128 = n12223 ^ n7353 ^ 1'b0 ;
  assign n19129 = n19128 ^ n12072 ^ 1'b0 ;
  assign n19130 = ~n5928 & n19129 ;
  assign n19131 = n19127 | n19130 ;
  assign n19132 = n2866 ^ n2107 ^ 1'b0 ;
  assign n19133 = n10590 | n19132 ;
  assign n19134 = n1914 & ~n11899 ;
  assign n19135 = n19133 & n19134 ;
  assign n19136 = n4350 & ~n10348 ;
  assign n19137 = n11519 & n19136 ;
  assign n19138 = n1405 & n19137 ;
  assign n19139 = ~n13339 & n19138 ;
  assign n19140 = n19135 & n19139 ;
  assign n19141 = n5012 ^ n4101 ^ 1'b0 ;
  assign n19142 = n19141 ^ n15180 ^ 1'b0 ;
  assign n19143 = ~x65 & n14211 ;
  assign n19144 = n5718 & n6053 ;
  assign n19145 = n1159 | n9730 ;
  assign n19146 = n7527 & ~n8123 ;
  assign n19147 = ~n1521 & n4354 ;
  assign n19148 = ~n4354 & n19147 ;
  assign n19149 = n3451 | n19148 ;
  assign n19150 = n3451 & ~n19149 ;
  assign n19151 = n951 | n1571 ;
  assign n19152 = n951 & ~n19151 ;
  assign n19153 = n19152 ^ n2001 ^ 1'b0 ;
  assign n19154 = n19150 | n19153 ;
  assign n19155 = n4244 & ~n10521 ;
  assign n19156 = ~n4244 & n19155 ;
  assign n19157 = n18464 ^ n8954 ^ 1'b0 ;
  assign n19158 = n19156 | n19157 ;
  assign n19159 = n7228 | n16561 ;
  assign n19160 = n16561 & ~n19159 ;
  assign n19161 = n672 | n2106 ;
  assign n19162 = n2106 & ~n19161 ;
  assign n19163 = n10936 & ~n19162 ;
  assign n19164 = ~n10936 & n19163 ;
  assign n19165 = n11416 | n17814 ;
  assign n19166 = n19164 | n19165 ;
  assign n19167 = n19160 & ~n19166 ;
  assign n19168 = n19158 | n19167 ;
  assign n19169 = n19154 & ~n19168 ;
  assign n19170 = n10637 ^ n1605 ^ 1'b0 ;
  assign n19171 = n11295 & n17579 ;
  assign n19172 = ~n17721 & n19171 ;
  assign n19173 = ~x84 & n10965 ;
  assign n19174 = n19173 ^ n5692 ^ 1'b0 ;
  assign n19175 = n3325 & ~n8969 ;
  assign n19176 = n2725 & ~n19175 ;
  assign n19177 = ~n9353 & n19176 ;
  assign n19178 = n3922 & ~n5148 ;
  assign n19179 = n2037 & n19178 ;
  assign n19180 = n1693 | n19179 ;
  assign n19181 = n4521 & n19180 ;
  assign n19182 = n18725 ^ n16421 ^ 1'b0 ;
  assign n19183 = n19181 & n19182 ;
  assign n19184 = ~n2274 & n16861 ;
  assign n19185 = n13370 ^ n3186 ^ 1'b0 ;
  assign n19186 = ~n10744 & n19185 ;
  assign n19193 = ~n1159 & n11862 ;
  assign n19194 = n4122 & n19193 ;
  assign n19195 = n19194 ^ n6662 ^ 1'b0 ;
  assign n19188 = n5382 ^ n3275 ^ 1'b0 ;
  assign n19189 = x215 & ~n19188 ;
  assign n19190 = n4455 ^ n320 ^ 1'b0 ;
  assign n19191 = n19189 & n19190 ;
  assign n19187 = n17591 ^ n7256 ^ 1'b0 ;
  assign n19192 = n19191 ^ n19187 ^ 1'b0 ;
  assign n19196 = n19195 ^ n19192 ^ 1'b0 ;
  assign n19197 = n1269 & n3692 ;
  assign n19198 = n5573 & n6854 ;
  assign n19199 = n13473 ^ n532 ^ 1'b0 ;
  assign n19200 = ~n4314 & n5059 ;
  assign n19201 = n2254 & n19200 ;
  assign n19202 = n12241 & ~n19201 ;
  assign n19203 = n19202 ^ n3468 ^ 1'b0 ;
  assign n19204 = n12775 & ~n19203 ;
  assign n19205 = ~n7864 & n16879 ;
  assign n19206 = n8427 | n10555 ;
  assign n19207 = n19206 ^ n1883 ^ 1'b0 ;
  assign n19208 = n19207 ^ n1070 ^ 1'b0 ;
  assign n19209 = n3124 ^ n2841 ^ 1'b0 ;
  assign n19210 = n14871 & ~n18615 ;
  assign n19211 = ~n19209 & n19210 ;
  assign n19212 = n3501 | n12711 ;
  assign n19213 = n19212 ^ n10081 ^ 1'b0 ;
  assign n19214 = n14397 ^ n12770 ^ 1'b0 ;
  assign n19215 = n8890 & n12141 ;
  assign n19216 = n19215 ^ n14643 ^ n12141 ;
  assign n19217 = ( ~n4932 & n19214 ) | ( ~n4932 & n19216 ) | ( n19214 & n19216 ) ;
  assign n19218 = n7569 & ~n7727 ;
  assign n19219 = n6108 & n11829 ;
  assign n19220 = ~n19218 & n19219 ;
  assign n19221 = n5618 & n7788 ;
  assign n19222 = ~n12268 & n19221 ;
  assign n19223 = n11868 & ~n13317 ;
  assign n19224 = n19223 ^ n18481 ^ 1'b0 ;
  assign n19225 = n2496 & ~n6389 ;
  assign n19226 = n4880 & n19225 ;
  assign n19227 = ~n5540 & n19226 ;
  assign n19228 = n3266 | n19227 ;
  assign n19229 = n19228 ^ n5779 ^ 1'b0 ;
  assign n19230 = n8738 ^ n7342 ^ 1'b0 ;
  assign n19231 = n18418 ^ n18117 ^ 1'b0 ;
  assign n19232 = n11884 ^ n3577 ^ 1'b0 ;
  assign n19233 = n11522 ^ n10265 ^ 1'b0 ;
  assign n19234 = n12787 ^ n7009 ^ n978 ;
  assign n19235 = n536 & ~n12270 ;
  assign n19236 = n7070 | n10348 ;
  assign n19237 = n13732 ^ n6644 ^ 1'b0 ;
  assign n19238 = n4564 & ~n19237 ;
  assign n19239 = n1809 & ~n1843 ;
  assign n19240 = x154 | n6061 ;
  assign n19241 = n19240 ^ n9304 ^ 1'b0 ;
  assign n19242 = n1803 & n19241 ;
  assign n19243 = n19242 ^ n1207 ^ 1'b0 ;
  assign n19244 = n5462 ^ n3477 ^ 1'b0 ;
  assign n19245 = n19243 & n19244 ;
  assign n19246 = n4573 | n11611 ;
  assign n19247 = n2116 & ~n19246 ;
  assign n19248 = n19247 ^ n8913 ^ 1'b0 ;
  assign n19249 = n5159 & n19248 ;
  assign n19250 = n6446 ^ x232 ^ 1'b0 ;
  assign n19251 = n4393 | n13317 ;
  assign n19252 = n5384 & ~n19251 ;
  assign n19253 = ( n956 & ~n2185 ) | ( n956 & n19252 ) | ( ~n2185 & n19252 ) ;
  assign n19254 = ~n3630 & n8465 ;
  assign n19255 = n19254 ^ n2223 ^ 1'b0 ;
  assign n19261 = n5507 & ~n6745 ;
  assign n19256 = ~n3224 & n6889 ;
  assign n19257 = n19256 ^ n1710 ^ 1'b0 ;
  assign n19258 = n12734 ^ n8584 ^ 1'b0 ;
  assign n19259 = ~n19257 & n19258 ;
  assign n19260 = n18571 & n19259 ;
  assign n19262 = n19261 ^ n19260 ^ 1'b0 ;
  assign n19263 = ~x70 & n1277 ;
  assign n19264 = n19263 ^ n12767 ^ 1'b0 ;
  assign n19265 = ~n8345 & n18760 ;
  assign n19266 = n4655 & ~n19265 ;
  assign n19267 = ~n7148 & n11304 ;
  assign n19268 = n19267 ^ n5654 ^ 1'b0 ;
  assign n19269 = ~n5613 & n9440 ;
  assign n19270 = ( n3175 & ~n15995 ) | ( n3175 & n19269 ) | ( ~n15995 & n19269 ) ;
  assign n19271 = ~n2842 & n13778 ;
  assign n19272 = n19271 ^ n5670 ^ 1'b0 ;
  assign n19273 = n15532 & ~n19272 ;
  assign n19274 = n19273 ^ n5427 ^ 1'b0 ;
  assign n19275 = n8336 & ~n19274 ;
  assign n19276 = n4460 & n7622 ;
  assign n19278 = n10422 ^ n3647 ^ n1826 ;
  assign n19277 = ~n1865 & n7312 ;
  assign n19279 = n19278 ^ n19277 ^ 1'b0 ;
  assign n19280 = n19276 & n19279 ;
  assign n19281 = n19280 ^ n3071 ^ 1'b0 ;
  assign n19282 = n9726 ^ x177 ^ 1'b0 ;
  assign n19283 = n7820 & n19282 ;
  assign n19284 = n19283 ^ n4874 ^ 1'b0 ;
  assign n19285 = n3158 | n19284 ;
  assign n19286 = n7720 & n16429 ;
  assign n19287 = n17203 ^ x176 ^ 1'b0 ;
  assign n19288 = n3637 ^ n1611 ^ 1'b0 ;
  assign n19289 = n4863 ^ n387 ^ 1'b0 ;
  assign n19290 = ~n3458 & n19289 ;
  assign n19291 = n1404 | n19290 ;
  assign n19292 = n7317 & n7459 ;
  assign n19293 = n9387 & n19292 ;
  assign n19294 = n11857 ^ n1533 ^ 1'b0 ;
  assign n19295 = n1731 & ~n19294 ;
  assign n19296 = n19295 ^ n6961 ^ n3891 ;
  assign n19297 = n19296 ^ n1524 ^ 1'b0 ;
  assign n19298 = ( ~n2135 & n2660 ) | ( ~n2135 & n19297 ) | ( n2660 & n19297 ) ;
  assign n19299 = n6939 & n19298 ;
  assign n19303 = n7105 ^ n6999 ^ 1'b0 ;
  assign n19300 = n2269 & ~n6015 ;
  assign n19301 = n19300 ^ n7314 ^ 1'b0 ;
  assign n19302 = n3796 & n19301 ;
  assign n19304 = n19303 ^ n19302 ^ n2392 ;
  assign n19305 = n10081 ^ n2737 ^ 1'b0 ;
  assign n19306 = n809 ^ n648 ^ 1'b0 ;
  assign n19307 = n3791 ^ n2406 ^ 1'b0 ;
  assign n19308 = ~n3086 & n9910 ;
  assign n19309 = n2072 & n19308 ;
  assign n19310 = n19309 ^ n924 ^ 1'b0 ;
  assign n19311 = n395 & n19310 ;
  assign n19312 = n19311 ^ n320 ^ 1'b0 ;
  assign n19313 = n3610 & ~n15614 ;
  assign n19314 = n19313 ^ n683 ^ 1'b0 ;
  assign n19315 = n7769 & ~n19314 ;
  assign n19317 = n3325 & n14652 ;
  assign n19316 = n1684 & n5861 ;
  assign n19318 = n19317 ^ n19316 ^ 1'b0 ;
  assign n19319 = n16067 & ~n19318 ;
  assign n19320 = x17 & ~n593 ;
  assign n19321 = n19320 ^ n1836 ^ 1'b0 ;
  assign n19322 = n5360 & n11584 ;
  assign n19323 = ~n2642 & n11050 ;
  assign n19324 = n1658 & n19323 ;
  assign n19325 = n19324 ^ x113 ^ 1'b0 ;
  assign n19326 = n16692 & ~n19325 ;
  assign n19327 = n19326 ^ n18392 ^ 1'b0 ;
  assign n19328 = n1172 | n13507 ;
  assign n19331 = n7036 ^ n4501 ^ 1'b0 ;
  assign n19332 = n8254 | n19331 ;
  assign n19333 = n13771 | n19332 ;
  assign n19334 = n8570 | n19333 ;
  assign n19329 = n13968 ^ x2 ^ 1'b0 ;
  assign n19330 = n14007 | n19329 ;
  assign n19335 = n19334 ^ n19330 ^ 1'b0 ;
  assign n19336 = ~n1745 & n1899 ;
  assign n19337 = n11517 & n19336 ;
  assign n19338 = n18084 & n19337 ;
  assign n19339 = ~n9380 & n17247 ;
  assign n19340 = n12745 & n19339 ;
  assign n19341 = n19340 ^ n16026 ^ 1'b0 ;
  assign n19342 = n5148 & n14463 ;
  assign n19343 = n19342 ^ n788 ^ 1'b0 ;
  assign n19344 = n5994 & ~n19343 ;
  assign n19348 = x226 & ~n6297 ;
  assign n19349 = n19348 ^ n579 ^ 1'b0 ;
  assign n19345 = ~n4930 & n8642 ;
  assign n19346 = n19345 ^ n1883 ^ 1'b0 ;
  assign n19347 = n4485 | n19346 ;
  assign n19350 = n19349 ^ n19347 ^ 1'b0 ;
  assign n19351 = n19350 ^ n5535 ^ x226 ;
  assign n19352 = n3669 & ~n3973 ;
  assign n19353 = ~n1298 & n19352 ;
  assign n19354 = ~n5097 & n19353 ;
  assign n19355 = n13230 & ~n19354 ;
  assign n19356 = n19355 ^ n6030 ^ 1'b0 ;
  assign n19357 = ~n8637 & n15874 ;
  assign n19358 = n19357 ^ n17244 ^ 1'b0 ;
  assign n19359 = n7737 ^ n4294 ^ 1'b0 ;
  assign n19360 = n18141 | n19359 ;
  assign n19361 = n1985 & n7345 ;
  assign n19362 = n19361 ^ n12594 ^ 1'b0 ;
  assign n19363 = ~n7593 & n17566 ;
  assign n19364 = n2542 | n19363 ;
  assign n19365 = n1899 ^ n833 ^ 1'b0 ;
  assign n19366 = n19364 & ~n19365 ;
  assign n19367 = n19366 ^ n2179 ^ 1'b0 ;
  assign n19368 = n11234 & ~n19367 ;
  assign n19369 = n8692 ^ n6741 ^ 1'b0 ;
  assign n19370 = n5723 & ~n19369 ;
  assign n19371 = ~n4186 & n6555 ;
  assign n19372 = ~n2740 & n19371 ;
  assign n19373 = n1727 | n4112 ;
  assign n19374 = n19373 ^ n415 ^ 1'b0 ;
  assign n19375 = n7679 & ~n10030 ;
  assign n19376 = ~n7679 & n19375 ;
  assign n19377 = ~n733 & n2443 ;
  assign n19378 = n733 & n19377 ;
  assign n19379 = ~n9406 & n19378 ;
  assign n19380 = ~n3902 & n19379 ;
  assign n19381 = n19380 ^ n9436 ^ 1'b0 ;
  assign n19382 = n19376 | n19381 ;
  assign n19383 = ~n8281 & n19382 ;
  assign n19384 = n12758 | n14770 ;
  assign n19385 = n9905 | n19384 ;
  assign n19386 = ~n1690 & n13225 ;
  assign n19387 = n19386 ^ n8840 ^ 1'b0 ;
  assign n19388 = ~n9959 & n19387 ;
  assign n19389 = ~n967 & n6071 ;
  assign n19390 = n8039 & n19389 ;
  assign n19391 = ~n19388 & n19390 ;
  assign n19392 = n18609 ^ n13651 ^ 1'b0 ;
  assign n19393 = n4395 ^ n2314 ^ 1'b0 ;
  assign n19394 = n8795 & n19393 ;
  assign n19395 = n4903 & n6651 ;
  assign n19396 = n7756 ^ n2074 ^ 1'b0 ;
  assign n19397 = n2906 | n10018 ;
  assign n19398 = n14277 | n19397 ;
  assign n19399 = n2420 | n9654 ;
  assign n19400 = n8740 | n19399 ;
  assign n19401 = n1175 | n1799 ;
  assign n19402 = n1175 & ~n19401 ;
  assign n19403 = n3741 & ~n19402 ;
  assign n19404 = ~n3741 & n19403 ;
  assign n19405 = n4099 | n13876 ;
  assign n19406 = n19404 | n19405 ;
  assign n19407 = n19406 ^ n19175 ^ 1'b0 ;
  assign n19408 = n7407 ^ n2186 ^ 1'b0 ;
  assign n19409 = n11891 & ~n19408 ;
  assign n19410 = x127 & n18519 ;
  assign n19411 = n9580 ^ n8624 ^ 1'b0 ;
  assign n19412 = n1451 | n19411 ;
  assign n19413 = n4331 & n7667 ;
  assign n19414 = ~n15627 & n19413 ;
  assign n19415 = ~n2629 & n9869 ;
  assign n19416 = n7685 & n19415 ;
  assign n19417 = n6499 ^ n2947 ^ 1'b0 ;
  assign n19418 = n13099 & ~n19417 ;
  assign n19419 = n19418 ^ n8617 ^ n5808 ;
  assign n19420 = n10875 ^ n7638 ^ 1'b0 ;
  assign n19421 = n387 & n6540 ;
  assign n19422 = n838 & n19421 ;
  assign n19423 = n8352 & ~n17412 ;
  assign n19424 = n1829 & ~n15999 ;
  assign n19425 = n19424 ^ n5448 ^ 1'b0 ;
  assign n19426 = ~n618 & n1370 ;
  assign n19427 = ~n575 & n19426 ;
  assign n19431 = ~n2191 & n6355 ;
  assign n19432 = n19431 ^ n4109 ^ 1'b0 ;
  assign n19429 = n6780 | n9380 ;
  assign n19430 = ~n18457 & n19429 ;
  assign n19433 = n19432 ^ n19430 ^ 1'b0 ;
  assign n19428 = n8517 & ~n15354 ;
  assign n19434 = n19433 ^ n19428 ^ 1'b0 ;
  assign n19435 = ~n7822 & n12338 ;
  assign n19436 = n3499 ^ n1638 ^ 1'b0 ;
  assign n19437 = n9006 ^ n6935 ^ 1'b0 ;
  assign n19438 = n19437 ^ n8992 ^ 1'b0 ;
  assign n19439 = n4803 ^ n1824 ^ 1'b0 ;
  assign n19440 = n3249 & n5454 ;
  assign n19441 = n6138 ^ n2411 ^ 1'b0 ;
  assign n19442 = ~n19440 & n19441 ;
  assign n19443 = ~n1571 & n19442 ;
  assign n19444 = n19443 ^ n3331 ^ 1'b0 ;
  assign n19445 = n19439 & ~n19444 ;
  assign n19446 = n5696 ^ n1928 ^ n1704 ;
  assign n19447 = n19446 ^ n832 ^ 1'b0 ;
  assign n19448 = ~n2099 & n19447 ;
  assign n19449 = ~n2389 & n19448 ;
  assign n19450 = n19449 ^ n6179 ^ 1'b0 ;
  assign n19451 = n18492 ^ n11751 ^ 1'b0 ;
  assign n19452 = n5622 & ~n19451 ;
  assign n19453 = n6496 ^ n3237 ^ 1'b0 ;
  assign n19454 = ~n1399 & n19453 ;
  assign n19455 = ~n5094 & n19454 ;
  assign n19456 = n5859 ^ n1656 ^ 1'b0 ;
  assign n19457 = n19455 | n19456 ;
  assign n19458 = n6644 & ~n8384 ;
  assign n19459 = n19458 ^ n19033 ^ n14658 ;
  assign n19460 = n2543 & ~n10686 ;
  assign n19461 = n1111 & n2089 ;
  assign n19464 = n2953 & n12334 ;
  assign n19462 = n10849 ^ x219 ^ 1'b0 ;
  assign n19463 = ~n8428 & n19462 ;
  assign n19465 = n19464 ^ n19463 ^ 1'b0 ;
  assign n19466 = n14431 | n19465 ;
  assign n19467 = n19461 | n19466 ;
  assign n19468 = n19467 ^ n13819 ^ 1'b0 ;
  assign n19469 = ~n3329 & n8173 ;
  assign n19470 = n11433 ^ n2310 ^ 1'b0 ;
  assign n19471 = n19470 ^ n19302 ^ 1'b0 ;
  assign n19472 = n19469 & n19471 ;
  assign n19473 = n1673 | n10334 ;
  assign n19474 = n6151 | n19473 ;
  assign n19475 = ( n522 & ~n5597 ) | ( n522 & n19474 ) | ( ~n5597 & n19474 ) ;
  assign n19476 = n685 & ~n2099 ;
  assign n19477 = n19476 ^ n12206 ^ 1'b0 ;
  assign n19478 = n6302 & ~n19477 ;
  assign n19479 = n1293 & ~n3159 ;
  assign n19480 = n17887 ^ n7179 ^ 1'b0 ;
  assign n19481 = n19479 & ~n19480 ;
  assign n19482 = n5931 & ~n17311 ;
  assign n19483 = n9135 & n19482 ;
  assign n19484 = n3514 | n11282 ;
  assign n19485 = n19484 ^ n15289 ^ 1'b0 ;
  assign n19486 = n13252 & n19485 ;
  assign n19487 = n8796 ^ n269 ^ 1'b0 ;
  assign n19488 = x52 & n19487 ;
  assign n19489 = n9341 ^ n1106 ^ 1'b0 ;
  assign n19490 = ~n3973 & n19489 ;
  assign n19491 = ~n9781 & n19490 ;
  assign n19492 = ~n19490 & n19491 ;
  assign n19493 = n16640 ^ n14354 ^ 1'b0 ;
  assign n19494 = n3784 | n19493 ;
  assign n19497 = n3542 | n4032 ;
  assign n19498 = n19497 ^ n8010 ^ 1'b0 ;
  assign n19499 = n6590 & n19498 ;
  assign n19500 = ~n663 & n19499 ;
  assign n19495 = n13418 | n17085 ;
  assign n19496 = n5996 & ~n19495 ;
  assign n19501 = n19500 ^ n19496 ^ 1'b0 ;
  assign n19502 = n461 & ~n4685 ;
  assign n19503 = n3100 ^ n259 ^ 1'b0 ;
  assign n19504 = ~n13055 & n19503 ;
  assign n19505 = n1710 | n6333 ;
  assign n19506 = n2990 & ~n19505 ;
  assign n19507 = n5627 ^ n1102 ^ 1'b0 ;
  assign n19508 = n14841 ^ n2423 ^ 1'b0 ;
  assign n19509 = n19508 ^ n7247 ^ 1'b0 ;
  assign n19510 = n6498 ^ n4433 ^ 1'b0 ;
  assign n19511 = n1419 | n19510 ;
  assign n19512 = n18284 & ~n19511 ;
  assign n19513 = ~n18141 & n19512 ;
  assign n19515 = ~n4418 & n5398 ;
  assign n19514 = n968 & ~n14608 ;
  assign n19516 = n19515 ^ n19514 ^ 1'b0 ;
  assign n19517 = x130 & n3533 ;
  assign n19518 = n16132 & n19517 ;
  assign n19519 = n19518 ^ n6178 ^ 1'b0 ;
  assign n19520 = n4059 | n5670 ;
  assign n19521 = n6879 ^ n720 ^ 1'b0 ;
  assign n19522 = n14171 ^ n4281 ^ 1'b0 ;
  assign n19523 = n18415 ^ x173 ^ 1'b0 ;
  assign n19524 = n19523 ^ n2870 ^ 1'b0 ;
  assign n19525 = n6250 & n6511 ;
  assign n19526 = n19525 ^ n6372 ^ 1'b0 ;
  assign n19527 = n1126 & ~n19526 ;
  assign n19528 = n461 & ~n19527 ;
  assign n19529 = n19528 ^ x99 ^ 1'b0 ;
  assign n19530 = n10718 & ~n13867 ;
  assign n19531 = ~n6340 & n18932 ;
  assign n19532 = n1706 | n2138 ;
  assign n19533 = n19532 ^ n3480 ^ 1'b0 ;
  assign n19534 = n4506 | n19533 ;
  assign n19535 = n13506 ^ n10350 ^ 1'b0 ;
  assign n19536 = n13228 & ~n19535 ;
  assign n19537 = n12185 & ~n14197 ;
  assign n19538 = n19537 ^ n5998 ^ 1'b0 ;
  assign n19539 = n12080 ^ n2173 ^ 1'b0 ;
  assign n19540 = n19538 & ~n19539 ;
  assign n19541 = ~n5656 & n19540 ;
  assign n19542 = n19541 ^ n10563 ^ 1'b0 ;
  assign n19543 = ~n1227 & n5182 ;
  assign n19544 = n19543 ^ n4054 ^ 1'b0 ;
  assign n19545 = n19542 & ~n19544 ;
  assign n19546 = n9449 & n19545 ;
  assign n19547 = n10754 & n19546 ;
  assign n19548 = n8696 ^ n7121 ^ 1'b0 ;
  assign n19549 = n16627 ^ n3118 ^ 1'b0 ;
  assign n19550 = n11242 & n12789 ;
  assign n19551 = ~n18284 & n19550 ;
  assign n19552 = n12305 ^ n9564 ^ 1'b0 ;
  assign n19553 = n19552 ^ n1559 ^ 1'b0 ;
  assign n19554 = n6754 ^ n1181 ^ 1'b0 ;
  assign n19555 = n5512 & n19554 ;
  assign n19556 = n15395 & n19555 ;
  assign n19557 = n19556 ^ n5452 ^ 1'b0 ;
  assign n19558 = n11945 & ~n19557 ;
  assign n19559 = n6018 & n8468 ;
  assign n19560 = n19559 ^ n4041 ^ 1'b0 ;
  assign n19561 = n10436 & ~n19560 ;
  assign n19563 = n4836 & ~n10924 ;
  assign n19564 = n19563 ^ n2393 ^ 1'b0 ;
  assign n19562 = n6528 | n13103 ;
  assign n19565 = n19564 ^ n19562 ^ 1'b0 ;
  assign n19566 = ~n1195 & n2277 ;
  assign n19567 = n19565 & n19566 ;
  assign n19568 = n6486 ^ n1236 ^ 1'b0 ;
  assign n19569 = n4516 & n7019 ;
  assign n19570 = ~n1675 & n19569 ;
  assign n19571 = n19570 ^ n11345 ^ 1'b0 ;
  assign n19572 = ~n9608 & n19571 ;
  assign n19573 = n6199 | n14072 ;
  assign n19574 = n19573 ^ n2720 ^ 1'b0 ;
  assign n19575 = n13052 ^ n5956 ^ 1'b0 ;
  assign n19576 = x110 & ~n14978 ;
  assign n19577 = n19575 & n19576 ;
  assign n19578 = ~n11671 & n16889 ;
  assign n19579 = n6106 & n19555 ;
  assign n19580 = n18289 & n19579 ;
  assign n19581 = n6087 | n9461 ;
  assign n19582 = ~n3321 & n12420 ;
  assign n19583 = n19582 ^ n14288 ^ 1'b0 ;
  assign n19584 = n12592 ^ n2778 ^ 1'b0 ;
  assign n19585 = n19583 & ~n19584 ;
  assign n19586 = n4086 ^ n4075 ^ 1'b0 ;
  assign n19587 = n5240 ^ n2423 ^ 1'b0 ;
  assign n19588 = n19586 | n19587 ;
  assign n19589 = n809 ^ x253 ^ 1'b0 ;
  assign n19590 = n5645 ^ n5636 ^ 1'b0 ;
  assign n19591 = n16989 | n19590 ;
  assign n19592 = n19591 ^ n8932 ^ 1'b0 ;
  assign n19593 = n4467 & ~n8358 ;
  assign n19594 = n1117 & n2475 ;
  assign n19595 = ~n18876 & n19594 ;
  assign n19596 = ~n959 & n13268 ;
  assign n19597 = ~n3429 & n19596 ;
  assign n19598 = n7097 & ~n19597 ;
  assign n19599 = n19598 ^ n8448 ^ 1'b0 ;
  assign n19600 = n8742 & n12381 ;
  assign n19601 = n19600 ^ n4960 ^ 1'b0 ;
  assign n19602 = n10092 ^ n3886 ^ 1'b0 ;
  assign n19603 = n12694 | n19602 ;
  assign n19604 = n19603 ^ n2311 ^ 1'b0 ;
  assign n19607 = n423 & n2185 ;
  assign n19608 = n19607 ^ n2891 ^ 1'b0 ;
  assign n19605 = n7528 ^ n3210 ^ 1'b0 ;
  assign n19606 = n5994 & n19605 ;
  assign n19609 = n19608 ^ n19606 ^ 1'b0 ;
  assign n19610 = n2187 | n19609 ;
  assign n19611 = n9816 ^ n3740 ^ 1'b0 ;
  assign n19612 = n1698 | n19611 ;
  assign n19613 = n6207 & n19612 ;
  assign n19614 = n19610 | n19613 ;
  assign n19615 = n10520 ^ n8773 ^ 1'b0 ;
  assign n19616 = n13139 ^ n5828 ^ 1'b0 ;
  assign n19617 = n14924 & n19616 ;
  assign n19618 = n15179 ^ n436 ^ 1'b0 ;
  assign n19619 = ~n8164 & n19618 ;
  assign n19620 = n13301 ^ n8181 ^ 1'b0 ;
  assign n19621 = n14554 ^ n6054 ^ 1'b0 ;
  assign n19622 = n19621 ^ n11373 ^ 1'b0 ;
  assign n19623 = n1901 & n6682 ;
  assign n19624 = n3774 ^ n3694 ^ 1'b0 ;
  assign n19625 = n19623 | n19624 ;
  assign n19626 = n14124 & ~n19625 ;
  assign n19627 = n1522 & n19626 ;
  assign n19629 = n2463 & ~n2818 ;
  assign n19628 = n1047 & n6162 ;
  assign n19630 = n19629 ^ n19628 ^ 1'b0 ;
  assign n19632 = n6876 & ~n9539 ;
  assign n19633 = n19632 ^ n1400 ^ 1'b0 ;
  assign n19631 = n2778 & ~n3532 ;
  assign n19634 = n19633 ^ n19631 ^ 1'b0 ;
  assign n19635 = n19634 ^ n9741 ^ 1'b0 ;
  assign n19636 = n10048 ^ n3641 ^ 1'b0 ;
  assign n19637 = n13521 & n19636 ;
  assign n19639 = n12716 & n17172 ;
  assign n19640 = n19639 ^ n11357 ^ 1'b0 ;
  assign n19641 = ~n956 & n19640 ;
  assign n19642 = n19641 ^ n10843 ^ 1'b0 ;
  assign n19643 = n663 & ~n19642 ;
  assign n19638 = n10167 & ~n15897 ;
  assign n19644 = n19643 ^ n19638 ^ 1'b0 ;
  assign n19645 = n5814 | n19644 ;
  assign n19646 = n3333 | n19645 ;
  assign n19651 = n5504 ^ n1793 ^ 1'b0 ;
  assign n19652 = n1068 | n19651 ;
  assign n19647 = n12691 ^ n4682 ^ 1'b0 ;
  assign n19648 = ~n11074 & n19647 ;
  assign n19649 = ~n16619 & n19648 ;
  assign n19650 = x143 & n19649 ;
  assign n19653 = n19652 ^ n19650 ^ 1'b0 ;
  assign n19654 = n14511 ^ x89 ^ 1'b0 ;
  assign n19655 = n14304 | n19654 ;
  assign n19656 = x0 & n3621 ;
  assign n19657 = n3908 & n5968 ;
  assign n19658 = ~n5968 & n19657 ;
  assign n19659 = x28 & ~n19658 ;
  assign n19660 = ~x28 & n19659 ;
  assign n19661 = n11666 & ~n19660 ;
  assign n19662 = n19660 & n19661 ;
  assign n19663 = n19662 ^ n11454 ^ 1'b0 ;
  assign n19664 = ~n15884 & n19663 ;
  assign n19665 = ~n5232 & n19664 ;
  assign n19666 = n1885 ^ n1846 ^ 1'b0 ;
  assign n19667 = n4946 & n19666 ;
  assign n19668 = n19667 ^ n8644 ^ 1'b0 ;
  assign n19669 = n4396 ^ n2215 ^ 1'b0 ;
  assign n19670 = ~x151 & n8364 ;
  assign n19671 = n14159 & n19670 ;
  assign n19672 = n19671 ^ n9911 ^ 1'b0 ;
  assign n19673 = n403 | n19672 ;
  assign n19674 = ~n597 & n3069 ;
  assign n19675 = ~n18905 & n19674 ;
  assign n19676 = n1080 | n8531 ;
  assign n19677 = n19676 ^ n2954 ^ 1'b0 ;
  assign n19678 = n4375 & ~n19677 ;
  assign n19679 = n10974 ^ n8553 ^ 1'b0 ;
  assign n19680 = n4821 & ~n16702 ;
  assign n19681 = ~n4927 & n6313 ;
  assign n19682 = n19681 ^ n2987 ^ 1'b0 ;
  assign n19683 = n6211 ^ n1485 ^ 1'b0 ;
  assign n19684 = n9174 | n19683 ;
  assign n19685 = n1630 | n19684 ;
  assign n19686 = n19685 ^ n4101 ^ 1'b0 ;
  assign n19687 = n5223 | n19686 ;
  assign n19688 = n725 & ~n4766 ;
  assign n19689 = ~n12695 & n19688 ;
  assign n19690 = n2296 & ~n16733 ;
  assign n19691 = n19690 ^ n1029 ^ 1'b0 ;
  assign n19692 = n19691 ^ n1575 ^ 1'b0 ;
  assign n19693 = n897 & n19692 ;
  assign n19694 = ~n1239 & n3895 ;
  assign n19695 = n6382 & ~n7865 ;
  assign n19696 = ~n9126 & n19695 ;
  assign n19697 = n10278 | n19696 ;
  assign n19698 = ~n4433 & n14401 ;
  assign n19700 = n461 & n9339 ;
  assign n19701 = n19700 ^ n8827 ^ 1'b0 ;
  assign n19702 = n19701 ^ n6614 ^ 1'b0 ;
  assign n19699 = n2906 | n14375 ;
  assign n19703 = n19702 ^ n19699 ^ 1'b0 ;
  assign n19704 = n15425 ^ n5355 ^ 1'b0 ;
  assign n19705 = n10918 & n12961 ;
  assign n19706 = ~n1159 & n4529 ;
  assign n19707 = n19705 & n19706 ;
  assign n19708 = n4677 & ~n14953 ;
  assign n19709 = n6411 & ~n14445 ;
  assign n19710 = n19709 ^ n9444 ^ 1'b0 ;
  assign n19711 = ~n329 & n19710 ;
  assign n19712 = n3371 & n19711 ;
  assign n19713 = n17736 ^ n10160 ^ 1'b0 ;
  assign n19714 = n19712 | n19713 ;
  assign n19715 = n2725 & n17182 ;
  assign n19716 = n14971 ^ n10035 ^ n3872 ;
  assign n19717 = n15515 ^ n10303 ^ 1'b0 ;
  assign n19719 = ~n401 & n12030 ;
  assign n19718 = ( n2380 & n11751 ) | ( n2380 & ~n17379 ) | ( n11751 & ~n17379 ) ;
  assign n19720 = n19719 ^ n19718 ^ 1'b0 ;
  assign n19721 = n8872 ^ n1812 ^ 1'b0 ;
  assign n19722 = n5106 & n19721 ;
  assign n19723 = n5669 ^ n3431 ^ 1'b0 ;
  assign n19724 = n3575 & n19723 ;
  assign n19725 = ( n8162 & n19722 ) | ( n8162 & ~n19724 ) | ( n19722 & ~n19724 ) ;
  assign n19726 = n12468 ^ n3111 ^ 1'b0 ;
  assign n19727 = n1273 & ~n4715 ;
  assign n19728 = n19727 ^ n7407 ^ 1'b0 ;
  assign n19729 = n17014 | n19728 ;
  assign n19730 = n7809 & ~n19729 ;
  assign n19731 = n9860 ^ n6886 ^ 1'b0 ;
  assign n19732 = n1540 & n19075 ;
  assign n19733 = ~n5032 & n19732 ;
  assign n19734 = n3120 ^ n2181 ^ 1'b0 ;
  assign n19735 = n3248 & ~n5879 ;
  assign n19736 = ~n2175 & n8947 ;
  assign n19737 = n11591 ^ n637 ^ 1'b0 ;
  assign n19738 = n19736 & n19737 ;
  assign n19739 = ~n5626 & n19738 ;
  assign n19740 = n19735 & n19739 ;
  assign n19741 = n838 & n6629 ;
  assign n19742 = n19741 ^ n4066 ^ 1'b0 ;
  assign n19743 = n19742 ^ n12030 ^ 1'b0 ;
  assign n19744 = n4271 | n19743 ;
  assign n19745 = n7501 & ~n12013 ;
  assign n19746 = n19744 & n19745 ;
  assign n19747 = n12723 | n19746 ;
  assign n19748 = x61 | n15540 ;
  assign n19749 = n9382 | n19748 ;
  assign n19750 = n4122 ^ n3903 ^ 1'b0 ;
  assign n19751 = n6950 | n10267 ;
  assign n19752 = n17255 & ~n19751 ;
  assign n19753 = n3982 & n10744 ;
  assign n19754 = n311 & ~n7466 ;
  assign n19755 = n2623 | n11847 ;
  assign n19756 = ~n8320 & n9135 ;
  assign n19757 = n17395 | n19756 ;
  assign n19758 = n19757 ^ n7838 ^ 1'b0 ;
  assign n19759 = n19758 ^ n2495 ^ 1'b0 ;
  assign n19760 = n10118 & ~n19759 ;
  assign n19761 = ~n10094 & n16160 ;
  assign n19762 = n19761 ^ n7275 ^ 1'b0 ;
  assign n19763 = n19762 ^ n6255 ^ 1'b0 ;
  assign n19764 = n4705 & ~n5890 ;
  assign n19765 = ~n5032 & n7863 ;
  assign n19766 = n19765 ^ n18206 ^ n9913 ;
  assign n19767 = n4919 | n10924 ;
  assign n19768 = n19767 ^ n2140 ^ 1'b0 ;
  assign n19769 = n12241 & ~n19768 ;
  assign n19770 = ~n9279 & n19769 ;
  assign n19771 = n11654 ^ n9446 ^ n8990 ;
  assign n19772 = n19771 ^ n526 ^ 1'b0 ;
  assign n19773 = n14689 ^ n2804 ^ 1'b0 ;
  assign n19774 = n8020 & n19773 ;
  assign n19775 = ( n1154 & n1366 ) | ( n1154 & n2423 ) | ( n1366 & n2423 ) ;
  assign n19776 = n19775 ^ n4570 ^ 1'b0 ;
  assign n19777 = ~n15918 & n19776 ;
  assign n19778 = n18148 & n19777 ;
  assign n19779 = ~n11268 & n19778 ;
  assign n19787 = ~n1295 & n5330 ;
  assign n19788 = n1295 & n19787 ;
  assign n19784 = n643 & n744 ;
  assign n19785 = ~n643 & n19784 ;
  assign n19782 = n1850 & n6557 ;
  assign n19783 = ~n6557 & n19782 ;
  assign n19786 = n19785 ^ n19783 ^ 1'b0 ;
  assign n19789 = n19788 ^ n19786 ^ n11052 ;
  assign n19780 = n12738 ^ n1673 ^ 1'b0 ;
  assign n19781 = n14479 & ~n19780 ;
  assign n19790 = n19789 ^ n19781 ^ 1'b0 ;
  assign n19791 = n3097 & ~n19790 ;
  assign n19794 = n1075 & n2854 ;
  assign n19792 = n14373 ^ n2546 ^ 1'b0 ;
  assign n19793 = n3811 | n19792 ;
  assign n19795 = n19794 ^ n19793 ^ 1'b0 ;
  assign n19796 = n6784 & ~n19795 ;
  assign n19797 = n1354 & n19796 ;
  assign n19798 = n4647 & ~n19797 ;
  assign n19799 = n717 & ~n6039 ;
  assign n19800 = n19799 ^ n9764 ^ 1'b0 ;
  assign n19801 = n5991 | n11797 ;
  assign n19802 = ~n1656 & n19801 ;
  assign n19803 = ~n3855 & n19802 ;
  assign n19804 = n18734 ^ n15827 ^ 1'b0 ;
  assign n19806 = n5029 ^ n275 ^ 1'b0 ;
  assign n19807 = n8010 & n19806 ;
  assign n19808 = n12572 & n19807 ;
  assign n19805 = n12990 ^ n6311 ^ 1'b0 ;
  assign n19809 = n19808 ^ n19805 ^ n4854 ;
  assign n19810 = n13793 ^ n7789 ^ 1'b0 ;
  assign n19811 = n7189 | n19810 ;
  assign n19812 = n2162 | n16770 ;
  assign n19813 = n13372 & ~n19812 ;
  assign n19814 = n10986 ^ n3069 ^ 1'b0 ;
  assign n19815 = n19352 & n19814 ;
  assign n19816 = n18644 & n19815 ;
  assign n19820 = n7100 ^ n1082 ^ 1'b0 ;
  assign n19817 = n2397 & n3865 ;
  assign n19818 = n5066 & n19817 ;
  assign n19819 = n19818 ^ n8244 ^ 1'b0 ;
  assign n19821 = n19820 ^ n19819 ^ 1'b0 ;
  assign n19822 = ~x23 & n19821 ;
  assign n19823 = n3608 & n19017 ;
  assign n19824 = ~n16928 & n19823 ;
  assign n19825 = ~n8564 & n10000 ;
  assign n19826 = n7785 & n19825 ;
  assign n19827 = n11859 | n19826 ;
  assign n19828 = n9929 & ~n19827 ;
  assign n19829 = ~n8516 & n15142 ;
  assign n19830 = n18604 ^ n18309 ^ 1'b0 ;
  assign n19831 = ~n4294 & n14778 ;
  assign n19832 = n18751 ^ n18339 ^ 1'b0 ;
  assign n19833 = n2707 & ~n2846 ;
  assign n19834 = ~n5366 & n19833 ;
  assign n19835 = n6093 & ~n7723 ;
  assign n19836 = x202 | n7545 ;
  assign n19837 = ~n2431 & n19836 ;
  assign n19838 = n19835 & ~n19837 ;
  assign n19839 = n19838 ^ n13850 ^ 1'b0 ;
  assign n19840 = n7680 ^ n2021 ^ 1'b0 ;
  assign n19841 = ~n2760 & n5784 ;
  assign n19842 = n7438 | n19841 ;
  assign n19843 = n19840 | n19842 ;
  assign n19844 = ~n939 & n19843 ;
  assign n19845 = n19844 ^ n1890 ^ 1'b0 ;
  assign n19846 = n19137 ^ n16284 ^ 1'b0 ;
  assign n19847 = n1018 | n19846 ;
  assign n19848 = n1985 & n10046 ;
  assign n19849 = n3049 | n19848 ;
  assign n19850 = n19849 ^ n9361 ^ 1'b0 ;
  assign n19851 = n14041 ^ n6584 ^ 1'b0 ;
  assign n19852 = n6681 & n19851 ;
  assign n19853 = n19852 ^ n10443 ^ 1'b0 ;
  assign n19854 = n1233 & n4917 ;
  assign n19855 = n7179 & ~n19854 ;
  assign n19856 = n19855 ^ n12743 ^ 1'b0 ;
  assign n19857 = n8913 ^ n5650 ^ x60 ;
  assign n19858 = n14602 ^ n12981 ^ 1'b0 ;
  assign n19859 = n3221 & ~n6162 ;
  assign n19860 = ~n3221 & n19859 ;
  assign n19861 = n19860 ^ n17163 ^ 1'b0 ;
  assign n19862 = ~n19858 & n19861 ;
  assign n19863 = n19858 & n19862 ;
  assign n19864 = n6737 & ~n11991 ;
  assign n19865 = n14350 & n19864 ;
  assign n19866 = n13043 ^ n9578 ^ n3412 ;
  assign n19867 = ~n1354 & n3698 ;
  assign n19868 = n19867 ^ n9154 ^ 1'b0 ;
  assign n19869 = n2223 | n19868 ;
  assign n19870 = n18432 ^ n13348 ^ 1'b0 ;
  assign n19871 = n1505 ^ n648 ^ 1'b0 ;
  assign n19872 = n19871 ^ n9208 ^ n5401 ;
  assign n19873 = x57 & ~n6794 ;
  assign n19874 = n4488 ^ n3415 ^ 1'b0 ;
  assign n19875 = ~n13768 & n19874 ;
  assign n19876 = n7785 ^ n1028 ^ 1'b0 ;
  assign n19877 = n19875 & n19876 ;
  assign n19878 = n6735 & ~n19877 ;
  assign n19879 = n14374 ^ n1308 ^ 1'b0 ;
  assign n19883 = n19000 ^ n12255 ^ 1'b0 ;
  assign n19880 = ~n930 & n9153 ;
  assign n19881 = ~n6972 & n19880 ;
  assign n19882 = n13422 & ~n19881 ;
  assign n19884 = n19883 ^ n19882 ^ 1'b0 ;
  assign n19885 = x228 & n6231 ;
  assign n19886 = n19885 ^ n10089 ^ 1'b0 ;
  assign n19887 = n16367 ^ n10523 ^ 1'b0 ;
  assign n19888 = n3964 & ~n4780 ;
  assign n19889 = n19888 ^ n9894 ^ 1'b0 ;
  assign n19890 = n3477 ^ n519 ^ 1'b0 ;
  assign n19891 = n7349 & n19890 ;
  assign n19892 = n17307 | n19891 ;
  assign n19893 = n14997 ^ n14708 ^ 1'b0 ;
  assign n19894 = n3656 | n14502 ;
  assign n19895 = n19894 ^ n16418 ^ 1'b0 ;
  assign n19896 = n14093 ^ n13012 ^ 1'b0 ;
  assign n19897 = ~n1499 & n12680 ;
  assign n19903 = n2394 & ~n10663 ;
  assign n19904 = ~n2394 & n19903 ;
  assign n19898 = n3307 & ~n8314 ;
  assign n19899 = ~n3307 & n19898 ;
  assign n19900 = x204 & ~n12032 ;
  assign n19901 = n19900 ^ n1658 ^ 1'b0 ;
  assign n19902 = ~n19899 & n19901 ;
  assign n19905 = n19904 ^ n19902 ^ 1'b0 ;
  assign n19906 = n5060 ^ n4971 ^ 1'b0 ;
  assign n19907 = n13570 & ~n19906 ;
  assign n19908 = n19907 ^ n10452 ^ 1'b0 ;
  assign n19909 = n9065 & ~n10220 ;
  assign n19910 = n19909 ^ n16621 ^ 1'b0 ;
  assign n19911 = n19910 ^ n19591 ^ 1'b0 ;
  assign n19912 = n19911 ^ n9105 ^ 1'b0 ;
  assign n19913 = n19908 & n19912 ;
  assign n19915 = n10875 ^ n7206 ^ 1'b0 ;
  assign n19914 = n1981 & n14654 ;
  assign n19916 = n19915 ^ n19914 ^ 1'b0 ;
  assign n19917 = n5665 | n9991 ;
  assign n19918 = ~n1190 & n8449 ;
  assign n19919 = n19918 ^ n1964 ^ 1'b0 ;
  assign n19920 = n9197 & n19024 ;
  assign n19921 = n19920 ^ n18219 ^ 1'b0 ;
  assign n19922 = ~x85 & n10817 ;
  assign n19923 = n3731 | n18732 ;
  assign n19924 = n18196 | n19923 ;
  assign n19925 = ~n6330 & n19924 ;
  assign n19926 = n1395 & n16399 ;
  assign n19927 = n19926 ^ n18353 ^ 1'b0 ;
  assign n19928 = ~n749 & n1608 ;
  assign n19929 = n19928 ^ n16594 ^ 1'b0 ;
  assign n19930 = n4117 | n7657 ;
  assign n19931 = n19930 ^ n1518 ^ 1'b0 ;
  assign n19932 = ~n4873 & n5484 ;
  assign n19933 = n19932 ^ n728 ^ 1'b0 ;
  assign n19934 = n3440 & n12121 ;
  assign n19935 = n16134 & n19934 ;
  assign n19936 = ~n1775 & n6517 ;
  assign n19937 = n1495 & ~n3333 ;
  assign n19938 = n3059 & n19937 ;
  assign n19939 = n10877 & ~n19938 ;
  assign n19940 = n19652 ^ n6700 ^ 1'b0 ;
  assign n19941 = n9111 ^ n283 ^ 1'b0 ;
  assign n19942 = n5765 & n19941 ;
  assign n19943 = n5908 & n10827 ;
  assign n19944 = n19942 & n19943 ;
  assign n19945 = n19944 ^ n16055 ^ 1'b0 ;
  assign n19946 = n4940 | n17754 ;
  assign n19947 = n6236 & ~n19946 ;
  assign n19948 = n19947 ^ n19824 ^ 1'b0 ;
  assign n19949 = n5857 | n13248 ;
  assign n19950 = n19949 ^ n747 ^ 1'b0 ;
  assign n19951 = n9578 & ~n19950 ;
  assign n19952 = n418 ^ n337 ^ 1'b0 ;
  assign n19953 = n415 & ~n19952 ;
  assign n19954 = n19124 ^ n18519 ^ 1'b0 ;
  assign n19955 = n19954 ^ x81 ^ 1'b0 ;
  assign n19956 = n10145 & ~n19955 ;
  assign n19957 = ( n754 & ~n2275 ) | ( n754 & n3697 ) | ( ~n2275 & n3697 ) ;
  assign n19958 = n10018 & ~n15088 ;
  assign n19959 = ( n17726 & n19957 ) | ( n17726 & ~n19958 ) | ( n19957 & ~n19958 ) ;
  assign n19961 = n1181 & ~n3718 ;
  assign n19962 = n3718 & n19961 ;
  assign n19963 = n13721 | n19962 ;
  assign n19964 = n19963 ^ n6150 ^ 1'b0 ;
  assign n19965 = n7636 & ~n11668 ;
  assign n19966 = ~n19964 & n19965 ;
  assign n19960 = n9690 | n11568 ;
  assign n19967 = n19966 ^ n19960 ^ 1'b0 ;
  assign n19968 = ~n5897 & n8475 ;
  assign n19969 = n1641 & n5767 ;
  assign n19971 = ~n7643 & n9836 ;
  assign n19972 = ~n4329 & n19971 ;
  assign n19973 = n8096 ^ n1393 ^ 1'b0 ;
  assign n19974 = n19972 | n19973 ;
  assign n19970 = ~n6948 & n10646 ;
  assign n19975 = n19974 ^ n19970 ^ 1'b0 ;
  assign n19976 = n4712 ^ n3099 ^ 1'b0 ;
  assign n19977 = n3334 | n19976 ;
  assign n19978 = ~n3462 & n9793 ;
  assign n19979 = n11543 & n19978 ;
  assign n19980 = n16090 ^ n10404 ^ 1'b0 ;
  assign n19981 = ~n2072 & n14205 ;
  assign n19982 = n19980 & n19981 ;
  assign n19983 = n5484 | n7816 ;
  assign n19984 = n19983 ^ n15217 ^ 1'b0 ;
  assign n19985 = n6710 & n9194 ;
  assign n19986 = x248 & n19985 ;
  assign n19987 = n19986 ^ n11738 ^ 1'b0 ;
  assign n19988 = n8957 & n17540 ;
  assign n19989 = n19988 ^ n9854 ^ 1'b0 ;
  assign n19990 = n8392 & n19989 ;
  assign n19991 = n19990 ^ n13093 ^ 1'b0 ;
  assign n19993 = ~n2283 & n2669 ;
  assign n19994 = n19993 ^ n18068 ^ 1'b0 ;
  assign n19995 = n8198 ^ n6633 ^ 1'b0 ;
  assign n19996 = n19994 & ~n19995 ;
  assign n19992 = n18835 ^ n16076 ^ 1'b0 ;
  assign n19997 = n19996 ^ n19992 ^ 1'b0 ;
  assign n19998 = n6516 ^ n4222 ^ 1'b0 ;
  assign n19999 = n6637 & ~n19998 ;
  assign n20000 = ~n11196 & n19999 ;
  assign n20001 = n11304 & n17754 ;
  assign n20002 = n20000 | n20001 ;
  assign n20003 = n20002 ^ n1910 ^ 1'b0 ;
  assign n20007 = n15566 ^ n1324 ^ 1'b0 ;
  assign n20004 = n3959 | n4301 ;
  assign n20005 = n3199 & ~n17506 ;
  assign n20006 = n20004 & n20005 ;
  assign n20008 = n20007 ^ n20006 ^ 1'b0 ;
  assign n20009 = n4728 & ~n9350 ;
  assign n20010 = ~n16351 & n20009 ;
  assign n20011 = n20010 ^ n2630 ^ 1'b0 ;
  assign n20012 = n8289 ^ n4828 ^ 1'b0 ;
  assign n20013 = n3984 | n4965 ;
  assign n20014 = ~n4747 & n20013 ;
  assign n20015 = ~n12397 & n20014 ;
  assign n20016 = n20015 ^ n16206 ^ n2589 ;
  assign n20017 = n7248 & n12576 ;
  assign n20018 = n10314 | n18053 ;
  assign n20019 = n20018 ^ n5082 ^ 1'b0 ;
  assign n20020 = ~x42 & n20019 ;
  assign n20021 = n16767 & n20020 ;
  assign n20022 = n11768 ^ n3086 ^ n2079 ;
  assign n20023 = n20022 ^ n12134 ^ 1'b0 ;
  assign n20024 = n8192 & ~n14871 ;
  assign n20025 = n20024 ^ n18788 ^ 1'b0 ;
  assign n20026 = x174 & n13741 ;
  assign n20027 = n20026 ^ n1510 ^ 1'b0 ;
  assign n20028 = n5157 | n10556 ;
  assign n20029 = ~n681 & n3869 ;
  assign n20030 = ~n4834 & n20029 ;
  assign n20031 = n20030 ^ n4553 ^ 1'b0 ;
  assign n20032 = n728 & n1847 ;
  assign n20033 = n20032 ^ n2861 ^ 1'b0 ;
  assign n20034 = n3053 ^ n1826 ^ 1'b0 ;
  assign n20035 = n20033 & ~n20034 ;
  assign n20036 = n1601 & ~n15891 ;
  assign n20037 = n5031 & n20036 ;
  assign n20038 = n2920 & ~n14144 ;
  assign n20039 = ~n2920 & n20038 ;
  assign n20040 = n3248 & n20039 ;
  assign n20041 = n9672 ^ n4562 ^ 1'b0 ;
  assign n20042 = n20040 & n20041 ;
  assign n20043 = n2399 & n20042 ;
  assign n20044 = n20037 | n20043 ;
  assign n20045 = n20037 & ~n20044 ;
  assign n20046 = n6783 & ~n20045 ;
  assign n20047 = n20045 & n20046 ;
  assign n20048 = n1727 ^ n1637 ^ 1'b0 ;
  assign n20049 = ~n20047 & n20048 ;
  assign n20062 = n2368 & ~n11557 ;
  assign n20063 = ~n2368 & n20062 ;
  assign n20064 = n4913 & n20063 ;
  assign n20065 = ~n10513 & n20064 ;
  assign n20066 = n10513 & n20065 ;
  assign n20055 = x134 & ~n366 ;
  assign n20056 = ~x134 & n20055 ;
  assign n20057 = n3336 | n20056 ;
  assign n20058 = n3336 & ~n20057 ;
  assign n20059 = n1232 | n2770 ;
  assign n20060 = n20058 & ~n20059 ;
  assign n20061 = n12154 | n20060 ;
  assign n20067 = n20066 ^ n20061 ^ 1'b0 ;
  assign n20050 = n2393 ^ n779 ^ 1'b0 ;
  assign n20051 = n5105 | n20050 ;
  assign n20052 = n20050 & ~n20051 ;
  assign n20053 = n380 & ~n5775 ;
  assign n20054 = ~n20052 & n20053 ;
  assign n20068 = n20067 ^ n20054 ^ 1'b0 ;
  assign n20069 = n20049 & ~n20068 ;
  assign n20071 = n4425 | n5118 ;
  assign n20072 = n3318 & ~n20071 ;
  assign n20070 = n12238 & n15348 ;
  assign n20073 = n20072 ^ n20070 ^ 1'b0 ;
  assign n20074 = n17304 ^ n15444 ^ 1'b0 ;
  assign n20075 = n13447 & ~n20074 ;
  assign n20076 = n14184 & n20075 ;
  assign n20077 = n20076 ^ n2863 ^ 1'b0 ;
  assign n20078 = n10240 & n17073 ;
  assign n20079 = n7135 ^ n3501 ^ 1'b0 ;
  assign n20080 = n8387 | n9793 ;
  assign n20081 = n9137 & ~n20080 ;
  assign n20082 = n4755 ^ n3395 ^ 1'b0 ;
  assign n20083 = n1793 & n20082 ;
  assign n20084 = n20083 ^ n3891 ^ 1'b0 ;
  assign n20085 = n309 | n11271 ;
  assign n20086 = ~n20084 & n20085 ;
  assign n20087 = n8755 ^ n8546 ^ 1'b0 ;
  assign n20088 = n5742 & ~n20087 ;
  assign n20089 = ~n16993 & n20088 ;
  assign n20090 = n3880 ^ n3089 ^ 1'b0 ;
  assign n20091 = ~n2720 & n11207 ;
  assign n20092 = n2026 | n12531 ;
  assign n20093 = n722 & ~n10222 ;
  assign n20094 = n20093 ^ n3049 ^ 1'b0 ;
  assign n20095 = n13630 & n20094 ;
  assign n20096 = n20092 & n20095 ;
  assign n20097 = n2117 | n11488 ;
  assign n20098 = n9630 & ~n20097 ;
  assign n20099 = n20098 ^ n8169 ^ 1'b0 ;
  assign n20100 = n20099 ^ n9060 ^ 1'b0 ;
  assign n20102 = n6756 & n14866 ;
  assign n20103 = n13252 & n20102 ;
  assign n20101 = n1094 & n8580 ;
  assign n20104 = n20103 ^ n20101 ^ 1'b0 ;
  assign n20105 = n4506 ^ n460 ^ 1'b0 ;
  assign n20106 = ~n12744 & n20105 ;
  assign n20107 = n3891 ^ n1186 ^ 1'b0 ;
  assign n20108 = n4932 & n20107 ;
  assign n20109 = n5265 | n7275 ;
  assign n20110 = n20109 ^ n7845 ^ 1'b0 ;
  assign n20112 = n1521 | n5155 ;
  assign n20113 = n7777 | n20112 ;
  assign n20114 = ~n18260 & n20113 ;
  assign n20115 = n20114 ^ n8074 ^ 1'b0 ;
  assign n20111 = n4384 & n17039 ;
  assign n20116 = n20115 ^ n20111 ^ 1'b0 ;
  assign n20117 = n20116 ^ n6601 ^ 1'b0 ;
  assign n20118 = n20110 & n20117 ;
  assign n20120 = n2599 & n12397 ;
  assign n20119 = n1540 & n5903 ;
  assign n20121 = n20120 ^ n20119 ^ 1'b0 ;
  assign n20122 = ~n2849 & n3759 ;
  assign n20125 = ~n1622 & n2093 ;
  assign n20124 = n327 | n4199 ;
  assign n20123 = n14612 ^ n7028 ^ 1'b0 ;
  assign n20126 = n20125 ^ n20124 ^ n20123 ;
  assign n20127 = n10564 ^ n2474 ^ 1'b0 ;
  assign n20128 = n6804 & ~n20127 ;
  assign n20129 = n20128 ^ n14250 ^ 1'b0 ;
  assign n20130 = n18243 & n20129 ;
  assign n20131 = x130 & ~n4913 ;
  assign n20132 = n8846 & n20131 ;
  assign n20133 = n535 & ~n7732 ;
  assign n20134 = n4385 ^ n3869 ^ 1'b0 ;
  assign n20135 = n9609 & ~n20134 ;
  assign n20136 = n20135 ^ n13109 ^ 1'b0 ;
  assign n20137 = n20133 | n20136 ;
  assign n20138 = n20132 & ~n20137 ;
  assign n20139 = n17969 ^ n12412 ^ 1'b0 ;
  assign n20140 = n6146 ^ n5468 ^ 1'b0 ;
  assign n20141 = n7248 ^ n1622 ^ 1'b0 ;
  assign n20142 = n9345 ^ n1298 ^ 1'b0 ;
  assign n20143 = n20142 ^ n17800 ^ 1'b0 ;
  assign n20144 = n20141 & n20143 ;
  assign n20145 = n15458 ^ n12932 ^ n4819 ;
  assign n20146 = n20145 ^ n19437 ^ 1'b0 ;
  assign n20147 = n6070 & n20146 ;
  assign n20148 = n5020 & ~n15841 ;
  assign n20149 = n2524 & n20148 ;
  assign n20150 = n7508 & n20149 ;
  assign n20151 = n15463 & n17269 ;
  assign n20152 = ~n2957 & n16101 ;
  assign n20153 = n13852 & n20152 ;
  assign n20154 = n19464 ^ n8319 ^ 1'b0 ;
  assign n20155 = n19736 & n20154 ;
  assign n20156 = n12559 ^ n2364 ^ 1'b0 ;
  assign n20157 = n13301 & n20156 ;
  assign n20158 = n20157 ^ n4145 ^ 1'b0 ;
  assign n20159 = ~n19689 & n20158 ;
  assign n20160 = ~n20155 & n20159 ;
  assign n20161 = n7516 ^ n820 ^ 1'b0 ;
  assign n20162 = n1854 & n6220 ;
  assign n20163 = n797 & n3046 ;
  assign n20164 = n20163 ^ n14845 ^ 1'b0 ;
  assign n20165 = n6145 ^ n1525 ^ 1'b0 ;
  assign n20166 = n20164 | n20165 ;
  assign n20167 = n20162 & ~n20166 ;
  assign n20168 = n7544 & n20167 ;
  assign n20169 = n8617 ^ n2846 ^ 1'b0 ;
  assign n20170 = n18658 ^ n3392 ^ 1'b0 ;
  assign n20171 = n4695 & ~n7046 ;
  assign n20172 = ~n10317 & n20171 ;
  assign n20173 = n11014 ^ n4178 ^ 1'b0 ;
  assign n20174 = ( ~n5433 & n13740 ) | ( ~n5433 & n20173 ) | ( n13740 & n20173 ) ;
  assign n20175 = n11261 ^ n8305 ^ 1'b0 ;
  assign n20176 = n6360 & n20175 ;
  assign n20177 = n4031 | n6618 ;
  assign n20178 = n20177 ^ n1487 ^ 1'b0 ;
  assign n20179 = n720 | n20178 ;
  assign n20180 = n1920 & ~n16785 ;
  assign n20181 = n20180 ^ n2153 ^ 1'b0 ;
  assign n20182 = n4701 & n20181 ;
  assign n20183 = n10865 & n20182 ;
  assign n20184 = n1969 & ~n3520 ;
  assign n20185 = n20184 ^ n4493 ^ 1'b0 ;
  assign n20186 = n629 | n20185 ;
  assign n20187 = ~n3059 & n8250 ;
  assign n20188 = ~n20186 & n20187 ;
  assign n20189 = n1602 & n18276 ;
  assign n20190 = ( n9921 & n17921 ) | ( n9921 & ~n20189 ) | ( n17921 & ~n20189 ) ;
  assign n20191 = ( n740 & n2838 ) | ( n740 & n10488 ) | ( n2838 & n10488 ) ;
  assign n20192 = n20191 ^ n12850 ^ 1'b0 ;
  assign n20193 = n17908 | n20192 ;
  assign n20194 = n9580 ^ n4238 ^ n3107 ;
  assign n20195 = n11538 | n20194 ;
  assign n20203 = n426 | n11119 ;
  assign n20196 = n918 & ~n1513 ;
  assign n20197 = ~n918 & n20196 ;
  assign n20198 = n535 & ~n1021 ;
  assign n20199 = n2892 | n3035 ;
  assign n20200 = n3035 & ~n20199 ;
  assign n20201 = ~n20198 & n20200 ;
  assign n20202 = ~n20197 & n20201 ;
  assign n20204 = n20203 ^ n20202 ^ 1'b0 ;
  assign n20205 = n18820 ^ n8727 ^ 1'b0 ;
  assign n20206 = n5050 & n20205 ;
  assign n20208 = n3610 ^ n3116 ^ 1'b0 ;
  assign n20207 = n3652 & ~n14652 ;
  assign n20209 = n20208 ^ n20207 ^ 1'b0 ;
  assign n20210 = ~n9358 & n20209 ;
  assign n20211 = n20123 ^ n2785 ^ 1'b0 ;
  assign n20212 = n1937 & ~n10620 ;
  assign n20213 = n20212 ^ n1566 ^ 1'b0 ;
  assign n20214 = n20213 ^ n10967 ^ 1'b0 ;
  assign n20215 = n20211 | n20214 ;
  assign n20216 = n4325 ^ n2615 ^ 1'b0 ;
  assign n20217 = n713 | n20216 ;
  assign n20218 = n12945 & ~n20217 ;
  assign n20219 = n9803 ^ n4382 ^ 1'b0 ;
  assign n20220 = ~n7974 & n20219 ;
  assign n20221 = ~n956 & n20220 ;
  assign n20222 = n20221 ^ n8162 ^ 1'b0 ;
  assign n20223 = n2466 ^ n2427 ^ 1'b0 ;
  assign n20224 = n19560 ^ n12305 ^ 1'b0 ;
  assign n20225 = n20223 | n20224 ;
  assign n20226 = n4897 | n5286 ;
  assign n20227 = n20225 & ~n20226 ;
  assign n20228 = ( ~n1490 & n2910 ) | ( ~n1490 & n4271 ) | ( n2910 & n4271 ) ;
  assign n20229 = n3833 ^ n2306 ^ 1'b0 ;
  assign n20230 = n20229 ^ n1419 ^ 1'b0 ;
  assign n20231 = n20228 & ~n20230 ;
  assign n20232 = n8900 ^ n8663 ^ n2357 ;
  assign n20233 = ( n4413 & ~n5750 ) | ( n4413 & n20232 ) | ( ~n5750 & n20232 ) ;
  assign n20234 = x93 | n17853 ;
  assign n20235 = n1099 | n19029 ;
  assign n20236 = n20235 ^ n14919 ^ 1'b0 ;
  assign n20237 = n7126 & ~n14182 ;
  assign n20238 = ( n6020 & n7467 ) | ( n6020 & n13393 ) | ( n7467 & n13393 ) ;
  assign n20239 = n12787 ^ n3895 ^ 1'b0 ;
  assign n20240 = n6596 ^ n2587 ^ 1'b0 ;
  assign n20241 = n2842 & n3578 ;
  assign n20242 = n20241 ^ n5438 ^ 1'b0 ;
  assign n20243 = n14993 | n20242 ;
  assign n20244 = n4243 & ~n5399 ;
  assign n20245 = n20243 & n20244 ;
  assign n20246 = n13520 & ~n20245 ;
  assign n20247 = n20246 ^ n1523 ^ 1'b0 ;
  assign n20248 = n430 & n3948 ;
  assign n20251 = n3561 ^ n2221 ^ 1'b0 ;
  assign n20249 = n10016 & n11754 ;
  assign n20250 = n20249 ^ n10963 ^ 1'b0 ;
  assign n20252 = n20251 ^ n20250 ^ n19095 ;
  assign n20254 = n2510 | n3683 ;
  assign n20255 = n4543 | n20254 ;
  assign n20256 = n20255 ^ n9342 ^ n6539 ;
  assign n20253 = n6662 ^ n6041 ^ 1'b0 ;
  assign n20257 = n20256 ^ n20253 ^ 1'b0 ;
  assign n20258 = n20257 ^ n14605 ^ 1'b0 ;
  assign n20259 = n602 & ~n14885 ;
  assign n20260 = n1606 | n5927 ;
  assign n20261 = n20260 ^ n2239 ^ 1'b0 ;
  assign n20263 = n9875 ^ n7430 ^ 1'b0 ;
  assign n20264 = n9458 & n20263 ;
  assign n20262 = n5047 & ~n10392 ;
  assign n20265 = n20264 ^ n20262 ^ 1'b0 ;
  assign n20269 = n5413 ^ n4586 ^ 1'b0 ;
  assign n20270 = n438 & ~n20269 ;
  assign n20266 = n7419 ^ n5624 ^ 1'b0 ;
  assign n20267 = n9976 & ~n20266 ;
  assign n20268 = n8336 & n20267 ;
  assign n20271 = n20270 ^ n20268 ^ 1'b0 ;
  assign n20272 = n5534 ^ n602 ^ 1'b0 ;
  assign n20273 = n15298 & ~n16303 ;
  assign n20274 = n20273 ^ n15265 ^ 1'b0 ;
  assign n20275 = ~n9208 & n20274 ;
  assign n20276 = n14853 & ~n18041 ;
  assign n20277 = n5015 | n18591 ;
  assign n20278 = n10306 & ~n20277 ;
  assign n20279 = n20278 ^ n5990 ^ 1'b0 ;
  assign n20280 = ~n6050 & n10456 ;
  assign n20281 = n20280 ^ n17554 ^ 1'b0 ;
  assign n20282 = n6165 ^ x75 ^ 1'b0 ;
  assign n20283 = ~n1056 & n20282 ;
  assign n20284 = n1572 & ~n3561 ;
  assign n20285 = n20283 & ~n20284 ;
  assign n20286 = ~n2374 & n11808 ;
  assign n20287 = n5574 & ~n7064 ;
  assign n20288 = ~n20142 & n20287 ;
  assign n20289 = n6727 & ~n11258 ;
  assign n20290 = n5332 & n12809 ;
  assign n20291 = n3217 ^ n2374 ^ 1'b0 ;
  assign n20292 = n2135 | n9250 ;
  assign n20293 = ( x34 & n809 ) | ( x34 & ~n9990 ) | ( n809 & ~n9990 ) ;
  assign n20294 = n5197 | n20293 ;
  assign n20295 = ~n9446 & n11068 ;
  assign n20299 = n15325 ^ n2267 ^ 1'b0 ;
  assign n20296 = n15507 ^ n7066 ^ 1'b0 ;
  assign n20297 = n1634 & ~n20296 ;
  assign n20298 = ~n15741 & n20297 ;
  assign n20300 = n20299 ^ n20298 ^ 1'b0 ;
  assign n20301 = n1528 & ~n20300 ;
  assign n20302 = n4684 | n11434 ;
  assign n20303 = n16312 & n20302 ;
  assign n20304 = n20303 ^ n16403 ^ 1'b0 ;
  assign n20305 = n1139 & n20304 ;
  assign n20306 = n20305 ^ n1793 ^ 1'b0 ;
  assign n20307 = n18134 ^ n1710 ^ 1'b0 ;
  assign n20308 = n18700 ^ n11709 ^ 1'b0 ;
  assign n20309 = n5398 & n12559 ;
  assign n20310 = n6267 ^ n564 ^ 1'b0 ;
  assign n20311 = n3718 ^ n2706 ^ 1'b0 ;
  assign n20312 = n20310 & n20311 ;
  assign n20313 = n556 & n3368 ;
  assign n20314 = n20313 ^ n1728 ^ 1'b0 ;
  assign n20315 = n20027 ^ n966 ^ 1'b0 ;
  assign n20316 = ~n3314 & n7789 ;
  assign n20317 = n5293 & n11544 ;
  assign n20318 = n2286 & n20317 ;
  assign n20319 = n13800 | n14047 ;
  assign n20320 = ~x21 & n6186 ;
  assign n20321 = n20320 ^ n15429 ^ 1'b0 ;
  assign n20323 = n19805 ^ n9287 ^ 1'b0 ;
  assign n20324 = n399 & ~n20323 ;
  assign n20322 = x153 | n4010 ;
  assign n20325 = n20324 ^ n20322 ^ 1'b0 ;
  assign n20326 = ~n4454 & n13235 ;
  assign n20327 = n20326 ^ n18036 ^ 1'b0 ;
  assign n20328 = n11461 ^ x101 ^ 1'b0 ;
  assign n20329 = n1184 & ~n15088 ;
  assign n20330 = n4595 & ~n16218 ;
  assign n20331 = n7762 ^ n3641 ^ 1'b0 ;
  assign n20332 = n7773 ^ n6490 ^ 1'b0 ;
  assign n20333 = n10192 & n20332 ;
  assign n20334 = ~n2212 & n20333 ;
  assign n20335 = n2034 & ~n15407 ;
  assign n20336 = n5283 & ~n6250 ;
  assign n20337 = ( ~n4660 & n5304 ) | ( ~n4660 & n17539 ) | ( n5304 & n17539 ) ;
  assign n20338 = n20337 ^ n12671 ^ 1'b0 ;
  assign n20339 = ~n2293 & n5475 ;
  assign n20340 = n20339 ^ n2782 ^ 1'b0 ;
  assign n20341 = n9116 & n20340 ;
  assign n20342 = n8508 & n16101 ;
  assign n20343 = n12983 & n20342 ;
  assign n20344 = n13570 ^ n2897 ^ 1'b0 ;
  assign n20345 = n20344 ^ n19089 ^ n11469 ;
  assign n20346 = n3896 & n16152 ;
  assign n20347 = n9011 ^ n5433 ^ 1'b0 ;
  assign n20348 = n10381 & n20347 ;
  assign n20349 = ~n8150 & n14497 ;
  assign n20350 = ~n6198 & n9163 ;
  assign n20351 = n7845 ^ n4172 ^ 1'b0 ;
  assign n20352 = n20351 ^ n7704 ^ 1'b0 ;
  assign n20353 = n5141 & ~n20352 ;
  assign n20354 = n5413 & n20353 ;
  assign n20355 = ~n2164 & n20354 ;
  assign n20356 = n17894 ^ n7241 ^ 1'b0 ;
  assign n20357 = n3964 & ~n20356 ;
  assign n20358 = ( ~n956 & n4857 ) | ( ~n956 & n10141 ) | ( n4857 & n10141 ) ;
  assign n20359 = n871 & n3408 ;
  assign n20360 = n3118 & ~n14451 ;
  assign n20361 = n13679 & n20360 ;
  assign n20362 = n15096 ^ n5500 ^ 1'b0 ;
  assign n20363 = n6797 & n7726 ;
  assign n20364 = n20363 ^ n420 ^ 1'b0 ;
  assign n20365 = n20362 & ~n20364 ;
  assign n20366 = n20365 ^ n13303 ^ 1'b0 ;
  assign n20367 = n20366 ^ n1747 ^ 1'b0 ;
  assign n20368 = n17140 & ~n20367 ;
  assign n20369 = x250 & ~n9280 ;
  assign n20370 = n4548 ^ n2199 ^ n2026 ;
  assign n20371 = n20369 & n20370 ;
  assign n20372 = x93 & n286 ;
  assign n20373 = n787 & ~n3269 ;
  assign n20374 = n20373 ^ n3257 ^ 1'b0 ;
  assign n20375 = n8823 ^ n8675 ^ 1'b0 ;
  assign n20376 = n10041 & ~n20375 ;
  assign n20377 = n19897 | n20376 ;
  assign n20378 = n11481 | n20377 ;
  assign n20379 = n11287 & ~n14635 ;
  assign n20380 = n20379 ^ n9771 ^ 1'b0 ;
  assign n20381 = n552 & ~n11908 ;
  assign n20382 = n20381 ^ n14593 ^ 1'b0 ;
  assign n20383 = n18162 ^ n8888 ^ 1'b0 ;
  assign n20384 = n10525 & n20383 ;
  assign n20385 = n20384 ^ n15445 ^ 1'b0 ;
  assign n20386 = n19674 ^ n14861 ^ 1'b0 ;
  assign n20387 = n8628 & n20386 ;
  assign n20388 = n10996 ^ n1264 ^ 1'b0 ;
  assign n20389 = n10902 & n20388 ;
  assign n20390 = n3112 & ~n10279 ;
  assign n20391 = n736 & n20390 ;
  assign n20392 = n6118 | n19807 ;
  assign n20393 = n3432 & ~n8025 ;
  assign n20394 = n20393 ^ n7362 ^ 1'b0 ;
  assign n20395 = n8963 & ~n12531 ;
  assign n20396 = n20395 ^ n709 ^ 1'b0 ;
  assign n20397 = n3585 & ~n15912 ;
  assign n20398 = n415 & ~n12161 ;
  assign n20399 = n20398 ^ n5852 ^ 1'b0 ;
  assign n20400 = n15878 ^ n2663 ^ 1'b0 ;
  assign n20401 = n17352 | n20400 ;
  assign n20402 = n16085 ^ n4577 ^ 1'b0 ;
  assign n20404 = n18858 ^ n1637 ^ 1'b0 ;
  assign n20405 = n12438 & n20404 ;
  assign n20403 = n8312 & ~n10406 ;
  assign n20406 = n20405 ^ n20403 ^ 1'b0 ;
  assign n20407 = n19722 ^ x111 ^ 1'b0 ;
  assign n20408 = ~n1961 & n20407 ;
  assign n20409 = n9025 ^ n1898 ^ 1'b0 ;
  assign n20410 = ~n11567 & n20409 ;
  assign n20411 = ~n14769 & n20410 ;
  assign n20412 = n1352 ^ x160 ^ 1'b0 ;
  assign n20413 = n3733 & n20412 ;
  assign n20414 = n1118 & n20413 ;
  assign n20415 = n8397 & ~n20414 ;
  assign n20416 = ~x199 & n20415 ;
  assign n20417 = n19856 ^ n5452 ^ 1'b0 ;
  assign n20418 = n1421 | n20417 ;
  assign n20419 = n1758 & n9976 ;
  assign n20420 = n20419 ^ n2632 ^ 1'b0 ;
  assign n20421 = n7068 | n16127 ;
  assign n20422 = n20421 ^ n17294 ^ 1'b0 ;
  assign n20423 = n2689 & n10767 ;
  assign n20424 = ~n5310 & n8027 ;
  assign n20425 = n20424 ^ n10039 ^ 1'b0 ;
  assign n20426 = n9801 ^ n9267 ^ 1'b0 ;
  assign n20427 = ( n956 & n7749 ) | ( n956 & ~n17445 ) | ( n7749 & ~n17445 ) ;
  assign n20428 = n20427 ^ n4671 ^ 1'b0 ;
  assign n20429 = n11119 | n13286 ;
  assign n20430 = n12504 | n20429 ;
  assign n20431 = n809 & ~n20430 ;
  assign n20432 = n20431 ^ n2394 ^ 1'b0 ;
  assign n20433 = ~n3948 & n20432 ;
  assign n20434 = n4124 ^ n1706 ^ 1'b0 ;
  assign n20435 = ~n6790 & n10840 ;
  assign n20436 = n13145 & n20435 ;
  assign n20437 = n1351 & ~n10886 ;
  assign n20438 = n1427 | n20437 ;
  assign n20439 = n20438 ^ n11356 ^ 1'b0 ;
  assign n20440 = n5484 | n8387 ;
  assign n20441 = n15974 & ~n20440 ;
  assign n20444 = n2082 | n5627 ;
  assign n20445 = n8139 | n20444 ;
  assign n20446 = n20445 ^ n16375 ^ 1'b0 ;
  assign n20447 = n1071 & ~n20446 ;
  assign n20442 = n478 | n12536 ;
  assign n20443 = n8445 & ~n20442 ;
  assign n20448 = n20447 ^ n20443 ^ 1'b0 ;
  assign n20449 = n16246 | n17906 ;
  assign n20450 = n20449 ^ n10751 ^ 1'b0 ;
  assign n20451 = n9174 ^ n1967 ^ 1'b0 ;
  assign n20452 = n2883 & ~n20451 ;
  assign n20453 = n11740 ^ n9290 ^ 1'b0 ;
  assign n20454 = n6694 & n19007 ;
  assign n20455 = n2296 & n13062 ;
  assign n20456 = n20455 ^ n7544 ^ 1'b0 ;
  assign n20457 = n4232 | n5897 ;
  assign n20458 = n14922 ^ n10877 ^ 1'b0 ;
  assign n20459 = n13372 ^ n10123 ^ 1'b0 ;
  assign n20460 = n12793 | n20166 ;
  assign n20462 = ~n12763 & n14845 ;
  assign n20463 = ~n4500 & n20462 ;
  assign n20461 = n6553 & ~n14045 ;
  assign n20464 = n20463 ^ n20461 ^ 1'b0 ;
  assign n20465 = ~n1745 & n14407 ;
  assign n20466 = n20465 ^ n15317 ^ 1'b0 ;
  assign n20467 = n19036 ^ n3143 ^ 1'b0 ;
  assign n20468 = n2593 & n20467 ;
  assign n20469 = n10334 ^ n2403 ^ 1'b0 ;
  assign n20470 = n15945 & n20469 ;
  assign n20471 = ~n918 & n1344 ;
  assign n20472 = n7428 & n10908 ;
  assign n20473 = ~n1404 & n4293 ;
  assign n20474 = n20473 ^ x134 ^ 1'b0 ;
  assign n20475 = n9974 | n20474 ;
  assign n20476 = ~n4496 & n20475 ;
  assign n20477 = n20476 ^ n1694 ^ 1'b0 ;
  assign n20478 = ~n13705 & n20477 ;
  assign n20479 = ~n13761 & n20478 ;
  assign n20480 = n351 | n6625 ;
  assign n20481 = n5692 | n9867 ;
  assign n20482 = n17304 | n20481 ;
  assign n20483 = n6570 & n13868 ;
  assign n20484 = n3532 | n9420 ;
  assign n20485 = n614 & ~n20484 ;
  assign n20486 = n6085 | n20485 ;
  assign n20487 = x188 & n20486 ;
  assign n20488 = ~n2185 & n20487 ;
  assign n20489 = n2858 ^ x11 ^ 1'b0 ;
  assign n20490 = n17821 & ~n20489 ;
  assign n20491 = n5676 ^ n5485 ^ 1'b0 ;
  assign n20492 = n20491 ^ n8816 ^ 1'b0 ;
  assign n20493 = n17895 | n20492 ;
  assign n20494 = ~n6401 & n7220 ;
  assign n20495 = n502 & n17119 ;
  assign n20496 = n20495 ^ n8992 ^ 1'b0 ;
  assign n20497 = n20496 ^ n5457 ^ 1'b0 ;
  assign n20498 = n5440 ^ n4354 ^ n366 ;
  assign n20499 = n3343 & ~n20498 ;
  assign n20500 = n1696 & n4741 ;
  assign n20501 = ~n15396 & n20500 ;
  assign n20502 = n17172 ^ n2333 ^ 1'b0 ;
  assign n20503 = n10599 | n20502 ;
  assign n20504 = n5056 | n5690 ;
  assign n20505 = n20504 ^ n3744 ^ 1'b0 ;
  assign n20506 = n20505 ^ n15416 ^ n8351 ;
  assign n20507 = n4149 | n20506 ;
  assign n20508 = n20507 ^ n9954 ^ 1'b0 ;
  assign n20509 = n4302 & n16621 ;
  assign n20510 = n12204 ^ n8223 ^ 1'b0 ;
  assign n20511 = ~n20509 & n20510 ;
  assign n20512 = n1304 & n15447 ;
  assign n20515 = n2295 ^ n669 ^ 1'b0 ;
  assign n20513 = ~n9142 & n14493 ;
  assign n20514 = ~n15912 & n20513 ;
  assign n20516 = n20515 ^ n20514 ^ 1'b0 ;
  assign n20517 = n2650 ^ n2099 ^ 1'b0 ;
  assign n20518 = ~n3521 & n20517 ;
  assign n20519 = n20518 ^ n3383 ^ 1'b0 ;
  assign n20520 = n20519 ^ n13133 ^ 1'b0 ;
  assign n20521 = n3476 & n20520 ;
  assign n20522 = n4294 & n20521 ;
  assign n20523 = n16144 & n20522 ;
  assign n20524 = n19601 & n20523 ;
  assign n20525 = n11744 & n16463 ;
  assign n20526 = x186 & ~n6031 ;
  assign n20527 = n5357 & ~n9210 ;
  assign n20528 = n20526 | n20527 ;
  assign n20529 = n6065 & ~n20528 ;
  assign n20530 = n3117 | n12893 ;
  assign n20531 = n7252 & ~n20530 ;
  assign n20532 = n4848 | n10394 ;
  assign n20533 = n17486 ^ n16736 ^ 1'b0 ;
  assign n20534 = n12860 | n20189 ;
  assign n20535 = n1023 & n8864 ;
  assign n20536 = n476 | n20535 ;
  assign n20537 = n20535 & ~n20536 ;
  assign n20538 = n1012 & ~n5643 ;
  assign n20539 = ~n20537 & n20538 ;
  assign n20540 = ~n5712 & n20539 ;
  assign n20541 = ~n1544 & n4367 ;
  assign n20542 = n1544 & n20541 ;
  assign n20543 = n8827 | n20542 ;
  assign n20544 = n8827 & ~n20543 ;
  assign n20545 = n6551 & n11816 ;
  assign n20546 = ~n11816 & n20545 ;
  assign n20547 = ~n16973 & n20546 ;
  assign n20548 = n20547 ^ n6744 ^ 1'b0 ;
  assign n20549 = ~n20544 & n20548 ;
  assign n20550 = ~n20151 & n20549 ;
  assign n20551 = n20540 & n20550 ;
  assign n20552 = ~n10024 & n16175 ;
  assign n20553 = n20552 ^ n7604 ^ 1'b0 ;
  assign n20554 = n3333 ^ n1104 ^ 1'b0 ;
  assign n20555 = n8827 | n20554 ;
  assign n20556 = n887 & ~n20555 ;
  assign n20557 = n4370 | n4451 ;
  assign n20558 = n15393 & ~n20557 ;
  assign n20559 = n20558 ^ n19197 ^ 1'b0 ;
  assign n20560 = n1162 & n10221 ;
  assign n20561 = n20560 ^ n12583 ^ 1'b0 ;
  assign n20562 = n11573 & ~n20561 ;
  assign n20563 = n7732 ^ n3028 ^ 1'b0 ;
  assign n20564 = n18180 & ~n20563 ;
  assign n20565 = n19564 & n20564 ;
  assign n20566 = n1782 & n3116 ;
  assign n20567 = n12675 ^ n11453 ^ 1'b0 ;
  assign n20568 = n16312 & n20567 ;
  assign n20569 = n19814 ^ n14122 ^ 1'b0 ;
  assign n20570 = n2127 & ~n9312 ;
  assign n20571 = n20570 ^ n1775 ^ 1'b0 ;
  assign n20572 = ~n12470 & n20571 ;
  assign n20573 = n20572 ^ n19030 ^ 1'b0 ;
  assign n20574 = n11346 & n20573 ;
  assign n20575 = n17488 ^ n5818 ^ 1'b0 ;
  assign n20576 = x122 & ~n20575 ;
  assign n20577 = ~n3343 & n18284 ;
  assign n20578 = n19625 & n20577 ;
  assign n20579 = ~n13403 & n15494 ;
  assign n20580 = ~n15781 & n20579 ;
  assign n20581 = ~n989 & n11689 ;
  assign n20582 = n509 & n20581 ;
  assign n20583 = n18123 ^ n5720 ^ 1'b0 ;
  assign n20584 = n20582 & n20583 ;
  assign n20585 = ( n894 & n6597 ) | ( n894 & ~n18157 ) | ( n6597 & ~n18157 ) ;
  assign n20586 = n9203 & n16911 ;
  assign n20587 = ~x155 & n20586 ;
  assign n20588 = n12848 | n20587 ;
  assign n20589 = n16648 ^ n8548 ^ 1'b0 ;
  assign n20590 = n1217 & ~n9165 ;
  assign n20591 = n20590 ^ n11873 ^ 1'b0 ;
  assign n20592 = n8750 ^ n1521 ^ 1'b0 ;
  assign n20593 = n11893 ^ n2743 ^ n2307 ;
  assign n20594 = n20592 | n20593 ;
  assign n20595 = n11928 ^ x115 ^ 1'b0 ;
  assign n20596 = n966 & ~n20595 ;
  assign n20597 = n7020 ^ n6647 ^ 1'b0 ;
  assign n20598 = ~n13830 & n19505 ;
  assign n20599 = ~n4833 & n20598 ;
  assign n20600 = ~n3516 & n19305 ;
  assign n20601 = ~n11295 & n20600 ;
  assign n20602 = n9234 | n20601 ;
  assign n20604 = n4185 & n8820 ;
  assign n20605 = n20604 ^ n8484 ^ 1'b0 ;
  assign n20606 = n20605 ^ n732 ^ 1'b0 ;
  assign n20603 = x100 & ~n7652 ;
  assign n20607 = n20606 ^ n20603 ^ 1'b0 ;
  assign n20608 = n10039 ^ n1159 ^ 1'b0 ;
  assign n20609 = n17218 ^ x98 ^ 1'b0 ;
  assign n20610 = n1678 & n19303 ;
  assign n20611 = n20610 ^ n17689 ^ 1'b0 ;
  assign n20612 = n14375 ^ n444 ^ 1'b0 ;
  assign n20613 = n12972 & n14348 ;
  assign n20615 = n1291 | n5447 ;
  assign n20614 = x24 & n14135 ;
  assign n20616 = n20615 ^ n20614 ^ 1'b0 ;
  assign n20617 = x182 | n20616 ;
  assign n20618 = n20206 ^ n5171 ^ 1'b0 ;
  assign n20619 = n1944 & n20618 ;
  assign n20620 = n19141 ^ n14589 ^ 1'b0 ;
  assign n20621 = n15411 & ~n20620 ;
  assign n20622 = n2517 & n20621 ;
  assign n20623 = n8933 ^ n2855 ^ 1'b0 ;
  assign n20624 = n14069 ^ n5619 ^ 1'b0 ;
  assign n20625 = n1679 & n3140 ;
  assign n20626 = ~n452 & n20625 ;
  assign n20627 = n5650 & ~n20626 ;
  assign n20628 = ~n8686 & n20627 ;
  assign n20629 = x182 | n6985 ;
  assign n20630 = n9256 & ~n11171 ;
  assign n20631 = x138 & n6281 ;
  assign n20632 = n20631 ^ n14214 ^ 1'b0 ;
  assign n20633 = n625 | n1632 ;
  assign n20634 = n625 & ~n20633 ;
  assign n20635 = n11731 & ~n20634 ;
  assign n20636 = n20635 ^ n10136 ^ 1'b0 ;
  assign n20637 = n17020 ^ n12385 ^ 1'b0 ;
  assign n20638 = n12849 & n20637 ;
  assign n20639 = n18800 ^ n6874 ^ n4222 ;
  assign n20640 = n5006 & n14598 ;
  assign n20641 = ~n10844 & n20640 ;
  assign n20642 = n16424 & ~n17010 ;
  assign n20643 = n14580 ^ n1619 ^ 1'b0 ;
  assign n20644 = ~n4955 & n20643 ;
  assign n20645 = ~n5895 & n20644 ;
  assign n20646 = n20645 ^ n11968 ^ 1'b0 ;
  assign n20647 = n512 | n4396 ;
  assign n20648 = ~n15582 & n20647 ;
  assign n20649 = n10469 | n12509 ;
  assign n20650 = x173 & ~n10623 ;
  assign n20651 = ( n5707 & n10077 ) | ( n5707 & n16401 ) | ( n10077 & n16401 ) ;
  assign n20652 = n20651 ^ n14972 ^ 1'b0 ;
  assign n20653 = n11891 & n20652 ;
  assign n20654 = n20653 ^ n7400 ^ 1'b0 ;
  assign n20655 = n20650 & n20654 ;
  assign n20656 = n6663 ^ n6267 ^ 1'b0 ;
  assign n20657 = n9568 & n20656 ;
  assign n20658 = n3107 | n5207 ;
  assign n20659 = n10997 & ~n20658 ;
  assign n20660 = n7430 & ~n7839 ;
  assign n20661 = n20659 & n20660 ;
  assign n20662 = n12412 & n20661 ;
  assign n20663 = n5408 | n10950 ;
  assign n20664 = n7076 & n11992 ;
  assign n20672 = n273 | n1160 ;
  assign n20668 = n1564 & n7475 ;
  assign n20669 = n20668 ^ n8718 ^ 1'b0 ;
  assign n20670 = n10300 & n20669 ;
  assign n20671 = n20670 ^ n10725 ^ 1'b0 ;
  assign n20673 = n20672 ^ n20671 ^ 1'b0 ;
  assign n20674 = ~n2868 & n20673 ;
  assign n20675 = n18088 & n20674 ;
  assign n20665 = n955 & ~n5788 ;
  assign n20666 = ~n9717 & n20665 ;
  assign n20667 = x200 | n20666 ;
  assign n20676 = n20675 ^ n20667 ^ 1'b0 ;
  assign n20677 = ( n3102 & ~n7779 ) | ( n3102 & n20676 ) | ( ~n7779 & n20676 ) ;
  assign n20678 = n4063 | n12882 ;
  assign n20679 = n2990 | n20678 ;
  assign n20680 = n16636 ^ n8969 ^ 1'b0 ;
  assign n20681 = n20556 | n20680 ;
  assign n20682 = n6355 & n19508 ;
  assign n20683 = ~n16754 & n20682 ;
  assign n20684 = n20683 ^ n1697 ^ 1'b0 ;
  assign n20685 = n2357 & n7197 ;
  assign n20686 = n5821 & n20685 ;
  assign n20687 = n20686 ^ n7069 ^ 1'b0 ;
  assign n20688 = n3633 ^ n3210 ^ 1'b0 ;
  assign n20689 = n14103 | n18541 ;
  assign n20690 = n4389 | n8127 ;
  assign n20691 = n13109 & n20690 ;
  assign n20692 = n13101 ^ n10108 ^ 1'b0 ;
  assign n20693 = n3562 & n20692 ;
  assign n20694 = n20693 ^ n17521 ^ 1'b0 ;
  assign n20695 = n3477 | n16357 ;
  assign n20696 = x219 & n20695 ;
  assign n20697 = n20696 ^ n809 ^ 1'b0 ;
  assign n20698 = n2221 & ~n20697 ;
  assign n20699 = ~n12251 & n20698 ;
  assign n20700 = x81 & ~n11792 ;
  assign n20701 = n15011 ^ n1410 ^ 1'b0 ;
  assign n20702 = n5350 & n6266 ;
  assign n20703 = ~n5883 & n9226 ;
  assign n20704 = n14799 ^ n12872 ^ 1'b0 ;
  assign n20705 = n9309 ^ n8681 ^ 1'b0 ;
  assign n20706 = n8560 ^ n3263 ^ 1'b0 ;
  assign n20707 = n20705 | n20706 ;
  assign n20708 = n9713 ^ n9539 ^ 1'b0 ;
  assign n20709 = n3446 | n20708 ;
  assign n20710 = n20709 ^ n2135 ^ 1'b0 ;
  assign n20711 = n17713 ^ n2296 ^ 1'b0 ;
  assign n20712 = ~n4175 & n20711 ;
  assign n20713 = ~n11705 & n16308 ;
  assign n20714 = n2597 & ~n7444 ;
  assign n20715 = ( n8092 & n11650 ) | ( n8092 & n20714 ) | ( n11650 & n20714 ) ;
  assign n20716 = n19940 & ~n20715 ;
  assign n20719 = x170 & ~n13539 ;
  assign n20720 = n20719 ^ n8722 ^ 1'b0 ;
  assign n20717 = n10218 ^ n3030 ^ 1'b0 ;
  assign n20718 = n10048 & ~n20717 ;
  assign n20721 = n20720 ^ n20718 ^ 1'b0 ;
  assign n20722 = n5004 & n8811 ;
  assign n20723 = n10555 | n20722 ;
  assign n20724 = n12519 | n20723 ;
  assign n20725 = n20724 ^ n5433 ^ 1'b0 ;
  assign n20726 = n20725 ^ n8474 ^ 1'b0 ;
  assign n20727 = n6243 & n20726 ;
  assign n20728 = n5702 | n14355 ;
  assign n20729 = n10972 | n20728 ;
  assign n20730 = n20729 ^ n327 ^ 1'b0 ;
  assign n20731 = n20727 | n20730 ;
  assign n20732 = n10092 | n11964 ;
  assign n20733 = n20732 ^ n12697 ^ n8097 ;
  assign n20734 = n17751 ^ n9109 ^ 1'b0 ;
  assign n20735 = ~n4119 & n12891 ;
  assign n20736 = n2627 & ~n3971 ;
  assign n20737 = ~n5287 & n20736 ;
  assign n20738 = x151 | n20737 ;
  assign n20739 = ~n959 & n9688 ;
  assign n20740 = n20738 & n20739 ;
  assign n20741 = n13157 & n20194 ;
  assign n20742 = n15101 ^ n5420 ^ n552 ;
  assign n20743 = n20742 ^ n14882 ^ n3065 ;
  assign n20744 = ~n5875 & n9256 ;
  assign n20745 = n20744 ^ n19107 ^ 1'b0 ;
  assign n20746 = n2897 & n3556 ;
  assign n20747 = n17109 & n20746 ;
  assign n20748 = n20232 ^ n4791 ^ 1'b0 ;
  assign n20749 = n8558 | n11176 ;
  assign n20750 = n955 & n20749 ;
  assign n20751 = n20750 ^ n2338 ^ 1'b0 ;
  assign n20752 = ~n1955 & n7500 ;
  assign n20753 = n20752 ^ n15731 ^ 1'b0 ;
  assign n20754 = n20751 | n20753 ;
  assign n20755 = n18289 ^ n9620 ^ 1'b0 ;
  assign n20756 = ~n4580 & n5344 ;
  assign n20757 = n20756 ^ n6468 ^ 1'b0 ;
  assign n20758 = n2310 & ~n5399 ;
  assign n20759 = ~n17984 & n20758 ;
  assign n20760 = ( n10968 & n18119 ) | ( n10968 & n20627 ) | ( n18119 & n20627 ) ;
  assign n20761 = n2707 | n18437 ;
  assign n20762 = n1529 & ~n4627 ;
  assign n20763 = ~n9815 & n20762 ;
  assign n20764 = n5694 & ~n20763 ;
  assign n20765 = n1275 & ~n12594 ;
  assign n20766 = ~n1275 & n20765 ;
  assign n20767 = n20764 | n20766 ;
  assign n20768 = n1299 | n20767 ;
  assign n20769 = n4769 & ~n5452 ;
  assign n20770 = n10198 ^ n8024 ^ 1'b0 ;
  assign n20771 = n8541 & n20770 ;
  assign n20772 = n20771 ^ n17344 ^ 1'b0 ;
  assign n20773 = n602 & n3069 ;
  assign n20774 = ~n1646 & n3754 ;
  assign n20775 = n20773 | n20774 ;
  assign n20776 = n1368 & ~n7339 ;
  assign n20777 = n3447 & ~n7710 ;
  assign n20778 = ~n20776 & n20777 ;
  assign n20779 = n357 | n20778 ;
  assign n20780 = n20779 ^ n3452 ^ 1'b0 ;
  assign n20781 = n2279 ^ n2085 ^ n551 ;
  assign n20782 = x25 | n20781 ;
  assign n20783 = n20780 | n20782 ;
  assign n20784 = n7832 ^ n1810 ^ 1'b0 ;
  assign n20785 = n16368 & n20784 ;
  assign n20786 = n19985 ^ n8029 ^ 1'b0 ;
  assign n20787 = n3862 & n14981 ;
  assign n20788 = n18800 ^ n4608 ^ 1'b0 ;
  assign n20789 = ~n950 & n15842 ;
  assign n20790 = ~n9012 & n20789 ;
  assign n20791 = n11891 | n20790 ;
  assign n20792 = ~n2712 & n5197 ;
  assign n20793 = n2828 & n4154 ;
  assign n20794 = n20793 ^ n7800 ^ 1'b0 ;
  assign n20795 = n18640 ^ n3442 ^ 1'b0 ;
  assign n20796 = n8835 & n20795 ;
  assign n20797 = n8530 & ~n14007 ;
  assign n20798 = n20797 ^ n20772 ^ 1'b0 ;
  assign n20799 = n2749 | n20798 ;
  assign n20800 = n16032 ^ n14023 ^ 1'b0 ;
  assign n20801 = n6884 & n19007 ;
  assign n20802 = n20801 ^ n18086 ^ 1'b0 ;
  assign n20803 = n7039 & n7331 ;
  assign n20804 = n20802 & n20803 ;
  assign n20805 = n9660 ^ n797 ^ 1'b0 ;
  assign n20806 = ~n6900 & n11394 ;
  assign n20807 = n5955 & n9385 ;
  assign n20808 = n17706 & n20807 ;
  assign n20809 = ~n2768 & n5823 ;
  assign n20810 = ~n1184 & n5573 ;
  assign n20811 = n20810 ^ n18063 ^ 1'b0 ;
  assign n20812 = n20811 ^ n15401 ^ 1'b0 ;
  assign n20813 = n1843 & n20812 ;
  assign n20814 = n12762 ^ n10118 ^ 1'b0 ;
  assign n20815 = ~n14993 & n20814 ;
  assign n20816 = ~n5128 & n6817 ;
  assign n20817 = n20816 ^ n1240 ^ 1'b0 ;
  assign n20818 = ~n8470 & n10488 ;
  assign n20819 = n17150 ^ n3485 ^ 1'b0 ;
  assign n20820 = n3751 | n4423 ;
  assign n20821 = n20820 ^ n5809 ^ 1'b0 ;
  assign n20822 = n20819 | n20821 ;
  assign n20823 = n1139 & n6693 ;
  assign n20824 = n6247 & n20823 ;
  assign n20825 = x43 & n4340 ;
  assign n20826 = n5877 & ~n20825 ;
  assign n20827 = n20824 & n20826 ;
  assign n20828 = n18353 ^ n4799 ^ 1'b0 ;
  assign n20829 = n4573 | n20828 ;
  assign n20830 = ( n923 & n2037 ) | ( n923 & ~n12627 ) | ( n2037 & ~n12627 ) ;
  assign n20831 = n6198 ^ n2505 ^ 1'b0 ;
  assign n20832 = n10004 | n20831 ;
  assign n20833 = n2325 ^ n1267 ^ 1'b0 ;
  assign n20834 = n20832 | n20833 ;
  assign n20836 = n15193 ^ n7670 ^ 1'b0 ;
  assign n20835 = n5100 ^ n800 ^ 1'b0 ;
  assign n20837 = n20836 ^ n20835 ^ n3125 ;
  assign n20838 = n772 & n20837 ;
  assign n20839 = x65 & n4944 ;
  assign n20843 = n6876 & n14060 ;
  assign n20844 = n271 & n20843 ;
  assign n20840 = n6416 & ~n18954 ;
  assign n20841 = ~n9449 & n20840 ;
  assign n20842 = n6629 & n20841 ;
  assign n20845 = n20844 ^ n20842 ^ 1'b0 ;
  assign n20846 = n10385 ^ n3226 ^ 1'b0 ;
  assign n20847 = n8608 & n20846 ;
  assign n20848 = ~n14005 & n20847 ;
  assign n20849 = n12151 ^ n3181 ^ 1'b0 ;
  assign n20850 = n9607 & n20849 ;
  assign n20851 = n16681 ^ n12080 ^ n9503 ;
  assign n20852 = n327 | n1272 ;
  assign n20853 = n327 & ~n20852 ;
  assign n20854 = n3153 | n20853 ;
  assign n20855 = n1112 & n13044 ;
  assign n20856 = n20854 | n20855 ;
  assign n20857 = n10658 & ~n20856 ;
  assign n20858 = n11235 ^ n5633 ^ 1'b0 ;
  assign n20862 = n6700 ^ n4049 ^ 1'b0 ;
  assign n20859 = n11165 ^ n327 ^ 1'b0 ;
  assign n20860 = n20859 ^ n265 ^ 1'b0 ;
  assign n20861 = ~n7544 & n20860 ;
  assign n20863 = n20862 ^ n20861 ^ n6747 ;
  assign n20864 = n4144 ^ n4101 ^ 1'b0 ;
  assign n20865 = n7395 & n11435 ;
  assign n20866 = n851 & n20865 ;
  assign n20867 = n10024 ^ n7392 ^ n337 ;
  assign n20868 = ~n1061 & n20867 ;
  assign n20869 = n20868 ^ n3745 ^ 1'b0 ;
  assign n20870 = x157 & n15071 ;
  assign n20872 = n395 | n871 ;
  assign n20873 = n20872 ^ x187 ^ 1'b0 ;
  assign n20871 = n5691 | n11972 ;
  assign n20874 = n20873 ^ n20871 ^ n1845 ;
  assign n20875 = n11613 ^ n1857 ^ 1'b0 ;
  assign n20876 = n1641 & n20875 ;
  assign n20877 = ~n800 & n1608 ;
  assign n20882 = ~n1291 & n14323 ;
  assign n20878 = n872 & ~n8674 ;
  assign n20879 = n4154 & n20878 ;
  assign n20880 = n12795 & ~n20879 ;
  assign n20881 = ~x130 & n20880 ;
  assign n20883 = n20882 ^ n20881 ^ 1'b0 ;
  assign n20884 = n6031 ^ n1077 ^ 1'b0 ;
  assign n20885 = n9239 ^ n6938 ^ 1'b0 ;
  assign n20886 = n2828 & ~n6961 ;
  assign n20887 = n9067 & n20886 ;
  assign n20888 = n15361 | n20887 ;
  assign n20889 = n11322 ^ x3 ^ 1'b0 ;
  assign n20890 = n860 & ~n5034 ;
  assign n20891 = n5851 & n20890 ;
  assign n20892 = n4370 ^ n2689 ^ 1'b0 ;
  assign n20893 = n20892 ^ n7371 ^ 1'b0 ;
  assign n20894 = n16952 | n20893 ;
  assign n20895 = n8608 ^ n8128 ^ 1'b0 ;
  assign n20896 = n3924 ^ x61 ^ 1'b0 ;
  assign n20897 = n1819 & ~n19309 ;
  assign n20898 = ~n3272 & n20897 ;
  assign n20899 = n11810 ^ n7437 ^ 1'b0 ;
  assign n20900 = ~n15814 & n20899 ;
  assign n20901 = n397 & n11891 ;
  assign n20902 = n20901 ^ n12804 ^ 1'b0 ;
  assign n20903 = n15780 ^ n3366 ^ n2008 ;
  assign n20904 = n20903 ^ n7189 ^ 1'b0 ;
  assign n20905 = x86 & n20904 ;
  assign n20906 = n19179 & n20905 ;
  assign n20907 = n20906 ^ n13186 ^ 1'b0 ;
  assign n20908 = x112 & n11618 ;
  assign n20909 = n4389 ^ n3637 ^ 1'b0 ;
  assign n20910 = n18949 ^ n2557 ^ 1'b0 ;
  assign n20911 = ~n20909 & n20910 ;
  assign n20912 = n672 & n14392 ;
  assign n20913 = n20912 ^ n15565 ^ 1'b0 ;
  assign n20914 = n17614 | n20913 ;
  assign n20917 = ( n2393 & ~n2793 ) | ( n2393 & n5286 ) | ( ~n2793 & n5286 ) ;
  assign n20918 = n20917 ^ n9964 ^ 1'b0 ;
  assign n20915 = n8722 ^ n3981 ^ 1'b0 ;
  assign n20916 = n20915 ^ n4390 ^ 1'b0 ;
  assign n20919 = n20918 ^ n20916 ^ 1'b0 ;
  assign n20920 = n15641 ^ n2926 ^ 1'b0 ;
  assign n20921 = n4734 | n18925 ;
  assign n20922 = n5203 & ~n20921 ;
  assign n20923 = n7132 ^ x231 ^ 1'b0 ;
  assign n20924 = n20923 ^ n12765 ^ 1'b0 ;
  assign n20926 = x152 & ~n14102 ;
  assign n20925 = ~n13169 & n18428 ;
  assign n20927 = n20926 ^ n20925 ^ 1'b0 ;
  assign n20928 = ~n955 & n18956 ;
  assign n20929 = n3167 & ~n20928 ;
  assign n20930 = n2632 | n15744 ;
  assign n20931 = n20930 ^ n9576 ^ 1'b0 ;
  assign n20932 = n6524 & n20931 ;
  assign n20933 = ~n14524 & n20932 ;
  assign n20934 = n5781 ^ n5620 ^ n482 ;
  assign n20935 = n1286 | n7062 ;
  assign n20936 = n1451 & ~n20935 ;
  assign n20937 = n5475 & n20936 ;
  assign n20938 = n2368 ^ x121 ^ 1'b0 ;
  assign n20939 = n6125 ^ n2076 ^ 1'b0 ;
  assign n20940 = ~n20217 & n20939 ;
  assign n20941 = n12126 & n20940 ;
  assign n20942 = n395 | n20941 ;
  assign n20945 = n271 & n967 ;
  assign n20946 = n20945 ^ n8406 ^ 1'b0 ;
  assign n20943 = n17631 ^ n5896 ^ 1'b0 ;
  assign n20944 = x53 & n20943 ;
  assign n20947 = n20946 ^ n20944 ^ 1'b0 ;
  assign n20948 = n11720 & ~n20947 ;
  assign n20949 = n6882 & n6963 ;
  assign n20950 = n20949 ^ n2769 ^ 1'b0 ;
  assign n20951 = n5283 ^ n1709 ^ 1'b0 ;
  assign n20952 = n8642 ^ n7047 ^ 1'b0 ;
  assign n20953 = n11329 ^ x110 ^ 1'b0 ;
  assign n20954 = ~n10150 & n20953 ;
  assign n20955 = n8742 & n20954 ;
  assign n20956 = n11356 & n20955 ;
  assign n20957 = ( ~n10626 & n11502 ) | ( ~n10626 & n20956 ) | ( n11502 & n20956 ) ;
  assign n20958 = n17633 ^ n12192 ^ 1'b0 ;
  assign n20959 = n16780 & ~n17340 ;
  assign n20960 = n620 & n5672 ;
  assign n20961 = n20960 ^ n630 ^ 1'b0 ;
  assign n20962 = x230 & ~n20961 ;
  assign n20963 = n20962 ^ n4554 ^ 1'b0 ;
  assign n20964 = n1442 & ~n20963 ;
  assign n20965 = ~n5068 & n5159 ;
  assign n20966 = n10332 & ~n20965 ;
  assign n20967 = n8646 ^ n2670 ^ 1'b0 ;
  assign n20968 = ~x178 & n20967 ;
  assign n20969 = ~n6089 & n15928 ;
  assign n20970 = n5748 & ~n12136 ;
  assign n20971 = n20970 ^ n3790 ^ 1'b0 ;
  assign n20972 = n4515 | n14694 ;
  assign n20973 = n13669 & ~n20972 ;
  assign n20974 = ~n2955 & n12785 ;
  assign n20975 = n14647 & n20974 ;
  assign n20976 = ~n5072 & n20975 ;
  assign n20977 = ~n10394 & n10780 ;
  assign n20978 = n20650 ^ n15507 ^ 1'b0 ;
  assign n20979 = n1926 | n20978 ;
  assign n20982 = n7792 ^ n4888 ^ 1'b0 ;
  assign n20983 = n20982 ^ n3308 ^ 1'b0 ;
  assign n20980 = n7474 ^ n288 ^ 1'b0 ;
  assign n20981 = n9495 & n20980 ;
  assign n20984 = n20983 ^ n20981 ^ 1'b0 ;
  assign n20985 = ~n430 & n11938 ;
  assign n20986 = n20985 ^ n7526 ^ 1'b0 ;
  assign n20987 = n20982 & ~n20986 ;
  assign n20988 = n3239 & n7098 ;
  assign n20989 = n10563 | n20988 ;
  assign n20990 = n16861 & ~n20989 ;
  assign n20991 = n4084 & ~n4720 ;
  assign n20992 = n14106 ^ x77 ^ 1'b0 ;
  assign n20993 = n20992 ^ n7971 ^ 1'b0 ;
  assign n20994 = n20993 ^ n20153 ^ 1'b0 ;
  assign n20995 = x252 & ~n7868 ;
  assign n20996 = ~x76 & n20995 ;
  assign n20997 = n20996 ^ n5950 ^ 1'b0 ;
  assign n20998 = n2593 & ~n7864 ;
  assign n20999 = n16608 ^ n666 ^ 1'b0 ;
  assign n21002 = n2764 & ~n11891 ;
  assign n21003 = n21002 ^ x250 ^ 1'b0 ;
  assign n21004 = n4409 & ~n21003 ;
  assign n21000 = n6421 ^ n4276 ^ 1'b0 ;
  assign n21001 = ~n7883 & n21000 ;
  assign n21005 = n21004 ^ n21001 ^ 1'b0 ;
  assign n21006 = n7748 ^ n1116 ^ 1'b0 ;
  assign n21007 = n12805 ^ n10016 ^ 1'b0 ;
  assign n21008 = n10993 & n21007 ;
  assign n21009 = n8611 & ~n14422 ;
  assign n21010 = n21009 ^ n3548 ^ 1'b0 ;
  assign n21011 = n298 | n1625 ;
  assign n21012 = n21011 ^ n8644 ^ 1'b0 ;
  assign n21013 = n10988 & ~n21012 ;
  assign n21014 = n7569 ^ n5195 ^ 1'b0 ;
  assign n21015 = n354 & n21014 ;
  assign n21016 = n21015 ^ n12161 ^ 1'b0 ;
  assign n21017 = n3994 & n21016 ;
  assign n21018 = n3814 | n4104 ;
  assign n21019 = n2500 & ~n4606 ;
  assign n21020 = n21019 ^ n3911 ^ 1'b0 ;
  assign n21021 = n6427 ^ n4119 ^ 1'b0 ;
  assign n21022 = n3217 & ~n21021 ;
  assign n21023 = n4328 & ~n16656 ;
  assign n21024 = ~n21022 & n21023 ;
  assign n21025 = ~n16130 & n21024 ;
  assign n21026 = n9830 | n19976 ;
  assign n21027 = n6966 & ~n9407 ;
  assign n21028 = n21027 ^ n13053 ^ 1'b0 ;
  assign n21029 = ~n21026 & n21028 ;
  assign n21030 = ~n5798 & n6507 ;
  assign n21031 = n21030 ^ n13001 ^ n2183 ;
  assign n21032 = n16612 ^ n3336 ^ 1'b0 ;
  assign n21033 = n12498 ^ n1873 ^ 1'b0 ;
  assign n21034 = n5382 & ~n12795 ;
  assign n21035 = n16362 | n19728 ;
  assign n21036 = n21035 ^ n7925 ^ 1'b0 ;
  assign n21040 = x172 & n3174 ;
  assign n21037 = n4119 & n16150 ;
  assign n21038 = n21037 ^ x245 ^ 1'b0 ;
  assign n21039 = n6478 & n21038 ;
  assign n21041 = n21040 ^ n21039 ^ 1'b0 ;
  assign n21042 = ~n1680 & n1845 ;
  assign n21043 = n21042 ^ n14379 ^ 1'b0 ;
  assign n21044 = ( n919 & ~n6450 ) | ( n919 & n21043 ) | ( ~n6450 & n21043 ) ;
  assign n21045 = n4370 & ~n18833 ;
  assign n21046 = ~n8205 & n13102 ;
  assign n21047 = ~n13192 & n21046 ;
  assign n21048 = n3003 & n3913 ;
  assign n21049 = n21047 & n21048 ;
  assign n21050 = n6972 & n20898 ;
  assign n21051 = n8170 & ~n17268 ;
  assign n21052 = n1613 & n21051 ;
  assign n21053 = ~n6647 & n8228 ;
  assign n21054 = ~n786 & n21053 ;
  assign n21055 = n6403 & ~n9186 ;
  assign n21056 = n11158 & ~n19424 ;
  assign n21057 = ~n9439 & n13820 ;
  assign n21059 = n2035 ^ n354 ^ 1'b0 ;
  assign n21058 = n7400 ^ n6123 ^ 1'b0 ;
  assign n21060 = n21059 ^ n21058 ^ 1'b0 ;
  assign n21061 = ~n19568 & n21060 ;
  assign n21063 = n9380 ^ n2502 ^ 1'b0 ;
  assign n21062 = n2354 & n9940 ;
  assign n21064 = n21063 ^ n21062 ^ 1'b0 ;
  assign n21065 = n2903 | n7410 ;
  assign n21066 = n21065 ^ n12449 ^ 1'b0 ;
  assign n21067 = n21064 | n21066 ;
  assign n21068 = n12527 ^ n3325 ^ 1'b0 ;
  assign n21069 = n3143 & n21068 ;
  assign n21070 = n18900 & n21069 ;
  assign n21071 = ~n21069 & n21070 ;
  assign n21072 = n7940 ^ n6815 ^ 1'b0 ;
  assign n21073 = n16435 & ~n21072 ;
  assign n21074 = n21073 ^ x57 ^ 1'b0 ;
  assign n21075 = n21074 ^ n11339 ^ 1'b0 ;
  assign n21076 = n12395 ^ n1217 ^ 1'b0 ;
  assign n21077 = n10798 & ~n15665 ;
  assign n21078 = n1314 | n7228 ;
  assign n21079 = n5213 & ~n21078 ;
  assign n21080 = n21079 ^ n8608 ^ 1'b0 ;
  assign n21081 = n10408 & n15393 ;
  assign n21082 = n21081 ^ n1499 ^ 1'b0 ;
  assign n21083 = n3970 ^ n2062 ^ 1'b0 ;
  assign n21084 = n20139 ^ n3744 ^ 1'b0 ;
  assign n21085 = ~n5305 & n10800 ;
  assign n21086 = n18611 & n21085 ;
  assign n21087 = ~n1219 & n12519 ;
  assign n21088 = n3755 & n11004 ;
  assign n21089 = ~n355 & n5199 ;
  assign n21090 = ~n2760 & n21089 ;
  assign n21091 = n21090 ^ n19800 ^ 1'b0 ;
  assign n21092 = n4469 & ~n12818 ;
  assign n21093 = ~n21091 & n21092 ;
  assign n21094 = n8008 & n13398 ;
  assign n21095 = n21094 ^ n16470 ^ 1'b0 ;
  assign n21096 = n7533 ^ n5073 ^ 1'b0 ;
  assign n21097 = n21096 ^ n1050 ^ 1'b0 ;
  assign n21098 = n6392 ^ n930 ^ 1'b0 ;
  assign n21099 = n21097 | n21098 ;
  assign n21100 = n21099 ^ n4801 ^ 1'b0 ;
  assign n21101 = n5624 | n7204 ;
  assign n21102 = n1173 | n21101 ;
  assign n21103 = n2110 & n21102 ;
  assign n21104 = n19187 & n21103 ;
  assign n21105 = n3920 & ~n9052 ;
  assign n21106 = ~n956 & n10133 ;
  assign n21107 = ~n10133 & n21106 ;
  assign n21108 = n20705 ^ n2728 ^ 1'b0 ;
  assign n21109 = n8236 | n21108 ;
  assign n21110 = n21109 ^ n17453 ^ 1'b0 ;
  assign n21111 = n21110 ^ n16120 ^ n12859 ;
  assign n21112 = n3126 & ~n9111 ;
  assign n21113 = ~n12893 & n21112 ;
  assign n21114 = n18387 ^ n9266 ^ 1'b0 ;
  assign n21115 = n21113 | n21114 ;
  assign n21116 = n11918 ^ n2842 ^ 1'b0 ;
  assign n21117 = n21116 ^ n1877 ^ 1'b0 ;
  assign n21118 = ( ~n6696 & n8847 ) | ( ~n6696 & n9415 ) | ( n8847 & n9415 ) ;
  assign n21119 = n15241 ^ n5192 ^ 1'b0 ;
  assign n21120 = n18243 & n21119 ;
  assign n21121 = n3397 | n7456 ;
  assign n21122 = n3905 ^ n1093 ^ 1'b0 ;
  assign n21123 = n6034 & ~n8195 ;
  assign n21124 = ~n1602 & n21123 ;
  assign n21125 = n3230 & n3263 ;
  assign n21126 = n8388 & n21125 ;
  assign n21127 = n21124 & n21126 ;
  assign n21128 = n11343 ^ n5679 ^ n486 ;
  assign n21129 = n15138 ^ n9254 ^ 1'b0 ;
  assign n21130 = n4720 | n21129 ;
  assign n21131 = n11565 ^ x123 ^ 1'b0 ;
  assign n21132 = n423 & ~n21131 ;
  assign n21133 = n9143 & n21132 ;
  assign n21134 = n21133 ^ n14842 ^ 1'b0 ;
  assign n21135 = ~n5700 & n10527 ;
  assign n21136 = n8921 & n21135 ;
  assign n21137 = n5931 ^ n1046 ^ 1'b0 ;
  assign n21138 = n13813 ^ n1857 ^ 1'b0 ;
  assign n21139 = n2450 & ~n21138 ;
  assign n21140 = n17846 | n19078 ;
  assign n21141 = ~n5926 & n21140 ;
  assign n21142 = n21141 ^ n10179 ^ 1'b0 ;
  assign n21143 = n10484 ^ n9978 ^ 1'b0 ;
  assign n21144 = n1847 & ~n21143 ;
  assign n21154 = n18716 | n19446 ;
  assign n21153 = n1978 ^ n1111 ^ 1'b0 ;
  assign n21145 = ~n6762 & n15124 ;
  assign n21146 = n1736 & ~n10972 ;
  assign n21147 = n21146 ^ n13914 ^ 1'b0 ;
  assign n21148 = n21145 | n21147 ;
  assign n21149 = n16319 ^ n1499 ^ 1'b0 ;
  assign n21150 = n1967 | n21149 ;
  assign n21151 = n21150 ^ n16499 ^ 1'b0 ;
  assign n21152 = ~n21148 & n21151 ;
  assign n21155 = n21154 ^ n21153 ^ n21152 ;
  assign n21156 = n3017 | n5031 ;
  assign n21157 = n7605 & ~n21156 ;
  assign n21158 = n1499 & ~n14580 ;
  assign n21159 = ~n6381 & n11808 ;
  assign n21160 = ~n2939 & n21159 ;
  assign n21161 = n17111 ^ n15463 ^ 1'b0 ;
  assign n21162 = n21161 ^ n5097 ^ x233 ;
  assign n21163 = n4678 | n7049 ;
  assign n21164 = n8709 | n21163 ;
  assign n21165 = n8553 & ~n13635 ;
  assign n21166 = ~n9739 & n12533 ;
  assign n21167 = n21166 ^ n562 ^ 1'b0 ;
  assign n21168 = x135 & n10039 ;
  assign n21169 = n4737 & ~n7227 ;
  assign n21170 = n21169 ^ n18502 ^ 1'b0 ;
  assign n21171 = n13656 | n21170 ;
  assign n21172 = n1249 & ~n7102 ;
  assign n21173 = n21172 ^ n11241 ^ 1'b0 ;
  assign n21174 = n1622 | n6469 ;
  assign n21175 = n14005 ^ n3879 ^ 1'b0 ;
  assign n21176 = n5484 & ~n12208 ;
  assign n21177 = n21176 ^ n1175 ^ 1'b0 ;
  assign n21178 = n3013 & n12159 ;
  assign n21179 = n4314 | n7111 ;
  assign n21180 = ~n15656 & n15829 ;
  assign n21181 = n9803 | n21180 ;
  assign n21182 = n5670 & n10678 ;
  assign n21183 = n2412 & ~n21182 ;
  assign n21184 = n21183 ^ n9284 ^ 1'b0 ;
  assign n21185 = x226 & ~n10990 ;
  assign n21186 = n884 & n11272 ;
  assign n21187 = n4920 & ~n20183 ;
  assign n21188 = ~n4955 & n11635 ;
  assign n21189 = n19041 ^ n5746 ^ 1'b0 ;
  assign n21190 = n7017 & n12962 ;
  assign n21191 = n21190 ^ n3801 ^ 1'b0 ;
  assign n21192 = n6008 | n21191 ;
  assign n21193 = n21192 ^ n754 ^ 1'b0 ;
  assign n21194 = ~n1507 & n13795 ;
  assign n21195 = ~n1485 & n16449 ;
  assign n21196 = ~n15436 & n21195 ;
  assign n21197 = ( n4118 & ~n9313 ) | ( n4118 & n10612 ) | ( ~n9313 & n10612 ) ;
  assign n21198 = n10240 & n12190 ;
  assign n21199 = n5339 & n7874 ;
  assign n21200 = n780 & n21199 ;
  assign n21201 = n21200 ^ n10082 ^ 1'b0 ;
  assign n21202 = n10016 & ~n21201 ;
  assign n21203 = n5225 ^ n4711 ^ 1'b0 ;
  assign n21204 = ~n3871 & n21203 ;
  assign n21205 = n21204 ^ n14344 ^ 1'b0 ;
  assign n21206 = n11854 ^ n7822 ^ 1'b0 ;
  assign n21207 = n17449 | n21206 ;
  assign n21208 = n3272 | n3381 ;
  assign n21209 = n2443 & n21208 ;
  assign n21210 = n9152 & ~n12636 ;
  assign n21211 = n5152 & n21210 ;
  assign n21212 = n3402 | n21211 ;
  assign n21213 = n15668 & ~n16711 ;
  assign n21214 = ~x191 & n21213 ;
  assign n21215 = n4831 | n5125 ;
  assign n21216 = n2370 | n21215 ;
  assign n21217 = ~n7384 & n12652 ;
  assign n21218 = n21217 ^ n17614 ^ 1'b0 ;
  assign n21219 = n9376 ^ n4949 ^ 1'b0 ;
  assign n21220 = n4006 & ~n21219 ;
  assign n21221 = n19036 ^ n7411 ^ 1'b0 ;
  assign n21222 = n11483 & ~n11566 ;
  assign n21223 = n11252 ^ n3445 ^ 1'b0 ;
  assign n21224 = n20532 | n21223 ;
  assign n21225 = n6471 | n21224 ;
  assign n21226 = n21222 | n21225 ;
  assign n21227 = n9223 | n21226 ;
  assign n21228 = n21221 | n21227 ;
  assign n21229 = n4328 & n17375 ;
  assign n21230 = n21229 ^ n10551 ^ 1'b0 ;
  assign n21231 = n5375 | n21230 ;
  assign n21232 = n3283 ^ x227 ^ 1'b0 ;
  assign n21233 = n3619 & n21232 ;
  assign n21234 = n261 | n11514 ;
  assign n21235 = n21234 ^ n1587 ^ 1'b0 ;
  assign n21236 = n6402 & ~n11239 ;
  assign n21237 = n21236 ^ n6049 ^ 1'b0 ;
  assign n21238 = n4319 & ~n5166 ;
  assign n21239 = n21238 ^ n13186 ^ 1'b0 ;
  assign n21240 = n10066 | n21239 ;
  assign n21241 = n5828 ^ n3940 ^ 1'b0 ;
  assign n21242 = n10098 ^ n5504 ^ 1'b0 ;
  assign n21243 = n21242 ^ n16055 ^ 1'b0 ;
  assign n21244 = n2018 & n21243 ;
  assign n21245 = n1291 | n1299 ;
  assign n21246 = n21245 ^ n2765 ^ 1'b0 ;
  assign n21247 = n481 ^ n461 ^ 1'b0 ;
  assign n21248 = n21246 & ~n21247 ;
  assign n21249 = n1464 | n5583 ;
  assign n21250 = n18133 & ~n21249 ;
  assign n21251 = n1523 & ~n18104 ;
  assign n21252 = n15624 & ~n21251 ;
  assign n21253 = n21252 ^ n6582 ^ 1'b0 ;
  assign n21254 = n4130 ^ n2979 ^ 1'b0 ;
  assign n21255 = n1988 | n21254 ;
  assign n21256 = ~n9860 & n21255 ;
  assign n21257 = n13663 ^ n3534 ^ 1'b0 ;
  assign n21258 = n18638 ^ n3189 ^ 1'b0 ;
  assign n21259 = n5307 & n21258 ;
  assign n21260 = ~x113 & x178 ;
  assign n21261 = n3495 ^ n1330 ^ 1'b0 ;
  assign n21262 = n15644 ^ n12440 ^ 1'b0 ;
  assign n21263 = n426 & ~n21262 ;
  assign n21264 = n21263 ^ n13893 ^ 1'b0 ;
  assign n21265 = n4398 ^ n3880 ^ 1'b0 ;
  assign n21266 = n7643 ^ n2833 ^ 1'b0 ;
  assign n21267 = n21266 ^ n14825 ^ 1'b0 ;
  assign n21268 = n21265 & ~n21267 ;
  assign n21269 = n7121 & n21268 ;
  assign n21270 = n10269 ^ n6945 ^ 1'b0 ;
  assign n21271 = n6296 & n21142 ;
  assign n21272 = n11964 & ~n18632 ;
  assign n21273 = n17332 ^ n16209 ^ n2968 ;
  assign n21274 = n15543 ^ n13694 ^ 1'b0 ;
  assign n21275 = ~n7942 & n18527 ;
  assign n21277 = n8970 ^ n3739 ^ 1'b0 ;
  assign n21276 = n11427 | n17902 ;
  assign n21278 = n21277 ^ n21276 ^ 1'b0 ;
  assign n21279 = n3890 | n21278 ;
  assign n21280 = n21279 ^ n4606 ^ 1'b0 ;
  assign n21281 = n8855 & ~n21251 ;
  assign n21282 = n5509 & n7743 ;
  assign n21283 = n3270 & ~n21282 ;
  assign n21284 = ~n20905 & n21283 ;
  assign n21285 = x193 & n302 ;
  assign n21286 = ~x193 & n21285 ;
  assign n21287 = ~n1658 & n2765 ;
  assign n21288 = n21286 & n21287 ;
  assign n21289 = n18253 | n21288 ;
  assign n21290 = n18253 & ~n21289 ;
  assign n21291 = ~n17298 & n21290 ;
  assign n21292 = n1344 & n3908 ;
  assign n21293 = n21292 ^ n4087 ^ 1'b0 ;
  assign n21294 = x182 & n21293 ;
  assign n21295 = ~n21291 & n21294 ;
  assign n21296 = ~n11865 & n14272 ;
  assign n21297 = n9545 ^ n7529 ^ 1'b0 ;
  assign n21298 = n20469 ^ n11374 ^ 1'b0 ;
  assign n21299 = n2698 & n21298 ;
  assign n21300 = ~n21297 & n21299 ;
  assign n21301 = n1328 & ~n7170 ;
  assign n21302 = n21301 ^ n715 ^ 1'b0 ;
  assign n21303 = n21302 ^ n1028 ^ 1'b0 ;
  assign n21304 = n6934 ^ n6637 ^ 1'b0 ;
  assign n21305 = ~n17062 & n21304 ;
  assign n21306 = n18491 ^ n9184 ^ 1'b0 ;
  assign n21307 = n12083 & ~n21306 ;
  assign n21308 = n19059 ^ n2591 ^ 1'b0 ;
  assign n21309 = n18114 & ~n21308 ;
  assign n21310 = n1310 ^ x230 ^ 1'b0 ;
  assign n21311 = n21310 ^ n4653 ^ 1'b0 ;
  assign n21312 = ~n1951 & n7771 ;
  assign n21313 = ~n21311 & n21312 ;
  assign n21314 = ~n1488 & n8964 ;
  assign n21315 = n6743 ^ n2366 ^ 1'b0 ;
  assign n21316 = n6076 & n11963 ;
  assign n21317 = n21315 & n21316 ;
  assign n21318 = n3407 & n5938 ;
  assign n21319 = n21318 ^ n16420 ^ 1'b0 ;
  assign n21320 = ~n15037 & n21319 ;
  assign n21321 = n9913 ^ n546 ^ 1'b0 ;
  assign n21322 = n5047 & ~n19680 ;
  assign n21323 = n21321 & n21322 ;
  assign n21324 = n11937 ^ n1111 ^ 1'b0 ;
  assign n21325 = n1470 | n21324 ;
  assign n21326 = n7349 ^ n2185 ^ 1'b0 ;
  assign n21327 = n21325 | n21326 ;
  assign n21328 = n3142 ^ n2417 ^ 1'b0 ;
  assign n21329 = n21328 ^ n1184 ^ 1'b0 ;
  assign n21330 = ~n18038 & n21329 ;
  assign n21331 = n21327 & n21330 ;
  assign n21332 = n1742 & ~n8233 ;
  assign n21333 = ~n7021 & n8123 ;
  assign n21334 = n6032 ^ n535 ^ 1'b0 ;
  assign n21335 = ~n3614 & n21334 ;
  assign n21336 = n5861 | n21335 ;
  assign n21337 = n1028 | n3774 ;
  assign n21338 = n2786 | n21337 ;
  assign n21339 = ~n4523 & n6431 ;
  assign n21340 = n21338 & ~n21339 ;
  assign n21341 = n8435 ^ n7108 ^ 1'b0 ;
  assign n21342 = n15719 | n21341 ;
  assign n21343 = n17283 & n21342 ;
  assign n21344 = ~x157 & n7007 ;
  assign n21345 = n8658 | n13554 ;
  assign n21346 = n21345 ^ n13892 ^ 1'b0 ;
  assign n21347 = ~n1909 & n16269 ;
  assign n21348 = n9562 & n21347 ;
  assign n21349 = n9254 | n12859 ;
  assign n21350 = n3199 & ~n11116 ;
  assign n21351 = n2786 | n6278 ;
  assign n21352 = n21351 ^ n10550 ^ 1'b0 ;
  assign n21353 = n12140 | n21352 ;
  assign n21354 = n12223 & ~n21353 ;
  assign n21355 = n1325 & ~n18049 ;
  assign n21356 = n21355 ^ n7841 ^ 1'b0 ;
  assign n21357 = n296 & n21356 ;
  assign n21358 = n21357 ^ n20811 ^ 1'b0 ;
  assign n21359 = n12702 & n14472 ;
  assign n21360 = n16208 ^ n10630 ^ 1'b0 ;
  assign n21361 = n10814 & n21360 ;
  assign n21362 = n6425 & n21361 ;
  assign n21363 = n21362 ^ n16034 ^ 1'b0 ;
  assign n21364 = n11511 ^ n6198 ^ 1'b0 ;
  assign n21365 = n21363 | n21364 ;
  assign n21366 = n8014 & n21042 ;
  assign n21367 = n21366 ^ n361 ^ 1'b0 ;
  assign n21368 = n14024 | n21367 ;
  assign n21369 = n6792 & ~n18896 ;
  assign n21370 = n21368 & n21369 ;
  assign n21371 = n2987 & ~n14380 ;
  assign n21372 = ~n17432 & n20568 ;
  assign n21373 = n5870 & n21372 ;
  assign n21374 = x163 | n6592 ;
  assign n21378 = n7216 ^ n349 ^ 1'b0 ;
  assign n21379 = n6649 & n21378 ;
  assign n21375 = ~n551 & n8875 ;
  assign n21376 = n21375 ^ n8572 ^ 1'b0 ;
  assign n21377 = n445 & n21376 ;
  assign n21380 = n21379 ^ n21377 ^ 1'b0 ;
  assign n21381 = ~n17311 & n21380 ;
  assign n21382 = n16564 ^ n11291 ^ 1'b0 ;
  assign n21383 = ~n6571 & n14170 ;
  assign n21384 = n12585 ^ n6372 ^ 1'b0 ;
  assign n21385 = n21384 ^ n9816 ^ 1'b0 ;
  assign n21386 = ~n3219 & n9234 ;
  assign n21387 = n21386 ^ n14395 ^ 1'b0 ;
  assign n21388 = n3902 & ~n10666 ;
  assign n21389 = n21388 ^ n6307 ^ 1'b0 ;
  assign n21390 = n21387 & n21389 ;
  assign n21391 = n2824 & n12071 ;
  assign n21392 = n21391 ^ n2718 ^ 1'b0 ;
  assign n21393 = ( ~n21064 & n21390 ) | ( ~n21064 & n21392 ) | ( n21390 & n21392 ) ;
  assign n21394 = n3270 & ~n5286 ;
  assign n21395 = ~n10972 & n21394 ;
  assign n21397 = n9176 ^ n4637 ^ 1'b0 ;
  assign n21396 = n10044 & n12652 ;
  assign n21398 = n21397 ^ n21396 ^ 1'b0 ;
  assign n21399 = n11096 ^ n392 ^ 1'b0 ;
  assign n21400 = n21128 ^ n16483 ^ 1'b0 ;
  assign n21401 = n594 | n21400 ;
  assign n21402 = n11945 & n18872 ;
  assign n21409 = n3774 | n4444 ;
  assign n21410 = n21409 ^ n6931 ^ 1'b0 ;
  assign n21411 = n1503 & n5207 ;
  assign n21412 = n21410 & n21411 ;
  assign n21413 = n21412 ^ n3116 ^ 1'b0 ;
  assign n21403 = n2938 & n10708 ;
  assign n21404 = ~n9711 & n21403 ;
  assign n21405 = n2629 | n14635 ;
  assign n21406 = n7510 | n21405 ;
  assign n21407 = n11207 & ~n21406 ;
  assign n21408 = n21404 | n21407 ;
  assign n21414 = n21413 ^ n21408 ^ 1'b0 ;
  assign n21415 = n5197 & ~n7527 ;
  assign n21416 = n1442 & n21415 ;
  assign n21417 = n21416 ^ n16783 ^ 1'b0 ;
  assign n21418 = ~n1135 & n4075 ;
  assign n21419 = n6442 ^ n881 ^ 1'b0 ;
  assign n21420 = n11915 & ~n13225 ;
  assign n21421 = ( ~n8300 & n21419 ) | ( ~n8300 & n21420 ) | ( n21419 & n21420 ) ;
  assign n21422 = n13000 ^ n7968 ^ 1'b0 ;
  assign n21423 = n492 & n21422 ;
  assign n21424 = n14974 ^ n5660 ^ 1'b0 ;
  assign n21425 = n6517 & n21424 ;
  assign n21426 = n5600 & ~n16931 ;
  assign n21427 = n16927 ^ n4509 ^ 1'b0 ;
  assign n21428 = n7508 & n19121 ;
  assign n21429 = n11543 & n21428 ;
  assign n21430 = n7971 & n9575 ;
  assign n21431 = n21430 ^ n8928 ^ 1'b0 ;
  assign n21432 = n3123 & n21431 ;
  assign n21433 = n7769 & n18510 ;
  assign n21434 = n4012 | n21433 ;
  assign n21435 = n3928 & ~n15692 ;
  assign n21436 = n6054 & ~n13325 ;
  assign n21437 = n4172 ^ n1291 ^ 1'b0 ;
  assign n21438 = n8088 | n21437 ;
  assign n21439 = n6752 & n14084 ;
  assign n21440 = n21439 ^ n14510 ^ 1'b0 ;
  assign n21441 = n2440 & n6014 ;
  assign n21442 = n7634 & n21441 ;
  assign n21443 = n10699 ^ n6722 ^ 1'b0 ;
  assign n21444 = n13617 ^ n673 ^ 1'b0 ;
  assign n21445 = n18609 & ~n21444 ;
  assign n21446 = n12959 ^ n4283 ^ 1'b0 ;
  assign n21447 = n16572 & n21446 ;
  assign n21448 = x148 & ~n15507 ;
  assign n21449 = ~n7098 & n17283 ;
  assign n21450 = n9367 ^ n1409 ^ 1'b0 ;
  assign n21451 = n21450 ^ x248 ^ 1'b0 ;
  assign n21452 = ( n1646 & n10863 ) | ( n1646 & n17379 ) | ( n10863 & n17379 ) ;
  assign n21453 = n6020 & ~n20232 ;
  assign n21454 = ~n6020 & n21453 ;
  assign n21455 = n21454 ^ n3091 ^ 1'b0 ;
  assign n21456 = ~n17464 & n21455 ;
  assign n21457 = ~n19488 & n21456 ;
  assign n21458 = ~x142 & n13535 ;
  assign n21459 = n6001 | n21080 ;
  assign n21460 = n11345 & ~n15827 ;
  assign n21464 = n5069 ^ n4021 ^ 1'b0 ;
  assign n21465 = n2744 & n21464 ;
  assign n21461 = n2423 & ~n4538 ;
  assign n21462 = n21461 ^ n1974 ^ 1'b0 ;
  assign n21463 = ~n347 & n21462 ;
  assign n21466 = n21465 ^ n21463 ^ 1'b0 ;
  assign n21467 = n21304 ^ n18059 ^ 1'b0 ;
  assign n21468 = n3974 & ~n21467 ;
  assign n21469 = n2885 & ~n17448 ;
  assign n21470 = n4982 & n9906 ;
  assign n21471 = n955 & n11789 ;
  assign n21472 = n21471 ^ n3462 ^ 1'b0 ;
  assign n21474 = n7746 ^ n6617 ^ 1'b0 ;
  assign n21473 = ~n10584 & n11397 ;
  assign n21475 = n21474 ^ n21473 ^ 1'b0 ;
  assign n21476 = ( n557 & n3908 ) | ( n557 & ~n9479 ) | ( n3908 & ~n9479 ) ;
  assign n21477 = n8456 | n19428 ;
  assign n21478 = n21476 & ~n21477 ;
  assign n21479 = n8669 | n10201 ;
  assign n21480 = n21479 ^ n14538 ^ 1'b0 ;
  assign n21481 = n681 | n11327 ;
  assign n21482 = n21481 ^ n17738 ^ 1'b0 ;
  assign n21483 = n6112 ^ n495 ^ 1'b0 ;
  assign n21484 = n21483 ^ n6033 ^ 1'b0 ;
  assign n21485 = n8223 ^ n7567 ^ 1'b0 ;
  assign n21486 = ~n21484 & n21485 ;
  assign n21487 = ( ~n6574 & n21482 ) | ( ~n6574 & n21486 ) | ( n21482 & n21486 ) ;
  assign n21488 = n21480 & n21487 ;
  assign n21489 = n10530 ^ n9580 ^ 1'b0 ;
  assign n21490 = n11858 ^ n10780 ^ 1'b0 ;
  assign n21491 = n15235 | n18716 ;
  assign n21492 = n10491 | n21491 ;
  assign n21493 = n19691 | n21492 ;
  assign n21494 = n951 | n12535 ;
  assign n21495 = n19241 ^ n8207 ^ 1'b0 ;
  assign n21496 = n21495 ^ n17045 ^ n2564 ;
  assign n21497 = n4690 | n5626 ;
  assign n21498 = n2074 & ~n2295 ;
  assign n21499 = n21498 ^ n14498 ^ n8728 ;
  assign n21500 = n9528 ^ n3069 ^ 1'b0 ;
  assign n21501 = n5095 ^ n2404 ^ x236 ;
  assign n21502 = ~n661 & n3256 ;
  assign n21503 = n8915 ^ n335 ^ 1'b0 ;
  assign n21504 = n10739 ^ n2544 ^ 1'b0 ;
  assign n21505 = n21504 ^ n10983 ^ 1'b0 ;
  assign n21506 = n21505 ^ n3789 ^ n838 ;
  assign n21507 = n1955 & ~n15820 ;
  assign n21508 = n8103 ^ n5409 ^ n2550 ;
  assign n21509 = n6602 ^ n1559 ^ 1'b0 ;
  assign n21510 = n4693 & ~n10344 ;
  assign n21511 = ~n21509 & n21510 ;
  assign n21512 = ~n14717 & n21511 ;
  assign n21513 = ~n1810 & n21512 ;
  assign n21514 = n5859 & ~n6553 ;
  assign n21515 = n10955 & n21514 ;
  assign n21516 = n11073 & n21515 ;
  assign n21517 = ~n1890 & n7026 ;
  assign n21518 = n21517 ^ n18768 ^ 1'b0 ;
  assign n21519 = n1272 | n1922 ;
  assign n21520 = n13438 ^ n1248 ^ 1'b0 ;
  assign n21521 = n8706 & ~n21520 ;
  assign n21522 = n21521 ^ n3404 ^ 1'b0 ;
  assign n21523 = n14229 & n21522 ;
  assign n21524 = n21519 & n21523 ;
  assign n21525 = n18251 ^ n11818 ^ 1'b0 ;
  assign n21526 = n1819 & ~n13133 ;
  assign n21527 = n21526 ^ n6900 ^ 1'b0 ;
  assign n21528 = n810 | n21527 ;
  assign n21529 = n9354 & ~n21528 ;
  assign n21530 = n7805 | n21529 ;
  assign n21531 = n14514 & n14755 ;
  assign n21532 = n13321 & n21531 ;
  assign n21533 = n6879 & n15851 ;
  assign n21534 = n2716 & ~n13524 ;
  assign n21536 = n9244 ^ n4260 ^ 1'b0 ;
  assign n21537 = n12795 & n21536 ;
  assign n21538 = ~n19115 & n21537 ;
  assign n21535 = n7136 | n9051 ;
  assign n21539 = n21538 ^ n21535 ^ 1'b0 ;
  assign n21540 = n3065 ^ n1808 ^ 1'b0 ;
  assign n21541 = n7326 & n21540 ;
  assign n21542 = n2350 & n3729 ;
  assign n21543 = n1540 | n21542 ;
  assign n21544 = n11133 ^ n8532 ^ 1'b0 ;
  assign n21545 = n12142 ^ n2571 ^ 1'b0 ;
  assign n21546 = n21545 ^ n13359 ^ 1'b0 ;
  assign n21547 = ~n19264 & n21546 ;
  assign n21548 = ~n3067 & n8412 ;
  assign n21549 = n21548 ^ n13385 ^ n11599 ;
  assign n21550 = n14675 ^ n3966 ^ 1'b0 ;
  assign n21551 = ~n8503 & n21550 ;
  assign n21552 = ~n10859 & n21551 ;
  assign n21553 = n21552 ^ n1195 ^ 1'b0 ;
  assign n21554 = ~n503 & n2885 ;
  assign n21555 = n8638 | n21554 ;
  assign n21556 = n6825 | n16050 ;
  assign n21557 = n17003 ^ n1896 ^ 1'b0 ;
  assign n21558 = n1548 | n21557 ;
  assign n21559 = n9010 & ~n21558 ;
  assign n21560 = n21559 ^ n17329 ^ 1'b0 ;
  assign n21562 = n420 & n15705 ;
  assign n21563 = ~n2011 & n21562 ;
  assign n21561 = n5891 & n19790 ;
  assign n21564 = n21563 ^ n21561 ^ 1'b0 ;
  assign n21565 = n13749 & n21564 ;
  assign n21566 = n15733 & n21565 ;
  assign n21567 = ~n407 & n4483 ;
  assign n21568 = n21567 ^ n15900 ^ 1'b0 ;
  assign n21569 = n7014 & n8474 ;
  assign n21570 = n21437 & n21569 ;
  assign n21571 = n1397 & ~n11210 ;
  assign n21572 = n1941 & ~n10080 ;
  assign n21573 = ~n21038 & n21572 ;
  assign n21574 = n21571 | n21573 ;
  assign n21575 = n15652 ^ n3549 ^ 1'b0 ;
  assign n21576 = n2768 ^ n696 ^ 1'b0 ;
  assign n21577 = n1339 & ~n21576 ;
  assign n21578 = n21577 ^ n9541 ^ n5748 ;
  assign n21579 = n2900 ^ n2348 ^ 1'b0 ;
  assign n21580 = n18128 | n21579 ;
  assign n21581 = n21580 ^ n13389 ^ 1'b0 ;
  assign n21582 = n298 & ~n21581 ;
  assign n21583 = n21582 ^ n14693 ^ 1'b0 ;
  assign n21584 = n2239 & ~n2343 ;
  assign n21585 = n5314 & n21584 ;
  assign n21586 = ~n9563 & n21585 ;
  assign n21587 = n10400 ^ n8765 ^ 1'b0 ;
  assign n21588 = n21586 | n21587 ;
  assign n21589 = n12838 ^ n3568 ^ 1'b0 ;
  assign n21590 = ~n13082 & n21589 ;
  assign n21591 = n21588 & n21590 ;
  assign n21592 = ( n8963 & n11345 ) | ( n8963 & ~n13383 ) | ( n11345 & ~n13383 ) ;
  assign n21593 = n14323 & n20820 ;
  assign n21594 = n8122 ^ x232 ^ 1'b0 ;
  assign n21595 = n9522 & n21594 ;
  assign n21596 = n21595 ^ n16439 ^ 1'b0 ;
  assign n21597 = n9518 & n21596 ;
  assign n21598 = n2063 & ~n21597 ;
  assign n21599 = n18311 | n21598 ;
  assign n21600 = x62 & n8597 ;
  assign n21601 = n21600 ^ n13821 ^ 1'b0 ;
  assign n21602 = n8059 ^ n337 ^ 1'b0 ;
  assign n21603 = n2531 & ~n21602 ;
  assign n21604 = n8655 & n11235 ;
  assign n21605 = ~n21603 & n21604 ;
  assign n21606 = n21605 ^ n15337 ^ 1'b0 ;
  assign n21607 = ~n14122 & n20837 ;
  assign n21608 = n3575 | n10130 ;
  assign n21609 = ~x248 & n3707 ;
  assign n21610 = n21608 & ~n21609 ;
  assign n21611 = n5932 ^ n5472 ^ 1'b0 ;
  assign n21612 = n21611 ^ n5823 ^ 1'b0 ;
  assign n21613 = x201 & ~n10774 ;
  assign n21614 = ( n14799 & n15552 ) | ( n14799 & ~n21613 ) | ( n15552 & ~n21613 ) ;
  assign n21615 = n2997 & ~n3438 ;
  assign n21616 = n2735 & n19235 ;
  assign n21617 = ~n7097 & n21616 ;
  assign n21618 = n21617 ^ n18293 ^ n1866 ;
  assign n21619 = ~n2145 & n3713 ;
  assign n21620 = n6944 & n21619 ;
  assign n21621 = n1337 | n21620 ;
  assign n21622 = ~n4298 & n21621 ;
  assign n21623 = n21622 ^ n18180 ^ 1'b0 ;
  assign n21624 = n2652 & n7967 ;
  assign n21625 = n21624 ^ n3397 ^ 1'b0 ;
  assign n21626 = n21625 ^ n1295 ^ 1'b0 ;
  assign n21627 = n3189 & n7882 ;
  assign n21628 = n21627 ^ n20236 ^ 1'b0 ;
  assign n21629 = n10674 ^ n4091 ^ 1'b0 ;
  assign n21630 = n19775 & ~n21629 ;
  assign n21631 = n21630 ^ n6001 ^ 1'b0 ;
  assign n21632 = n1120 & ~n20469 ;
  assign n21635 = n16403 ^ n2362 ^ 1'b0 ;
  assign n21633 = n17652 & ~n18253 ;
  assign n21634 = n9455 & n21633 ;
  assign n21636 = n21635 ^ n21634 ^ 1'b0 ;
  assign n21637 = n21636 ^ n8553 ^ 1'b0 ;
  assign n21638 = n5157 | n21637 ;
  assign n21639 = n19313 & ~n21638 ;
  assign n21640 = n5928 & n21639 ;
  assign n21643 = ~n9747 & n10264 ;
  assign n21644 = n1227 & n21643 ;
  assign n21645 = ( n12087 & n13668 ) | ( n12087 & ~n21644 ) | ( n13668 & ~n21644 ) ;
  assign n21641 = n15737 & ~n17531 ;
  assign n21642 = n5371 & n21641 ;
  assign n21646 = n21645 ^ n21642 ^ 1'b0 ;
  assign n21647 = n10708 ^ n10226 ^ n4625 ;
  assign n21648 = n5798 | n21647 ;
  assign n21649 = n2378 & ~n7504 ;
  assign n21650 = n1505 & n21649 ;
  assign n21651 = n294 | n21650 ;
  assign n21652 = n21651 ^ x65 ^ 1'b0 ;
  assign n21653 = n4627 | n7628 ;
  assign n21654 = n21653 ^ n9799 ^ 1'b0 ;
  assign n21655 = n6522 ^ n3974 ^ 1'b0 ;
  assign n21656 = n8661 & n21655 ;
  assign n21657 = n11004 ^ n9983 ^ 1'b0 ;
  assign n21658 = n7708 & ~n21657 ;
  assign n21660 = x9 | n11221 ;
  assign n21659 = n8617 | n9059 ;
  assign n21661 = n21660 ^ n21659 ^ n9109 ;
  assign n21662 = n4551 & n21661 ;
  assign n21663 = x139 | n20790 ;
  assign n21664 = n600 | n2066 ;
  assign n21665 = n9472 & ~n21664 ;
  assign n21666 = n9388 & n19644 ;
  assign n21667 = n5423 ^ n4804 ^ 1'b0 ;
  assign n21668 = n10699 & ~n13725 ;
  assign n21669 = n8959 ^ n7996 ^ n1575 ;
  assign n21670 = n21669 ^ n3968 ^ 1'b0 ;
  assign n21671 = ~n1160 & n6775 ;
  assign n21672 = n13237 ^ n4375 ^ 1'b0 ;
  assign n21673 = n4652 & n21672 ;
  assign n21674 = n10281 | n14989 ;
  assign n21675 = n17965 | n21674 ;
  assign n21676 = n12200 ^ n7098 ^ 1'b0 ;
  assign n21677 = n12795 & n19832 ;
  assign n21678 = ~n21676 & n21677 ;
  assign n21679 = n13835 | n18464 ;
  assign n21680 = n5364 | n21679 ;
  assign n21681 = n6448 & n8750 ;
  assign n21682 = n1116 ^ x194 ^ 1'b0 ;
  assign n21688 = n13153 ^ n12329 ^ 1'b0 ;
  assign n21687 = n12189 & n18432 ;
  assign n21689 = n21688 ^ n21687 ^ 1'b0 ;
  assign n21683 = ~n4178 & n7744 ;
  assign n21684 = n21683 ^ n6529 ^ 1'b0 ;
  assign n21685 = n21684 ^ n11543 ^ 1'b0 ;
  assign n21686 = n6527 | n21685 ;
  assign n21690 = n21689 ^ n21686 ^ 1'b0 ;
  assign n21691 = n10017 ^ n8811 ^ 1'b0 ;
  assign n21692 = n12297 & n21691 ;
  assign n21693 = n2172 | n10924 ;
  assign n21694 = ~n2278 & n21693 ;
  assign n21695 = n21694 ^ n8489 ^ 1'b0 ;
  assign n21696 = n21692 | n21695 ;
  assign n21697 = n4540 & n7268 ;
  assign n21698 = n5573 & n12695 ;
  assign n21699 = ~n4097 & n21698 ;
  assign n21700 = n21699 ^ n13616 ^ 1'b0 ;
  assign n21702 = n585 | n5489 ;
  assign n21703 = n21702 ^ n2179 ^ 1'b0 ;
  assign n21701 = n7818 & ~n15820 ;
  assign n21704 = n21703 ^ n21701 ^ 1'b0 ;
  assign n21705 = n860 & ~n6179 ;
  assign n21706 = n3223 & n21705 ;
  assign n21707 = n16137 ^ n9005 ^ 1'b0 ;
  assign n21708 = n6369 | n21707 ;
  assign n21709 = n1424 & ~n20700 ;
  assign n21710 = n21708 & n21709 ;
  assign n21712 = n13439 ^ n3825 ^ 1'b0 ;
  assign n21713 = n8059 | n21712 ;
  assign n21714 = n3412 & ~n21713 ;
  assign n21711 = ~n4075 & n5778 ;
  assign n21715 = n21714 ^ n21711 ^ 1'b0 ;
  assign n21716 = n21715 ^ n7818 ^ 1'b0 ;
  assign n21717 = n6172 ^ n4751 ^ 1'b0 ;
  assign n21718 = n16130 | n21717 ;
  assign n21721 = n13173 ^ n4938 ^ 1'b0 ;
  assign n21722 = n7431 & n21721 ;
  assign n21719 = n5737 ^ n4726 ^ 1'b0 ;
  assign n21720 = ~n5384 & n21719 ;
  assign n21723 = n21722 ^ n21720 ^ 1'b0 ;
  assign n21724 = n9600 ^ n2990 ^ 1'b0 ;
  assign n21725 = n1654 ^ n968 ^ 1'b0 ;
  assign n21726 = ~n4573 & n10771 ;
  assign n21727 = ~n19807 & n21726 ;
  assign n21728 = n10100 ^ n6200 ^ n271 ;
  assign n21729 = n20988 ^ n6998 ^ 1'b0 ;
  assign n21730 = n10697 ^ n7401 ^ 1'b0 ;
  assign n21731 = ~n516 & n6784 ;
  assign n21732 = n6346 ^ x1 ^ 1'b0 ;
  assign n21733 = n1467 | n21732 ;
  assign n21734 = n10239 & ~n21733 ;
  assign n21735 = ~n4399 & n21734 ;
  assign n21736 = ~n3747 & n21735 ;
  assign n21737 = n3468 | n6544 ;
  assign n21738 = n15789 & ~n21737 ;
  assign n21739 = n3520 & n15842 ;
  assign n21740 = ~n4188 & n16181 ;
  assign n21741 = n17101 ^ n3941 ^ 1'b0 ;
  assign n21742 = n2127 & ~n5121 ;
  assign n21743 = ~n15434 & n21742 ;
  assign n21744 = n14308 ^ n6322 ^ 1'b0 ;
  assign n21745 = n5105 ^ n1077 ^ 1'b0 ;
  assign n21746 = n4270 & n14421 ;
  assign n21747 = n2055 ^ n502 ^ 1'b0 ;
  assign n21748 = n5398 & ~n21747 ;
  assign n21749 = x144 & ~n9428 ;
  assign n21750 = n16057 & n21749 ;
  assign n21751 = n13012 ^ n12707 ^ 1'b0 ;
  assign n21752 = n18440 | n19383 ;
  assign n21753 = n17806 | n21752 ;
  assign n21754 = n14440 ^ n3411 ^ 1'b0 ;
  assign n21755 = n6715 ^ n1400 ^ 1'b0 ;
  assign n21756 = n21755 ^ n19272 ^ 1'b0 ;
  assign n21757 = n4772 & ~n19265 ;
  assign n21758 = n21756 & n21757 ;
  assign n21759 = n17230 ^ n4986 ^ 1'b0 ;
  assign n21760 = n12239 & n19907 ;
  assign n21761 = ~n8379 & n21760 ;
  assign n21762 = n7337 ^ n1037 ^ 1'b0 ;
  assign n21763 = n12948 & ~n21762 ;
  assign n21764 = n10800 & ~n13949 ;
  assign n21765 = n16783 | n21764 ;
  assign n21766 = n21765 ^ n17838 ^ 1'b0 ;
  assign n21767 = n14991 ^ n7429 ^ 1'b0 ;
  assign n21768 = n3533 & ~n21767 ;
  assign n21769 = n21768 ^ n4031 ^ 1'b0 ;
  assign n21770 = n7475 & n12887 ;
  assign n21771 = n21770 ^ n3466 ^ 1'b0 ;
  assign n21772 = n21674 ^ n9188 ^ 1'b0 ;
  assign n21773 = ~n1696 & n21772 ;
  assign n21774 = n1793 ^ n607 ^ 1'b0 ;
  assign n21775 = n14866 ^ n2057 ^ 1'b0 ;
  assign n21776 = n8328 | n16624 ;
  assign n21777 = x226 & n6322 ;
  assign n21778 = n21777 ^ n15589 ^ 1'b0 ;
  assign n21779 = ~n2225 & n21778 ;
  assign n21780 = x1 & ~n320 ;
  assign n21781 = n15579 ^ n12048 ^ 1'b0 ;
  assign n21782 = n13045 & ~n21781 ;
  assign n21783 = n21782 ^ n19058 ^ n2866 ;
  assign n21784 = n3796 ^ x142 ^ 1'b0 ;
  assign n21785 = n21783 | n21784 ;
  assign n21786 = n10753 & n15049 ;
  assign n21787 = n18134 & n18410 ;
  assign n21788 = n3308 & n21787 ;
  assign n21789 = n5898 ^ n1805 ^ 1'b0 ;
  assign n21790 = ~n2711 & n21789 ;
  assign n21791 = n19054 ^ n733 ^ 1'b0 ;
  assign n21792 = x132 & ~n4276 ;
  assign n21793 = ~n21791 & n21792 ;
  assign n21794 = n21793 ^ n16767 ^ 1'b0 ;
  assign n21795 = n11916 ^ n2089 ^ 1'b0 ;
  assign n21796 = n11864 & n21795 ;
  assign n21797 = n21796 ^ n4345 ^ 1'b0 ;
  assign n21798 = n21794 & ~n21797 ;
  assign n21799 = n7427 ^ n6904 ^ 1'b0 ;
  assign n21800 = ~n8957 & n21799 ;
  assign n21801 = n14852 & n21800 ;
  assign n21802 = ~n9985 & n21801 ;
  assign n21803 = ~n7897 & n17669 ;
  assign n21804 = n4826 ^ n4010 ^ 1'b0 ;
  assign n21805 = n7876 & ~n21804 ;
  assign n21806 = n2665 & n6879 ;
  assign n21807 = n21806 ^ n10310 ^ 1'b0 ;
  assign n21808 = n2668 | n11597 ;
  assign n21809 = n16238 & ~n21808 ;
  assign n21810 = ~n1696 & n13029 ;
  assign n21811 = ~n16022 & n21810 ;
  assign n21812 = n21809 & n21811 ;
  assign n21813 = n1108 & ~n3216 ;
  assign n21814 = n14187 | n21813 ;
  assign n21815 = n21814 ^ n903 ^ 1'b0 ;
  assign n21816 = n21815 ^ n4655 ^ 1'b0 ;
  assign n21817 = n6886 & n10306 ;
  assign n21818 = n21817 ^ n12697 ^ 1'b0 ;
  assign n21819 = n11979 | n19885 ;
  assign n21820 = n6827 & n10462 ;
  assign n21821 = n512 & ~n8753 ;
  assign n21822 = ~n8912 & n21821 ;
  assign n21823 = n6431 & n21822 ;
  assign n21825 = n1405 & n5798 ;
  assign n21826 = n1370 & n21825 ;
  assign n21824 = n2283 & n11431 ;
  assign n21827 = n21826 ^ n21824 ^ 1'b0 ;
  assign n21828 = n5642 ^ n1299 ^ 1'b0 ;
  assign n21829 = n21827 & n21828 ;
  assign n21830 = n899 & ~n8345 ;
  assign n21831 = n21830 ^ n15011 ^ 1'b0 ;
  assign n21832 = ~n21124 & n21831 ;
  assign n21833 = n1159 & n3333 ;
  assign n21834 = n9791 & n17590 ;
  assign n21835 = n21834 ^ n4502 ^ 1'b0 ;
  assign n21836 = n7631 ^ n5692 ^ 1'b0 ;
  assign n21837 = n21835 | n21836 ;
  assign n21838 = n2610 ^ n1740 ^ 1'b0 ;
  assign n21839 = ~n16887 & n21838 ;
  assign n21840 = n8233 | n10585 ;
  assign n21841 = n17467 & ~n21840 ;
  assign n21842 = n15067 & n21841 ;
  assign n21843 = n13062 | n21842 ;
  assign n21844 = n1339 ^ x113 ^ 1'b0 ;
  assign n21845 = n4106 ^ n752 ^ 1'b0 ;
  assign n21846 = n9284 & n21845 ;
  assign n21847 = ~n2276 & n21846 ;
  assign n21848 = n1330 ^ n903 ^ 1'b0 ;
  assign n21849 = n17062 & n21848 ;
  assign n21850 = n5385 & n8148 ;
  assign n21851 = n21850 ^ n14647 ^ 1'b0 ;
  assign n21852 = n21851 ^ n13189 ^ 1'b0 ;
  assign n21853 = n11673 | n21852 ;
  assign n21854 = n21853 ^ n17690 ^ 1'b0 ;
  assign n21855 = n2855 & n5675 ;
  assign n21856 = ~n13498 & n21855 ;
  assign n21857 = ~n14491 & n21522 ;
  assign n21858 = n12535 & ~n18422 ;
  assign n21859 = ( ~n6307 & n9071 ) | ( ~n6307 & n19805 ) | ( n9071 & n19805 ) ;
  assign n21860 = n3212 & ~n3667 ;
  assign n21861 = n21860 ^ n2539 ^ 1'b0 ;
  assign n21862 = n4460 & ~n21861 ;
  assign n21863 = ~n15263 & n17820 ;
  assign n21864 = n10488 ^ n9596 ^ 1'b0 ;
  assign n21865 = n18926 ^ n9559 ^ 1'b0 ;
  assign n21866 = n4970 ^ n3089 ^ 1'b0 ;
  assign n21867 = n18971 & ~n21866 ;
  assign n21868 = n21867 ^ n1770 ^ 1'b0 ;
  assign n21869 = ~n21352 & n21868 ;
  assign n21870 = n1085 & n3710 ;
  assign n21871 = n21870 ^ n7054 ^ 1'b0 ;
  assign n21872 = n5555 ^ n1672 ^ 1'b0 ;
  assign n21873 = n6990 & ~n21872 ;
  assign n21874 = ( n3982 & ~n4173 ) | ( n3982 & n14279 ) | ( ~n4173 & n14279 ) ;
  assign n21875 = n19486 ^ n7994 ^ 1'b0 ;
  assign n21876 = n4290 & ~n21875 ;
  assign n21877 = n5987 & n18617 ;
  assign n21878 = n5026 & ~n17788 ;
  assign n21879 = n21878 ^ n3126 ^ 1'b0 ;
  assign n21880 = n9380 & ~n20420 ;
  assign n21881 = n3808 & n21880 ;
  assign n21882 = n18650 ^ n1814 ^ 1'b0 ;
  assign n21883 = n1935 & ~n8803 ;
  assign n21884 = n21883 ^ n2772 ^ 1'b0 ;
  assign n21885 = n21884 ^ n9643 ^ 1'b0 ;
  assign n21886 = n8094 ^ n7281 ^ n964 ;
  assign n21887 = n3143 & n21886 ;
  assign n21888 = n3473 ^ n1656 ^ 1'b0 ;
  assign n21889 = n5563 | n21888 ;
  assign n21890 = n9653 & n14240 ;
  assign n21891 = n13786 & n21890 ;
  assign n21892 = n3177 & ~n18206 ;
  assign n21893 = n6878 & ~n21892 ;
  assign n21894 = n6764 ^ n5023 ^ 1'b0 ;
  assign n21895 = n15963 & ~n21894 ;
  assign n21896 = n1252 & n6372 ;
  assign n21897 = ~n6372 & n21896 ;
  assign n21898 = n1339 | n21897 ;
  assign n21899 = n17067 & ~n21898 ;
  assign n21900 = n3850 | n5396 ;
  assign n21901 = n2142 | n21900 ;
  assign n21902 = n16823 ^ n7243 ^ 1'b0 ;
  assign n21903 = n15161 & n21902 ;
  assign n21904 = n6541 & n14316 ;
  assign n21905 = ~n7732 & n21904 ;
  assign n21906 = n8545 & n17094 ;
  assign n21907 = n9893 & n21906 ;
  assign n21908 = n18120 & n19264 ;
  assign n21909 = n5371 & n10233 ;
  assign n21910 = ( n2426 & ~n13222 ) | ( n2426 & n21909 ) | ( ~n13222 & n21909 ) ;
  assign n21911 = n6506 | n18456 ;
  assign n21912 = n6413 & n18431 ;
  assign n21913 = n21912 ^ n6343 ^ 1'b0 ;
  assign n21914 = ~n8341 & n16206 ;
  assign n21915 = n13787 & n21914 ;
  assign n21916 = n14247 ^ n2274 ^ 1'b0 ;
  assign n21917 = n13062 & n21916 ;
  assign n21918 = n14635 ^ n12037 ^ 1'b0 ;
  assign n21919 = n10725 & ~n13971 ;
  assign n21920 = n4420 | n21919 ;
  assign n21921 = n790 & ~n21920 ;
  assign n21922 = n858 & n7991 ;
  assign n21923 = n21922 ^ n9364 ^ 1'b0 ;
  assign n21924 = n5253 ^ n671 ^ 1'b0 ;
  assign n21925 = n8792 & ~n16709 ;
  assign n21926 = n17930 & ~n21925 ;
  assign n21927 = n21926 ^ n14842 ^ 1'b0 ;
  assign n21928 = n4289 ^ n2962 ^ 1'b0 ;
  assign n21929 = n9620 | n18668 ;
  assign n21930 = ~n1691 & n21929 ;
  assign n21931 = n5948 | n21930 ;
  assign n21932 = n11650 ^ n10030 ^ 1'b0 ;
  assign n21933 = n715 | n11928 ;
  assign n21934 = n1790 & ~n21933 ;
  assign n21935 = n21932 & ~n21934 ;
  assign n21936 = n9361 ^ n2373 ^ 1'b0 ;
  assign n21937 = n3985 ^ n3536 ^ 1'b0 ;
  assign n21938 = n1690 | n21937 ;
  assign n21939 = n7126 | n9329 ;
  assign n21940 = n3711 | n21939 ;
  assign n21941 = n21938 & ~n21940 ;
  assign n21942 = n21941 ^ x108 ^ 1'b0 ;
  assign n21943 = n21936 | n21942 ;
  assign n21944 = ~n5715 & n5923 ;
  assign n21945 = n6895 | n10199 ;
  assign n21946 = n1773 | n21945 ;
  assign n21947 = n5223 | n20855 ;
  assign n21948 = n21947 ^ n3036 ^ 1'b0 ;
  assign n21949 = n3308 ^ n1135 ^ 1'b0 ;
  assign n21950 = n3988 & n21949 ;
  assign n21951 = n2836 | n5203 ;
  assign n21952 = n5203 & ~n21951 ;
  assign n21953 = n21952 ^ n732 ^ 1'b0 ;
  assign n21954 = n21950 & n21953 ;
  assign n21955 = n18748 ^ n1835 ^ 1'b0 ;
  assign n21957 = n13890 ^ n2213 ^ n2195 ;
  assign n21956 = n12572 ^ n3895 ^ 1'b0 ;
  assign n21958 = n21957 ^ n21956 ^ 1'b0 ;
  assign n21959 = n6006 & ~n21958 ;
  assign n21960 = n21959 ^ n10514 ^ 1'b0 ;
  assign n21961 = ~n13310 & n21960 ;
  assign n21962 = n14484 ^ n9806 ^ 1'b0 ;
  assign n21963 = ~n1951 & n4675 ;
  assign n21964 = n21963 ^ n3383 ^ 1'b0 ;
  assign n21966 = n963 | n13603 ;
  assign n21967 = n5443 & ~n21966 ;
  assign n21965 = ~n7155 & n7485 ;
  assign n21968 = n21967 ^ n21965 ^ 1'b0 ;
  assign n21969 = n21964 & n21968 ;
  assign n21970 = n3710 & ~n7136 ;
  assign n21971 = ~n21969 & n21970 ;
  assign n21972 = n20876 ^ n20284 ^ n666 ;
  assign n21973 = ( n2524 & n11456 ) | ( n2524 & ~n15894 ) | ( n11456 & ~n15894 ) ;
  assign n21974 = ~n7754 & n10993 ;
  assign n21975 = n21974 ^ n376 ^ 1'b0 ;
  assign n21976 = ~n21973 & n21975 ;
  assign n21977 = n14225 & ~n21750 ;
  assign n21978 = n11968 & n21977 ;
  assign n21979 = n9947 ^ n3284 ^ 1'b0 ;
  assign n21980 = n21979 ^ n13344 ^ n1700 ;
  assign n21981 = n8704 & ~n19753 ;
  assign n21982 = x245 & ~n15187 ;
  assign n21983 = n21982 ^ n1389 ^ 1'b0 ;
  assign n21984 = n5021 & ~n12586 ;
  assign n21985 = ~n5021 & n21984 ;
  assign n21986 = n21985 ^ n8568 ^ 1'b0 ;
  assign n21987 = n11961 ^ n4556 ^ 1'b0 ;
  assign n21988 = ~n21986 & n21987 ;
  assign n21989 = n1126 & n4329 ;
  assign n21990 = n2027 & ~n12718 ;
  assign n21991 = n21990 ^ n17009 ^ 1'b0 ;
  assign n21992 = n21989 & n21991 ;
  assign n22002 = n18984 ^ n438 ^ 1'b0 ;
  assign n21993 = n17698 ^ n822 ^ 1'b0 ;
  assign n21994 = n1242 & ~n21993 ;
  assign n21995 = n11938 & n21994 ;
  assign n21997 = n9304 ^ n3424 ^ 1'b0 ;
  assign n21998 = ~n2860 & n21997 ;
  assign n21996 = n3126 | n5136 ;
  assign n21999 = n21998 ^ n21996 ^ 1'b0 ;
  assign n22000 = n21999 ^ n18984 ^ n3888 ;
  assign n22001 = n21995 & ~n22000 ;
  assign n22003 = n22002 ^ n22001 ^ 1'b0 ;
  assign n22004 = n18289 ^ n9550 ^ x23 ;
  assign n22005 = n659 & n4348 ;
  assign n22008 = ~n4927 & n7653 ;
  assign n22009 = n1360 & n22008 ;
  assign n22006 = ~n4674 & n5287 ;
  assign n22007 = ~n4580 & n22006 ;
  assign n22010 = n22009 ^ n22007 ^ 1'b0 ;
  assign n22011 = n15786 & n22010 ;
  assign n22012 = x31 & n1667 ;
  assign n22013 = n7442 | n20277 ;
  assign n22014 = n13247 | n22013 ;
  assign n22015 = ~n1654 & n10048 ;
  assign n22016 = n18056 & n22015 ;
  assign n22017 = n22016 ^ n3591 ^ 1'b0 ;
  assign n22018 = n3397 & ~n22017 ;
  assign n22019 = n6081 | n18783 ;
  assign n22020 = n22019 ^ n14324 ^ 1'b0 ;
  assign n22021 = n15456 | n17892 ;
  assign n22022 = n21735 | n22021 ;
  assign n22023 = x223 & n4553 ;
  assign n22024 = ~x223 & n22023 ;
  assign n22025 = n8727 ^ n6041 ^ 1'b0 ;
  assign n22026 = n22024 & n22025 ;
  assign n22027 = n5137 & ~n22026 ;
  assign n22028 = n10871 & n22027 ;
  assign n22029 = ~n22027 & n22028 ;
  assign n22030 = n2883 | n4207 ;
  assign n22031 = ~n1657 & n5877 ;
  assign n22032 = n8846 ^ n4970 ^ 1'b0 ;
  assign n22033 = n1429 & n14497 ;
  assign n22034 = n8809 ^ n7984 ^ n415 ;
  assign n22035 = n3568 & n9688 ;
  assign n22036 = n10766 ^ n7968 ^ 1'b0 ;
  assign n22037 = n22035 & ~n22036 ;
  assign n22049 = n3941 & n15050 ;
  assign n22038 = n9094 ^ n4605 ^ 1'b0 ;
  assign n22045 = n7613 ^ n2801 ^ 1'b0 ;
  assign n22041 = n13524 ^ n10877 ^ 1'b0 ;
  assign n22042 = n22041 ^ n1501 ^ 1'b0 ;
  assign n22043 = n22042 ^ n19278 ^ 1'b0 ;
  assign n22044 = n22043 ^ n2948 ^ x129 ;
  assign n22046 = n22045 ^ n22044 ^ 1'b0 ;
  assign n22039 = n15598 ^ n8619 ^ 1'b0 ;
  assign n22040 = n10864 | n22039 ;
  assign n22047 = n22046 ^ n22040 ^ 1'b0 ;
  assign n22048 = n22038 & ~n22047 ;
  assign n22050 = n22049 ^ n22048 ^ 1'b0 ;
  assign n22051 = n975 & ~n13054 ;
  assign n22052 = ~n11108 & n11926 ;
  assign n22053 = ( ~n6455 & n10400 ) | ( ~n6455 & n14375 ) | ( n10400 & n14375 ) ;
  assign n22054 = n10914 & n17624 ;
  assign n22055 = n16335 & n22054 ;
  assign n22056 = n4461 & n8740 ;
  assign n22057 = ~x73 & n22056 ;
  assign n22058 = n22055 | n22057 ;
  assign n22059 = n460 & ~n22058 ;
  assign n22060 = n18457 ^ n11685 ^ 1'b0 ;
  assign n22061 = n1052 & n21612 ;
  assign n22062 = n22061 ^ n11082 ^ 1'b0 ;
  assign n22063 = n16007 ^ n10864 ^ n3833 ;
  assign n22064 = n8885 & n22063 ;
  assign n22065 = n22064 ^ n5802 ^ 1'b0 ;
  assign n22066 = n13870 & n18751 ;
  assign n22067 = n22065 & n22066 ;
  assign n22068 = n1100 & n4009 ;
  assign n22069 = n9926 & n22068 ;
  assign n22070 = n21778 & n22069 ;
  assign n22071 = n19437 ^ n15867 ^ 1'b0 ;
  assign n22072 = n6112 ^ n6051 ^ 1'b0 ;
  assign n22073 = n1928 & ~n22072 ;
  assign n22074 = n22073 ^ n14053 ^ 1'b0 ;
  assign n22075 = n9260 ^ n1544 ^ 1'b0 ;
  assign n22076 = ~n6278 & n22075 ;
  assign n22077 = n12579 & n22076 ;
  assign n22078 = n22077 ^ n12033 ^ 1'b0 ;
  assign n22079 = n22078 ^ n14854 ^ n14103 ;
  assign n22080 = n2097 & n15597 ;
  assign n22081 = n22080 ^ n7675 ^ 1'b0 ;
  assign n22082 = n6858 ^ n4113 ^ 1'b0 ;
  assign n22083 = n8670 & ~n22082 ;
  assign n22084 = ~n9410 & n19507 ;
  assign n22085 = ~n1553 & n19718 ;
  assign n22086 = n917 | n3176 ;
  assign n22087 = n3176 & ~n22086 ;
  assign n22088 = n2119 & ~n9051 ;
  assign n22089 = n22087 & n22088 ;
  assign n22090 = ~n1914 & n22089 ;
  assign n22091 = n22090 ^ n14361 ^ 1'b0 ;
  assign n22092 = ~n10021 & n14938 ;
  assign n22093 = n6838 | n7398 ;
  assign n22094 = n22092 & ~n22093 ;
  assign n22095 = n4731 ^ n954 ^ 1'b0 ;
  assign n22096 = ( n1738 & ~n3754 ) | ( n1738 & n4323 ) | ( ~n3754 & n4323 ) ;
  assign n22097 = n22096 ^ n18070 ^ 1'b0 ;
  assign n22098 = ~n22095 & n22097 ;
  assign n22099 = n5331 ^ n2892 ^ 1'b0 ;
  assign n22100 = n19124 ^ n12703 ^ 1'b0 ;
  assign n22101 = ~n4546 & n22100 ;
  assign n22102 = n12265 ^ n2486 ^ 1'b0 ;
  assign n22103 = n4437 ^ n2642 ^ 1'b0 ;
  assign n22104 = ~n512 & n22103 ;
  assign n22105 = n5472 & n22104 ;
  assign n22106 = n10559 ^ n2257 ^ 1'b0 ;
  assign n22107 = n12733 & ~n22106 ;
  assign n22108 = ~n22105 & n22107 ;
  assign n22109 = n15904 ^ n7513 ^ 1'b0 ;
  assign n22110 = n2153 & n22109 ;
  assign n22113 = n786 & ~n3825 ;
  assign n22114 = n22113 ^ n13842 ^ 1'b0 ;
  assign n22111 = n2263 & n14352 ;
  assign n22112 = n19592 & n22111 ;
  assign n22115 = n22114 ^ n22112 ^ 1'b0 ;
  assign n22116 = n3827 & n15501 ;
  assign n22117 = n4108 | n5626 ;
  assign n22118 = n18485 | n22117 ;
  assign n22119 = n7509 | n19286 ;
  assign n22120 = ~n4024 & n5076 ;
  assign n22121 = n8456 | n14361 ;
  assign n22122 = n22121 ^ n3858 ^ 1'b0 ;
  assign n22124 = n3583 & n7805 ;
  assign n22123 = n1920 | n2505 ;
  assign n22125 = n22124 ^ n22123 ^ 1'b0 ;
  assign n22126 = n1537 & ~n12636 ;
  assign n22127 = n22126 ^ n3258 ^ 1'b0 ;
  assign n22128 = ~n4753 & n6822 ;
  assign n22129 = n21356 ^ n3546 ^ 1'b0 ;
  assign n22130 = n2001 ^ n476 ^ 1'b0 ;
  assign n22131 = n15440 & ~n22130 ;
  assign n22132 = x251 & n22131 ;
  assign n22133 = ~n22129 & n22132 ;
  assign n22134 = n22128 & ~n22133 ;
  assign n22135 = n3554 | n18849 ;
  assign n22136 = n22135 ^ n801 ^ 1'b0 ;
  assign n22137 = n6015 & n10610 ;
  assign n22138 = n22137 ^ n16908 ^ 1'b0 ;
  assign n22139 = n22136 & ~n22138 ;
  assign n22140 = ~x11 & n15280 ;
  assign n22141 = n3741 & n22140 ;
  assign n22142 = ~n7149 & n12793 ;
  assign n22143 = n22142 ^ n12853 ^ 1'b0 ;
  assign n22144 = ~n8830 & n9759 ;
  assign n22145 = n6371 ^ n913 ^ 1'b0 ;
  assign n22146 = n5079 & n7446 ;
  assign n22147 = ~n9919 & n11680 ;
  assign n22148 = n22146 & n22147 ;
  assign n22149 = n12901 | n20587 ;
  assign n22150 = n22149 ^ n2769 ^ 1'b0 ;
  assign n22151 = n4249 & n10298 ;
  assign n22152 = x67 & n22151 ;
  assign n22153 = n18960 | n22152 ;
  assign n22154 = n22153 ^ n12633 ^ n9569 ;
  assign n22155 = n9063 | n11809 ;
  assign n22160 = n6511 ^ n3575 ^ 1'b0 ;
  assign n22161 = n8677 | n22160 ;
  assign n22162 = n22161 ^ n2735 ^ 1'b0 ;
  assign n22163 = ~n2403 & n22162 ;
  assign n22156 = n6448 ^ n4974 ^ 1'b0 ;
  assign n22157 = ~n3884 & n22156 ;
  assign n22158 = ~n1815 & n22157 ;
  assign n22159 = n12061 & ~n22158 ;
  assign n22164 = n22163 ^ n22159 ^ 1'b0 ;
  assign n22167 = n3720 & n14504 ;
  assign n22168 = ~n4219 & n22167 ;
  assign n22169 = ( n8359 & n20437 ) | ( n8359 & n22168 ) | ( n20437 & n22168 ) ;
  assign n22165 = n9269 ^ n8424 ^ 1'b0 ;
  assign n22166 = n4487 & ~n22165 ;
  assign n22170 = n22169 ^ n22166 ^ 1'b0 ;
  assign n22171 = n3065 & n13542 ;
  assign n22172 = ~n936 & n22171 ;
  assign n22173 = n9789 | n22172 ;
  assign n22174 = n4647 | n10630 ;
  assign n22175 = n22174 ^ n12235 ^ 1'b0 ;
  assign n22176 = n486 | n22175 ;
  assign n22179 = n1728 | n2576 ;
  assign n22180 = n21482 | n22179 ;
  assign n22177 = n4910 & n12386 ;
  assign n22178 = n854 & ~n22177 ;
  assign n22181 = n22180 ^ n22178 ^ 1'b0 ;
  assign n22182 = n17325 ^ n13439 ^ 1'b0 ;
  assign n22183 = n3362 & n13314 ;
  assign n22184 = n9068 ^ n7164 ^ 1'b0 ;
  assign n22185 = n2289 | n22184 ;
  assign n22188 = n8442 & ~n12120 ;
  assign n22186 = ~n3197 & n3886 ;
  assign n22187 = n20607 & n22186 ;
  assign n22189 = n22188 ^ n22187 ^ 1'b0 ;
  assign n22190 = x120 & n1972 ;
  assign n22191 = ~n1972 & n22190 ;
  assign n22192 = ~n631 & n1299 ;
  assign n22193 = n631 & n22192 ;
  assign n22194 = n9651 | n22193 ;
  assign n22195 = n22191 & ~n22194 ;
  assign n22196 = ( n5539 & n15489 ) | ( n5539 & ~n22195 ) | ( n15489 & ~n22195 ) ;
  assign n22197 = ( n11264 & n15686 ) | ( n11264 & ~n16728 ) | ( n15686 & ~n16728 ) ;
  assign n22198 = n12982 & ~n22197 ;
  assign n22199 = n22197 & n22198 ;
  assign n22200 = n22196 | n22199 ;
  assign n22201 = n22196 & ~n22200 ;
  assign n22202 = n17518 ^ n4708 ^ 1'b0 ;
  assign n22203 = n5575 & n22202 ;
  assign n22204 = n10864 ^ n4005 ^ 1'b0 ;
  assign n22205 = n6149 | n22204 ;
  assign n22206 = n3945 & n9522 ;
  assign n22207 = n22206 ^ n15675 ^ 1'b0 ;
  assign n22208 = n12610 & n22207 ;
  assign n22209 = n1221 ^ x151 ^ 1'b0 ;
  assign n22210 = n11353 & n22209 ;
  assign n22211 = n657 | n4622 ;
  assign n22212 = n3824 | n22211 ;
  assign n22213 = n8663 ^ n6655 ^ 1'b0 ;
  assign n22214 = n22212 & n22213 ;
  assign n22215 = ~n7738 & n22214 ;
  assign n22216 = n14241 & n22215 ;
  assign n22217 = n16659 ^ n1160 ^ 1'b0 ;
  assign n22218 = n12562 | n17816 ;
  assign n22219 = n22218 ^ n10988 ^ 1'b0 ;
  assign n22220 = x54 & ~n6076 ;
  assign n22221 = n11306 ^ n279 ^ 1'b0 ;
  assign n22222 = n6400 | n12061 ;
  assign n22223 = n22222 ^ n12506 ^ 1'b0 ;
  assign n22224 = n21038 & ~n22223 ;
  assign n22225 = ~n4099 & n10164 ;
  assign n22226 = ~n10106 & n22225 ;
  assign n22227 = n22226 ^ n12077 ^ 1'b0 ;
  assign n22228 = n18835 ^ n1291 ^ 1'b0 ;
  assign n22229 = n7126 | n11356 ;
  assign n22230 = n22229 ^ n11708 ^ 1'b0 ;
  assign n22231 = n6960 ^ n948 ^ 1'b0 ;
  assign n22232 = n8209 | n20125 ;
  assign n22233 = x15 & x130 ;
  assign n22234 = ~n9517 & n22233 ;
  assign n22235 = n8602 ^ n5892 ^ 1'b0 ;
  assign n22236 = ~n4333 & n6897 ;
  assign n22237 = n22236 ^ n13187 ^ 1'b0 ;
  assign n22238 = n22237 ^ n11241 ^ 1'b0 ;
  assign n22239 = ~n3915 & n21892 ;
  assign n22240 = ~n9210 & n17694 ;
  assign n22241 = n20527 & n22240 ;
  assign n22242 = ~n1343 & n17620 ;
  assign n22243 = n20514 & n22242 ;
  assign n22246 = ~n4936 & n7695 ;
  assign n22244 = n3456 ^ n2997 ^ 1'b0 ;
  assign n22245 = n5925 & ~n22244 ;
  assign n22247 = n22246 ^ n22245 ^ 1'b0 ;
  assign n22248 = n17207 & n22247 ;
  assign n22252 = n6030 | n10663 ;
  assign n22253 = n22252 ^ n4602 ^ 1'b0 ;
  assign n22249 = n5564 & n7419 ;
  assign n22250 = n14529 & n22249 ;
  assign n22251 = n22250 ^ n19448 ^ 1'b0 ;
  assign n22254 = n22253 ^ n22251 ^ n1926 ;
  assign n22256 = n5855 ^ n1172 ^ 1'b0 ;
  assign n22255 = n9143 & ~n11341 ;
  assign n22257 = n22256 ^ n22255 ^ 1'b0 ;
  assign n22258 = n8092 ^ n7190 ^ 1'b0 ;
  assign n22259 = n9018 ^ n903 ^ 1'b0 ;
  assign n22260 = ~n7381 & n22259 ;
  assign n22262 = ~n5540 & n10418 ;
  assign n22261 = ~n11960 & n22006 ;
  assign n22263 = n22262 ^ n22261 ^ 1'b0 ;
  assign n22264 = n5614 ^ n2001 ^ 1'b0 ;
  assign n22265 = n22264 ^ n17026 ^ 1'b0 ;
  assign n22266 = n1720 | n5603 ;
  assign n22267 = n7515 & n18092 ;
  assign n22268 = n2770 & n22267 ;
  assign n22269 = n22266 & ~n22268 ;
  assign n22270 = n11979 ^ n10150 ^ 1'b0 ;
  assign n22271 = ~n1757 & n19065 ;
  assign n22272 = n1948 & n8023 ;
  assign n22273 = n11653 | n13343 ;
  assign n22274 = n22272 & ~n22273 ;
  assign n22275 = n2730 ^ n956 ^ 1'b0 ;
  assign n22276 = x251 & ~n22275 ;
  assign n22277 = n22276 ^ n2311 ^ 1'b0 ;
  assign n22278 = n5665 & n6178 ;
  assign n22279 = n22278 ^ n8274 ^ 1'b0 ;
  assign n22280 = n22279 ^ n21145 ^ 1'b0 ;
  assign n22285 = ~n4914 & n5168 ;
  assign n22286 = ~n3707 & n22285 ;
  assign n22287 = n4502 | n22286 ;
  assign n22288 = n22287 ^ n3697 ^ 1'b0 ;
  assign n22289 = n22288 ^ n19974 ^ 1'b0 ;
  assign n22281 = n18730 ^ n8964 ^ 1'b0 ;
  assign n22282 = n257 & ~n1139 ;
  assign n22283 = n22282 ^ n956 ^ 1'b0 ;
  assign n22284 = n22281 | n22283 ;
  assign n22290 = n22289 ^ n22284 ^ n18741 ;
  assign n22291 = n1093 & n8733 ;
  assign n22292 = n8175 ^ n2673 ^ 1'b0 ;
  assign n22293 = ( n4473 & ~n4811 ) | ( n4473 & n22292 ) | ( ~n4811 & n22292 ) ;
  assign n22294 = ( n3862 & n6691 ) | ( n3862 & n17736 ) | ( n6691 & n17736 ) ;
  assign n22295 = n2774 | n8792 ;
  assign n22296 = n22294 | n22295 ;
  assign n22297 = n5265 & ~n5571 ;
  assign n22298 = n5571 & n22297 ;
  assign n22299 = n3437 & n22298 ;
  assign n22300 = n322 | n3397 ;
  assign n22301 = n22300 ^ n1511 ^ 1'b0 ;
  assign n22302 = n5166 | n22301 ;
  assign n22303 = n22299 & ~n22302 ;
  assign n22304 = n22296 & n22303 ;
  assign n22305 = n14477 | n16905 ;
  assign n22306 = ~n1477 & n16712 ;
  assign n22307 = n6663 ^ n1098 ^ 1'b0 ;
  assign n22308 = n21387 & ~n22307 ;
  assign n22309 = n6025 ^ n2109 ^ 1'b0 ;
  assign n22310 = ~n1160 & n22309 ;
  assign n22311 = ~n9895 & n13617 ;
  assign n22312 = n22311 ^ n13696 ^ 1'b0 ;
  assign n22313 = ( n3331 & n22310 ) | ( n3331 & n22312 ) | ( n22310 & n22312 ) ;
  assign n22314 = n4258 & ~n22313 ;
  assign n22315 = n22314 ^ n15633 ^ 1'b0 ;
  assign n22316 = n6325 & n21675 ;
  assign n22319 = x41 & n11196 ;
  assign n22317 = n6997 ^ n3270 ^ 1'b0 ;
  assign n22318 = n22317 ^ n13319 ^ 1'b0 ;
  assign n22320 = n22319 ^ n22318 ^ 1'b0 ;
  assign n22321 = ~n13848 & n16002 ;
  assign n22322 = n15106 & n22321 ;
  assign n22323 = n8212 & ~n9485 ;
  assign n22324 = n7459 ^ n5482 ^ 1'b0 ;
  assign n22325 = n22323 & n22324 ;
  assign n22326 = n7851 ^ n3824 ^ 1'b0 ;
  assign n22327 = n10619 & n17384 ;
  assign n22328 = n22327 ^ n9449 ^ 1'b0 ;
  assign n22329 = n1402 ^ x11 ^ 1'b0 ;
  assign n22330 = n926 & n22329 ;
  assign n22331 = n22328 & n22330 ;
  assign n22332 = ~n6372 & n21799 ;
  assign n22333 = n2613 | n11486 ;
  assign n22334 = n19652 ^ n15007 ^ 1'b0 ;
  assign n22335 = n10400 & n22334 ;
  assign n22336 = n8118 | n12695 ;
  assign n22337 = n16867 & n20141 ;
  assign n22338 = n22336 & n22337 ;
  assign n22339 = n14506 | n14575 ;
  assign n22340 = n7494 | n22339 ;
  assign n22341 = n5728 ^ n512 ^ 1'b0 ;
  assign n22342 = ~n623 & n6162 ;
  assign n22343 = n9340 & n22342 ;
  assign n22344 = n22343 ^ n2013 ^ 1'b0 ;
  assign n22345 = ~n21495 & n22344 ;
  assign n22347 = n5399 ^ n4242 ^ 1'b0 ;
  assign n22348 = n5923 | n22347 ;
  assign n22346 = n3931 | n11083 ;
  assign n22349 = n22348 ^ n22346 ^ 1'b0 ;
  assign n22350 = n5763 ^ n3343 ^ 1'b0 ;
  assign n22351 = n4063 | n22350 ;
  assign n22352 = n22351 ^ n2247 ^ 1'b0 ;
  assign n22353 = n380 & ~n1126 ;
  assign n22354 = ~n395 & n22353 ;
  assign n22355 = n22352 & ~n22354 ;
  assign n22356 = n22355 ^ n13125 ^ 1'b0 ;
  assign n22357 = n2575 & n8076 ;
  assign n22358 = n15513 & n22357 ;
  assign n22359 = n3999 & n5292 ;
  assign n22360 = n18185 & n22359 ;
  assign n22361 = ~n1481 & n20809 ;
  assign n22362 = n11886 & ~n22361 ;
  assign n22363 = n22362 ^ n10954 ^ 1'b0 ;
  assign n22364 = ( n1089 & n3896 ) | ( n1089 & n3903 ) | ( n3896 & n3903 ) ;
  assign n22365 = n22364 ^ n6981 ^ 1'b0 ;
  assign n22366 = n6331 ^ n4005 ^ 1'b0 ;
  assign n22367 = n5151 ^ n4720 ^ 1'b0 ;
  assign n22368 = n22366 | n22367 ;
  assign n22369 = n15743 & ~n22368 ;
  assign n22370 = n7745 ^ n6570 ^ n6290 ;
  assign n22371 = n22370 ^ n16069 ^ 1'b0 ;
  assign n22372 = n8093 & ~n22371 ;
  assign n22373 = n7206 & ~n18737 ;
  assign n22374 = n5620 | n6339 ;
  assign n22375 = n22374 ^ n11989 ^ 1'b0 ;
  assign n22376 = ( n3288 & ~n20622 ) | ( n3288 & n22375 ) | ( ~n20622 & n22375 ) ;
  assign n22377 = n6255 | n22376 ;
  assign n22378 = n1405 | n3328 ;
  assign n22379 = x222 & ~n22378 ;
  assign n22380 = n22379 ^ n3911 ^ 1'b0 ;
  assign n22381 = ~n3376 & n22380 ;
  assign n22382 = n22381 ^ n2451 ^ 1'b0 ;
  assign n22383 = n10936 ^ n6647 ^ 1'b0 ;
  assign n22384 = n5032 & n22383 ;
  assign n22385 = ~n1608 & n4660 ;
  assign n22386 = n4833 ^ n3778 ^ 1'b0 ;
  assign n22387 = n5516 | n22386 ;
  assign n22388 = n22387 ^ n7039 ^ 1'b0 ;
  assign n22389 = ~n22385 & n22388 ;
  assign n22390 = n12225 ^ n9427 ^ n7792 ;
  assign n22391 = n1025 | n2054 ;
  assign n22392 = n8967 & n10387 ;
  assign n22393 = ( n16109 & n18947 ) | ( n16109 & ~n22392 ) | ( n18947 & ~n22392 ) ;
  assign n22398 = ~n405 & n3171 ;
  assign n22399 = n22398 ^ n6548 ^ 1'b0 ;
  assign n22394 = n3493 & ~n10018 ;
  assign n22395 = n7034 ^ n3213 ^ 1'b0 ;
  assign n22396 = n22394 & ~n22395 ;
  assign n22397 = n2806 & ~n22396 ;
  assign n22400 = n22399 ^ n22397 ^ 1'b0 ;
  assign n22401 = n4899 ^ n1419 ^ 1'b0 ;
  assign n22402 = ~n3353 & n5101 ;
  assign n22403 = n22402 ^ n7378 ^ 1'b0 ;
  assign n22404 = n7549 | n22403 ;
  assign n22405 = n22401 | n22404 ;
  assign n22406 = n12467 & ~n22405 ;
  assign n22410 = n2910 ^ n1195 ^ 1'b0 ;
  assign n22407 = n5112 & ~n12559 ;
  assign n22408 = ( ~n630 & n1031 ) | ( ~n630 & n22407 ) | ( n1031 & n22407 ) ;
  assign n22409 = n1451 & ~n22408 ;
  assign n22411 = n22410 ^ n22409 ^ 1'b0 ;
  assign n22412 = n7277 ^ n580 ^ 1'b0 ;
  assign n22413 = n12494 ^ x155 ^ 1'b0 ;
  assign n22414 = ~n15745 & n22413 ;
  assign n22415 = n13717 ^ n11276 ^ 1'b0 ;
  assign n22416 = ~n1028 & n6253 ;
  assign n22417 = n22416 ^ n880 ^ 1'b0 ;
  assign n22418 = n22134 | n22417 ;
  assign n22419 = n22418 ^ n16778 ^ 1'b0 ;
  assign n22420 = n527 & ~n17542 ;
  assign n22421 = n22420 ^ n3986 ^ 1'b0 ;
  assign n22422 = n3189 & n4175 ;
  assign n22423 = n3477 | n4396 ;
  assign n22424 = n22422 & ~n22423 ;
  assign n22425 = n4104 & ~n11069 ;
  assign n22426 = n17634 & ~n22425 ;
  assign n22427 = n22424 & n22426 ;
  assign n22428 = n4851 ^ n3678 ^ 1'b0 ;
  assign n22429 = n7995 & n22428 ;
  assign n22430 = n1172 & n8768 ;
  assign n22431 = ~n1573 & n22430 ;
  assign n22432 = ~n22017 & n22431 ;
  assign n22433 = n1397 & n2527 ;
  assign n22434 = n22433 ^ n8033 ^ 1'b0 ;
  assign n22435 = n12353 | n22434 ;
  assign n22436 = n22435 ^ n19054 ^ 1'b0 ;
  assign n22437 = n22318 | n22436 ;
  assign n22438 = n5197 | n13725 ;
  assign n22439 = n22438 ^ n12848 ^ 1'b0 ;
  assign n22440 = n10857 | n15531 ;
  assign n22441 = n10563 ^ n4749 ^ 1'b0 ;
  assign n22442 = n713 | n733 ;
  assign n22443 = n733 & ~n22442 ;
  assign n22444 = n14341 | n22443 ;
  assign n22445 = n14341 & ~n22444 ;
  assign n22446 = n20644 & n22445 ;
  assign n22447 = ~n6834 & n8417 ;
  assign n22448 = n22447 ^ n1639 ^ 1'b0 ;
  assign n22449 = x130 & n22448 ;
  assign n22450 = ~x181 & n22449 ;
  assign n22451 = n11266 | n22450 ;
  assign n22452 = n8604 | n22451 ;
  assign n22453 = n16303 & n22452 ;
  assign n22454 = n2463 ^ n397 ^ 1'b0 ;
  assign n22455 = n903 | n2787 ;
  assign n22456 = n17853 & ~n22455 ;
  assign n22457 = ~n7249 & n9643 ;
  assign n22458 = n1521 & ~n10178 ;
  assign n22459 = n6165 ^ n3255 ^ 1'b0 ;
  assign n22460 = x98 & ~n22459 ;
  assign n22461 = ~n10220 & n10511 ;
  assign n22462 = n4079 | n20556 ;
  assign n22463 = ( x26 & ~n13568 ) | ( x26 & n14401 ) | ( ~n13568 & n14401 ) ;
  assign n22464 = n2975 & n9001 ;
  assign n22465 = n5750 & n22464 ;
  assign n22466 = n16832 & n22465 ;
  assign n22467 = n21886 ^ n16396 ^ n5559 ;
  assign n22468 = n15233 & n22467 ;
  assign n22469 = n1679 & ~n4027 ;
  assign n22470 = ~n20248 & n21379 ;
  assign n22471 = ~x61 & n6703 ;
  assign n22472 = n8925 & n22471 ;
  assign n22473 = n6311 & ~n22065 ;
  assign n22474 = ~n14818 & n22473 ;
  assign n22475 = n12288 ^ n8613 ^ n1521 ;
  assign n22476 = ~n22474 & n22475 ;
  assign n22478 = n8907 | n13884 ;
  assign n22477 = n2122 | n7483 ;
  assign n22479 = n22478 ^ n22477 ^ 1'b0 ;
  assign n22482 = n941 | n11356 ;
  assign n22480 = n1980 ^ n1061 ^ 1'b0 ;
  assign n22481 = n22480 ^ n9052 ^ n2765 ;
  assign n22483 = n22482 ^ n22481 ^ 1'b0 ;
  assign n22484 = n754 & n22483 ;
  assign n22485 = ~n1117 & n3959 ;
  assign n22486 = n22485 ^ n6337 ^ 1'b0 ;
  assign n22487 = n8737 & ~n22486 ;
  assign n22488 = ~n2403 & n9152 ;
  assign n22489 = ~n7115 & n22488 ;
  assign n22490 = n14632 | n22489 ;
  assign n22491 = n22490 ^ n10144 ^ 1'b0 ;
  assign n22492 = n21684 ^ n3879 ^ 1'b0 ;
  assign n22493 = n4979 ^ n423 ^ 1'b0 ;
  assign n22494 = n10440 & ~n22493 ;
  assign n22495 = n9869 ^ n4954 ^ 1'b0 ;
  assign n22496 = n1977 | n20647 ;
  assign n22498 = n8747 & n9163 ;
  assign n22497 = n5891 & ~n15618 ;
  assign n22499 = n22498 ^ n22497 ^ 1'b0 ;
  assign n22500 = n13166 ^ n1836 ^ 1'b0 ;
  assign n22501 = n444 & n22500 ;
  assign n22502 = n16024 & n22501 ;
  assign n22503 = n17465 ^ n9588 ^ 1'b0 ;
  assign n22504 = n10861 | n22503 ;
  assign n22505 = n1302 | n7016 ;
  assign n22506 = ~n21934 & n22505 ;
  assign n22507 = n13355 ^ n4541 ^ 1'b0 ;
  assign n22508 = n540 & ~n1820 ;
  assign n22509 = ( x61 & ~n1353 ) | ( x61 & n22508 ) | ( ~n1353 & n22508 ) ;
  assign n22511 = n1291 | n3250 ;
  assign n22510 = n2899 & n2928 ;
  assign n22512 = n22511 ^ n22510 ^ 1'b0 ;
  assign n22513 = n22509 & n22512 ;
  assign n22515 = n10967 | n19109 ;
  assign n22516 = n22515 ^ n11809 ^ 1'b0 ;
  assign n22514 = n13313 & n16817 ;
  assign n22517 = n22516 ^ n22514 ^ 1'b0 ;
  assign n22518 = n18212 ^ x251 ^ 1'b0 ;
  assign n22519 = n1314 & ~n3324 ;
  assign n22520 = ~n1828 & n6553 ;
  assign n22521 = n643 & ~n4291 ;
  assign n22522 = ~n3182 & n6738 ;
  assign n22523 = n22521 & n22522 ;
  assign n22524 = n21480 ^ n9097 ^ 1'b0 ;
  assign n22525 = n11400 ^ n709 ^ 1'b0 ;
  assign n22526 = n4634 & n6681 ;
  assign n22527 = n14632 | n22526 ;
  assign n22528 = ( ~n8324 & n22428 ) | ( ~n8324 & n22527 ) | ( n22428 & n22527 ) ;
  assign n22529 = ~n8314 & n12726 ;
  assign n22530 = ~n967 & n22529 ;
  assign n22531 = n11237 | n22530 ;
  assign n22532 = ~n1240 & n9906 ;
  assign n22533 = ~n8939 & n22532 ;
  assign n22534 = n22533 ^ n6526 ^ n1075 ;
  assign n22535 = ~n1068 & n9018 ;
  assign n22536 = n22535 ^ n6346 ^ 1'b0 ;
  assign n22537 = n20923 & ~n22536 ;
  assign n22538 = n15866 ^ n13657 ^ 1'b0 ;
  assign n22539 = n7124 | n22538 ;
  assign n22540 = n4938 & ~n18905 ;
  assign n22541 = n22540 ^ n4366 ^ 1'b0 ;
  assign n22542 = n1236 ^ x130 ^ 1'b0 ;
  assign n22543 = n1826 ^ n273 ^ 1'b0 ;
  assign n22544 = n6408 | n22543 ;
  assign n22545 = n341 | n22544 ;
  assign n22546 = n698 & ~n22545 ;
  assign n22547 = ~n2536 & n3577 ;
  assign n22548 = ~n3670 & n22547 ;
  assign n22549 = n11738 | n22548 ;
  assign n22550 = n22549 ^ n18507 ^ 1'b0 ;
  assign n22551 = n8217 & ~n11476 ;
  assign n22552 = ~n16160 & n22551 ;
  assign n22553 = n963 | n6368 ;
  assign n22554 = n22552 & ~n22553 ;
  assign n22555 = n4095 & n4402 ;
  assign n22556 = n1094 | n10797 ;
  assign n22557 = n5079 & ~n19938 ;
  assign n22558 = n22556 & ~n22557 ;
  assign n22559 = n3378 & ~n18917 ;
  assign n22560 = n22559 ^ n8528 ^ 1'b0 ;
  assign n22561 = n19925 ^ n4238 ^ 1'b0 ;
  assign n22562 = n20841 ^ n5211 ^ 1'b0 ;
  assign n22563 = n22562 ^ n14863 ^ n2901 ;
  assign n22564 = n19730 ^ n6621 ^ 1'b0 ;
  assign n22565 = n22563 & ~n22564 ;
  assign n22566 = n9029 ^ n6442 ^ 1'b0 ;
  assign n22567 = n1054 & ~n22566 ;
  assign n22568 = n5715 & n9495 ;
  assign n22569 = n4204 & n22568 ;
  assign n22570 = ( ~n10438 & n22567 ) | ( ~n10438 & n22569 ) | ( n22567 & n22569 ) ;
  assign n22571 = n3862 ^ n3397 ^ 1'b0 ;
  assign n22572 = n2485 | n22571 ;
  assign n22573 = n4328 | n22572 ;
  assign n22574 = n4524 & ~n21825 ;
  assign n22575 = n22574 ^ n3152 ^ 1'b0 ;
  assign n22576 = n10331 & n14922 ;
  assign n22577 = n22576 ^ n10130 ^ n9367 ;
  assign n22578 = n22577 ^ n13882 ^ n11110 ;
  assign n22579 = n10953 & ~n22578 ;
  assign n22580 = n15846 ^ n10595 ^ 1'b0 ;
  assign n22581 = n8843 & ~n22580 ;
  assign n22582 = ~n11496 & n14629 ;
  assign n22583 = ~n22581 & n22582 ;
  assign n22584 = n13222 & ~n18422 ;
  assign n22585 = ~n8560 & n13356 ;
  assign n22586 = n1507 & n22585 ;
  assign n22587 = n20915 ^ n401 ^ 1'b0 ;
  assign n22588 = ~n22586 & n22587 ;
  assign n22591 = ( n2935 & n4673 ) | ( n2935 & n4841 ) | ( n4673 & n4841 ) ;
  assign n22592 = n22591 ^ n3257 ^ 1'b0 ;
  assign n22589 = n1622 & ~n19040 ;
  assign n22590 = ~n1622 & n22589 ;
  assign n22593 = n22592 ^ n22590 ^ 1'b0 ;
  assign n22594 = n22593 ^ n2546 ^ 1'b0 ;
  assign n22595 = n895 | n6950 ;
  assign n22596 = n22595 ^ n16861 ^ 1'b0 ;
  assign n22597 = n22594 & ~n22596 ;
  assign n22598 = ~n13386 & n22597 ;
  assign n22599 = x88 | n10561 ;
  assign n22600 = n11377 ^ n4802 ^ 1'b0 ;
  assign n22601 = ~n1638 & n22600 ;
  assign n22602 = x47 & n3533 ;
  assign n22603 = ~x228 & n22602 ;
  assign n22604 = n8281 ^ n6002 ^ 1'b0 ;
  assign n22605 = n22603 | n22604 ;
  assign n22606 = n1507 & ~n11616 ;
  assign n22607 = n22606 ^ n11119 ^ 1'b0 ;
  assign n22608 = n5712 & ~n16989 ;
  assign n22609 = n22608 ^ n4500 ^ 1'b0 ;
  assign n22610 = n22609 ^ n8727 ^ n4347 ;
  assign n22611 = n7688 ^ n700 ^ 1'b0 ;
  assign n22612 = n1256 & ~n19712 ;
  assign n22613 = n22612 ^ n19803 ^ 1'b0 ;
  assign n22614 = n9032 & ~n22613 ;
  assign n22615 = n15825 ^ n7580 ^ 1'b0 ;
  assign n22616 = n1339 | n22615 ;
  assign n22617 = ~n11682 & n19213 ;
  assign n22618 = n12189 & ~n13400 ;
  assign n22619 = n2366 | n3906 ;
  assign n22620 = n6184 | n22619 ;
  assign n22621 = n3074 | n22620 ;
  assign n22622 = n22621 ^ n5695 ^ 1'b0 ;
  assign n22623 = ~n2062 & n22622 ;
  assign n22624 = n16410 ^ n15854 ^ 1'b0 ;
  assign n22625 = n16322 ^ n14980 ^ n9624 ;
  assign n22626 = n1742 | n4209 ;
  assign n22627 = n7572 ^ n3342 ^ 1'b0 ;
  assign n22628 = ~n22626 & n22627 ;
  assign n22629 = n13949 | n16783 ;
  assign n22630 = n3216 ^ n1670 ^ n1198 ;
  assign n22631 = n6644 & ~n22630 ;
  assign n22632 = ~n19710 & n22631 ;
  assign n22633 = n8139 ^ n5002 ^ 1'b0 ;
  assign n22634 = n10459 & n22317 ;
  assign n22635 = n15692 & n22634 ;
  assign n22636 = n22635 ^ n895 ^ 1'b0 ;
  assign n22637 = n12948 & ~n22636 ;
  assign n22638 = n7461 & ~n13911 ;
  assign n22639 = ~n13635 & n22638 ;
  assign n22640 = n4040 & ~n7500 ;
  assign n22641 = n22640 ^ n7936 ^ 1'b0 ;
  assign n22642 = n8312 & ~n22641 ;
  assign n22643 = ~n6297 & n14858 ;
  assign n22644 = ~n22642 & n22643 ;
  assign n22645 = n8233 ^ n5394 ^ 1'b0 ;
  assign n22646 = n1348 | n5381 ;
  assign n22647 = n4871 ^ n3801 ^ 1'b0 ;
  assign n22648 = n5507 & ~n20498 ;
  assign n22649 = n20082 ^ n13331 ^ 1'b0 ;
  assign n22650 = n22648 | n22649 ;
  assign n22651 = n5692 | n16377 ;
  assign n22652 = n22651 ^ n1539 ^ 1'b0 ;
  assign n22653 = n3437 ^ n3174 ^ 1'b0 ;
  assign n22654 = n13547 & n22653 ;
  assign n22655 = n5405 & n9397 ;
  assign n22657 = ~n538 & n6054 ;
  assign n22658 = n22657 ^ n22063 ^ n7051 ;
  assign n22656 = n2042 | n5408 ;
  assign n22659 = n22658 ^ n22656 ^ 1'b0 ;
  assign n22660 = n13532 ^ n285 ^ 1'b0 ;
  assign n22661 = n8554 & n22660 ;
  assign n22664 = ( ~n4821 & n5791 ) | ( ~n4821 & n14436 ) | ( n5791 & n14436 ) ;
  assign n22662 = ~n9752 & n13173 ;
  assign n22663 = n22662 ^ n13775 ^ 1'b0 ;
  assign n22665 = n22664 ^ n22663 ^ n3982 ;
  assign n22670 = n5403 ^ n3136 ^ 1'b0 ;
  assign n22671 = n7347 | n22670 ;
  assign n22666 = ~n1965 & n9222 ;
  assign n22667 = n22666 ^ n4220 ^ 1'b0 ;
  assign n22668 = n5673 & n22667 ;
  assign n22669 = n8332 & n22668 ;
  assign n22672 = n22671 ^ n22669 ^ n6409 ;
  assign n22673 = n17488 ^ n5021 ^ 1'b0 ;
  assign n22674 = n22672 | n22673 ;
  assign n22675 = ~n9590 & n14981 ;
  assign n22676 = n12586 & n22675 ;
  assign n22677 = n22676 ^ n8776 ^ 1'b0 ;
  assign n22678 = ~n17790 & n22677 ;
  assign n22679 = n14852 ^ n4979 ^ 1'b0 ;
  assign n22680 = ~n728 & n22679 ;
  assign n22681 = n9793 ^ n5369 ^ 1'b0 ;
  assign n22682 = n22680 & n22681 ;
  assign n22683 = n6941 | n11119 ;
  assign n22684 = n22683 ^ n6381 ^ 1'b0 ;
  assign n22685 = n22684 ^ n1111 ^ 1'b0 ;
  assign n22686 = n22682 & n22685 ;
  assign n22687 = n11705 ^ n5265 ^ 1'b0 ;
  assign n22688 = ~n15800 & n22687 ;
  assign n22689 = ~n8146 & n8627 ;
  assign n22690 = n22689 ^ n11912 ^ 1'b0 ;
  assign n22691 = n9695 ^ n8474 ^ 1'b0 ;
  assign n22692 = n723 & n22691 ;
  assign n22693 = n22692 ^ n14356 ^ n3065 ;
  assign n22694 = n3065 ^ n2379 ^ 1'b0 ;
  assign n22695 = n7428 ^ n3480 ^ 1'b0 ;
  assign n22696 = n12911 & ~n22695 ;
  assign n22697 = n22696 ^ n9371 ^ 1'b0 ;
  assign n22698 = n6647 ^ n4408 ^ 1'b0 ;
  assign n22699 = ~n10886 & n22698 ;
  assign n22700 = n22699 ^ n4122 ^ 1'b0 ;
  assign n22701 = n10757 | n21113 ;
  assign n22702 = n4850 & n22002 ;
  assign n22703 = n10014 ^ n1076 ^ 1'b0 ;
  assign n22704 = n22702 & n22703 ;
  assign n22705 = ( n1286 & n2752 ) | ( n1286 & ~n5781 ) | ( n2752 & ~n5781 ) ;
  assign n22706 = n13157 & n14981 ;
  assign n22707 = n2455 & ~n2670 ;
  assign n22708 = n22707 ^ n16062 ^ 1'b0 ;
  assign n22709 = n2629 & n22708 ;
  assign n22710 = n5146 ^ n4574 ^ 1'b0 ;
  assign n22711 = n11237 | n22710 ;
  assign n22712 = n22711 ^ n7421 ^ 1'b0 ;
  assign n22713 = ~n18900 & n22712 ;
  assign n22714 = n17905 ^ n11226 ^ 1'b0 ;
  assign n22715 = n12429 & n16102 ;
  assign n22716 = n4413 | n22017 ;
  assign n22717 = n22715 | n22716 ;
  assign n22718 = n10715 ^ n6443 ^ n1181 ;
  assign n22719 = n14652 ^ n8333 ^ n1533 ;
  assign n22720 = n2351 & ~n22719 ;
  assign n22721 = n1890 | n3856 ;
  assign n22722 = n2216 ^ n1360 ^ 1'b0 ;
  assign n22723 = n5595 | n22722 ;
  assign n22724 = ~n8890 & n12963 ;
  assign n22725 = ~n14895 & n22724 ;
  assign n22726 = n875 & ~n22725 ;
  assign n22727 = n13863 ^ n10777 ^ 1'b0 ;
  assign n22728 = n3127 & n22727 ;
  assign n22729 = x106 & ~n22728 ;
  assign n22730 = n9060 & ~n22729 ;
  assign n22731 = n22730 ^ n9902 ^ 1'b0 ;
  assign n22732 = ~n562 & n17804 ;
  assign n22733 = n1387 & n22732 ;
  assign n22734 = ~n13820 & n16208 ;
  assign n22735 = n22733 & n22734 ;
  assign n22736 = ~n2578 & n22482 ;
  assign n22737 = n8657 ^ n2438 ^ 1'b0 ;
  assign n22738 = ~n3381 & n22737 ;
  assign n22739 = n6006 & n13066 ;
  assign n22740 = n9223 & n22739 ;
  assign n22741 = ( n7527 & n9682 ) | ( n7527 & n22740 ) | ( n9682 & n22740 ) ;
  assign n22742 = n1540 & ~n5700 ;
  assign n22743 = n22742 ^ n5133 ^ 1'b0 ;
  assign n22744 = n710 & n8097 ;
  assign n22746 = n2974 ^ n2547 ^ 1'b0 ;
  assign n22747 = ( n546 & n1568 ) | ( n546 & n22746 ) | ( n1568 & n22746 ) ;
  assign n22748 = n22747 ^ n10306 ^ 1'b0 ;
  assign n22745 = n18835 & n20285 ;
  assign n22749 = n22748 ^ n22745 ^ 1'b0 ;
  assign n22750 = ~x244 & n21293 ;
  assign n22751 = n4414 ^ n1815 ^ 1'b0 ;
  assign n22752 = ~n22750 & n22751 ;
  assign n22753 = ~n14613 & n22752 ;
  assign n22756 = n10070 ^ n3383 ^ 1'b0 ;
  assign n22754 = n8006 ^ n4256 ^ 1'b0 ;
  assign n22755 = n5529 & n22754 ;
  assign n22757 = n22756 ^ n22755 ^ n2669 ;
  assign n22758 = n6677 | n22757 ;
  assign n22759 = n16293 & n17836 ;
  assign n22760 = n10771 | n20801 ;
  assign n22761 = n22760 ^ n10076 ^ n1399 ;
  assign n22762 = n6283 & n22761 ;
  assign n22763 = n3073 & n7634 ;
  assign n22764 = n15214 & n22763 ;
  assign n22765 = n19316 & ~n22764 ;
  assign n22766 = n22765 ^ n9351 ^ 1'b0 ;
  assign n22767 = n4903 ^ n3920 ^ 1'b0 ;
  assign n22768 = n22766 & ~n22767 ;
  assign n22769 = n22768 ^ n21882 ^ 1'b0 ;
  assign n22770 = n5978 ^ n1684 ^ 1'b0 ;
  assign n22771 = n2955 | n18534 ;
  assign n22772 = n17015 ^ n13348 ^ 1'b0 ;
  assign n22773 = n10993 & n13538 ;
  assign n22774 = n22773 ^ n5824 ^ 1'b0 ;
  assign n22775 = n1507 & ~n7984 ;
  assign n22776 = ~n9503 & n22775 ;
  assign n22777 = n22776 ^ n15436 ^ 1'b0 ;
  assign n22778 = ~n22774 & n22777 ;
  assign n22779 = n1321 & ~n17073 ;
  assign n22780 = n12118 & ~n15007 ;
  assign n22781 = ( n6724 & ~n18895 ) | ( n6724 & n22076 ) | ( ~n18895 & n22076 ) ;
  assign n22782 = n22781 ^ n16807 ^ 1'b0 ;
  assign n22783 = n2761 | n20174 ;
  assign n22784 = n6213 ^ n2361 ^ 1'b0 ;
  assign n22785 = n7466 ^ n5503 ^ 1'b0 ;
  assign n22786 = n15224 & ~n22785 ;
  assign n22787 = n9988 ^ n6375 ^ 1'b0 ;
  assign n22788 = n1903 & n5806 ;
  assign n22789 = n22788 ^ n8068 ^ 1'b0 ;
  assign n22790 = n1152 | n12346 ;
  assign n22791 = n6012 | n22790 ;
  assign n22792 = n22789 & n22791 ;
  assign n22793 = ~n16206 & n22792 ;
  assign n22794 = n6740 ^ n315 ^ 1'b0 ;
  assign n22795 = n22794 ^ n19175 ^ 1'b0 ;
  assign n22796 = n4024 & ~n4051 ;
  assign n22797 = n11851 ^ n10477 ^ 1'b0 ;
  assign n22798 = n6962 ^ n4661 ^ 1'b0 ;
  assign n22799 = n6189 | n21435 ;
  assign n22800 = n22798 & ~n22799 ;
  assign n22801 = n2289 | n11007 ;
  assign n22802 = ~n11013 & n22801 ;
  assign n22803 = n18599 ^ n11508 ^ 1'b0 ;
  assign n22804 = n22181 ^ n1859 ^ 1'b0 ;
  assign n22805 = n2939 & ~n19735 ;
  assign n22806 = n13717 ^ x14 ^ 1'b0 ;
  assign n22807 = n22805 & ~n22806 ;
  assign n22808 = ( ~n3740 & n3901 ) | ( ~n3740 & n4776 ) | ( n3901 & n4776 ) ;
  assign n22809 = n3852 ^ n1931 ^ 1'b0 ;
  assign n22810 = n3083 | n6333 ;
  assign n22811 = n19622 | n22810 ;
  assign n22812 = n15187 ^ n7259 ^ 1'b0 ;
  assign n22813 = n11331 | n22812 ;
  assign n22814 = ( n9929 & n14889 ) | ( n9929 & ~n22813 ) | ( n14889 & ~n22813 ) ;
  assign n22815 = n2358 | n10539 ;
  assign n22817 = ~n2106 & n2507 ;
  assign n22818 = n22817 ^ n7940 ^ 1'b0 ;
  assign n22819 = n4313 | n22818 ;
  assign n22820 = n715 | n22819 ;
  assign n22816 = n21432 & n21810 ;
  assign n22821 = n22820 ^ n22816 ^ 1'b0 ;
  assign n22822 = n505 & n3694 ;
  assign n22823 = n22822 ^ n6058 ^ 1'b0 ;
  assign n22824 = ~n4130 & n22823 ;
  assign n22825 = n22824 ^ n6771 ^ 1'b0 ;
  assign n22826 = ~n1283 & n2629 ;
  assign n22827 = n3666 & n22826 ;
  assign n22829 = ~n2270 & n9304 ;
  assign n22828 = x81 & ~n6764 ;
  assign n22830 = n22829 ^ n22828 ^ 1'b0 ;
  assign n22831 = n7915 | n22830 ;
  assign n22832 = n22831 ^ x248 ^ 1'b0 ;
  assign n22833 = n22832 ^ n7261 ^ 1'b0 ;
  assign n22834 = n13863 | n17947 ;
  assign n22838 = n3798 | n4605 ;
  assign n22836 = n5955 ^ n3768 ^ 1'b0 ;
  assign n22837 = ~n22401 & n22836 ;
  assign n22839 = n22838 ^ n22837 ^ 1'b0 ;
  assign n22835 = n7915 ^ n6496 ^ 1'b0 ;
  assign n22840 = n22839 ^ n22835 ^ n3342 ;
  assign n22841 = n21799 ^ n2187 ^ 1'b0 ;
  assign n22842 = n12887 ^ n3917 ^ 1'b0 ;
  assign n22843 = ~n2589 & n7358 ;
  assign n22844 = ~n22842 & n22843 ;
  assign n22845 = ~n1217 & n6954 ;
  assign n22846 = n3458 | n3751 ;
  assign n22847 = ( ~n10433 & n20454 ) | ( ~n10433 & n22846 ) | ( n20454 & n22846 ) ;
  assign n22848 = n8165 & ~n13619 ;
  assign n22849 = n22848 ^ n1443 ^ 1'b0 ;
  assign n22850 = n4506 | n22849 ;
  assign n22851 = ~n16911 & n22850 ;
  assign n22852 = ~n8997 & n22851 ;
  assign n22853 = x250 & ~n608 ;
  assign n22854 = n608 & n22853 ;
  assign n22855 = n1831 & ~n22854 ;
  assign n22856 = n22854 & n22855 ;
  assign n22857 = n2406 & n22856 ;
  assign n22858 = n444 & ~n4382 ;
  assign n22859 = ~n444 & n22858 ;
  assign n22860 = n10758 & ~n22859 ;
  assign n22861 = n22857 & n22860 ;
  assign n22862 = ~n1630 & n22861 ;
  assign n22863 = n9438 | n22862 ;
  assign n22864 = ~n3998 & n13626 ;
  assign n22865 = n3998 & n22864 ;
  assign n22866 = n22863 & ~n22865 ;
  assign n22867 = ~n22863 & n22866 ;
  assign n22868 = n3926 & n21492 ;
  assign n22869 = n10140 ^ n1381 ^ 1'b0 ;
  assign n22870 = n13523 ^ n5916 ^ 1'b0 ;
  assign n22871 = n4351 & n8016 ;
  assign n22872 = ~n6368 & n22871 ;
  assign n22873 = n700 & n7691 ;
  assign n22874 = n22873 ^ n22819 ^ 1'b0 ;
  assign n22875 = n22874 ^ n5885 ^ 1'b0 ;
  assign n22876 = n2307 & ~n22875 ;
  assign n22877 = n12729 | n22876 ;
  assign n22878 = n1507 ^ n963 ^ 1'b0 ;
  assign n22879 = n12389 | n22878 ;
  assign n22880 = n10126 & n22879 ;
  assign n22881 = ~n9892 & n16285 ;
  assign n22882 = ~n7136 & n11815 ;
  assign n22885 = ~n2793 & n3880 ;
  assign n22883 = ( n2895 & n3308 ) | ( n2895 & ~n3621 ) | ( n3308 & ~n3621 ) ;
  assign n22884 = n5496 & ~n22883 ;
  assign n22886 = n22885 ^ n22884 ^ 1'b0 ;
  assign n22887 = n5347 | n7199 ;
  assign n22888 = x64 & ~n9351 ;
  assign n22889 = ~n22887 & n22888 ;
  assign n22890 = ~x220 & n7739 ;
  assign n22891 = n18119 & n22890 ;
  assign n22892 = n6574 ^ n5457 ^ 1'b0 ;
  assign n22893 = n22891 | n22892 ;
  assign n22894 = n16019 | n20805 ;
  assign n22895 = n5316 ^ n3597 ^ n1588 ;
  assign n22896 = ~n3933 & n22895 ;
  assign n22897 = n22896 ^ n3270 ^ 1'b0 ;
  assign n22898 = n6750 & n14406 ;
  assign n22899 = n2392 & n8571 ;
  assign n22900 = n22898 | n22899 ;
  assign n22901 = ~n6118 & n8553 ;
  assign n22902 = n10000 & n14587 ;
  assign n22903 = n14303 & n22902 ;
  assign n22904 = n8208 & ~n20820 ;
  assign n22905 = n22904 ^ n3128 ^ 1'b0 ;
  assign n22906 = ~n2566 & n9797 ;
  assign n22907 = n9362 & n17159 ;
  assign n22908 = n5673 & n19207 ;
  assign n22909 = n22908 ^ n6872 ^ 1'b0 ;
  assign n22910 = n10487 | n22909 ;
  assign n22911 = n9072 | n22910 ;
  assign n22912 = n964 | n22911 ;
  assign n22913 = n12204 ^ n7194 ^ 1'b0 ;
  assign n22914 = n9109 & ~n22913 ;
  assign n22915 = ~n8435 & n22914 ;
  assign n22916 = n2085 & n7212 ;
  assign n22917 = n3567 ^ n3423 ^ 1'b0 ;
  assign n22918 = n818 & ~n22917 ;
  assign n22919 = n22916 & n22918 ;
  assign n22920 = n18770 & ~n22919 ;
  assign n22921 = n16728 & n22920 ;
  assign n22922 = n2686 | n4705 ;
  assign n22923 = n17168 & ~n21919 ;
  assign n22924 = x211 & n9402 ;
  assign n22925 = n22924 ^ n13929 ^ 1'b0 ;
  assign n22926 = n859 & n4454 ;
  assign n22927 = ( n11213 & n22925 ) | ( n11213 & ~n22926 ) | ( n22925 & ~n22926 ) ;
  assign n22928 = ~n3158 & n20687 ;
  assign n22929 = ( n366 & ~n12686 ) | ( n366 & n21407 ) | ( ~n12686 & n21407 ) ;
  assign n22930 = n1885 ^ n1027 ^ 1'b0 ;
  assign n22931 = n2760 & n8875 ;
  assign n22932 = n22931 ^ n974 ^ 1'b0 ;
  assign n22933 = n6584 | n13317 ;
  assign n22934 = n22932 | n22933 ;
  assign n22935 = n22934 ^ n10002 ^ 1'b0 ;
  assign n22936 = n9345 | n22935 ;
  assign n22937 = n4213 & n15909 ;
  assign n22938 = n19445 ^ n13798 ^ 1'b0 ;
  assign n22939 = n8283 | n13965 ;
  assign n22940 = n10164 | n17130 ;
  assign n22942 = n17095 ^ n1435 ^ 1'b0 ;
  assign n22943 = ~n18990 & n22942 ;
  assign n22941 = n5926 | n22387 ;
  assign n22944 = n22943 ^ n22941 ^ 1'b0 ;
  assign n22945 = ~n2697 & n9001 ;
  assign n22946 = n4172 & ~n19747 ;
  assign n22947 = ~n4451 & n22946 ;
  assign n22948 = n22947 ^ n21265 ^ n2725 ;
  assign n22949 = ~n1630 & n22948 ;
  assign n22950 = ~n10886 & n22949 ;
  assign n22951 = n1685 & ~n7569 ;
  assign n22952 = n22951 ^ n5144 ^ 1'b0 ;
  assign n22953 = x170 & ~n1503 ;
  assign n22954 = n22953 ^ n14481 ^ 1'b0 ;
  assign n22955 = n2006 & n12250 ;
  assign n22956 = n15436 ^ n4214 ^ 1'b0 ;
  assign n22957 = n15193 | n22956 ;
  assign n22958 = n1130 | n2668 ;
  assign n22959 = n4107 | n22958 ;
  assign n22960 = n3915 & n9978 ;
  assign n22961 = n1441 & n8708 ;
  assign n22962 = n22961 ^ x123 ^ 1'b0 ;
  assign n22963 = n18877 & ~n22962 ;
  assign n22964 = n2632 | n3419 ;
  assign n22965 = n22964 ^ n11462 ^ n1199 ;
  assign n22966 = n16297 ^ n10169 ^ 1'b0 ;
  assign n22967 = n1871 | n22966 ;
  assign n22968 = ( n3601 & ~n13273 ) | ( n3601 & n16174 ) | ( ~n13273 & n16174 ) ;
  assign n22969 = n22968 ^ n13644 ^ 1'b0 ;
  assign n22970 = n7421 | n22969 ;
  assign n22971 = n8704 & n13155 ;
  assign n22972 = n22971 ^ n3408 ^ 1'b0 ;
  assign n22973 = n15388 & ~n22972 ;
  assign n22974 = n10981 & ~n15302 ;
  assign n22975 = n22974 ^ n8760 ^ 1'b0 ;
  assign n22977 = n3676 | n8242 ;
  assign n22976 = n3227 & n6145 ;
  assign n22978 = n22977 ^ n22976 ^ 1'b0 ;
  assign n22979 = n16627 ^ n15054 ^ 1'b0 ;
  assign n22980 = n7100 | n22979 ;
  assign n22981 = n679 & ~n22980 ;
  assign n22982 = n467 & n11964 ;
  assign n22983 = n11074 & ~n22982 ;
  assign n22984 = n5896 | n13742 ;
  assign n22993 = n781 | n11945 ;
  assign n22988 = x65 & n978 ;
  assign n22989 = n22988 ^ n3359 ^ 1'b0 ;
  assign n22990 = n22989 ^ n11482 ^ 1'b0 ;
  assign n22991 = n5237 & n22990 ;
  assign n22985 = n2180 & n6945 ;
  assign n22986 = n1395 & n22985 ;
  assign n22987 = n1366 | n22986 ;
  assign n22992 = n22991 ^ n22987 ^ 1'b0 ;
  assign n22994 = n22993 ^ n22992 ^ n926 ;
  assign n22995 = n275 | n20194 ;
  assign n22996 = n18606 ^ x19 ^ 1'b0 ;
  assign n22997 = n22068 ^ n6172 ^ 1'b0 ;
  assign n22998 = ~n808 & n3746 ;
  assign n22999 = ~n15651 & n22998 ;
  assign n23000 = n3989 | n4400 ;
  assign n23001 = ~n22999 & n23000 ;
  assign n23002 = n16140 ^ n2527 ^ 1'b0 ;
  assign n23003 = n21111 & ~n23002 ;
  assign n23004 = n5907 & n5928 ;
  assign n23005 = n9279 | n23004 ;
  assign n23006 = ~n7051 & n10682 ;
  assign n23007 = n3995 & n7753 ;
  assign n23008 = n23006 & n23007 ;
  assign n23009 = n13051 & ~n23008 ;
  assign n23010 = n23009 ^ n7061 ^ 1'b0 ;
  assign n23011 = n741 | n20799 ;
  assign n23012 = n14639 ^ n4238 ^ n1736 ;
  assign n23013 = n1569 | n23012 ;
  assign n23014 = n22288 ^ n10305 ^ 1'b0 ;
  assign n23015 = ~n4694 & n13884 ;
  assign n23016 = n20555 | n23015 ;
  assign n23017 = n23016 ^ n8767 ^ 1'b0 ;
  assign n23018 = n8390 & ~n23017 ;
  assign n23019 = ~n5376 & n7352 ;
  assign n23020 = n562 & n23019 ;
  assign n23021 = n12914 ^ n4490 ^ n2264 ;
  assign n23022 = n23021 ^ n18157 ^ x53 ;
  assign n23023 = n6560 | n18608 ;
  assign n23024 = ~n1952 & n2786 ;
  assign n23025 = n22889 ^ n9880 ^ 1'b0 ;
  assign n23026 = n6409 ^ n981 ^ 1'b0 ;
  assign n23027 = n8054 | n23026 ;
  assign n23028 = ~n696 & n6496 ;
  assign n23029 = ~n14198 & n23028 ;
  assign n23030 = n5715 | n23029 ;
  assign n23031 = n23027 & n23030 ;
  assign n23032 = n23031 ^ n10296 ^ 1'b0 ;
  assign n23033 = n23032 ^ n13149 ^ 1'b0 ;
  assign n23034 = ~x226 & n23033 ;
  assign n23035 = ~n8005 & n10491 ;
  assign n23036 = n23035 ^ n3324 ^ 1'b0 ;
  assign n23037 = n7844 & ~n23036 ;
  assign n23038 = n18070 ^ n2113 ^ 1'b0 ;
  assign n23039 = n2472 | n2922 ;
  assign n23040 = n10658 ^ n5864 ^ 1'b0 ;
  assign n23041 = n23039 & n23040 ;
  assign n23042 = n6207 ^ n3171 ^ 1'b0 ;
  assign n23043 = n16399 & n23042 ;
  assign n23044 = n23043 ^ n387 ^ 1'b0 ;
  assign n23045 = n10371 & ~n22035 ;
  assign n23046 = n15664 ^ n3466 ^ 1'b0 ;
  assign n23047 = n12429 ^ n1538 ^ 1'b0 ;
  assign n23048 = ~n23046 & n23047 ;
  assign n23049 = n23048 ^ n3078 ^ 1'b0 ;
  assign n23050 = n19421 & ~n23049 ;
  assign n23051 = n1463 & ~n2116 ;
  assign n23052 = ~n17549 & n23051 ;
  assign n23053 = n23052 ^ n11532 ^ 1'b0 ;
  assign n23054 = ~n10259 & n16102 ;
  assign n23055 = n22746 & n23054 ;
  assign n23056 = x10 & ~n11519 ;
  assign n23057 = n23056 ^ n14168 ^ 1'b0 ;
  assign n23058 = n3901 & ~n17447 ;
  assign n23059 = n1880 | n23058 ;
  assign n23060 = n10552 ^ n3621 ^ 1'b0 ;
  assign n23061 = n6295 & ~n14170 ;
  assign n23062 = n23061 ^ n21685 ^ 1'b0 ;
  assign n23063 = n3389 ^ n3027 ^ 1'b0 ;
  assign n23064 = n4493 | n17056 ;
  assign n23065 = n4714 | n22073 ;
  assign n23066 = n6026 & ~n11775 ;
  assign n23067 = n23065 & n23066 ;
  assign n23068 = n3888 | n10991 ;
  assign n23069 = n23068 ^ n9331 ^ 1'b0 ;
  assign n23070 = n22226 ^ n5744 ^ x81 ;
  assign n23071 = n9627 | n9741 ;
  assign n23072 = n20007 ^ n8854 ^ 1'b0 ;
  assign n23073 = n22570 & n23072 ;
  assign n23074 = n1324 & n23073 ;
  assign n23075 = n17357 ^ n13113 ^ 1'b0 ;
  assign n23076 = n12749 & ~n23075 ;
  assign n23077 = ~n8190 & n8223 ;
  assign n23078 = n20134 ^ n8089 ^ n2541 ;
  assign n23079 = n659 | n3675 ;
  assign n23080 = n19523 & ~n23079 ;
  assign n23081 = n6651 & n9769 ;
  assign n23082 = ~n4238 & n23081 ;
  assign n23083 = n23080 & n23082 ;
  assign n23084 = n5799 | n8205 ;
  assign n23085 = n1243 | n1546 ;
  assign n23086 = n1546 & ~n23085 ;
  assign n23087 = n5568 & ~n23086 ;
  assign n23088 = n23086 & n23087 ;
  assign n23089 = n23088 ^ n15546 ^ 1'b0 ;
  assign n23090 = n23084 & ~n23089 ;
  assign n23091 = n294 | n15640 ;
  assign n23092 = n9158 & ~n23091 ;
  assign n23093 = n17349 | n23092 ;
  assign n23094 = n23090 | n23093 ;
  assign n23095 = ~n10183 & n20832 ;
  assign n23096 = n12972 ^ n1066 ^ 1'b0 ;
  assign n23097 = n9386 & n23096 ;
  assign n23098 = ( n2333 & n4409 ) | ( n2333 & n11694 ) | ( n4409 & n11694 ) ;
  assign n23099 = n17186 ^ n15005 ^ 1'b0 ;
  assign n23100 = n7022 & ~n23099 ;
  assign n23101 = n3013 | n5173 ;
  assign n23102 = ~n21093 & n23101 ;
  assign n23103 = ~n23100 & n23102 ;
  assign n23104 = n3759 ^ n1770 ^ 1'b0 ;
  assign n23105 = n13330 & ~n23104 ;
  assign n23106 = n8729 & n12849 ;
  assign n23107 = n1435 | n9018 ;
  assign n23108 = ~n729 & n1131 ;
  assign n23109 = ~n1131 & n23108 ;
  assign n23110 = n372 & n1054 ;
  assign n23111 = ~n1054 & n23110 ;
  assign n23112 = n1251 & n23111 ;
  assign n23113 = ~n7130 & n23112 ;
  assign n23114 = n797 & ~n934 ;
  assign n23115 = n934 & n23114 ;
  assign n23116 = n3314 & ~n7400 ;
  assign n23117 = ~n3314 & n23116 ;
  assign n23118 = n23115 | n23117 ;
  assign n23119 = n23113 | n23118 ;
  assign n23120 = ~n23109 & n23119 ;
  assign n23121 = n23109 & n23120 ;
  assign n23122 = n15487 ^ n7246 ^ 1'b0 ;
  assign n23123 = n2391 | n4154 ;
  assign n23124 = n23123 ^ n16308 ^ 1'b0 ;
  assign n23125 = n6494 ^ n5300 ^ 1'b0 ;
  assign n23126 = n11945 & n23125 ;
  assign n23127 = n23126 ^ n405 ^ 1'b0 ;
  assign n23128 = ~n12536 & n23127 ;
  assign n23129 = n23128 ^ n521 ^ 1'b0 ;
  assign n23130 = ~n1018 & n13943 ;
  assign n23131 = x58 & ~n7716 ;
  assign n23132 = n23131 ^ n7204 ^ 1'b0 ;
  assign n23133 = n23132 ^ n18782 ^ n4664 ;
  assign n23134 = n2772 & ~n4695 ;
  assign n23135 = n2179 & n23134 ;
  assign n23136 = n23135 ^ n4414 ^ 1'b0 ;
  assign n23137 = n16219 ^ n3143 ^ 1'b0 ;
  assign n23138 = n23137 ^ n4478 ^ 1'b0 ;
  assign n23139 = n9592 | n18870 ;
  assign n23140 = n3939 | n5419 ;
  assign n23141 = n23140 ^ n564 ^ 1'b0 ;
  assign n23142 = ~n977 & n8939 ;
  assign n23143 = n23142 ^ n1485 ^ 1'b0 ;
  assign n23144 = n11258 ^ n6842 ^ 1'b0 ;
  assign n23145 = n23144 ^ n14773 ^ 1'b0 ;
  assign n23146 = ~n19070 & n23145 ;
  assign n23147 = n11469 ^ n981 ^ 1'b0 ;
  assign n23148 = n6288 & ~n23147 ;
  assign n23149 = n17018 ^ n6039 ^ n5838 ;
  assign n23150 = n22364 ^ n6933 ^ 1'b0 ;
  assign n23151 = ~n17695 & n23150 ;
  assign n23152 = ~n23149 & n23151 ;
  assign n23153 = ~n4048 & n23152 ;
  assign n23154 = n2376 | n14490 ;
  assign n23155 = ( x23 & ~n14652 ) | ( x23 & n15172 ) | ( ~n14652 & n15172 ) ;
  assign n23156 = n8283 ^ n6840 ^ 1'b0 ;
  assign n23157 = n1018 & ~n23156 ;
  assign n23158 = n23157 ^ n381 ^ 1'b0 ;
  assign n23159 = n13913 | n21627 ;
  assign n23160 = n23159 ^ n4584 ^ 1'b0 ;
  assign n23161 = ~n23158 & n23160 ;
  assign n23162 = n296 ^ x56 ^ 1'b0 ;
  assign n23163 = ~n6969 & n16129 ;
  assign n23164 = ~n23162 & n23163 ;
  assign n23165 = ~x245 & n13075 ;
  assign n23166 = ~n6710 & n13009 ;
  assign n23167 = n23166 ^ n3796 ^ 1'b0 ;
  assign n23168 = ~x93 & n1111 ;
  assign n23169 = x93 & n23168 ;
  assign n23170 = n3765 & n23169 ;
  assign n23171 = ~n832 & n23170 ;
  assign n23172 = n832 & n23171 ;
  assign n23173 = n1906 & ~n5542 ;
  assign n23174 = n16258 & n23173 ;
  assign n23175 = x23 & ~n23174 ;
  assign n23176 = n23174 & n23175 ;
  assign n23177 = n5590 & ~n23176 ;
  assign n23178 = n23176 & n23177 ;
  assign n23179 = n7583 & ~n23178 ;
  assign n23180 = n23178 & n23179 ;
  assign n23181 = n23172 | n23180 ;
  assign n23182 = n23172 & ~n23181 ;
  assign n23183 = n22647 & ~n23182 ;
  assign n23184 = ( n13360 & n23167 ) | ( n13360 & ~n23183 ) | ( n23167 & ~n23183 ) ;
  assign n23185 = n13613 ^ n10513 ^ 1'b0 ;
  assign n23186 = n21944 & ~n22808 ;
  assign n23187 = n11385 & n23186 ;
  assign n23188 = n5266 ^ n2737 ^ 1'b0 ;
  assign n23189 = ~n10022 & n23188 ;
  assign n23190 = n23189 ^ n3973 ^ 1'b0 ;
  assign n23191 = ~n19924 & n23190 ;
  assign n23192 = ~n12310 & n16130 ;
  assign n23194 = n6823 ^ x113 ^ 1'b0 ;
  assign n23193 = n15081 ^ n746 ^ 1'b0 ;
  assign n23195 = n23194 ^ n23193 ^ n14481 ;
  assign n23198 = n20194 ^ n7706 ^ 1'b0 ;
  assign n23199 = ~n10314 & n23198 ;
  assign n23196 = n1970 | n15814 ;
  assign n23197 = n13175 & ~n23196 ;
  assign n23200 = n23199 ^ n23197 ^ 1'b0 ;
  assign n23201 = n4274 ^ n1304 ^ 1'b0 ;
  assign n23202 = n21682 ^ n18405 ^ 1'b0 ;
  assign n23205 = n1528 & ~n3158 ;
  assign n23206 = n1059 & n23205 ;
  assign n23203 = n10397 & n15224 ;
  assign n23204 = n23203 ^ n6198 ^ 1'b0 ;
  assign n23207 = n23206 ^ n23204 ^ 1'b0 ;
  assign n23208 = ~n1021 & n8947 ;
  assign n23209 = n583 & ~n1703 ;
  assign n23210 = ~n16941 & n23209 ;
  assign n23211 = n23210 ^ n17758 ^ 1'b0 ;
  assign n23212 = n23208 & n23211 ;
  assign n23213 = n23212 ^ n2505 ^ 1'b0 ;
  assign n23214 = ~n838 & n3242 ;
  assign n23215 = n6026 & ~n23214 ;
  assign n23216 = n23215 ^ n9786 ^ 1'b0 ;
  assign n23217 = n628 | n12576 ;
  assign n23218 = n10887 ^ n2057 ^ 1'b0 ;
  assign n23219 = n10396 & n23218 ;
  assign n23220 = n6296 ^ n527 ^ 1'b0 ;
  assign n23221 = n12170 & ~n23220 ;
  assign n23222 = n23221 ^ n8818 ^ 1'b0 ;
  assign n23223 = n4552 & n23222 ;
  assign n23224 = n4949 & n23223 ;
  assign n23225 = ( n4524 & n10915 ) | ( n4524 & ~n10965 ) | ( n10915 & ~n10965 ) ;
  assign n23226 = n2643 | n4578 ;
  assign n23227 = n3349 | n23226 ;
  assign n23228 = n23227 ^ n4324 ^ 1'b0 ;
  assign n23229 = n4253 & ~n11775 ;
  assign n23230 = n23228 & n23229 ;
  assign n23231 = ~n436 & n11808 ;
  assign n23232 = n23231 ^ n2500 ^ 1'b0 ;
  assign n23233 = n343 & n1042 ;
  assign n23234 = n23233 ^ n7625 ^ 1'b0 ;
  assign n23235 = ~n1245 & n22631 ;
  assign n23236 = n14324 & ~n16333 ;
  assign n23237 = n4678 & ~n17432 ;
  assign n23239 = n1877 & ~n20882 ;
  assign n23240 = n23239 ^ n1691 ^ 1'b0 ;
  assign n23238 = n4021 | n18754 ;
  assign n23241 = n23240 ^ n23238 ^ 1'b0 ;
  assign n23242 = n734 | n13899 ;
  assign n23243 = n10002 ^ n7066 ^ 1'b0 ;
  assign n23244 = n4084 & ~n23243 ;
  assign n23245 = n23244 ^ n11972 ^ 1'b0 ;
  assign n23246 = ~n6527 & n23245 ;
  assign n23247 = ~n2443 & n23246 ;
  assign n23248 = n5091 ^ n3046 ^ 1'b0 ;
  assign n23249 = n333 & n5583 ;
  assign n23250 = ~n5903 & n19035 ;
  assign n23251 = n6437 & n23250 ;
  assign n23252 = n23251 ^ n8901 ^ 1'b0 ;
  assign n23253 = n1393 & n7000 ;
  assign n23254 = n23253 ^ n2309 ^ 1'b0 ;
  assign n23255 = n3886 & ~n23206 ;
  assign n23256 = n23254 & n23255 ;
  assign n23257 = n18622 ^ n7627 ^ 1'b0 ;
  assign n23258 = ~n9432 & n23257 ;
  assign n23259 = n2667 & ~n15322 ;
  assign n23260 = ~n12579 & n23259 ;
  assign n23261 = n15235 | n23260 ;
  assign n23262 = n23261 ^ n6981 ^ 1'b0 ;
  assign n23263 = n7700 ^ n6250 ^ 1'b0 ;
  assign n23264 = n2116 | n14139 ;
  assign n23265 = n5120 & ~n5850 ;
  assign n23266 = ~n18555 & n23265 ;
  assign n23267 = n23266 ^ n2306 ^ 1'b0 ;
  assign n23268 = ~n18677 & n19107 ;
  assign n23269 = ~n15743 & n23268 ;
  assign n23270 = n4785 & n8613 ;
  assign n23272 = n2766 ^ n807 ^ 1'b0 ;
  assign n23273 = ~n966 & n23272 ;
  assign n23271 = n2582 & ~n18536 ;
  assign n23274 = n23273 ^ n23271 ^ 1'b0 ;
  assign n23275 = n345 & ~n1854 ;
  assign n23276 = n23275 ^ n15591 ^ 1'b0 ;
  assign n23277 = n2768 & n23276 ;
  assign n23278 = n4602 | n6036 ;
  assign n23279 = n1681 & ~n23278 ;
  assign n23280 = n23279 ^ n11299 ^ n3197 ;
  assign n23281 = n7693 | n23280 ;
  assign n23282 = n19462 ^ n10336 ^ 1'b0 ;
  assign n23283 = n23281 & ~n23282 ;
  assign n23284 = n11472 & n23283 ;
  assign n23285 = n9989 | n22312 ;
  assign n23286 = n3059 | n18148 ;
  assign n23287 = n21658 ^ n12115 ^ 1'b0 ;
  assign n23288 = ~n15216 & n23287 ;
  assign n23289 = n10123 ^ n5809 ^ 1'b0 ;
  assign n23290 = n5593 & ~n23097 ;
  assign n23291 = n23290 ^ n19253 ^ 1'b0 ;
  assign n23292 = n6516 & ~n13081 ;
  assign n23293 = n23292 ^ n503 ^ 1'b0 ;
  assign n23294 = n17907 ^ n3905 ^ 1'b0 ;
  assign n23295 = ~n21066 & n23294 ;
  assign n23296 = n3097 & n15516 ;
  assign n23297 = n5382 & n23296 ;
  assign n23298 = n2744 ^ n1272 ^ 1'b0 ;
  assign n23299 = n23297 | n23298 ;
  assign n23300 = n841 & n20582 ;
  assign n23301 = ~x222 & n1731 ;
  assign n23302 = n23300 & n23301 ;
  assign n23303 = n23302 ^ n17551 ^ 1'b0 ;
  assign n23304 = ~n3219 & n3551 ;
  assign n23305 = n23304 ^ n3527 ^ 1'b0 ;
  assign n23306 = n9894 & n10994 ;
  assign n23307 = ~n21356 & n23306 ;
  assign n23308 = n23307 ^ n3473 ^ 1'b0 ;
  assign n23309 = x19 & n4638 ;
  assign n23310 = n23309 ^ n2366 ^ 1'b0 ;
  assign n23311 = n23310 ^ n22740 ^ 1'b0 ;
  assign n23312 = n16752 ^ n7809 ^ 1'b0 ;
  assign n23313 = n729 & ~n2689 ;
  assign n23314 = ~n458 & n5073 ;
  assign n23315 = n6899 & n23314 ;
  assign n23316 = n23313 & n23315 ;
  assign n23317 = n18975 ^ n1221 ^ 1'b0 ;
  assign n23318 = ~n16387 & n23317 ;
  assign n23319 = n23318 ^ n12030 ^ 1'b0 ;
  assign n23320 = n2650 & n10460 ;
  assign n23321 = n11142 | n23320 ;
  assign n23322 = n23321 ^ n2078 ^ 1'b0 ;
  assign n23323 = n5551 & n23322 ;
  assign n23324 = ~n13268 & n23323 ;
  assign n23325 = n3402 & ~n5257 ;
  assign n23326 = n9679 ^ n8253 ^ 1'b0 ;
  assign n23327 = n23325 | n23326 ;
  assign n23328 = n4294 & n18228 ;
  assign n23329 = n2868 & n23328 ;
  assign n23330 = ~n1159 & n15696 ;
  assign n23331 = n23330 ^ n7887 ^ 1'b0 ;
  assign n23332 = n10375 & ~n21380 ;
  assign n23333 = n23332 ^ n1757 ^ 1'b0 ;
  assign n23334 = n11856 | n14400 ;
  assign n23335 = n9592 ^ n8309 ^ 1'b0 ;
  assign n23336 = ~n8655 & n23335 ;
  assign n23337 = n20450 | n23336 ;
  assign n23338 = ~n8151 & n12352 ;
  assign n23339 = n23338 ^ n923 ^ 1'b0 ;
  assign n23340 = n4812 ^ n3258 ^ 1'b0 ;
  assign n23341 = ~n5176 & n23340 ;
  assign n23342 = ~n1783 & n23341 ;
  assign n23343 = n6373 & n23342 ;
  assign n23344 = n9103 ^ n5622 ^ 1'b0 ;
  assign n23345 = n6146 & ~n12539 ;
  assign n23346 = n5798 & n23345 ;
  assign n23347 = n3542 & ~n4166 ;
  assign n23348 = n1847 & n23347 ;
  assign n23349 = n23348 ^ n22895 ^ 1'b0 ;
  assign n23350 = ~n11421 & n23349 ;
  assign n23351 = n3475 | n4554 ;
  assign n23352 = n10824 & ~n23351 ;
  assign n23353 = n2668 & n12081 ;
  assign n23356 = n2416 & ~n12260 ;
  assign n23354 = n2143 & ~n6376 ;
  assign n23355 = n12901 | n23354 ;
  assign n23357 = n23356 ^ n23355 ^ 1'b0 ;
  assign n23358 = n3116 & n20301 ;
  assign n23359 = n9464 ^ n5959 ^ n1608 ;
  assign n23360 = n7567 & ~n23359 ;
  assign n23361 = ~n4648 & n23360 ;
  assign n23362 = n23361 ^ n11107 ^ 1'b0 ;
  assign n23363 = n19527 ^ n3184 ^ 1'b0 ;
  assign n23364 = n4388 & ~n23363 ;
  assign n23365 = n4132 ^ n623 ^ 1'b0 ;
  assign n23366 = ~n20526 & n23365 ;
  assign n23367 = ~n2855 & n16101 ;
  assign n23368 = n23367 ^ n3648 ^ 1'b0 ;
  assign n23369 = n3189 & n23368 ;
  assign n23370 = n2869 | n18695 ;
  assign n23371 = n1020 | n23370 ;
  assign n23372 = ~n10050 & n23371 ;
  assign n23373 = n23372 ^ n14972 ^ 1'b0 ;
  assign n23374 = n1706 | n13437 ;
  assign n23375 = n7155 ^ n1967 ^ 1'b0 ;
  assign n23376 = n4421 & ~n23375 ;
  assign n23379 = n14302 & ~n20572 ;
  assign n23377 = n3795 | n6834 ;
  assign n23378 = n4857 | n23377 ;
  assign n23380 = n23379 ^ n23378 ^ 1'b0 ;
  assign n23381 = n6832 ^ n4424 ^ 1'b0 ;
  assign n23382 = ~n13273 & n23381 ;
  assign n23383 = n23382 ^ n4747 ^ 1'b0 ;
  assign n23387 = n538 | n11863 ;
  assign n23384 = n2185 & n15164 ;
  assign n23385 = n23384 ^ n6801 ^ 1'b0 ;
  assign n23386 = ~n9301 & n23385 ;
  assign n23388 = n23387 ^ n23386 ^ 1'b0 ;
  assign n23389 = ~n23383 & n23388 ;
  assign n23392 = n13506 & n14779 ;
  assign n23390 = n14323 ^ n5715 ^ 1'b0 ;
  assign n23391 = ~n17078 & n23390 ;
  assign n23393 = n23392 ^ n23391 ^ 1'b0 ;
  assign n23394 = n2728 & ~n6736 ;
  assign n23395 = n6736 & n23394 ;
  assign n23396 = n23395 ^ n13330 ^ 1'b0 ;
  assign n23397 = n9077 | n23396 ;
  assign n23398 = ~n10528 & n23397 ;
  assign n23399 = n3741 & n10705 ;
  assign n23400 = n6420 | n13113 ;
  assign n23403 = n1368 & n8622 ;
  assign n23401 = n3105 ^ x94 ^ 1'b0 ;
  assign n23402 = n23401 ^ n12850 ^ 1'b0 ;
  assign n23404 = n23403 ^ n23402 ^ 1'b0 ;
  assign n23405 = ~n1580 & n23404 ;
  assign n23406 = n1117 & n5082 ;
  assign n23407 = n23406 ^ n21304 ^ 1'b0 ;
  assign n23408 = n9832 & n23407 ;
  assign n23409 = n16939 & n23408 ;
  assign n23410 = n19452 ^ n1096 ^ 1'b0 ;
  assign n23411 = ~n726 & n3863 ;
  assign n23412 = n23411 ^ n17222 ^ 1'b0 ;
  assign n23413 = ~n2982 & n23412 ;
  assign n23414 = n694 & n11696 ;
  assign n23415 = ( ~n825 & n1202 ) | ( ~n825 & n3666 ) | ( n1202 & n3666 ) ;
  assign n23416 = n15248 | n16189 ;
  assign n23419 = n5893 & ~n6079 ;
  assign n23420 = ~n8228 & n23419 ;
  assign n23417 = n15675 | n16591 ;
  assign n23418 = ( n1888 & n18141 ) | ( n1888 & n23417 ) | ( n18141 & n23417 ) ;
  assign n23421 = n23420 ^ n23418 ^ 1'b0 ;
  assign n23422 = n23416 | n23421 ;
  assign n23423 = n20917 ^ n10440 ^ 1'b0 ;
  assign n23424 = n19538 ^ n6674 ^ 1'b0 ;
  assign n23425 = n5619 | n23424 ;
  assign n23426 = n23423 & n23425 ;
  assign n23427 = n23426 ^ n17285 ^ 1'b0 ;
  assign n23428 = n4065 ^ n3943 ^ 1'b0 ;
  assign n23429 = n14884 & n22755 ;
  assign n23430 = n4664 ^ n1893 ^ 1'b0 ;
  assign n23431 = n23430 ^ n3054 ^ 1'b0 ;
  assign n23432 = ~n5629 & n7076 ;
  assign n23433 = n19264 ^ n1337 ^ 1'b0 ;
  assign n23435 = ~n10935 & n13293 ;
  assign n23434 = n5138 & ~n9199 ;
  assign n23436 = n23435 ^ n23434 ^ 1'b0 ;
  assign n23437 = ~n16451 & n23436 ;
  assign n23438 = ~n9989 & n15101 ;
  assign n23439 = ~n3859 & n7802 ;
  assign n23440 = n23439 ^ n20457 ^ 1'b0 ;
  assign n23441 = n4771 ^ n2550 ^ 1'b0 ;
  assign n23442 = ~n14003 & n23441 ;
  assign n23443 = n290 & n8126 ;
  assign n23444 = n14876 & n23443 ;
  assign n23445 = n1152 & n1784 ;
  assign n23446 = ~n1152 & n23445 ;
  assign n23447 = n11782 & ~n23446 ;
  assign n23448 = ~n11782 & n23447 ;
  assign n23449 = n965 | n3836 ;
  assign n23450 = n11576 & ~n23449 ;
  assign n23451 = ~n2476 & n23450 ;
  assign n23452 = n23448 | n23451 ;
  assign n23453 = n23448 & ~n23452 ;
  assign n23454 = n667 & n5180 ;
  assign n23455 = n2089 ^ n273 ^ 1'b0 ;
  assign n23456 = n23454 & ~n23455 ;
  assign n23457 = ~n8451 & n23456 ;
  assign n23458 = n23457 ^ n19684 ^ 1'b0 ;
  assign n23459 = n4295 & ~n23458 ;
  assign n23460 = n2348 | n12176 ;
  assign n23461 = n23460 ^ n2527 ^ 1'b0 ;
  assign n23462 = ~n5429 & n18313 ;
  assign n23463 = n7644 ^ n2597 ^ 1'b0 ;
  assign n23464 = n23463 ^ n7376 ^ 1'b0 ;
  assign n23465 = n20616 | n23464 ;
  assign n23466 = n15250 | n16784 ;
  assign n23467 = n9762 | n23466 ;
  assign n23468 = n2153 ^ x184 ^ 1'b0 ;
  assign n23469 = n13588 | n23468 ;
  assign n23470 = n18508 ^ n7928 ^ 1'b0 ;
  assign n23471 = n22893 | n23470 ;
  assign n23472 = n18671 ^ n1815 ^ 1'b0 ;
  assign n23473 = n13656 ^ n9986 ^ n9360 ;
  assign n23474 = n23473 ^ n1643 ^ 1'b0 ;
  assign n23475 = n16649 & ~n23474 ;
  assign n23476 = n14610 ^ n14234 ^ 1'b0 ;
  assign n23477 = x124 & n23476 ;
  assign n23478 = n628 | n21688 ;
  assign n23479 = n12781 | n23478 ;
  assign n23480 = n2495 & ~n11938 ;
  assign n23481 = n2135 | n4022 ;
  assign n23482 = n23481 ^ n5779 ^ 1'b0 ;
  assign n23483 = n23480 & ~n23482 ;
  assign n23484 = ~n8654 & n23483 ;
  assign n23485 = n20812 & n23484 ;
  assign n23486 = n1463 & n2624 ;
  assign n23487 = ~n16705 & n18576 ;
  assign n23488 = n20132 ^ n15537 ^ 1'b0 ;
  assign n23489 = n15600 | n23488 ;
  assign n23490 = ~x1 & n2735 ;
  assign n23491 = n23490 ^ n2806 ^ 1'b0 ;
  assign n23492 = n12801 & n17182 ;
  assign n23493 = ~n23491 & n23492 ;
  assign n23494 = n12980 | n23493 ;
  assign n23495 = n19568 | n23494 ;
  assign n23496 = n18824 ^ n16759 ^ 1'b0 ;
  assign n23497 = n1217 & ~n23496 ;
  assign n23498 = n12720 | n23497 ;
  assign n23499 = n21841 ^ n19875 ^ n9339 ;
  assign n23500 = n1939 | n15380 ;
  assign n23501 = n1765 & ~n8709 ;
  assign n23502 = n23501 ^ n18686 ^ 1'b0 ;
  assign n23503 = n2153 & ~n23502 ;
  assign n23504 = n11912 ^ n10236 ^ 1'b0 ;
  assign n23505 = n17846 & ~n23504 ;
  assign n23506 = n13157 | n18888 ;
  assign n23507 = n647 & ~n7659 ;
  assign n23508 = n23507 ^ n10587 ^ 1'b0 ;
  assign n23509 = n23508 ^ n2175 ^ 1'b0 ;
  assign n23510 = n5031 | n23509 ;
  assign n23511 = n23510 ^ n16463 ^ 1'b0 ;
  assign n23512 = n23506 | n23511 ;
  assign n23513 = n21395 | n23512 ;
  assign n23514 = n1429 & ~n13228 ;
  assign n23515 = n10188 ^ n2824 ^ 1'b0 ;
  assign n23516 = n23515 ^ n15417 ^ 1'b0 ;
  assign n23517 = n21598 & ~n23516 ;
  assign n23518 = n3272 & ~n20527 ;
  assign n23519 = n23518 ^ n8001 ^ 1'b0 ;
  assign n23520 = n23519 ^ n19943 ^ 1'b0 ;
  assign n23521 = n3707 | n23520 ;
  assign n23522 = n1405 | n10528 ;
  assign n23523 = n14695 & ~n23522 ;
  assign n23524 = n3488 & n23523 ;
  assign n23525 = n9941 | n14929 ;
  assign n23526 = n6015 | n23525 ;
  assign n23527 = n23526 ^ n2546 ^ 1'b0 ;
  assign n23528 = n23524 | n23527 ;
  assign n23529 = n2438 | n11977 ;
  assign n23530 = n14076 | n16841 ;
  assign n23531 = n4812 | n5150 ;
  assign n23532 = n5150 & ~n23531 ;
  assign n23533 = ~n10607 & n23532 ;
  assign n23534 = n512 & ~n22700 ;
  assign n23535 = n3875 & ~n8747 ;
  assign n23536 = n6962 & n23535 ;
  assign n23537 = n1271 & n19100 ;
  assign n23538 = n23537 ^ n10746 ^ 1'b0 ;
  assign n23539 = ~n1684 & n20145 ;
  assign n23540 = n23538 | n23539 ;
  assign n23541 = n3862 & ~n5651 ;
  assign n23542 = n1018 & n6884 ;
  assign n23543 = n10958 ^ n1453 ^ x119 ;
  assign n23544 = n14528 ^ n2482 ^ 1'b0 ;
  assign n23545 = ~n11055 & n23544 ;
  assign n23546 = n5118 & n17451 ;
  assign n23547 = n5159 & n6774 ;
  assign n23548 = n8421 ^ n4524 ^ n3432 ;
  assign n23549 = ~n16050 & n23548 ;
  assign n23550 = n458 | n3386 ;
  assign n23551 = n6283 & ~n23550 ;
  assign n23552 = n18687 ^ n11618 ^ 1'b0 ;
  assign n23553 = n23551 | n23552 ;
  assign n23554 = n20164 ^ n5495 ^ 1'b0 ;
  assign n23555 = n22822 ^ n10817 ^ 1'b0 ;
  assign n23556 = ~n23554 & n23555 ;
  assign n23557 = n11727 ^ n9783 ^ 1'b0 ;
  assign n23558 = n5238 ^ n5082 ^ n3419 ;
  assign n23559 = n2820 & n16770 ;
  assign n23560 = n23559 ^ n5512 ^ 1'b0 ;
  assign n23561 = ~n3694 & n23560 ;
  assign n23562 = n12312 | n17947 ;
  assign n23563 = n23562 ^ n3514 ^ 1'b0 ;
  assign n23564 = ~n3531 & n9711 ;
  assign n23565 = ~n12800 & n23564 ;
  assign n23566 = ~n23563 & n23565 ;
  assign n23567 = ~n3559 & n19594 ;
  assign n23568 = n20469 & n22964 ;
  assign n23569 = n23568 ^ n2879 ^ 1'b0 ;
  assign n23570 = n8083 & ~n23569 ;
  assign n23571 = n9608 & n23570 ;
  assign n23572 = ~n8915 & n17266 ;
  assign n23573 = n7708 ^ n4810 ^ 1'b0 ;
  assign n23574 = ~n15997 & n23573 ;
  assign n23575 = ~x68 & n8895 ;
  assign n23577 = ~n3499 & n5639 ;
  assign n23576 = ~n4674 & n15681 ;
  assign n23578 = n23577 ^ n23576 ^ 1'b0 ;
  assign n23579 = n8621 & n17727 ;
  assign n23580 = ~n11648 & n23579 ;
  assign n23581 = n23580 ^ n5914 ^ 1'b0 ;
  assign n23582 = n2629 | n23581 ;
  assign n23583 = n8773 & n11171 ;
  assign n23584 = n23583 ^ n7326 ^ 1'b0 ;
  assign n23585 = n2602 & ~n7960 ;
  assign n23586 = n14041 & ~n23585 ;
  assign n23587 = ~n8963 & n23586 ;
  assign n23589 = n11034 & n22676 ;
  assign n23588 = n15077 | n21781 ;
  assign n23590 = n23589 ^ n23588 ^ 1'b0 ;
  assign n23591 = ~n23587 & n23590 ;
  assign n23592 = n4375 ^ n2723 ^ 1'b0 ;
  assign n23593 = n3690 & n23592 ;
  assign n23594 = n5564 ^ n1533 ^ 1'b0 ;
  assign n23595 = n23593 & n23594 ;
  assign n23596 = ~n23591 & n23595 ;
  assign n23597 = n17035 | n18861 ;
  assign n23598 = n8804 & ~n18216 ;
  assign n23599 = ~n1508 & n23598 ;
  assign n23600 = n7839 | n23599 ;
  assign n23601 = n23600 ^ n20133 ^ 1'b0 ;
  assign n23602 = n23601 ^ n452 ^ 1'b0 ;
  assign n23603 = n23092 ^ n4267 ^ n633 ;
  assign n23604 = n4279 & ~n20474 ;
  assign n23605 = n8036 & n18797 ;
  assign n23606 = ~n8193 & n23605 ;
  assign n23607 = n10630 & n23606 ;
  assign n23608 = n12531 ^ n12306 ^ 1'b0 ;
  assign n23609 = n1508 & n10397 ;
  assign n23610 = n23609 ^ n13297 ^ 1'b0 ;
  assign n23611 = n4459 | n23610 ;
  assign n23612 = n23611 ^ x53 ^ 1'b0 ;
  assign n23613 = n3224 & n8338 ;
  assign n23614 = n5007 & n16384 ;
  assign n23615 = ( n2340 & n6666 ) | ( n2340 & ~n13214 ) | ( n6666 & ~n13214 ) ;
  assign n23616 = n16083 | n16505 ;
  assign n23617 = n23615 & ~n23616 ;
  assign n23618 = n607 & n8626 ;
  assign n23619 = n8774 & n23618 ;
  assign n23620 = n5530 ^ n1159 ^ 1'b0 ;
  assign n23621 = n12912 ^ n1819 ^ 1'b0 ;
  assign n23622 = n23621 ^ n14947 ^ 1'b0 ;
  assign n23623 = n1226 & n12172 ;
  assign n23624 = n23623 ^ n9916 ^ 1'b0 ;
  assign n23625 = n23624 ^ n13160 ^ 1'b0 ;
  assign n23626 = n23622 & n23625 ;
  assign n23630 = ~n1724 & n4590 ;
  assign n23629 = ~n8127 & n8281 ;
  assign n23631 = n23630 ^ n23629 ^ 1'b0 ;
  assign n23632 = n1379 & ~n23631 ;
  assign n23633 = n23632 ^ n13347 ^ 1'b0 ;
  assign n23627 = n18399 ^ n5821 ^ 1'b0 ;
  assign n23628 = ~n11013 & n23627 ;
  assign n23634 = n23633 ^ n23628 ^ 1'b0 ;
  assign n23635 = n8495 & ~n23634 ;
  assign n23636 = n5195 & ~n9886 ;
  assign n23637 = x239 & n23636 ;
  assign n23638 = n23637 ^ n4911 ^ 1'b0 ;
  assign n23639 = n10124 & ~n23638 ;
  assign n23640 = n2195 & ~n7164 ;
  assign n23641 = n2019 | n9961 ;
  assign n23642 = n23640 | n23641 ;
  assign n23643 = n18418 ^ n2591 ^ 1'b0 ;
  assign n23644 = n4466 & n23643 ;
  assign n23645 = n19281 ^ n6804 ^ 1'b0 ;
  assign n23646 = n9607 & n11543 ;
  assign n23647 = n17626 ^ n15100 ^ 1'b0 ;
  assign n23648 = n14602 | n23647 ;
  assign n23649 = ~n6790 & n23648 ;
  assign n23650 = n23649 ^ n16979 ^ 1'b0 ;
  assign n23651 = n5302 & n14864 ;
  assign n23652 = n23651 ^ n4372 ^ 1'b0 ;
  assign n23653 = n12237 ^ n5379 ^ 1'b0 ;
  assign n23654 = n23653 ^ n2431 ^ 1'b0 ;
  assign n23655 = n23652 & n23654 ;
  assign n23656 = n23655 ^ n965 ^ 1'b0 ;
  assign n23657 = n10395 ^ n5779 ^ 1'b0 ;
  assign n23658 = n4985 & n6626 ;
  assign n23659 = n23658 ^ n17267 ^ 1'b0 ;
  assign n23660 = ~n23657 & n23659 ;
  assign n23661 = n6276 | n13852 ;
  assign n23662 = n19409 ^ n8811 ^ n1475 ;
  assign n23663 = ~n8421 & n12340 ;
  assign n23664 = n23663 ^ n5207 ^ 1'b0 ;
  assign n23665 = n3447 & n4364 ;
  assign n23666 = n14531 ^ n1237 ^ 1'b0 ;
  assign n23672 = ~n3451 & n4338 ;
  assign n23673 = ~n2475 & n23672 ;
  assign n23667 = ~n3707 & n17022 ;
  assign n23668 = n23667 ^ n12748 ^ 1'b0 ;
  assign n23669 = ~n7316 & n23668 ;
  assign n23670 = n23669 ^ n3073 ^ 1'b0 ;
  assign n23671 = n9041 & n23670 ;
  assign n23674 = n23673 ^ n23671 ^ n1390 ;
  assign n23675 = n12167 ^ n6134 ^ 1'b0 ;
  assign n23676 = n13311 & ~n23675 ;
  assign n23677 = n7403 & n23676 ;
  assign n23678 = n10794 ^ n9612 ^ 1'b0 ;
  assign n23679 = n23677 | n23678 ;
  assign n23680 = n1914 | n9175 ;
  assign n23681 = n15089 ^ n789 ^ 1'b0 ;
  assign n23682 = n23680 | n23681 ;
  assign n23683 = n7232 & ~n8481 ;
  assign n23684 = n22667 & ~n23683 ;
  assign n23685 = n10413 | n16102 ;
  assign n23686 = n8054 & ~n22917 ;
  assign n23687 = n23686 ^ n17732 ^ 1'b0 ;
  assign n23688 = n7021 | n23687 ;
  assign n23689 = n15989 ^ n15354 ^ n14818 ;
  assign n23690 = ~n11158 & n15434 ;
  assign n23691 = n3739 & n18206 ;
  assign n23692 = n728 & n15991 ;
  assign n23693 = n23692 ^ n909 ^ 1'b0 ;
  assign n23694 = n8675 & ~n10141 ;
  assign n23695 = n23694 ^ n11045 ^ 1'b0 ;
  assign n23696 = n4739 ^ x15 ^ 1'b0 ;
  assign n23697 = n844 & n23696 ;
  assign n23698 = n23695 & n23697 ;
  assign n23699 = n9394 & n10602 ;
  assign n23700 = ~n15471 & n23699 ;
  assign n23701 = n1588 | n11792 ;
  assign n23702 = n23700 & ~n23701 ;
  assign n23703 = ~n7383 & n8956 ;
  assign n23704 = n1018 | n10030 ;
  assign n23705 = n958 & ~n23704 ;
  assign n23706 = n23703 & n23705 ;
  assign n23707 = n4952 ^ n4417 ^ 1'b0 ;
  assign n23709 = n12506 ^ n2765 ^ 1'b0 ;
  assign n23710 = n3886 & n23709 ;
  assign n23708 = n3756 & ~n9221 ;
  assign n23711 = n23710 ^ n23708 ^ 1'b0 ;
  assign n23712 = n14504 ^ n1267 ^ 1'b0 ;
  assign n23713 = ~n1429 & n4466 ;
  assign n23714 = x123 & ~n15677 ;
  assign n23715 = n9397 & ~n18132 ;
  assign n23716 = ~n5733 & n23715 ;
  assign n23717 = n2990 & ~n19013 ;
  assign n23718 = n911 | n21062 ;
  assign n23721 = x175 & n18407 ;
  assign n23719 = n4291 & ~n22396 ;
  assign n23720 = n11659 | n23719 ;
  assign n23722 = n23721 ^ n23720 ^ 1'b0 ;
  assign n23723 = n23722 ^ n14863 ^ 1'b0 ;
  assign n23724 = n2376 & ~n23723 ;
  assign n23725 = n1178 & ~n2856 ;
  assign n23726 = ~n1178 & n23725 ;
  assign n23727 = n16815 | n23726 ;
  assign n23728 = n16815 & ~n23727 ;
  assign n23729 = ( n853 & n6419 ) | ( n853 & n7902 ) | ( n6419 & n7902 ) ;
  assign n23730 = n21609 ^ n18541 ^ 1'b0 ;
  assign n23731 = ~n23729 & n23730 ;
  assign n23733 = n8574 ^ n7867 ^ n1651 ;
  assign n23732 = n493 | n1332 ;
  assign n23734 = n23733 ^ n23732 ^ 1'b0 ;
  assign n23735 = n23734 ^ n8033 ^ 1'b0 ;
  assign n23736 = n12616 ^ n2438 ^ 1'b0 ;
  assign n23737 = n5686 & ~n23736 ;
  assign n23738 = n3705 & ~n4582 ;
  assign n23739 = n23738 ^ n17465 ^ 1'b0 ;
  assign n23740 = n8619 & ~n21435 ;
  assign n23741 = n19264 & n23740 ;
  assign n23742 = x24 & n832 ;
  assign n23743 = n9150 & n23742 ;
  assign n23744 = n7746 ^ n6264 ^ n2274 ;
  assign n23745 = ~n2260 & n3968 ;
  assign n23746 = n6348 & n23745 ;
  assign n23747 = n23744 | n23746 ;
  assign n23756 = n4297 & ~n5462 ;
  assign n23748 = n498 & ~n791 ;
  assign n23749 = n6473 ^ x75 ^ 1'b0 ;
  assign n23750 = n23749 ^ n3645 ^ 1'b0 ;
  assign n23751 = n23748 & n23750 ;
  assign n23752 = n10112 & n23751 ;
  assign n23753 = n5310 | n11441 ;
  assign n23754 = n23752 & ~n23753 ;
  assign n23755 = n2978 & ~n23754 ;
  assign n23757 = n23756 ^ n23755 ^ 1'b0 ;
  assign n23758 = n18501 & ~n23681 ;
  assign n23759 = n3026 ^ n2315 ^ 1'b0 ;
  assign n23760 = n801 & n22836 ;
  assign n23761 = n23760 ^ n14837 ^ 1'b0 ;
  assign n23762 = n6427 & n13210 ;
  assign n23763 = n23762 ^ n18360 ^ 1'b0 ;
  assign n23764 = n23763 ^ n1363 ^ 1'b0 ;
  assign n23765 = n23764 ^ n4080 ^ 1'b0 ;
  assign n23766 = ~n22137 & n23765 ;
  assign n23767 = n19801 ^ n11573 ^ 1'b0 ;
  assign n23771 = n12788 ^ n10965 ^ 1'b0 ;
  assign n23768 = n1744 & ~n16384 ;
  assign n23769 = n13156 & n23768 ;
  assign n23770 = ~n21273 & n23769 ;
  assign n23772 = n23771 ^ n23770 ^ 1'b0 ;
  assign n23773 = n3979 & ~n14825 ;
  assign n23774 = n4825 & ~n18141 ;
  assign n23775 = n23774 ^ n3326 ^ 1'b0 ;
  assign n23776 = n2451 & ~n23775 ;
  assign n23777 = x240 & ~n23776 ;
  assign n23778 = n2892 | n8964 ;
  assign n23779 = n23778 ^ n17159 ^ 1'b0 ;
  assign n23780 = ~n10965 & n15049 ;
  assign n23781 = n10422 & n23780 ;
  assign n23782 = n6461 | n17599 ;
  assign n23783 = n23782 ^ n16908 ^ 1'b0 ;
  assign n23784 = ~n23781 & n23783 ;
  assign n23785 = n9177 ^ n7655 ^ n5883 ;
  assign n23786 = n3575 | n23785 ;
  assign n23787 = n20838 ^ n1773 ^ 1'b0 ;
  assign n23788 = n23787 ^ n11765 ^ n6093 ;
  assign n23789 = n15786 | n19316 ;
  assign n23790 = n8162 | n14024 ;
  assign n23791 = n10300 | n23790 ;
  assign n23793 = ~n2803 & n5293 ;
  assign n23794 = ~n5293 & n23793 ;
  assign n23795 = n16580 & ~n23794 ;
  assign n23792 = n7321 & ~n17424 ;
  assign n23796 = n23795 ^ n23792 ^ 1'b0 ;
  assign n23797 = n9768 & ~n12163 ;
  assign n23798 = n23797 ^ n20514 ^ 1'b0 ;
  assign n23799 = n11914 | n23798 ;
  assign n23800 = n17578 ^ n5439 ^ 1'b0 ;
  assign n23801 = n1853 & n23800 ;
  assign n23802 = n1031 & n13899 ;
  assign n23803 = x120 & n2447 ;
  assign n23804 = n23802 & n23803 ;
  assign n23807 = n1023 & n13133 ;
  assign n23805 = n8876 | n14817 ;
  assign n23806 = n10464 & ~n23805 ;
  assign n23808 = n23807 ^ n23806 ^ 1'b0 ;
  assign n23813 = n17876 ^ n17126 ^ 1'b0 ;
  assign n23811 = ~n2293 & n13778 ;
  assign n23812 = n23811 ^ n1907 ^ 1'b0 ;
  assign n23814 = n23813 ^ n23812 ^ 1'b0 ;
  assign n23815 = n7994 & n23814 ;
  assign n23809 = n6402 & n14676 ;
  assign n23810 = n23809 ^ n15435 ^ 1'b0 ;
  assign n23816 = n23815 ^ n23810 ^ 1'b0 ;
  assign n23817 = n13509 & ~n17201 ;
  assign n23818 = n23817 ^ n14924 ^ 1'b0 ;
  assign n23819 = ~n8257 & n23818 ;
  assign n23820 = n6407 & ~n23819 ;
  assign n23821 = ~n1283 & n4080 ;
  assign n23822 = ~n19386 & n23821 ;
  assign n23823 = n20873 & ~n23822 ;
  assign n23824 = n23823 ^ n9907 ^ 1'b0 ;
  assign n23825 = n444 & ~n2700 ;
  assign n23826 = n9238 ^ n6261 ^ 1'b0 ;
  assign n23827 = n23825 & ~n23826 ;
  assign n23828 = ~n9133 & n13748 ;
  assign n23829 = ~n13222 & n23828 ;
  assign n23830 = n8098 & n19281 ;
  assign n23831 = n23830 ^ n2591 ^ 1'b0 ;
  assign n23832 = ~n13291 & n17092 ;
  assign n23833 = n8747 & n23832 ;
  assign n23834 = n6203 & n7019 ;
  assign n23835 = n23834 ^ n15216 ^ 1'b0 ;
  assign n23836 = n11571 | n18973 ;
  assign n23837 = n23835 & ~n23836 ;
  assign n23838 = n23837 ^ n18072 ^ 1'b0 ;
  assign n23839 = n22791 ^ n10915 ^ 1'b0 ;
  assign n23840 = n17338 ^ n15652 ^ 1'b0 ;
  assign n23841 = n2812 & n23840 ;
  assign n23842 = n23841 ^ n12753 ^ 1'b0 ;
  assign n23843 = n13283 ^ n12816 ^ 1'b0 ;
  assign n23844 = n16712 & ~n23843 ;
  assign n23845 = n19334 ^ n9212 ^ 1'b0 ;
  assign n23846 = n2716 | n23845 ;
  assign n23847 = n23846 ^ n9837 ^ 1'b0 ;
  assign n23848 = n4655 | n23847 ;
  assign n23849 = ~n3237 & n15260 ;
  assign n23850 = n7720 & n23849 ;
  assign n23851 = n10692 ^ n7098 ^ 1'b0 ;
  assign n23852 = n3405 & n23851 ;
  assign n23853 = ~n23850 & n23852 ;
  assign n23859 = n3872 & ~n11806 ;
  assign n23860 = ~n3039 & n23859 ;
  assign n23854 = n458 & n1901 ;
  assign n23855 = ~n4307 & n23854 ;
  assign n23856 = n22642 ^ n2057 ^ 1'b0 ;
  assign n23857 = ( n4385 & n23855 ) | ( n4385 & n23856 ) | ( n23855 & n23856 ) ;
  assign n23858 = n22161 & n23857 ;
  assign n23861 = n23860 ^ n23858 ^ 1'b0 ;
  assign n23862 = ( n10259 & ~n15399 ) | ( n10259 & n19990 ) | ( ~n15399 & n19990 ) ;
  assign n23863 = n4378 & n9415 ;
  assign n23864 = n23863 ^ n22926 ^ 1'b0 ;
  assign n23865 = n2055 | n3123 ;
  assign n23866 = n13789 & ~n23865 ;
  assign n23867 = n6694 & n12694 ;
  assign n23868 = ~n10898 & n23867 ;
  assign n23869 = n8202 | n23868 ;
  assign n23870 = n23869 ^ n18677 ^ 1'b0 ;
  assign n23871 = n14349 & n16504 ;
  assign n23872 = n1928 & n3687 ;
  assign n23873 = n23872 ^ n9191 ^ 1'b0 ;
  assign n23874 = n23871 & ~n23873 ;
  assign n23875 = n2572 & n4367 ;
  assign n23876 = n23875 ^ n4319 ^ 1'b0 ;
  assign n23877 = ~x204 & n23876 ;
  assign n23878 = n23877 ^ n8556 ^ 1'b0 ;
  assign n23879 = n387 & n8137 ;
  assign n23880 = ~n14646 & n23879 ;
  assign n23881 = n21459 ^ n7123 ^ 1'b0 ;
  assign n23882 = n9679 & n23881 ;
  assign n23884 = n6635 ^ n3939 ^ 1'b0 ;
  assign n23883 = ( n2166 & n2503 ) | ( n2166 & n6573 ) | ( n2503 & n6573 ) ;
  assign n23885 = n23884 ^ n23883 ^ 1'b0 ;
  assign n23886 = n2818 | n3996 ;
  assign n23887 = n23885 & ~n23886 ;
  assign n23888 = x144 & n23887 ;
  assign n23890 = n3143 ^ x35 ^ 1'b0 ;
  assign n23891 = n2082 & ~n23890 ;
  assign n23892 = n7748 & n23891 ;
  assign n23889 = n4619 & n17046 ;
  assign n23893 = n23892 ^ n23889 ^ 1'b0 ;
  assign n23894 = ~n3128 & n23893 ;
  assign n23895 = n6747 & ~n10267 ;
  assign n23896 = n3448 & n23895 ;
  assign n23897 = ~n12956 & n18389 ;
  assign n23898 = n19549 & n23897 ;
  assign n23899 = n20248 & ~n23898 ;
  assign n23900 = n6154 ^ n934 ^ 1'b0 ;
  assign n23901 = ~n5400 & n6998 ;
  assign n23902 = n23900 & n23901 ;
  assign n23904 = n2671 & ~n4671 ;
  assign n23905 = n23904 ^ n3181 ^ 1'b0 ;
  assign n23903 = n5853 & ~n5938 ;
  assign n23906 = n23905 ^ n23903 ^ 1'b0 ;
  assign n23907 = n4961 | n14978 ;
  assign n23908 = n23907 ^ n23207 ^ 1'b0 ;
  assign n23909 = ~n19017 & n20162 ;
  assign n23910 = n23909 ^ n7316 ^ 1'b0 ;
  assign n23911 = n21277 ^ n18233 ^ 1'b0 ;
  assign n23912 = ~n23910 & n23911 ;
  assign n23913 = n13054 ^ n4582 ^ 1'b0 ;
  assign n23914 = ~n580 & n23913 ;
  assign n23915 = ~n20809 & n23914 ;
  assign n23916 = n23915 ^ n4203 ^ 1'b0 ;
  assign n23917 = n1832 & ~n23916 ;
  assign n23918 = n9786 | n15519 ;
  assign n23919 = n23918 ^ n19017 ^ 1'b0 ;
  assign n23920 = n23917 & n23919 ;
  assign n23921 = n9471 | n15189 ;
  assign n23922 = n3360 | n4857 ;
  assign n23923 = n17821 ^ n14678 ^ 1'b0 ;
  assign n23924 = n23922 & ~n23923 ;
  assign n23926 = n8816 ^ n6117 ^ 1'b0 ;
  assign n23925 = n638 & n9632 ;
  assign n23927 = n23926 ^ n23925 ^ 1'b0 ;
  assign n23928 = n13651 ^ n9384 ^ 1'b0 ;
  assign n23929 = ~n1404 & n23928 ;
  assign n23930 = n23929 ^ n22570 ^ 1'b0 ;
  assign n23931 = n7440 & ~n12660 ;
  assign n23932 = n19896 & ~n23353 ;
  assign n23933 = n11658 ^ n5682 ^ 1'b0 ;
  assign n23934 = ~n23133 & n23933 ;
  assign n23935 = n23934 ^ n355 ^ 1'b0 ;
  assign n23936 = ~n5305 & n5444 ;
  assign n23937 = n1139 & n23936 ;
  assign n23938 = n446 & ~n17395 ;
  assign n23939 = n12860 ^ n4616 ^ 1'b0 ;
  assign n23940 = n18357 & n23939 ;
  assign n23942 = n734 & ~n19691 ;
  assign n23941 = n1573 | n21121 ;
  assign n23943 = n23942 ^ n23941 ^ 1'b0 ;
  assign n23944 = n2513 & ~n12458 ;
  assign n23945 = n12296 ^ n3866 ^ 1'b0 ;
  assign n23946 = n23944 & n23945 ;
  assign n23947 = n21002 ^ n13388 ^ 1'b0 ;
  assign n23948 = n5622 & n9423 ;
  assign n23949 = ~n3182 & n23948 ;
  assign n23950 = n3707 & n23949 ;
  assign n23952 = n7410 & n7587 ;
  assign n23951 = ~n6258 & n7818 ;
  assign n23953 = n23952 ^ n23951 ^ 1'b0 ;
  assign n23954 = n23950 & ~n23953 ;
  assign n23955 = n11012 ^ n6991 ^ 1'b0 ;
  assign n23956 = n5712 & ~n17283 ;
  assign n23957 = ~n529 & n1275 ;
  assign n23958 = n23956 & n23957 ;
  assign n23959 = n1642 & ~n13460 ;
  assign n23960 = n741 & ~n6083 ;
  assign n23961 = ( n7613 & n13315 ) | ( n7613 & ~n23960 ) | ( n13315 & ~n23960 ) ;
  assign n23962 = n23961 ^ n12952 ^ 1'b0 ;
  assign n23963 = n10042 | n23962 ;
  assign n23964 = n2812 & ~n3599 ;
  assign n23965 = n23964 ^ n10861 ^ 1'b0 ;
  assign n23966 = n23965 ^ n14324 ^ 1'b0 ;
  assign n23967 = n23966 ^ n2289 ^ 1'b0 ;
  assign n23968 = n3119 & ~n10160 ;
  assign n23969 = n12921 & ~n23968 ;
  assign n23970 = n3169 & n23969 ;
  assign n23971 = n14696 | n15726 ;
  assign n23972 = n23970 & ~n23971 ;
  assign n23973 = ~n6997 & n7032 ;
  assign n23974 = n4138 & n16432 ;
  assign n23975 = n15328 | n18956 ;
  assign n23978 = n4161 & n7960 ;
  assign n23976 = n11958 & n16777 ;
  assign n23977 = n23976 ^ n16657 ^ 1'b0 ;
  assign n23979 = n23978 ^ n23977 ^ 1'b0 ;
  assign n23980 = n6359 & n23979 ;
  assign n23981 = n19950 ^ n15666 ^ 1'b0 ;
  assign n23982 = n7467 & n23981 ;
  assign n23983 = n8211 & ~n16939 ;
  assign n23984 = n7181 | n23983 ;
  assign n23985 = n16062 & n23984 ;
  assign n23986 = n16397 | n23985 ;
  assign n23987 = x44 & ~n5587 ;
  assign n23988 = n22370 ^ n4219 ^ 1'b0 ;
  assign n23989 = n12432 ^ n7174 ^ 1'b0 ;
  assign n23990 = n7398 | n15014 ;
  assign n23991 = n23990 ^ n9690 ^ 1'b0 ;
  assign n23992 = n23991 ^ n11623 ^ 1'b0 ;
  assign n23993 = n23989 & ~n23992 ;
  assign n23994 = n2663 | n3043 ;
  assign n23995 = n7788 | n23994 ;
  assign n23996 = n14518 | n23995 ;
  assign n23997 = ( ~n729 & n23354 ) | ( ~n729 & n23996 ) | ( n23354 & n23996 ) ;
  assign n23998 = n8081 & n23997 ;
  assign n23999 = ~n3915 & n23998 ;
  assign n24001 = ~n3392 & n14068 ;
  assign n24002 = n863 & n24001 ;
  assign n24000 = n4946 & ~n7148 ;
  assign n24003 = n24002 ^ n24000 ^ 1'b0 ;
  assign n24005 = n13400 ^ n754 ^ 1'b0 ;
  assign n24006 = n5819 & ~n24005 ;
  assign n24004 = ~n8111 & n8453 ;
  assign n24007 = n24006 ^ n24004 ^ 1'b0 ;
  assign n24008 = n24003 & n24007 ;
  assign n24009 = n5525 & n24008 ;
  assign n24010 = ~n10108 & n10112 ;
  assign n24011 = n3277 | n24010 ;
  assign n24012 = n4149 | n7295 ;
  assign n24013 = n11171 | n24012 ;
  assign n24014 = x2 & ~n20982 ;
  assign n24015 = n6278 ^ n2665 ^ 1'b0 ;
  assign n24016 = n10467 | n24015 ;
  assign n24017 = n24016 ^ n904 ^ 1'b0 ;
  assign n24018 = n12369 | n24017 ;
  assign n24019 = ~n2715 & n12807 ;
  assign n24020 = n24018 & n24019 ;
  assign n24021 = n11586 ^ n1951 ^ 1'b0 ;
  assign n24022 = n16001 & ~n24021 ;
  assign n24023 = n1883 | n4054 ;
  assign n24024 = n562 | n24023 ;
  assign n24025 = n11862 & ~n24024 ;
  assign n24026 = n24022 & ~n24025 ;
  assign n24027 = n1727 & n24026 ;
  assign n24028 = n12094 ^ n5533 ^ 1'b0 ;
  assign n24029 = n11133 & n24028 ;
  assign n24030 = n24029 ^ n2627 ^ 1'b0 ;
  assign n24031 = n23828 ^ n17056 ^ n1181 ;
  assign n24032 = n24031 ^ n12385 ^ 1'b0 ;
  assign n24033 = n810 | n24032 ;
  assign n24034 = n5083 ^ x81 ^ 1'b0 ;
  assign n24035 = ~n1356 & n24034 ;
  assign n24036 = n18862 ^ n1785 ^ 1'b0 ;
  assign n24037 = n4574 & ~n8246 ;
  assign n24038 = n24037 ^ x7 ^ 1'b0 ;
  assign n24039 = n24038 ^ n6823 ^ 1'b0 ;
  assign n24040 = n16925 ^ n4538 ^ 1'b0 ;
  assign n24041 = x222 | n13810 ;
  assign n24042 = n15429 | n24041 ;
  assign n24043 = n24042 ^ n7915 ^ 1'b0 ;
  assign n24044 = n3527 | n4879 ;
  assign n24045 = n822 & ~n12980 ;
  assign n24046 = n24044 & n24045 ;
  assign n24047 = n21588 ^ n6935 ^ 1'b0 ;
  assign n24048 = n13455 ^ n8148 ^ 1'b0 ;
  assign n24049 = n527 & n17669 ;
  assign n24050 = n24049 ^ n1443 ^ 1'b0 ;
  assign n24051 = n15208 & ~n24050 ;
  assign n24052 = ( ~x86 & n17601 ) | ( ~x86 & n20156 ) | ( n17601 & n20156 ) ;
  assign n24053 = ~n9034 & n24052 ;
  assign n24054 = n24053 ^ n1920 ^ 1'b0 ;
  assign n24055 = n8082 ^ n7993 ^ 1'b0 ;
  assign n24056 = n9998 ^ n5252 ^ 1'b0 ;
  assign n24057 = n3203 & n24056 ;
  assign n24058 = x213 & n24057 ;
  assign n24059 = n24055 & n24058 ;
  assign n24060 = n4318 ^ n3027 ^ 1'b0 ;
  assign n24061 = n2034 & ~n2889 ;
  assign n24062 = ~n2034 & n24061 ;
  assign n24063 = n2287 & ~n24062 ;
  assign n24064 = n24062 & n24063 ;
  assign n24065 = n24064 ^ n11029 ^ 1'b0 ;
  assign n24066 = n24060 | n24065 ;
  assign n24067 = n24060 & ~n24066 ;
  assign n24069 = n2091 & n12200 ;
  assign n24070 = n5256 & n24069 ;
  assign n24068 = n10560 & n19429 ;
  assign n24071 = n24070 ^ n24068 ^ 1'b0 ;
  assign n24072 = ~n3561 & n11586 ;
  assign n24073 = n24072 ^ n18727 ^ 1'b0 ;
  assign n24074 = ~n1886 & n6868 ;
  assign n24075 = n24074 ^ n2133 ^ 1'b0 ;
  assign n24077 = ~n10393 & n14601 ;
  assign n24078 = n24077 ^ n15509 ^ 1'b0 ;
  assign n24079 = n5821 | n24078 ;
  assign n24076 = n5423 ^ x88 ^ 1'b0 ;
  assign n24080 = n24079 ^ n24076 ^ n1635 ;
  assign n24081 = x247 & ~n10363 ;
  assign n24082 = n19788 & n24081 ;
  assign n24083 = n22964 ^ n1199 ^ 1'b0 ;
  assign n24084 = ( n24079 & ~n24082 ) | ( n24079 & n24083 ) | ( ~n24082 & n24083 ) ;
  assign n24085 = ~n4072 & n16744 ;
  assign n24086 = n15531 & n24085 ;
  assign n24087 = n6154 & n9881 ;
  assign n24088 = n5082 ^ n2602 ^ 1'b0 ;
  assign n24089 = n18436 & ~n24088 ;
  assign n24090 = n20136 & n24089 ;
  assign n24091 = n5613 | n8038 ;
  assign n24092 = n22041 & ~n24091 ;
  assign n24093 = ( n5903 & n15753 ) | ( n5903 & n24092 ) | ( n15753 & n24092 ) ;
  assign n24094 = n7995 ^ n6452 ^ 1'b0 ;
  assign n24095 = n9991 & ~n10178 ;
  assign n24096 = n24094 & n24095 ;
  assign n24097 = n1677 & n24096 ;
  assign n24098 = n11983 ^ n3229 ^ n2664 ;
  assign n24099 = x143 & n21950 ;
  assign n24100 = n4731 | n24099 ;
  assign n24101 = n24100 ^ n6804 ^ 1'b0 ;
  assign n24102 = n1792 & n10798 ;
  assign n24103 = n24102 ^ n10467 ^ 1'b0 ;
  assign n24104 = n24103 ^ n8811 ^ 1'b0 ;
  assign n24105 = n14858 & ~n24104 ;
  assign n24106 = n21703 ^ n6568 ^ 1'b0 ;
  assign n24107 = ~n913 & n6246 ;
  assign n24108 = ~n743 & n24107 ;
  assign n24109 = n8014 ^ n2942 ^ 1'b0 ;
  assign n24110 = n8010 & n24109 ;
  assign n24111 = n307 & n1643 ;
  assign n24112 = n9324 ^ n4063 ^ 1'b0 ;
  assign n24113 = ~n6904 & n24112 ;
  assign n24114 = n19505 & n22925 ;
  assign n24115 = n15265 ^ n1651 ^ 1'b0 ;
  assign n24116 = n1810 & n9379 ;
  assign n24117 = ( n8111 & n11240 ) | ( n8111 & n24116 ) | ( n11240 & n24116 ) ;
  assign n24118 = n6954 & n13959 ;
  assign n24119 = n24118 ^ n17891 ^ 1'b0 ;
  assign n24120 = n15253 & ~n15438 ;
  assign n24121 = ~n24119 & n24120 ;
  assign n24122 = n24121 ^ n5580 ^ 1'b0 ;
  assign n24123 = n4769 & ~n7867 ;
  assign n24124 = n875 & n24123 ;
  assign n24125 = n17834 | n24124 ;
  assign n24126 = n24125 ^ x222 ^ 1'b0 ;
  assign n24127 = n1990 & n21200 ;
  assign n24128 = n10771 ^ n7320 ^ 1'b0 ;
  assign n24129 = n16215 | n24128 ;
  assign n24130 = n10764 & n17249 ;
  assign n24131 = n4954 & ~n11233 ;
  assign n24132 = n24131 ^ n22999 ^ 1'b0 ;
  assign n24133 = n24132 ^ n8933 ^ 1'b0 ;
  assign n24134 = n4859 | n24133 ;
  assign n24135 = n24134 ^ n11013 ^ 1'b0 ;
  assign n24136 = n4671 & n24135 ;
  assign n24137 = n10637 ^ n4653 ^ 1'b0 ;
  assign n24138 = n10593 ^ n6745 ^ 1'b0 ;
  assign n24139 = ~n10160 & n24138 ;
  assign n24140 = n3548 & ~n24092 ;
  assign n24141 = n11572 & ~n12342 ;
  assign n24142 = n20125 & n24141 ;
  assign n24143 = n16929 & ~n24142 ;
  assign n24144 = n5604 & n21320 ;
  assign n24145 = n635 & n24144 ;
  assign n24146 = n5658 | n9455 ;
  assign n24147 = n13317 & ~n24146 ;
  assign n24148 = ~n12118 & n24115 ;
  assign n24149 = ~n6473 & n7838 ;
  assign n24150 = n24149 ^ n14685 ^ 1'b0 ;
  assign n24151 = ( x115 & ~n18029 ) | ( x115 & n24150 ) | ( ~n18029 & n24150 ) ;
  assign n24152 = n11580 | n24151 ;
  assign n24153 = n1103 ^ n1031 ^ 1'b0 ;
  assign n24165 = n2870 | n3673 ;
  assign n24166 = n3673 & ~n24165 ;
  assign n24154 = n343 & n467 ;
  assign n24155 = ~n343 & n24154 ;
  assign n24156 = x65 & x241 ;
  assign n24157 = ~x241 & n24156 ;
  assign n24158 = x253 & ~n24157 ;
  assign n24159 = n24155 & n24158 ;
  assign n24160 = ~n1488 & n4586 ;
  assign n24161 = ~n4586 & n24160 ;
  assign n24162 = n1442 & ~n5880 ;
  assign n24163 = n24161 & n24162 ;
  assign n24164 = n24159 | n24163 ;
  assign n24167 = n24166 ^ n24164 ^ 1'b0 ;
  assign n24168 = n4549 & n7879 ;
  assign n24169 = n24168 ^ n16518 ^ 1'b0 ;
  assign n24170 = n12274 ^ n1684 ^ 1'b0 ;
  assign n24171 = n24169 & n24170 ;
  assign n24172 = n663 & n2112 ;
  assign n24173 = n9823 & n24172 ;
  assign n24174 = n24173 ^ n1580 ^ 1'b0 ;
  assign n24175 = n1700 & n16446 ;
  assign n24176 = ~n13145 & n24175 ;
  assign n24177 = n24176 ^ n16109 ^ 1'b0 ;
  assign n24178 = n20209 & n24177 ;
  assign n24179 = ~n5729 & n18477 ;
  assign n24180 = ~n4108 & n10602 ;
  assign n24181 = n3854 & n24180 ;
  assign n24182 = ~n2511 & n10632 ;
  assign n24183 = n7851 & n24182 ;
  assign n24184 = n12266 | n24183 ;
  assign n24185 = n1841 & n3257 ;
  assign n24186 = ~n22993 & n24185 ;
  assign n24187 = n24186 ^ n7423 ^ n5814 ;
  assign n24188 = n4660 | n4708 ;
  assign n24189 = n2778 & n24188 ;
  assign n24190 = n2250 & ~n8133 ;
  assign n24191 = n17528 & n22771 ;
  assign n24192 = n8692 ^ n5946 ^ 1'b0 ;
  assign n24193 = ~n4544 & n24192 ;
  assign n24194 = ~n3870 & n24193 ;
  assign n24195 = n24194 ^ n17902 ^ 1'b0 ;
  assign n24196 = ~n5790 & n21584 ;
  assign n24197 = n24196 ^ n17209 ^ 1'b0 ;
  assign n24198 = n13057 & n22612 ;
  assign n24202 = n15841 ^ n1689 ^ 1'b0 ;
  assign n24203 = n6972 & n24202 ;
  assign n24199 = n3336 & n7734 ;
  assign n24200 = ~n7164 & n24199 ;
  assign n24201 = n21851 & ~n24200 ;
  assign n24204 = n24203 ^ n24201 ^ 1'b0 ;
  assign n24205 = n16397 & ~n23588 ;
  assign n24206 = n9358 & n24205 ;
  assign n24207 = n23965 ^ n2922 ^ 1'b0 ;
  assign n24208 = ~x93 & n10540 ;
  assign n24209 = n5262 & ~n24208 ;
  assign n24210 = n1387 | n14853 ;
  assign n24211 = n6870 | n24210 ;
  assign n24212 = n24209 & n24211 ;
  assign n24213 = n24212 ^ n5030 ^ 1'b0 ;
  assign n24214 = ~n1064 & n16965 ;
  assign n24215 = n24214 ^ n20944 ^ 1'b0 ;
  assign n24216 = n19374 ^ n2819 ^ 1'b0 ;
  assign n24217 = n20337 ^ n7700 ^ 1'b0 ;
  assign n24218 = n9854 | n17332 ;
  assign n24219 = n7769 ^ n6375 ^ 1'b0 ;
  assign n24221 = n602 | n5980 ;
  assign n24222 = n24221 ^ n13982 ^ n7864 ;
  assign n24223 = n1621 | n24222 ;
  assign n24220 = ~n13329 & n20156 ;
  assign n24224 = n24223 ^ n24220 ^ n12116 ;
  assign n24225 = x251 | n1181 ;
  assign n24226 = n12154 & ~n24225 ;
  assign n24227 = n2042 ^ n994 ^ 1'b0 ;
  assign n24228 = n1809 & ~n24227 ;
  assign n24229 = n6523 & ~n7810 ;
  assign n24230 = n3324 | n12035 ;
  assign n24231 = n13242 | n24230 ;
  assign n24232 = n6145 & ~n6635 ;
  assign n24233 = n12334 ^ n442 ^ 1'b0 ;
  assign n24234 = n2319 & n24233 ;
  assign n24235 = ( x142 & ~n6962 ) | ( x142 & n24234 ) | ( ~n6962 & n24234 ) ;
  assign n24236 = n21004 & n21843 ;
  assign n24237 = n7698 & n24236 ;
  assign n24238 = n21495 ^ n20811 ^ 1'b0 ;
  assign n24239 = n11083 ^ n8956 ^ 1'b0 ;
  assign n24240 = n13607 | n24239 ;
  assign n24241 = n14668 ^ n1668 ^ 1'b0 ;
  assign n24242 = ( n7162 & n7251 ) | ( n7162 & ~n12268 ) | ( n7251 & ~n12268 ) ;
  assign n24243 = n1035 & ~n6327 ;
  assign n24244 = ( n10400 & ~n12975 ) | ( n10400 & n17285 ) | ( ~n12975 & n17285 ) ;
  assign n24245 = n2848 & n12314 ;
  assign n24246 = n24245 ^ n913 ^ 1'b0 ;
  assign n24247 = ~n8697 & n24246 ;
  assign n24248 = n24247 ^ n14072 ^ 1'b0 ;
  assign n24249 = n5865 | n24248 ;
  assign n24250 = n2944 | n3043 ;
  assign n24251 = n4914 & ~n24250 ;
  assign n24252 = n4501 & n17156 ;
  assign n24253 = n24251 & n24252 ;
  assign n24255 = n6493 & ~n12824 ;
  assign n24256 = ~n3349 & n24255 ;
  assign n24257 = ~n8365 & n24256 ;
  assign n24254 = ~n3796 & n19352 ;
  assign n24258 = n24257 ^ n24254 ^ 1'b0 ;
  assign n24259 = n19199 ^ n6403 ^ 1'b0 ;
  assign n24260 = n9057 & ~n24259 ;
  assign n24261 = n13950 ^ n6000 ^ 1'b0 ;
  assign n24262 = n23712 | n24261 ;
  assign n24263 = n11638 ^ n10203 ^ 1'b0 ;
  assign n24264 = n24263 ^ n6558 ^ 1'b0 ;
  assign n24265 = n12242 & n24264 ;
  assign n24266 = n17746 ^ n8956 ^ 1'b0 ;
  assign n24267 = x151 & ~n24266 ;
  assign n24268 = x149 & n18097 ;
  assign n24269 = n11312 & n24268 ;
  assign n24270 = n24269 ^ n6679 ^ 1'b0 ;
  assign n24271 = n20320 & ~n24270 ;
  assign n24272 = ~n24267 & n24271 ;
  assign n24273 = ~n4999 & n22527 ;
  assign n24274 = ~n6281 & n21728 ;
  assign n24275 = n3567 ^ n3274 ^ 1'b0 ;
  assign n24276 = n3272 & ~n7496 ;
  assign n24277 = n15183 & n24276 ;
  assign n24278 = n14888 ^ n8872 ^ 1'b0 ;
  assign n24279 = n19792 ^ n14594 ^ 1'b0 ;
  assign n24280 = x92 & ~n3171 ;
  assign n24282 = ~n2110 & n6651 ;
  assign n24283 = n24282 ^ n9327 ^ 1'b0 ;
  assign n24281 = n6038 & n8014 ;
  assign n24284 = n24283 ^ n24281 ^ 1'b0 ;
  assign n24285 = n14608 ^ n5325 ^ 1'b0 ;
  assign n24286 = n14812 ^ n8477 ^ 1'b0 ;
  assign n24287 = n10330 | n20595 ;
  assign n24288 = n24287 ^ n11140 ^ 1'b0 ;
  assign n24290 = ~n327 & n1780 ;
  assign n24291 = ~n11891 & n24290 ;
  assign n24292 = n5413 & ~n24291 ;
  assign n24289 = ~n1988 & n6200 ;
  assign n24293 = n24292 ^ n24289 ^ 1'b0 ;
  assign n24294 = n5021 & n24293 ;
  assign n24295 = x24 & ~n13983 ;
  assign n24296 = n24295 ^ n7753 ^ 1'b0 ;
  assign n24297 = n7929 ^ n872 ^ 1'b0 ;
  assign n24298 = n10038 & n24297 ;
  assign n24299 = x92 & ~n4796 ;
  assign n24300 = n16774 & n24299 ;
  assign n24301 = n6174 & ~n9307 ;
  assign n24302 = n786 & n24301 ;
  assign n24303 = ~n2731 & n24302 ;
  assign n24304 = n24303 ^ n5970 ^ 1'b0 ;
  assign n24305 = n1977 & ~n18782 ;
  assign n24306 = n18508 & n24305 ;
  assign n24308 = ~n734 & n13507 ;
  assign n24309 = n734 & n24308 ;
  assign n24307 = n2892 | n21016 ;
  assign n24310 = n24309 ^ n24307 ^ 1'b0 ;
  assign n24311 = n24070 ^ n3298 ^ 1'b0 ;
  assign n24312 = n24243 ^ n11661 ^ 1'b0 ;
  assign n24313 = n9975 & n19296 ;
  assign n24314 = ~n11244 & n24313 ;
  assign n24315 = n18833 | n19526 ;
  assign n24316 = n24315 ^ n9066 ^ 1'b0 ;
  assign n24317 = n10657 & ~n14661 ;
  assign n24318 = ~n18502 & n23979 ;
  assign n24319 = ~n2566 & n8341 ;
  assign n24320 = n18364 & ~n24319 ;
  assign n24324 = n12448 ^ n3284 ^ x51 ;
  assign n24321 = n17822 ^ n6259 ^ n5793 ;
  assign n24322 = n24321 ^ n9654 ^ 1'b0 ;
  assign n24323 = n1321 & n24322 ;
  assign n24325 = n24324 ^ n24323 ^ 1'b0 ;
  assign n24326 = n1148 & n21950 ;
  assign n24327 = ~n1148 & n24326 ;
  assign n24328 = n24327 ^ n7818 ^ 1'b0 ;
  assign n24329 = n18882 & ~n24328 ;
  assign n24330 = ~n5826 & n6326 ;
  assign n24331 = n12221 & n24330 ;
  assign n24332 = ~n7193 & n18459 ;
  assign n24333 = n20802 & n24332 ;
  assign n24335 = n2073 & n14686 ;
  assign n24336 = n24335 ^ n1423 ^ 1'b0 ;
  assign n24334 = n2089 & n4451 ;
  assign n24337 = n24336 ^ n24334 ^ 1'b0 ;
  assign n24338 = n10675 ^ n4491 ^ 1'b0 ;
  assign n24339 = n22905 ^ n2663 ^ 1'b0 ;
  assign n24340 = ~n6471 & n24339 ;
  assign n24341 = n4613 & ~n13822 ;
  assign n24342 = ~n8692 & n10706 ;
  assign n24343 = n15817 ^ n14914 ^ 1'b0 ;
  assign n24344 = n2972 & ~n21549 ;
  assign n24345 = n24344 ^ n1347 ^ 1'b0 ;
  assign n24347 = n14689 ^ n1052 ^ 1'b0 ;
  assign n24348 = n15447 & ~n24347 ;
  assign n24349 = ( n17285 & n24242 ) | ( n17285 & n24348 ) | ( n24242 & n24348 ) ;
  assign n24350 = ~n5393 & n24349 ;
  assign n24346 = ~n4598 & n23961 ;
  assign n24351 = n24350 ^ n24346 ^ 1'b0 ;
  assign n24352 = n16981 & ~n23526 ;
  assign n24353 = n1974 & ~n4579 ;
  assign n24354 = n4617 & ~n8756 ;
  assign n24355 = n10501 & ~n24354 ;
  assign n24356 = n7475 & n13308 ;
  assign n24357 = n24356 ^ n19261 ^ 1'b0 ;
  assign n24358 = n1360 ^ n895 ^ 1'b0 ;
  assign n24359 = n6859 & ~n24358 ;
  assign n24360 = ~n3305 & n11501 ;
  assign n24361 = n24360 ^ n9985 ^ 1'b0 ;
  assign n24362 = n24361 ^ n23094 ^ 1'b0 ;
  assign n24363 = ~n12938 & n24362 ;
  assign n24364 = ~n11675 & n13054 ;
  assign n24365 = x106 & n24364 ;
  assign n24366 = n6824 & n24365 ;
  assign n24367 = n22109 & ~n24366 ;
  assign n24368 = n4577 & n14593 ;
  assign n24369 = n16683 & n22660 ;
  assign n24370 = n5588 ^ n1037 ^ 1'b0 ;
  assign n24371 = n4257 & n12574 ;
  assign n24372 = n24370 & ~n24371 ;
  assign n24373 = n24369 & n24372 ;
  assign n24374 = n17366 ^ n5468 ^ 1'b0 ;
  assign n24375 = x68 & n11073 ;
  assign n24376 = ~n24374 & n24375 ;
  assign n24377 = n500 & n5796 ;
  assign n24378 = n4459 & n24377 ;
  assign n24379 = ~n8544 & n15095 ;
  assign n24380 = n24379 ^ n18195 ^ n772 ;
  assign n24381 = n4180 & ~n13657 ;
  assign n24382 = ~n2312 & n24381 ;
  assign n24383 = ~n4411 & n7608 ;
  assign n24384 = ~n8619 & n24383 ;
  assign n24385 = n22235 ^ n1977 ^ 1'b0 ;
  assign n24386 = ( n3511 & n8154 ) | ( n3511 & ~n9810 ) | ( n8154 & ~n9810 ) ;
  assign n24387 = n24386 ^ n6941 ^ 1'b0 ;
  assign n24388 = n5334 & n24387 ;
  assign n24389 = n6736 | n24388 ;
  assign n24390 = ~n2142 & n7970 ;
  assign n24391 = n14984 ^ n2531 ^ 1'b0 ;
  assign n24393 = n14352 ^ n482 ^ 1'b0 ;
  assign n24392 = ~x28 & n5356 ;
  assign n24394 = n24393 ^ n24392 ^ 1'b0 ;
  assign n24395 = n7482 & ~n18191 ;
  assign n24396 = n20505 & n24395 ;
  assign n24397 = n23497 & ~n24396 ;
  assign n24398 = n22893 ^ n21644 ^ 1'b0 ;
  assign n24399 = ~n3884 & n21377 ;
  assign n24400 = n24399 ^ n1573 ^ 1'b0 ;
  assign n24401 = n13325 ^ n1249 ^ 1'b0 ;
  assign n24402 = n24400 | n24401 ;
  assign n24403 = n5026 ^ n2310 ^ 1'b0 ;
  assign n24404 = ~n7571 & n24403 ;
  assign n24405 = n806 & n24404 ;
  assign n24408 = n24107 ^ n9052 ^ 1'b0 ;
  assign n24409 = n24408 ^ n13225 ^ 1'b0 ;
  assign n24406 = ~n417 & n4932 ;
  assign n24407 = n1809 & ~n24406 ;
  assign n24410 = n24409 ^ n24407 ^ 1'b0 ;
  assign n24411 = ( ~n7657 & n7982 ) | ( ~n7657 & n8295 ) | ( n7982 & n8295 ) ;
  assign n24412 = n24411 ^ n21857 ^ 1'b0 ;
  assign n24413 = n822 | n4714 ;
  assign n24414 = n24413 ^ n6039 ^ 1'b0 ;
  assign n24415 = n17979 & ~n24414 ;
  assign n24416 = n6370 & n24415 ;
  assign n24417 = n24416 ^ n18935 ^ 1'b0 ;
  assign n24418 = n9508 ^ n4582 ^ 1'b0 ;
  assign n24419 = n11696 ^ n8959 ^ 1'b0 ;
  assign n24420 = ~n4493 & n24419 ;
  assign n24421 = ( ~n4061 & n19954 ) | ( ~n4061 & n24420 ) | ( n19954 & n24420 ) ;
  assign n24422 = n1048 & ~n4783 ;
  assign n24423 = n10443 & n22305 ;
  assign n24424 = n14888 ^ n8963 ^ 1'b0 ;
  assign n24425 = n9609 & n24424 ;
  assign n24426 = n23802 ^ n4745 ^ 1'b0 ;
  assign n24427 = n24426 ^ x115 ^ 1'b0 ;
  assign n24428 = n608 | n2725 ;
  assign n24429 = n17593 & ~n24428 ;
  assign n24430 = n11207 & n24429 ;
  assign n24431 = x80 & n1644 ;
  assign n24432 = n24431 ^ n18216 ^ 1'b0 ;
  assign n24433 = x204 & ~n4095 ;
  assign n24434 = n24433 ^ n14991 ^ 1'b0 ;
  assign n24435 = n24434 ^ n9602 ^ 1'b0 ;
  assign n24436 = ~n1951 & n19921 ;
  assign n24437 = n24436 ^ n1321 ^ 1'b0 ;
  assign n24438 = n20238 | n24437 ;
  assign n24439 = n4416 | n24438 ;
  assign n24440 = n15075 ^ n1738 ^ 1'b0 ;
  assign n24441 = n13524 & n24440 ;
  assign n24442 = n5786 & n12804 ;
  assign n24443 = n14418 ^ n7391 ^ 1'b0 ;
  assign n24444 = ~n15081 & n24443 ;
  assign n24445 = n12356 & n24444 ;
  assign n24446 = n24445 ^ n16432 ^ 1'b0 ;
  assign n24447 = n6555 | n24446 ;
  assign n24448 = n24447 ^ n16163 ^ 1'b0 ;
  assign n24449 = n5985 | n13319 ;
  assign n24450 = ~n7058 & n7255 ;
  assign n24451 = ~n6494 & n24450 ;
  assign n24452 = n7940 & ~n24451 ;
  assign n24453 = n6851 & n13596 ;
  assign n24454 = n10813 ^ n6568 ^ 1'b0 ;
  assign n24455 = n4709 | n24454 ;
  assign n24456 = n1311 & ~n24455 ;
  assign n24457 = n3297 & n24456 ;
  assign n24458 = n24457 ^ n17846 ^ 1'b0 ;
  assign n24459 = n4862 ^ x151 ^ 1'b0 ;
  assign n24460 = n14289 ^ n512 ^ 1'b0 ;
  assign n24461 = n24459 & ~n24460 ;
  assign n24462 = n6106 & n24461 ;
  assign n24463 = n5904 | n23206 ;
  assign n24464 = n24463 ^ n10281 ^ 1'b0 ;
  assign n24465 = n2581 & ~n17455 ;
  assign n24466 = n13127 | n21733 ;
  assign n24467 = n24466 ^ n15436 ^ n12293 ;
  assign n24468 = n9717 | n24467 ;
  assign n24469 = n13443 ^ n6433 ^ 1'b0 ;
  assign n24470 = n15429 ^ n13129 ^ 1'b0 ;
  assign n24471 = n24470 ^ n20164 ^ 1'b0 ;
  assign n24472 = n3816 & ~n11175 ;
  assign n24473 = n24472 ^ n6102 ^ 1'b0 ;
  assign n24474 = n24471 & ~n24473 ;
  assign n24475 = n19593 ^ n16818 ^ 1'b0 ;
  assign n24476 = n18666 & n24475 ;
  assign n24477 = ~x220 & n365 ;
  assign n24478 = n18924 & n24477 ;
  assign n24479 = ~n14084 & n24478 ;
  assign n24480 = n15057 & n22021 ;
  assign n24481 = n24480 ^ n14241 ^ n3970 ;
  assign n24482 = n5357 | n7100 ;
  assign n24483 = n6964 & n24482 ;
  assign n24484 = n3140 & n24483 ;
  assign n24486 = ~n4207 & n8992 ;
  assign n24487 = n6904 & n24486 ;
  assign n24485 = n5440 | n9687 ;
  assign n24488 = n24487 ^ n24485 ^ 1'b0 ;
  assign n24489 = n18504 | n24488 ;
  assign n24490 = n24489 ^ n288 ^ 1'b0 ;
  assign n24491 = n7057 ^ n1227 ^ 1'b0 ;
  assign n24492 = n19892 & n24491 ;
  assign n24493 = n3102 & ~n24492 ;
  assign n24494 = n24493 ^ n17714 ^ 1'b0 ;
  assign n24495 = n2579 ^ n1689 ^ 1'b0 ;
  assign n24496 = n4431 & n24495 ;
  assign n24497 = ~n1772 & n24496 ;
  assign n24498 = ~n22901 & n24497 ;
  assign n24499 = n15601 & ~n20427 ;
  assign n24500 = n4408 & ~n5583 ;
  assign n24501 = n24500 ^ n2848 ^ 1'b0 ;
  assign n24502 = n24393 ^ n10886 ^ 1'b0 ;
  assign n24503 = n14826 & n15890 ;
  assign n24504 = ~n1634 & n24503 ;
  assign n24505 = n4393 | n5484 ;
  assign n24506 = n10325 | n24505 ;
  assign n24507 = n10081 & ~n24506 ;
  assign n24508 = n10790 ^ n4308 ^ 1'b0 ;
  assign n24510 = n4291 & n13820 ;
  assign n24509 = ~n6025 & n9438 ;
  assign n24511 = n24510 ^ n24509 ^ 1'b0 ;
  assign n24512 = n6685 & n17607 ;
  assign n24513 = n24512 ^ n12813 ^ 1'b0 ;
  assign n24514 = n12667 ^ n10712 ^ 1'b0 ;
  assign n24515 = n1103 & n24514 ;
  assign n24516 = n1038 & ~n24515 ;
  assign n24517 = n14093 ^ n4229 ^ 1'b0 ;
  assign n24518 = n18112 ^ n7713 ^ 1'b0 ;
  assign n24519 = n3009 & n22928 ;
  assign n24520 = n24519 ^ n6676 ^ 1'b0 ;
  assign n24521 = n17469 ^ n7223 ^ 1'b0 ;
  assign n24522 = n18201 & ~n24521 ;
  assign n24523 = x141 & n9416 ;
  assign n24524 = n21609 ^ n8978 ^ 1'b0 ;
  assign n24525 = n1599 | n24524 ;
  assign n24526 = ~n4493 & n24525 ;
  assign n24527 = n14327 & n16389 ;
  assign n24528 = n24527 ^ n3408 ^ 1'b0 ;
  assign n24529 = n4118 | n8281 ;
  assign n24530 = n3207 & n13267 ;
  assign n24531 = n11743 ^ n4803 ^ 1'b0 ;
  assign n24532 = n24530 & n24531 ;
  assign n24533 = n5774 & n24532 ;
  assign n24534 = ~n4267 & n18389 ;
  assign n24535 = n3465 | n5650 ;
  assign n24536 = n20097 & ~n24535 ;
  assign n24537 = n24536 ^ n13676 ^ n13445 ;
  assign n24538 = n18436 ^ n2210 ^ 1'b0 ;
  assign n24539 = n23627 | n24538 ;
  assign n24540 = ~n6756 & n13715 ;
  assign n24541 = n8626 ^ n8152 ^ n3834 ;
  assign n24542 = n14277 & n17582 ;
  assign n24543 = n24542 ^ n2018 ^ 1'b0 ;
  assign n24544 = n4466 & ~n11403 ;
  assign n24545 = n24544 ^ n9294 ^ 1'b0 ;
  assign n24546 = n11797 ^ n261 ^ 1'b0 ;
  assign n24547 = n19913 & ~n24523 ;
  assign n24548 = n6531 | n13252 ;
  assign n24549 = n4238 & ~n24548 ;
  assign n24550 = n1826 & n8120 ;
  assign n24551 = n4867 & ~n13515 ;
  assign n24557 = n7680 | n9251 ;
  assign n24552 = n23774 ^ n6929 ^ 1'b0 ;
  assign n24553 = x228 & n11214 ;
  assign n24554 = n24553 ^ x11 ^ 1'b0 ;
  assign n24555 = n24554 ^ n16996 ^ 1'b0 ;
  assign n24556 = n24552 | n24555 ;
  assign n24558 = n24557 ^ n24556 ^ 1'b0 ;
  assign n24559 = ~n320 & n24558 ;
  assign n24560 = n5597 & ~n12094 ;
  assign n24561 = ( ~n2853 & n11891 ) | ( ~n2853 & n17669 ) | ( n11891 & n17669 ) ;
  assign n24562 = n2576 | n4791 ;
  assign n24563 = n24561 | n24562 ;
  assign n24564 = n13523 ^ n2972 ^ 1'b0 ;
  assign n24565 = n16349 | n24564 ;
  assign n24566 = n24565 ^ n11591 ^ 1'b0 ;
  assign n24567 = n1767 & ~n24566 ;
  assign n24568 = n24567 ^ n15539 ^ 1'b0 ;
  assign n24569 = n20393 ^ n16751 ^ n3223 ;
  assign n24570 = ~n3906 & n22965 ;
  assign n24571 = n10315 ^ n7787 ^ 1'b0 ;
  assign n24572 = n6310 & ~n7693 ;
  assign n24573 = n589 | n24572 ;
  assign n24574 = n24573 ^ n10049 ^ 1'b0 ;
  assign n24582 = x3 & ~n1283 ;
  assign n24583 = ~x3 & n24582 ;
  assign n24584 = n770 | n1077 ;
  assign n24585 = n24583 & ~n24584 ;
  assign n24586 = x151 & ~n887 ;
  assign n24587 = n887 & n24586 ;
  assign n24588 = n24585 & ~n24587 ;
  assign n24589 = n620 & ~n1698 ;
  assign n24590 = ~n620 & n24589 ;
  assign n24591 = n9986 & n24590 ;
  assign n24592 = n1027 & ~n24591 ;
  assign n24593 = n24588 & ~n24592 ;
  assign n24594 = ~n621 & n24593 ;
  assign n24577 = x240 & n738 ;
  assign n24578 = ~x240 & n24577 ;
  assign n24579 = ~n820 & n6165 ;
  assign n24580 = n24578 & n24579 ;
  assign n24581 = n9793 | n24580 ;
  assign n24595 = n24594 ^ n24581 ^ 1'b0 ;
  assign n24597 = x247 & n532 ;
  assign n24598 = ~n532 & n24597 ;
  assign n24599 = n24598 ^ n1233 ^ 1'b0 ;
  assign n24596 = n5685 & ~n12477 ;
  assign n24600 = n24599 ^ n24596 ^ 1'b0 ;
  assign n24601 = n6067 | n24600 ;
  assign n24602 = n24595 & ~n24601 ;
  assign n24575 = n4092 & n6893 ;
  assign n24576 = n24575 ^ n21462 ^ 1'b0 ;
  assign n24603 = n24602 ^ n24576 ^ n5615 ;
  assign n24604 = n6250 & n11500 ;
  assign n24605 = n24604 ^ n13431 ^ 1'b0 ;
  assign n24606 = n8322 & ~n24605 ;
  assign n24607 = n2412 ^ n1843 ^ 1'b0 ;
  assign n24608 = n3776 & ~n24607 ;
  assign n24609 = n24608 ^ n4162 ^ 1'b0 ;
  assign n24610 = n24606 & ~n24609 ;
  assign n24611 = n1538 | n7003 ;
  assign n24612 = n24611 ^ n19218 ^ 1'b0 ;
  assign n24613 = n24612 ^ n448 ^ 1'b0 ;
  assign n24614 = n1707 & n14080 ;
  assign n24615 = n8960 & n24614 ;
  assign n24616 = n24615 ^ n8225 ^ 1'b0 ;
  assign n24617 = ~n6888 & n21240 ;
  assign n24618 = n24616 & n24617 ;
  assign n24621 = ~n821 & n18998 ;
  assign n24619 = n14193 ^ n7430 ^ n5920 ;
  assign n24620 = n458 | n24619 ;
  assign n24622 = n24621 ^ n24620 ^ 1'b0 ;
  assign n24623 = n24501 & n24622 ;
  assign n24624 = n24623 ^ n6262 ^ 1'b0 ;
  assign n24625 = n9323 & ~n9528 ;
  assign n24626 = n24625 ^ n12559 ^ 1'b0 ;
  assign n24627 = n3727 & n22109 ;
  assign n24628 = n16751 ^ n6325 ^ n4265 ;
  assign n24629 = n23886 ^ n17373 ^ 1'b0 ;
  assign n24630 = n7513 & n24629 ;
  assign n24631 = n17152 ^ n13776 ^ 1'b0 ;
  assign n24632 = n12559 ^ n5427 ^ 1'b0 ;
  assign n24633 = n23149 & n24632 ;
  assign n24634 = n6889 ^ n2968 ^ 1'b0 ;
  assign n24635 = ~n891 & n24634 ;
  assign n24636 = n1295 | n10950 ;
  assign n24637 = n5207 & ~n24636 ;
  assign n24638 = n24637 ^ n21173 ^ 1'b0 ;
  assign n24639 = n18074 ^ n10240 ^ 1'b0 ;
  assign n24640 = ~n2632 & n24639 ;
  assign n24641 = ~n1507 & n3065 ;
  assign n24642 = n24641 ^ n4894 ^ 1'b0 ;
  assign n24643 = n1506 & ~n6489 ;
  assign n24644 = n24643 ^ n10338 ^ n7494 ;
  assign n24645 = n24644 ^ n16340 ^ n4119 ;
  assign n24646 = n24645 ^ n4536 ^ 1'b0 ;
  assign n24647 = n19282 & ~n24646 ;
  assign n24648 = n19024 & n24647 ;
  assign n24649 = n24648 ^ n8687 ^ 1'b0 ;
  assign n24650 = n6432 | n8139 ;
  assign n24651 = n24650 ^ n4341 ^ 1'b0 ;
  assign n24652 = ~n3850 & n24651 ;
  assign n24653 = n15300 ^ n6948 ^ 1'b0 ;
  assign n24654 = n10602 & ~n24653 ;
  assign n24655 = n934 & n24654 ;
  assign n24656 = n20585 | n24655 ;
  assign n24657 = n10611 & n24656 ;
  assign n24658 = n8182 & n24657 ;
  assign n24659 = n24658 ^ n14365 ^ n5982 ;
  assign n24660 = n21038 & n24659 ;
  assign n24661 = n3725 | n11390 ;
  assign n24662 = n24661 ^ n16630 ^ 1'b0 ;
  assign n24663 = ~n816 & n24662 ;
  assign n24664 = n24663 ^ n4466 ^ 1'b0 ;
  assign n24665 = ~n6079 & n17588 ;
  assign n24666 = n16179 | n24665 ;
  assign n24667 = n4652 & n24666 ;
  assign n24668 = n5617 | n20162 ;
  assign n24669 = n24668 ^ n12270 ^ 1'b0 ;
  assign n24670 = n6146 ^ n859 ^ 1'b0 ;
  assign n24672 = n7223 & n14854 ;
  assign n24673 = n8184 & n24672 ;
  assign n24671 = ~n9889 & n18880 ;
  assign n24674 = n24673 ^ n24671 ^ 1'b0 ;
  assign n24675 = ~n16483 & n24674 ;
  assign n24676 = ~n24262 & n24675 ;
  assign n24677 = ~n5030 & n18160 ;
  assign n24678 = n23610 ^ n7910 ^ 1'b0 ;
  assign n24679 = n2761 & ~n24678 ;
  assign n24680 = n5283 & n6891 ;
  assign n24681 = ~n24679 & n24680 ;
  assign n24682 = ~n4183 & n15452 ;
  assign n24683 = n11469 & n24682 ;
  assign n24687 = n9815 ^ n6612 ^ 1'b0 ;
  assign n24684 = n6642 ^ n6432 ^ n2955 ;
  assign n24685 = n9803 & n24684 ;
  assign n24686 = ~n22967 & n24685 ;
  assign n24688 = n24687 ^ n24686 ^ 1'b0 ;
  assign n24689 = n19359 ^ n5634 ^ 1'b0 ;
  assign n24690 = n7796 & n24689 ;
  assign n24691 = ( n3408 & n9190 ) | ( n3408 & ~n24690 ) | ( n9190 & ~n24690 ) ;
  assign n24692 = n13056 ^ n3879 ^ 1'b0 ;
  assign n24693 = n15193 & n24692 ;
  assign n24694 = n9870 & n21172 ;
  assign n24695 = n557 & n4310 ;
  assign n24696 = n24695 ^ n14378 ^ 1'b0 ;
  assign n24697 = n7791 & ~n24696 ;
  assign n24698 = ~n9582 & n24697 ;
  assign n24699 = n24698 ^ n5347 ^ 1'b0 ;
  assign n24700 = n24694 | n24699 ;
  assign n24701 = n14329 & n23883 ;
  assign n24702 = n2523 & n24701 ;
  assign n24703 = n24702 ^ n20723 ^ 1'b0 ;
  assign n24704 = n7634 & ~n12060 ;
  assign n24705 = n9108 & ~n19054 ;
  assign n24706 = n24705 ^ n19980 ^ 1'b0 ;
  assign n24707 = n2814 ^ x27 ^ 1'b0 ;
  assign n24708 = ~n7536 & n12291 ;
  assign n24709 = ~n3604 & n18998 ;
  assign n24710 = n24709 ^ n17812 ^ 1'b0 ;
  assign n24711 = n7646 & ~n24710 ;
  assign n24712 = n5755 | n12863 ;
  assign n24713 = n24711 | n24712 ;
  assign n24714 = n17082 ^ n1321 ^ 1'b0 ;
  assign n24715 = n2119 & ~n2489 ;
  assign n24716 = n24715 ^ n15021 ^ 1'b0 ;
  assign n24717 = n3727 & n11230 ;
  assign n24718 = n2379 & n24717 ;
  assign n24719 = n24718 ^ n6948 ^ 1'b0 ;
  assign n24720 = n8833 | n15579 ;
  assign n24721 = n24720 ^ x164 ^ 1'b0 ;
  assign n24722 = n7493 ^ n5195 ^ n4971 ;
  assign n24723 = n6471 | n24722 ;
  assign n24724 = n24723 ^ n8334 ^ 1'b0 ;
  assign n24725 = n24724 ^ n4881 ^ 1'b0 ;
  assign n24726 = n5844 & n24725 ;
  assign n24727 = n5062 ^ n3046 ^ 1'b0 ;
  assign n24728 = n5907 & ~n24727 ;
  assign n24729 = ~n5485 & n24728 ;
  assign n24730 = n24729 ^ n7863 ^ 1'b0 ;
  assign n24731 = n1867 & n5350 ;
  assign n24732 = ~n14573 & n24731 ;
  assign n24733 = n7449 ^ n3801 ^ 1'b0 ;
  assign n24734 = n13273 ^ n417 ^ 1'b0 ;
  assign n24735 = n1980 & n24734 ;
  assign n24736 = n8376 | n10996 ;
  assign n24737 = n13303 ^ n4524 ^ 1'b0 ;
  assign n24738 = x16 & x233 ;
  assign n24739 = ~x233 & n24738 ;
  assign n24740 = x222 | n24739 ;
  assign n24741 = x222 & ~n24740 ;
  assign n24742 = n3333 & n24741 ;
  assign n24743 = n24742 ^ n4955 ^ 1'b0 ;
  assign n24744 = x196 & ~n535 ;
  assign n24745 = ~x196 & n24744 ;
  assign n24746 = n2684 & ~n24745 ;
  assign n24747 = ~n2684 & n24746 ;
  assign n24748 = ~n329 & n387 ;
  assign n24749 = n329 & n24748 ;
  assign n24750 = n395 | n24749 ;
  assign n24751 = n24749 & ~n24750 ;
  assign n24752 = x229 & ~n24751 ;
  assign n24753 = n24751 & n24752 ;
  assign n24754 = n6375 | n24753 ;
  assign n24755 = n6375 & ~n24754 ;
  assign n24756 = n24747 | n24755 ;
  assign n24757 = n24747 & ~n24756 ;
  assign n24758 = ~n3197 & n24757 ;
  assign n24759 = ~n5255 & n24758 ;
  assign n24760 = n5255 & n24759 ;
  assign n24761 = x20 & n281 ;
  assign n24762 = ~n281 & n24761 ;
  assign n24763 = x109 & n24762 ;
  assign n24764 = n3687 & n24763 ;
  assign n24765 = ~n294 & n1501 ;
  assign n24766 = n294 & n24765 ;
  assign n24767 = n24764 & ~n24766 ;
  assign n24768 = n2076 & n24767 ;
  assign n24769 = n4385 & ~n24768 ;
  assign n24770 = ~n4385 & n24769 ;
  assign n24771 = n24760 | n24770 ;
  assign n24772 = n24760 & ~n24771 ;
  assign n24773 = n24743 & ~n24772 ;
  assign n24774 = n24773 ^ n3229 ^ 1'b0 ;
  assign n24775 = n24774 ^ n8369 ^ 1'b0 ;
  assign n24776 = n17856 | n24775 ;
  assign n24777 = n1973 & ~n24776 ;
  assign n24778 = n18148 ^ n7003 ^ n1720 ;
  assign n24779 = n24777 & ~n24778 ;
  assign n24780 = n5389 & n24779 ;
  assign n24781 = n3957 | n6003 ;
  assign n24782 = n22458 ^ n21358 ^ 1'b0 ;
  assign n24783 = n24781 & n24782 ;
  assign n24784 = ~n1632 & n10852 ;
  assign n24785 = n6362 & n24784 ;
  assign n24786 = n24785 ^ n20344 ^ 1'b0 ;
  assign n24787 = n15193 & ~n24786 ;
  assign n24788 = n11697 ^ n1507 ^ 1'b0 ;
  assign n24789 = n2058 & ~n24788 ;
  assign n24790 = n15039 ^ n4577 ^ 1'b0 ;
  assign n24791 = ~n9916 & n24790 ;
  assign n24792 = ( n6152 & n8883 ) | ( n6152 & n21437 ) | ( n8883 & n21437 ) ;
  assign n24793 = n24792 ^ n3768 ^ 1'b0 ;
  assign n24794 = n19097 & ~n24793 ;
  assign n24795 = n425 & n1671 ;
  assign n24796 = ~n10328 & n24795 ;
  assign n24797 = n5435 | n24796 ;
  assign n24798 = n7753 & ~n9799 ;
  assign n24799 = n24798 ^ n16163 ^ 1'b0 ;
  assign n24800 = n2164 & ~n5372 ;
  assign n24801 = n24800 ^ n6140 ^ 1'b0 ;
  assign n24802 = n9455 | n16556 ;
  assign n24803 = n4406 | n12829 ;
  assign n24804 = n11014 | n18506 ;
  assign n24805 = n11458 | n24804 ;
  assign n24806 = n1602 & n4444 ;
  assign n24807 = ~n6116 & n24806 ;
  assign n24808 = ~n1685 & n24807 ;
  assign n24809 = n24808 ^ n13761 ^ 1'b0 ;
  assign n24810 = n4611 & ~n8559 ;
  assign n24811 = n14433 ^ n6442 ^ n3159 ;
  assign n24812 = n8008 & n18167 ;
  assign n24813 = n18159 ^ n12841 ^ 1'b0 ;
  assign n24814 = n8010 & n24813 ;
  assign n24816 = n3073 & n12577 ;
  assign n24815 = n17038 | n21099 ;
  assign n24817 = n24816 ^ n24815 ^ 1'b0 ;
  assign n24818 = n13046 ^ n2968 ^ 1'b0 ;
  assign n24819 = n19046 ^ n9295 ^ 1'b0 ;
  assign n24820 = ~n7404 & n9311 ;
  assign n24821 = n24820 ^ n5559 ^ 1'b0 ;
  assign n24822 = n24819 & ~n24821 ;
  assign n24823 = ~n8223 & n24822 ;
  assign n24824 = n24823 ^ n4822 ^ 1'b0 ;
  assign n24825 = n492 & ~n22118 ;
  assign n24826 = ~n3050 & n22519 ;
  assign n24827 = n23886 ^ n741 ^ 1'b0 ;
  assign n24828 = n14525 | n24827 ;
  assign n24829 = n2266 | n7756 ;
  assign n24830 = n24829 ^ n7189 ^ 1'b0 ;
  assign n24831 = n24830 ^ n21573 ^ n633 ;
  assign n24832 = n1869 & ~n20277 ;
  assign n24833 = n2326 & ~n5694 ;
  assign n24834 = n24833 ^ n20310 ^ 1'b0 ;
  assign n24835 = n24834 ^ n18075 ^ 1'b0 ;
  assign n24836 = n3801 & ~n24835 ;
  assign n24837 = n1027 & ~n10135 ;
  assign n24838 = n16777 ^ n6602 ^ 1'b0 ;
  assign n24839 = n24837 & n24838 ;
  assign n24840 = n21386 ^ n4024 ^ 1'b0 ;
  assign n24841 = n23645 & ~n24840 ;
  assign n24842 = n24841 ^ n21076 ^ 1'b0 ;
  assign n24843 = n1236 | n11266 ;
  assign n24844 = n337 | n24843 ;
  assign n24845 = n24844 ^ n12850 ^ 1'b0 ;
  assign n24846 = n4623 | n24845 ;
  assign n24847 = n5297 & ~n17106 ;
  assign n24848 = n12917 & n24847 ;
  assign n24849 = n21755 ^ n519 ^ 1'b0 ;
  assign n24850 = n24848 | n24849 ;
  assign n24851 = n3232 | n16898 ;
  assign n24852 = n15681 | n24851 ;
  assign n24853 = n15636 & ~n24792 ;
  assign n24854 = n7113 ^ n1336 ^ 1'b0 ;
  assign n24855 = x136 & ~n12816 ;
  assign n24856 = ~n23893 & n24855 ;
  assign n24857 = n24856 ^ n19621 ^ 1'b0 ;
  assign n24858 = n1012 & n2893 ;
  assign n24859 = ~n1012 & n24858 ;
  assign n24860 = n10591 & ~n24859 ;
  assign n24861 = ~n10591 & n24860 ;
  assign n24862 = n8881 | n24861 ;
  assign n24863 = n14938 & ~n24862 ;
  assign n24864 = ~n24857 & n24863 ;
  assign n24865 = ~n4962 & n12295 ;
  assign n24867 = ~n1686 & n9261 ;
  assign n24866 = n387 & ~n8237 ;
  assign n24868 = n24867 ^ n24866 ^ 1'b0 ;
  assign n24869 = n444 & ~n24868 ;
  assign n24870 = n4576 ^ n2861 ^ 1'b0 ;
  assign n24871 = n2610 & n24870 ;
  assign n24872 = ~n3649 & n5385 ;
  assign n24873 = ~n24871 & n24872 ;
  assign n24874 = n9171 & n18627 ;
  assign n24875 = n3545 & ~n4980 ;
  assign n24876 = n15903 ^ n12230 ^ 1'b0 ;
  assign n24877 = n14658 | n24876 ;
  assign n24878 = n10920 & ~n24877 ;
  assign n24879 = n3620 ^ n1249 ^ 1'b0 ;
  assign n24880 = n24879 ^ n22025 ^ 1'b0 ;
  assign n24881 = x132 & ~n2334 ;
  assign n24882 = n2959 & ~n24881 ;
  assign n24883 = n22538 ^ n2546 ^ 1'b0 ;
  assign n24884 = n2129 & n17755 ;
  assign n24885 = n2143 & n10144 ;
  assign n24886 = n24884 & n24885 ;
  assign n24887 = n688 & n1797 ;
  assign n24888 = n12193 ^ n3877 ^ 1'b0 ;
  assign n24889 = n5038 ^ n4967 ^ 1'b0 ;
  assign n24890 = n17975 & n19085 ;
  assign n24891 = n11149 & n24890 ;
  assign n24892 = ~n24889 & n24891 ;
  assign n24893 = ~n3043 & n15638 ;
  assign n24899 = n5110 & ~n16672 ;
  assign n24897 = n11851 ^ n4913 ^ 1'b0 ;
  assign n24894 = n19007 ^ n6790 ^ 1'b0 ;
  assign n24895 = n1906 & ~n24894 ;
  assign n24896 = n23885 & n24895 ;
  assign n24898 = n24897 ^ n24896 ^ 1'b0 ;
  assign n24900 = n24899 ^ n24898 ^ 1'b0 ;
  assign n24901 = n24893 & n24900 ;
  assign n24908 = n23892 ^ n6224 ^ 1'b0 ;
  assign n24909 = n17998 & n24908 ;
  assign n24910 = ~n24908 & n24909 ;
  assign n24902 = n4755 & n7529 ;
  assign n24903 = ~n7529 & n24902 ;
  assign n24904 = ~n1082 & n24903 ;
  assign n24905 = n22193 ^ n7667 ^ 1'b0 ;
  assign n24906 = n24904 & ~n24905 ;
  assign n24907 = ~n6829 & n24906 ;
  assign n24911 = n24910 ^ n24907 ^ 1'b0 ;
  assign n24912 = n1158 & n1743 ;
  assign n24913 = ~n1158 & n24912 ;
  assign n24914 = n10875 & ~n24913 ;
  assign n24915 = ~n14731 & n24914 ;
  assign n24916 = ~n24911 & n24915 ;
  assign n24917 = ( n13821 & ~n16706 ) | ( n13821 & n24916 ) | ( ~n16706 & n24916 ) ;
  assign n24918 = n3477 | n23165 ;
  assign n24919 = n24918 ^ n4375 ^ 1'b0 ;
  assign n24920 = ~n1082 & n16688 ;
  assign n24921 = n24920 ^ n15884 ^ 1'b0 ;
  assign n24922 = n13506 | n15715 ;
  assign n24923 = n16209 ^ n7984 ^ 1'b0 ;
  assign n24924 = n8801 ^ n3872 ^ 1'b0 ;
  assign n24926 = x29 & ~n11709 ;
  assign n24925 = n2743 | n3171 ;
  assign n24927 = n24926 ^ n24925 ^ 1'b0 ;
  assign n24928 = ~n22461 & n24927 ;
  assign n24929 = n12737 & n13290 ;
  assign n24930 = ~n20477 & n24929 ;
  assign n24931 = ~n3533 & n18045 ;
  assign n24932 = ~n13714 & n24638 ;
  assign n24933 = n928 & n23144 ;
  assign n24934 = n5625 & n24933 ;
  assign n24935 = ~n1656 & n2314 ;
  assign n24936 = n24935 ^ n10056 ^ 1'b0 ;
  assign n24937 = ~n3989 & n24936 ;
  assign n24938 = n10507 ^ n5154 ^ 1'b0 ;
  assign n24939 = n24545 ^ n12058 ^ 1'b0 ;
  assign n24940 = n6428 ^ x17 ^ 1'b0 ;
  assign n24941 = n8995 & n24940 ;
  assign n24942 = n5897 ^ x199 ^ 1'b0 ;
  assign n24943 = n8019 ^ n5012 ^ 1'b0 ;
  assign n24944 = n6836 | n24943 ;
  assign n24945 = n9923 & ~n24944 ;
  assign n24946 = ~n18441 & n22715 ;
  assign n24947 = ~n20868 & n24946 ;
  assign n24948 = n9012 & ~n24947 ;
  assign n24949 = n24948 ^ n10194 ^ 1'b0 ;
  assign n24950 = n2325 | n21121 ;
  assign n24951 = n18232 ^ n5991 ^ 1'b0 ;
  assign n24952 = n23977 ^ n6355 ^ 1'b0 ;
  assign n24953 = n2669 & n6300 ;
  assign n24954 = n24953 ^ n4546 ^ 1'b0 ;
  assign n24955 = n8182 | n16362 ;
  assign n24956 = n24955 ^ n16144 ^ 1'b0 ;
  assign n24957 = n6970 | n24956 ;
  assign n24958 = n24954 | n24957 ;
  assign n24959 = n18125 ^ n18061 ^ 1'b0 ;
  assign n24960 = ~n11792 & n21509 ;
  assign n24961 = n8517 & ~n24960 ;
  assign n24962 = n7947 & n16497 ;
  assign n24963 = n679 | n1790 ;
  assign n24964 = n5364 | n24963 ;
  assign n24965 = n5420 & ~n23551 ;
  assign n24966 = n14231 & n24965 ;
  assign n24967 = n10236 & ~n24966 ;
  assign n24968 = n4822 & ~n18741 ;
  assign n24969 = n6413 & ~n24968 ;
  assign n24970 = n5507 & ~n11570 ;
  assign n24971 = n24970 ^ n10523 ^ 1'b0 ;
  assign n24972 = n3402 & n24971 ;
  assign n24973 = n24972 ^ n24261 ^ 1'b0 ;
  assign n24974 = n3247 ^ n1596 ^ 1'b0 ;
  assign n24975 = ~n12735 & n24974 ;
  assign n24976 = n24975 ^ n10523 ^ n9665 ;
  assign n24977 = n24976 ^ n2801 ^ 1'b0 ;
  assign n24978 = n9892 ^ n4664 ^ n621 ;
  assign n24979 = x217 & ~n1133 ;
  assign n24980 = n12882 & n24979 ;
  assign n24981 = n21480 | n24980 ;
  assign n24982 = n24978 | n24981 ;
  assign n24983 = n3417 & ~n19511 ;
  assign n24984 = ~n1423 & n24983 ;
  assign n24985 = n17246 | n24984 ;
  assign n24986 = n24985 ^ n14986 ^ 1'b0 ;
  assign n24987 = n24986 ^ n11210 ^ 1'b0 ;
  assign n24988 = n1159 | n20414 ;
  assign n24989 = ~n16463 & n16506 ;
  assign n24990 = x181 & n4473 ;
  assign n24991 = n24990 ^ n5278 ^ 1'b0 ;
  assign n24992 = n4828 ^ n2660 ^ 1'b0 ;
  assign n24993 = ~n13589 & n24992 ;
  assign n24994 = ( ~n1361 & n1521 ) | ( ~n1361 & n24993 ) | ( n1521 & n24993 ) ;
  assign n24995 = n8530 ^ n1017 ^ 1'b0 ;
  assign n24996 = n5648 | n24995 ;
  assign n24997 = n14399 | n24996 ;
  assign n24998 = x34 & n22343 ;
  assign n25001 = n7588 | n14947 ;
  assign n25002 = n25001 ^ n817 ^ 1'b0 ;
  assign n25003 = n13354 & ~n25002 ;
  assign n24999 = n14022 ^ n7202 ^ 1'b0 ;
  assign n25000 = n24999 ^ n22872 ^ n2712 ;
  assign n25004 = n25003 ^ n25000 ^ 1'b0 ;
  assign n25005 = n2186 ^ x218 ^ 1'b0 ;
  assign n25006 = ~n6605 & n25005 ;
  assign n25007 = n3791 ^ n2237 ^ 1'b0 ;
  assign n25008 = n15580 | n22767 ;
  assign n25009 = n25007 & ~n25008 ;
  assign n25010 = ~n1791 & n25009 ;
  assign n25011 = n14417 | n17348 ;
  assign n25012 = n19311 | n25011 ;
  assign n25013 = n20997 ^ n18314 ^ 1'b0 ;
  assign n25015 = ( ~n15323 & n18314 ) | ( ~n15323 & n23341 ) | ( n18314 & n23341 ) ;
  assign n25014 = n6287 & ~n13491 ;
  assign n25016 = n25015 ^ n25014 ^ 1'b0 ;
  assign n25017 = n4122 & ~n12888 ;
  assign n25018 = n4606 & ~n7477 ;
  assign n25019 = n796 | n19138 ;
  assign n25020 = n21361 & ~n25019 ;
  assign n25022 = n6423 ^ n2148 ^ 1'b0 ;
  assign n25023 = n6617 | n25022 ;
  assign n25021 = n10070 | n13125 ;
  assign n25024 = n25023 ^ n25021 ^ 1'b0 ;
  assign n25025 = ~x191 & n8568 ;
  assign n25026 = n12360 ^ n6583 ^ 1'b0 ;
  assign n25027 = n6702 ^ n4466 ^ 1'b0 ;
  assign n25028 = n13941 & n25027 ;
  assign n25029 = n9024 & ~n9612 ;
  assign n25030 = n4521 & ~n8808 ;
  assign n25031 = ( ~n17378 & n17837 ) | ( ~n17378 & n25030 ) | ( n17837 & n25030 ) ;
  assign n25032 = n24507 | n25031 ;
  assign n25033 = n5908 & ~n7021 ;
  assign n25034 = n25033 ^ n19000 ^ 1'b0 ;
  assign n25035 = n4529 & ~n7128 ;
  assign n25036 = n7766 & n25035 ;
  assign n25037 = ~n6471 & n16798 ;
  assign n25038 = ~n509 & n25037 ;
  assign n25039 = n25036 & n25038 ;
  assign n25040 = ~n5220 & n13763 ;
  assign n25041 = n25040 ^ n24022 ^ 1'b0 ;
  assign n25042 = n19797 | n25041 ;
  assign n25043 = ~n20295 & n21848 ;
  assign n25044 = ~n4149 & n8223 ;
  assign n25045 = n25044 ^ n20292 ^ 1'b0 ;
  assign n25046 = n10413 | n10794 ;
  assign n25047 = n15212 ^ n5976 ^ 1'b0 ;
  assign n25048 = n21034 & ~n25047 ;
  assign n25049 = n2333 | n6491 ;
  assign n25050 = n25049 ^ n15584 ^ 1'b0 ;
  assign n25051 = ~n8771 & n11651 ;
  assign n25052 = n25051 ^ n9460 ^ 1'b0 ;
  assign n25053 = n25052 ^ n22316 ^ 1'b0 ;
  assign n25054 = n24444 ^ n3434 ^ 1'b0 ;
  assign n25055 = n3265 & n5688 ;
  assign n25056 = ~n25054 & n25055 ;
  assign n25057 = n14612 & ~n23159 ;
  assign n25058 = ~n19368 & n25057 ;
  assign n25059 = n11887 | n19819 ;
  assign n25060 = n25059 ^ n1508 ^ 1'b0 ;
  assign n25061 = n8277 ^ n1663 ^ 1'b0 ;
  assign n25062 = n11207 & ~n25061 ;
  assign n25063 = n11274 ^ n9508 ^ 1'b0 ;
  assign n25064 = n4923 | n25062 ;
  assign n25065 = ~n526 & n1947 ;
  assign n25066 = ~n3143 & n25065 ;
  assign n25067 = n4003 | n14187 ;
  assign n25068 = n25066 & ~n25067 ;
  assign n25069 = n19131 | n25068 ;
  assign n25070 = n8094 | n15094 ;
  assign n25071 = n10822 | n24868 ;
  assign n25072 = n3629 & n6882 ;
  assign n25073 = n11042 | n25072 ;
  assign n25079 = ~n6978 & n22567 ;
  assign n25080 = n6978 & n25079 ;
  assign n25081 = n3390 & n25080 ;
  assign n25074 = n3994 & n6442 ;
  assign n25075 = ~n6442 & n25074 ;
  assign n25076 = n20419 & ~n25075 ;
  assign n25077 = x178 & ~n25076 ;
  assign n25078 = n25076 & n25077 ;
  assign n25082 = n25081 ^ n25078 ^ n363 ;
  assign n25083 = n14675 ^ n6493 ^ 1'b0 ;
  assign n25084 = n7636 & n14848 ;
  assign n25085 = n25084 ^ n18921 ^ 1'b0 ;
  assign n25087 = n22861 ^ n18165 ^ 1'b0 ;
  assign n25086 = n633 & ~n21957 ;
  assign n25088 = n25087 ^ n25086 ^ 1'b0 ;
  assign n25089 = n4652 & n6994 ;
  assign n25090 = ~n5419 & n5929 ;
  assign n25091 = ( ~n18861 & n22161 ) | ( ~n18861 & n25090 ) | ( n22161 & n25090 ) ;
  assign n25093 = n5946 ^ n1275 ^ 1'b0 ;
  assign n25094 = n4475 | n25093 ;
  assign n25095 = n2021 | n25094 ;
  assign n25096 = n25095 ^ n2918 ^ 1'b0 ;
  assign n25092 = ~n5849 & n6780 ;
  assign n25097 = n25096 ^ n25092 ^ 1'b0 ;
  assign n25098 = n8195 | n9239 ;
  assign n25099 = n25098 ^ n17680 ^ 1'b0 ;
  assign n25100 = x115 | n12230 ;
  assign n25101 = n5031 & ~n5553 ;
  assign n25102 = n25101 ^ n16565 ^ 1'b0 ;
  assign n25103 = ~n16729 & n21630 ;
  assign n25104 = n7988 & ~n12506 ;
  assign n25105 = ~n512 & n25104 ;
  assign n25106 = n21617 ^ x226 ^ 1'b0 ;
  assign n25107 = n4475 & n15167 ;
  assign n25108 = n4671 | n11261 ;
  assign n25109 = n4671 & ~n25108 ;
  assign n25110 = n25109 ^ n9253 ^ 1'b0 ;
  assign n25111 = n2068 & ~n2889 ;
  assign n25112 = n2889 & n25111 ;
  assign n25113 = n11069 | n25112 ;
  assign n25114 = n11069 & ~n25113 ;
  assign n25115 = n9148 | n25114 ;
  assign n25116 = n25110 | n25115 ;
  assign n25117 = n1419 | n17935 ;
  assign n25118 = n5105 & n5810 ;
  assign n25119 = n20168 ^ n6413 ^ 1'b0 ;
  assign n25120 = n11668 ^ n399 ^ 1'b0 ;
  assign n25121 = n10488 ^ n7359 ^ 1'b0 ;
  assign n25122 = n11220 & ~n25121 ;
  assign n25123 = n21851 & ~n25122 ;
  assign n25124 = n3197 & ~n16861 ;
  assign n25125 = n1775 & ~n3399 ;
  assign n25126 = n25125 ^ n1195 ^ 1'b0 ;
  assign n25127 = n3881 ^ n1725 ^ 1'b0 ;
  assign n25128 = n11783 | n25127 ;
  assign n25129 = n6812 | n25128 ;
  assign n25130 = n1689 ^ n281 ^ 1'b0 ;
  assign n25131 = n25130 ^ n18856 ^ 1'b0 ;
  assign n25132 = ~n25129 & n25131 ;
  assign n25133 = n25132 ^ n11719 ^ 1'b0 ;
  assign n25134 = n4520 & ~n5029 ;
  assign n25135 = x128 & ~n25134 ;
  assign n25136 = n3181 & ~n4952 ;
  assign n25137 = n8709 ^ n3710 ^ 1'b0 ;
  assign n25138 = n4913 & n25137 ;
  assign n25139 = n13030 ^ n12708 ^ n9817 ;
  assign n25140 = n15987 ^ n452 ^ 1'b0 ;
  assign n25141 = n4660 | n25140 ;
  assign n25142 = n17830 ^ n508 ^ 1'b0 ;
  assign n25143 = n561 & n25142 ;
  assign n25144 = n13003 | n14885 ;
  assign n25145 = n4465 & ~n21436 ;
  assign n25146 = n25145 ^ n14093 ^ 1'b0 ;
  assign n25147 = n13265 ^ n643 ^ 1'b0 ;
  assign n25148 = ~n805 & n15736 ;
  assign n25149 = n25148 ^ x29 ^ 1'b0 ;
  assign n25150 = n21415 ^ n2655 ^ 1'b0 ;
  assign n25151 = x248 & n21775 ;
  assign n25152 = n19976 & n25151 ;
  assign n25153 = n16175 | n17327 ;
  assign n25154 = ~n5369 & n10809 ;
  assign n25155 = ~n10144 & n25154 ;
  assign n25156 = ~n14641 & n25155 ;
  assign n25157 = ~n9276 & n25156 ;
  assign n25158 = n9123 & ~n22001 ;
  assign n25159 = n25158 ^ n8369 ^ 1'b0 ;
  assign n25160 = ( n3111 & ~n9875 ) | ( n3111 & n15318 ) | ( ~n9875 & n15318 ) ;
  assign n25161 = ~n1560 & n4730 ;
  assign n25162 = n7858 ^ n3062 ^ 1'b0 ;
  assign n25163 = ~n15419 & n25162 ;
  assign n25164 = n2004 | n8064 ;
  assign n25165 = n22925 ^ x75 ^ 1'b0 ;
  assign n25166 = n25164 | n25165 ;
  assign n25167 = n13294 ^ n3597 ^ 1'b0 ;
  assign n25168 = n5938 | n25167 ;
  assign n25169 = n20264 & ~n25168 ;
  assign n25170 = n8010 | n25169 ;
  assign n25171 = ~n1378 & n3604 ;
  assign n25172 = n3795 | n19349 ;
  assign n25173 = ~n934 & n22648 ;
  assign n25174 = n25173 ^ n771 ^ 1'b0 ;
  assign n25175 = n8277 & n13222 ;
  assign n25176 = n5440 ^ n2604 ^ 1'b0 ;
  assign n25177 = n11069 | n16140 ;
  assign n25178 = n25177 ^ n12607 ^ 1'b0 ;
  assign n25179 = ~n11635 & n25178 ;
  assign n25181 = n5840 | n23029 ;
  assign n25182 = n345 | n25181 ;
  assign n25180 = n4189 | n17973 ;
  assign n25183 = n25182 ^ n25180 ^ 1'b0 ;
  assign n25184 = n14771 ^ n633 ^ 1'b0 ;
  assign n25185 = n25183 & ~n25184 ;
  assign n25186 = n25185 ^ n13671 ^ 1'b0 ;
  assign n25187 = n9251 & n10611 ;
  assign n25188 = n25187 ^ n3780 ^ 1'b0 ;
  assign n25189 = ~n703 & n25188 ;
  assign n25190 = n7367 | n24047 ;
  assign n25191 = n25190 ^ n24193 ^ 1'b0 ;
  assign n25192 = ( n1345 & n7477 ) | ( n1345 & ~n10039 ) | ( n7477 & ~n10039 ) ;
  assign n25193 = n6254 & ~n9252 ;
  assign n25194 = n25192 & n25193 ;
  assign n25195 = n19994 ^ n10697 ^ 1'b0 ;
  assign n25196 = ~n21012 & n25195 ;
  assign n25197 = n25196 ^ n10781 ^ 1'b0 ;
  assign n25198 = ~n5207 & n21542 ;
  assign n25199 = n927 & ~n6174 ;
  assign n25200 = ~n25198 & n25199 ;
  assign n25201 = n2757 | n10613 ;
  assign n25202 = ~n4026 & n25201 ;
  assign n25203 = ~n2441 & n8925 ;
  assign n25204 = n1832 & ~n9105 ;
  assign n25205 = ~x88 & n25204 ;
  assign n25206 = n8001 | n15362 ;
  assign n25207 = n25206 ^ n23423 ^ n23045 ;
  assign n25208 = n8840 & ~n25207 ;
  assign n25209 = ( n2891 & n6267 ) | ( n2891 & ~n7183 ) | ( n6267 & ~n7183 ) ;
  assign n25210 = ( n8773 & n21979 ) | ( n8773 & n25209 ) | ( n21979 & n25209 ) ;
  assign n25211 = n20431 ^ n7482 ^ 1'b0 ;
  assign n25212 = n17238 ^ n833 ^ 1'b0 ;
  assign n25213 = n1758 & ~n4502 ;
  assign n25214 = n25213 ^ n10021 ^ 1'b0 ;
  assign n25215 = ~n2296 & n18005 ;
  assign n25216 = n25214 & n25215 ;
  assign n25217 = n6333 ^ n5734 ^ 1'b0 ;
  assign n25218 = n10382 & ~n25217 ;
  assign n25219 = n25218 ^ n16317 ^ 1'b0 ;
  assign n25220 = n7977 | n25219 ;
  assign n25221 = n10416 ^ n6014 ^ 1'b0 ;
  assign n25222 = n1429 & n8290 ;
  assign n25223 = n17219 & ~n25222 ;
  assign n25224 = n3888 | n8978 ;
  assign n25225 = n3888 & ~n25224 ;
  assign n25226 = n4763 & n11068 ;
  assign n25227 = n19130 ^ n2550 ^ 1'b0 ;
  assign n25228 = n24895 | n25227 ;
  assign n25229 = n22678 ^ n9598 ^ 1'b0 ;
  assign n25230 = n2254 | n25229 ;
  assign n25231 = n7723 ^ n7568 ^ 1'b0 ;
  assign n25232 = n7400 & n25231 ;
  assign n25233 = n3414 | n25232 ;
  assign n25234 = n809 & n21737 ;
  assign n25235 = n25234 ^ n14283 ^ 1'b0 ;
  assign n25236 = ~n3139 & n25235 ;
  assign n25237 = n3207 ^ n1738 ^ 1'b0 ;
  assign n25238 = n1304 | n25237 ;
  assign n25239 = n25238 ^ n2849 ^ 1'b0 ;
  assign n25240 = n472 & n6162 ;
  assign n25241 = n19777 ^ n10717 ^ n720 ;
  assign n25242 = n19591 ^ n3599 ^ 1'b0 ;
  assign n25243 = ~n2793 & n25242 ;
  assign n25244 = ~n8655 & n15641 ;
  assign n25245 = n25244 ^ n20870 ^ 1'b0 ;
  assign n25246 = n25243 & ~n25245 ;
  assign n25247 = x75 & n19570 ;
  assign n25248 = n8010 ^ n3437 ^ 1'b0 ;
  assign n25249 = ~n7436 & n8738 ;
  assign n25250 = n5943 | n25249 ;
  assign n25251 = n25250 ^ n7548 ^ 1'b0 ;
  assign n25252 = n25248 & ~n25251 ;
  assign n25253 = n6053 & n25252 ;
  assign n25254 = n25253 ^ n14103 ^ 1'b0 ;
  assign n25255 = n21387 ^ n7501 ^ 1'b0 ;
  assign n25256 = ~n22678 & n25255 ;
  assign n25257 = n22671 ^ n1297 ^ 1'b0 ;
  assign n25258 = n14177 & ~n25257 ;
  assign n25259 = n14245 & ~n25258 ;
  assign n25260 = ~n1928 & n23876 ;
  assign n25261 = ~n15187 & n25260 ;
  assign n25262 = ~n5192 & n6208 ;
  assign n25263 = n6858 | n25262 ;
  assign n25264 = n4162 & n7255 ;
  assign n25265 = n7695 & ~n25264 ;
  assign n25266 = n12371 ^ n335 ^ 1'b0 ;
  assign n25267 = n17373 & ~n25266 ;
  assign n25268 = ~n25265 & n25267 ;
  assign n25272 = n527 & ~n1663 ;
  assign n25273 = n15085 & n25272 ;
  assign n25274 = n25273 ^ n21755 ^ n9420 ;
  assign n25269 = n1994 & n2768 ;
  assign n25270 = n15533 ^ n5784 ^ 1'b0 ;
  assign n25271 = ~n25269 & n25270 ;
  assign n25275 = n25274 ^ n25271 ^ 1'b0 ;
  assign n25276 = n16384 & ~n25275 ;
  assign n25277 = n2794 | n17219 ;
  assign n25278 = n6878 & ~n25277 ;
  assign n25279 = n12088 | n25278 ;
  assign n25280 = n25279 ^ n9947 ^ 1'b0 ;
  assign n25281 = n25280 ^ n15809 ^ 1'b0 ;
  assign n25282 = n13696 ^ n1046 ^ 1'b0 ;
  assign n25283 = n5969 ^ n1898 ^ 1'b0 ;
  assign n25284 = n23917 ^ n11454 ^ 1'b0 ;
  assign n25285 = n25283 & n25284 ;
  assign n25286 = n11758 ^ n3872 ^ 1'b0 ;
  assign n25287 = n10167 ^ n8351 ^ 1'b0 ;
  assign n25288 = ~n7807 & n25287 ;
  assign n25289 = n25288 ^ n11512 ^ 1'b0 ;
  assign n25290 = n15589 | n25289 ;
  assign n25291 = n25290 ^ n22556 ^ 1'b0 ;
  assign n25292 = ~n5775 & n23221 ;
  assign n25293 = n25292 ^ n1638 ^ 1'b0 ;
  assign n25294 = n11608 & n25293 ;
  assign n25295 = n25294 ^ n17453 ^ 1'b0 ;
  assign n25296 = n8474 & n20772 ;
  assign n25297 = n25295 & n25296 ;
  assign n25298 = ~x105 & n25297 ;
  assign n25299 = n2589 & ~n17090 ;
  assign n25300 = n4741 & n21014 ;
  assign n25301 = n25300 ^ n2854 ^ 1'b0 ;
  assign n25302 = ~n6769 & n25301 ;
  assign n25303 = n7856 & ~n15772 ;
  assign n25304 = n25303 ^ n11873 ^ 1'b0 ;
  assign n25305 = ~n8622 & n25304 ;
  assign n25306 = ~n25302 & n25305 ;
  assign n25307 = n10027 ^ n909 ^ 1'b0 ;
  assign n25308 = n9398 & ~n21103 ;
  assign n25309 = n5405 & n13676 ;
  assign n25310 = ~n2861 & n19796 ;
  assign n25311 = n3140 & n8195 ;
  assign n25312 = n10954 ^ n3423 ^ 1'b0 ;
  assign n25313 = n6225 & n25312 ;
  assign n25314 = n3854 & n25313 ;
  assign n25315 = n16610 | n25314 ;
  assign n25316 = n11856 & ~n25315 ;
  assign n25317 = n25311 & ~n25316 ;
  assign n25326 = ~n5363 & n6551 ;
  assign n25327 = n5363 & n25326 ;
  assign n25318 = n1158 & n2159 ;
  assign n25319 = ~n2159 & n25318 ;
  assign n25320 = n594 | n25319 ;
  assign n25321 = n594 & ~n25320 ;
  assign n25322 = x37 & ~n25321 ;
  assign n25323 = n25321 & n25322 ;
  assign n25324 = n14689 | n25323 ;
  assign n25325 = n25324 ^ n9565 ^ 1'b0 ;
  assign n25328 = n25327 ^ n25325 ^ 1'b0 ;
  assign n25329 = n10555 | n25328 ;
  assign n25330 = n7443 & ~n25329 ;
  assign n25331 = n25330 ^ n18420 ^ 1'b0 ;
  assign n25332 = n8198 | n10932 ;
  assign n25333 = n25332 ^ n5781 ^ 1'b0 ;
  assign n25334 = n3156 & n9801 ;
  assign n25335 = n25334 ^ n1608 ^ 1'b0 ;
  assign n25336 = n4788 & n25335 ;
  assign n25337 = n25336 ^ n7266 ^ 1'b0 ;
  assign n25338 = n8493 & n25337 ;
  assign n25339 = n1383 & n25338 ;
  assign n25340 = ~n25333 & n25339 ;
  assign n25341 = n15847 ^ n6167 ^ 1'b0 ;
  assign n25342 = n8619 & n25341 ;
  assign n25343 = n13296 & ~n25342 ;
  assign n25344 = ~n2928 & n21744 ;
  assign n25345 = n13603 ^ n5293 ^ 1'b0 ;
  assign n25346 = n25345 ^ n18496 ^ 1'b0 ;
  assign n25347 = n25344 | n25346 ;
  assign n25348 = n9051 ^ n5712 ^ n2752 ;
  assign n25349 = n25348 ^ n21613 ^ 1'b0 ;
  assign n25350 = n8755 & n13561 ;
  assign n25351 = n15904 | n25350 ;
  assign n25352 = n6976 & ~n25351 ;
  assign n25353 = n25352 ^ n7325 ^ 1'b0 ;
  assign n25354 = ~n4333 & n24114 ;
  assign n25355 = n25354 ^ n20647 ^ 1'b0 ;
  assign n25356 = ~n14301 & n17579 ;
  assign n25357 = ~x40 & n25356 ;
  assign n25358 = n25357 ^ n4972 ^ 1'b0 ;
  assign n25359 = n1512 & n12184 ;
  assign n25360 = n1782 | n7903 ;
  assign n25361 = n2650 & n25360 ;
  assign n25362 = n10192 & ~n21127 ;
  assign n25363 = ( x100 & n2427 ) | ( x100 & ~n7381 ) | ( n2427 & ~n7381 ) ;
  assign n25364 = n12193 & n14300 ;
  assign n25365 = n25364 ^ n13932 ^ 1'b0 ;
  assign n25366 = n461 & ~n25365 ;
  assign n25367 = ~n25363 & n25366 ;
  assign n25368 = n6440 & ~n8402 ;
  assign n25369 = n25367 & n25368 ;
  assign n25372 = n8928 ^ n6114 ^ 1'b0 ;
  assign n25373 = n3589 & n25372 ;
  assign n25370 = n4560 ^ n4328 ^ 1'b0 ;
  assign n25371 = n6999 & ~n25370 ;
  assign n25374 = n25373 ^ n25371 ^ 1'b0 ;
  assign n25375 = n12327 & ~n24507 ;
  assign n25376 = n17150 ^ n9212 ^ 1'b0 ;
  assign n25377 = n6062 ^ n3212 ^ 1'b0 ;
  assign n25378 = n4555 & n20692 ;
  assign n25379 = n25378 ^ n24366 ^ 1'b0 ;
  assign n25380 = n2237 & n12726 ;
  assign n25381 = ~n6542 & n25380 ;
  assign n25382 = n16236 & ~n25381 ;
  assign n25383 = n2664 ^ n1316 ^ 1'b0 ;
  assign n25384 = ~n1082 & n7557 ;
  assign n25385 = n25384 ^ n10488 ^ 1'b0 ;
  assign n25386 = n23234 & ~n25385 ;
  assign n25387 = ~n3128 & n11733 ;
  assign n25388 = n5861 ^ x93 ^ 1'b0 ;
  assign n25389 = n12816 | n25388 ;
  assign n25390 = n25389 ^ n6399 ^ 1'b0 ;
  assign n25391 = n15436 & ~n25390 ;
  assign n25392 = n11709 ^ n2589 ^ 1'b0 ;
  assign n25393 = n681 | n25392 ;
  assign n25394 = n14782 | n25393 ;
  assign n25395 = n25394 ^ n325 ^ 1'b0 ;
  assign n25396 = n25395 ^ n10273 ^ 1'b0 ;
  assign n25397 = ~n23420 & n25396 ;
  assign n25398 = ~n7666 & n12754 ;
  assign n25399 = n12024 & n20336 ;
  assign n25400 = n18212 & n25399 ;
  assign n25402 = n3103 ^ n2106 ^ x164 ;
  assign n25401 = n9320 ^ n4097 ^ 1'b0 ;
  assign n25403 = n25402 ^ n25401 ^ n18437 ;
  assign n25404 = n4862 | n5961 ;
  assign n25405 = n25404 ^ n21274 ^ 1'b0 ;
  assign n25406 = n12505 & ~n25405 ;
  assign n25407 = n552 & n821 ;
  assign n25408 = n1867 | n23697 ;
  assign n25409 = n25408 ^ n24792 ^ 1'b0 ;
  assign n25410 = n25407 & n25409 ;
  assign n25411 = n18779 ^ n782 ^ 1'b0 ;
  assign n25412 = n20001 ^ n15907 ^ 1'b0 ;
  assign n25416 = n16400 | n24653 ;
  assign n25417 = n25416 ^ n4555 ^ 1'b0 ;
  assign n25413 = n13441 ^ n4555 ^ 1'b0 ;
  assign n25414 = ~n19998 & n25413 ;
  assign n25415 = n25414 ^ n11371 ^ 1'b0 ;
  assign n25418 = n25417 ^ n25415 ^ 1'b0 ;
  assign n25419 = n8137 & n11814 ;
  assign n25420 = n12754 | n14492 ;
  assign n25421 = ~n1657 & n25420 ;
  assign n25422 = ~n4117 & n8365 ;
  assign n25423 = n10519 | n15622 ;
  assign n25424 = ~n4991 & n24360 ;
  assign n25425 = n3117 | n9371 ;
  assign n25426 = n313 & ~n25425 ;
  assign n25427 = n25426 ^ n9166 ^ 1'b0 ;
  assign n25428 = n16684 ^ n305 ^ 1'b0 ;
  assign n25429 = n25428 ^ n25197 ^ 1'b0 ;
  assign n25430 = n7706 & n25429 ;
  assign n25431 = n552 & n23274 ;
  assign n25436 = n10213 ^ n3620 ^ n978 ;
  assign n25432 = ~n1372 & n2667 ;
  assign n25433 = n13603 & n25432 ;
  assign n25434 = n16024 ^ n4590 ^ 1'b0 ;
  assign n25435 = n25433 | n25434 ;
  assign n25437 = n25436 ^ n25435 ^ 1'b0 ;
  assign n25438 = n17080 ^ n3057 ^ 1'b0 ;
  assign n25439 = n25437 & ~n25438 ;
  assign n25440 = n14668 ^ n2085 ^ 1'b0 ;
  assign n25441 = n25440 ^ n13763 ^ 1'b0 ;
  assign n25442 = ~n5116 & n7011 ;
  assign n25443 = ~n6574 & n9950 ;
  assign n25444 = n7011 ^ n747 ^ 1'b0 ;
  assign n25445 = n16007 & ~n25444 ;
  assign n25446 = n25445 ^ n2618 ^ 1'b0 ;
  assign n25447 = ~n25443 & n25446 ;
  assign n25448 = x251 & n5903 ;
  assign n25449 = n17251 ^ n7281 ^ n7174 ;
  assign n25450 = ~n5783 & n20664 ;
  assign n25451 = n25450 ^ n5765 ^ 1'b0 ;
  assign n25452 = n1969 | n5963 ;
  assign n25453 = n25452 ^ n1356 ^ 1'b0 ;
  assign n25454 = n4179 & n17897 ;
  assign n25455 = n1981 & ~n2348 ;
  assign n25456 = n25455 ^ n337 ^ 1'b0 ;
  assign n25457 = n1457 & n8901 ;
  assign n25458 = n25456 & n25457 ;
  assign n25459 = n25458 ^ n13627 ^ n4857 ;
  assign n25460 = n11570 ^ x81 ^ 1'b0 ;
  assign n25461 = n8750 & ~n25460 ;
  assign n25462 = n4080 | n7148 ;
  assign n25463 = n15745 ^ n5686 ^ 1'b0 ;
  assign n25464 = n3252 | n4753 ;
  assign n25465 = n21964 & n25464 ;
  assign n25466 = ~n23631 & n25465 ;
  assign n25467 = n9802 & ~n22813 ;
  assign n25468 = ~n8681 & n25467 ;
  assign n25469 = n25468 ^ n8517 ^ 1'b0 ;
  assign n25470 = ~n22092 & n23850 ;
  assign n25478 = n820 & n1757 ;
  assign n25479 = ~n1757 & n25478 ;
  assign n25480 = n6885 & n25479 ;
  assign n25481 = ~n6341 & n25480 ;
  assign n25482 = ~n2667 & n25481 ;
  assign n25483 = n2746 & ~n13588 ;
  assign n25484 = n13588 & n25483 ;
  assign n25485 = ~n1511 & n3690 ;
  assign n25486 = ~n3690 & n25485 ;
  assign n25487 = n25484 | n25486 ;
  assign n25488 = n25482 & ~n25487 ;
  assign n25489 = n3841 & n4084 ;
  assign n25490 = ~n25488 & n25489 ;
  assign n25491 = n25488 & n25490 ;
  assign n25471 = n5748 ^ n2728 ^ 1'b0 ;
  assign n25472 = n2990 & n3863 ;
  assign n25473 = ~n3863 & n25472 ;
  assign n25474 = n2433 & n25473 ;
  assign n25475 = ~n25471 & n25474 ;
  assign n25476 = n17038 & n25475 ;
  assign n25477 = n13323 | n25476 ;
  assign n25492 = n25491 ^ n25477 ^ 1'b0 ;
  assign n25493 = n13133 ^ n3020 ^ 1'b0 ;
  assign n25494 = n16799 & ~n25493 ;
  assign n25495 = n5990 & ~n12506 ;
  assign n25496 = n10306 & n25495 ;
  assign n25497 = n7876 & ~n14344 ;
  assign n25498 = n25497 ^ x231 ^ 1'b0 ;
  assign n25499 = n25498 ^ n12612 ^ 1'b0 ;
  assign n25500 = n8051 & n25499 ;
  assign n25501 = n3089 | n19591 ;
  assign n25502 = n3089 & ~n25501 ;
  assign n25503 = ~n1660 & n5119 ;
  assign n25504 = n25502 & n25503 ;
  assign n25505 = n15686 ^ n10128 ^ 1'b0 ;
  assign n25506 = n3817 & ~n25505 ;
  assign n25507 = n23802 & n25506 ;
  assign n25508 = ( n2761 & n10787 ) | ( n2761 & n24635 ) | ( n10787 & n24635 ) ;
  assign n25509 = ~n2232 & n13761 ;
  assign n25510 = n25508 & n25509 ;
  assign n25511 = n1252 & ~n20582 ;
  assign n25512 = ~x88 & n25511 ;
  assign n25513 = n25512 ^ n6296 ^ 1'b0 ;
  assign n25514 = n10993 & n25513 ;
  assign n25515 = n10601 ^ n5627 ^ 1'b0 ;
  assign n25516 = n17910 & ~n25515 ;
  assign n25517 = n25516 ^ n8760 ^ 1'b0 ;
  assign n25518 = n13913 ^ n5021 ^ n1111 ;
  assign n25519 = ~n801 & n2521 ;
  assign n25520 = n10790 & n25519 ;
  assign n25521 = n25520 ^ n10100 ^ 1'b0 ;
  assign n25522 = n25518 | n25521 ;
  assign n25523 = n24557 | n25522 ;
  assign n25524 = n1805 & ~n25523 ;
  assign n25525 = n15703 ^ n12273 ^ 1'b0 ;
  assign n25526 = n1535 ^ n1314 ^ 1'b0 ;
  assign n25527 = n1429 & n20905 ;
  assign n25528 = n25527 ^ n9389 ^ 1'b0 ;
  assign n25529 = n25528 ^ n2379 ^ 1'b0 ;
  assign n25530 = n6851 | n25529 ;
  assign n25531 = n5159 & ~n11820 ;
  assign n25532 = n19774 ^ n3879 ^ 1'b0 ;
  assign n25533 = n25531 & ~n25532 ;
  assign n25534 = n4841 & ~n10441 ;
  assign n25535 = n25534 ^ n5439 ^ 1'b0 ;
  assign n25536 = n2328 & n2466 ;
  assign n25537 = n9652 | n23473 ;
  assign n25538 = x93 & ~n2581 ;
  assign n25539 = ~n1718 & n25538 ;
  assign n25540 = n25539 ^ n1148 ^ 1'b0 ;
  assign n25541 = n14882 | n25540 ;
  assign n25542 = n2465 & n3855 ;
  assign n25543 = n25542 ^ n19439 ^ 1'b0 ;
  assign n25544 = n504 | n5100 ;
  assign n25545 = n1184 & ~n25544 ;
  assign n25546 = ~n25543 & n25545 ;
  assign n25547 = n19589 | n19911 ;
  assign n25548 = n25547 ^ n458 ^ 1'b0 ;
  assign n25549 = ~n2761 & n3093 ;
  assign n25550 = n25549 ^ n2201 ^ 1'b0 ;
  assign n25551 = x218 & ~n25550 ;
  assign n25552 = n25551 ^ n22601 ^ 1'b0 ;
  assign n25553 = n23390 & ~n25552 ;
  assign n25554 = n10012 | n19104 ;
  assign n25555 = n5099 ^ n2315 ^ 1'b0 ;
  assign n25556 = n11720 ^ n445 ^ 1'b0 ;
  assign n25557 = n25556 ^ n13084 ^ 1'b0 ;
  assign n25558 = x116 & ~n25557 ;
  assign n25559 = n16508 ^ n11591 ^ n6407 ;
  assign n25560 = ~n4821 & n25559 ;
  assign n25561 = n2611 | n22094 ;
  assign n25562 = n10643 & n17874 ;
  assign n25563 = n2122 & n8036 ;
  assign n25564 = n15191 & ~n25563 ;
  assign n25565 = n8995 ^ n6578 ^ 1'b0 ;
  assign n25566 = ~n25564 & n25565 ;
  assign n25567 = n19054 ^ n6089 ^ n2761 ;
  assign n25568 = x129 & ~n7664 ;
  assign n25569 = ~n2949 & n8570 ;
  assign n25570 = ~n13369 & n25569 ;
  assign n25571 = n25570 ^ n14187 ^ 1'b0 ;
  assign n25572 = n19222 ^ n1184 ^ 1'b0 ;
  assign n25573 = n3145 ^ n836 ^ 1'b0 ;
  assign n25574 = ~n7109 & n25573 ;
  assign n25575 = n11710 & ~n17410 ;
  assign n25576 = n1181 & ~n2861 ;
  assign n25577 = n895 & ~n3624 ;
  assign n25578 = n1777 & n25577 ;
  assign n25579 = n25576 & n25578 ;
  assign n25580 = n23758 & n25579 ;
  assign n25581 = n25580 ^ n14381 ^ 1'b0 ;
  assign n25582 = ~n1690 & n6564 ;
  assign n25583 = n9356 ^ n966 ^ 1'b0 ;
  assign n25584 = n1661 & n25583 ;
  assign n25585 = ~n397 & n25584 ;
  assign n25586 = n2342 & n12601 ;
  assign n25587 = n2221 & ~n25586 ;
  assign n25588 = n25585 & n25587 ;
  assign n25589 = n1125 | n17698 ;
  assign n25590 = n25589 ^ n6311 ^ 1'b0 ;
  assign n25591 = n25590 ^ n12767 ^ 1'b0 ;
  assign n25592 = n9078 | n16224 ;
  assign n25593 = n16697 | n25592 ;
  assign n25594 = n305 & n25593 ;
  assign n25595 = n9702 & n25594 ;
  assign n25596 = n13301 | n18619 ;
  assign n25597 = ~n18074 & n25564 ;
  assign n25598 = n25597 ^ n14826 ^ 1'b0 ;
  assign n25599 = n3549 | n25598 ;
  assign n25600 = n3420 | n21957 ;
  assign n25601 = n9803 | n25600 ;
  assign n25602 = n14563 ^ n5043 ^ 1'b0 ;
  assign n25603 = n25601 & n25602 ;
  assign n25604 = n19068 ^ n11862 ^ 1'b0 ;
  assign n25605 = n25604 ^ n17053 ^ 1'b0 ;
  assign n25606 = n6225 & ~n25605 ;
  assign n25607 = x155 & n4310 ;
  assign n25608 = n25607 ^ n1790 ^ 1'b0 ;
  assign n25609 = n20345 ^ n10880 ^ 1'b0 ;
  assign n25610 = n25608 & ~n25609 ;
  assign n25611 = n15773 & n20437 ;
  assign n25612 = ~n20437 & n25611 ;
  assign n25613 = n7802 & ~n12427 ;
  assign n25614 = n8708 & n25613 ;
  assign n25615 = n23813 ^ n6360 ^ 1'b0 ;
  assign n25616 = n641 & n12182 ;
  assign n25617 = n22158 ^ n1608 ^ 1'b0 ;
  assign n25618 = ~n1709 & n10857 ;
  assign n25619 = n25618 ^ n1713 ^ 1'b0 ;
  assign n25620 = n15286 & ~n23885 ;
  assign n25621 = n4014 & ~n25620 ;
  assign n25622 = ~n11376 & n25621 ;
  assign n25623 = n2336 | n16396 ;
  assign n25624 = n25623 ^ n21522 ^ 1'b0 ;
  assign n25625 = n7940 & n25624 ;
  assign n25626 = n23991 ^ n13388 ^ 1'b0 ;
  assign n25627 = n19464 & ~n25626 ;
  assign n25628 = n25397 ^ n15904 ^ 1'b0 ;
  assign n25630 = n946 & ~n2411 ;
  assign n25631 = n25630 ^ n17335 ^ n8127 ;
  assign n25629 = n13836 & ~n18678 ;
  assign n25632 = n25631 ^ n25629 ^ n11458 ;
  assign n25633 = ~n25628 & n25632 ;
  assign n25634 = n559 & n1857 ;
  assign n25635 = n2048 & n14198 ;
  assign n25636 = n25635 ^ n6463 ^ 1'b0 ;
  assign n25637 = n1190 & n19718 ;
  assign n25638 = n9013 & n25637 ;
  assign n25639 = n15504 & n25638 ;
  assign n25640 = ~n3357 & n7879 ;
  assign n25641 = n516 | n2348 ;
  assign n25642 = n25640 & ~n25641 ;
  assign n25643 = n5774 ^ n4156 ^ 1'b0 ;
  assign n25644 = n20229 ^ n7627 ^ 1'b0 ;
  assign n25645 = ~n2546 & n25644 ;
  assign n25646 = n16329 ^ n11082 ^ 1'b0 ;
  assign n25647 = n2351 & n14707 ;
  assign n25648 = n10701 ^ n8135 ^ 1'b0 ;
  assign n25649 = ~n25647 & n25648 ;
  assign n25650 = n25649 ^ n1499 ^ 1'b0 ;
  assign n25651 = n7968 ^ n3485 ^ 1'b0 ;
  assign n25652 = n2409 ^ n1658 ^ 1'b0 ;
  assign n25653 = n8654 | n25652 ;
  assign n25654 = n19939 ^ n10153 ^ 1'b0 ;
  assign n25655 = ~n25653 & n25654 ;
  assign n25656 = n10177 ^ n454 ^ 1'b0 ;
  assign n25657 = n25655 & ~n25656 ;
  assign n25658 = n8997 ^ n4347 ^ 1'b0 ;
  assign n25659 = n12242 & n25658 ;
  assign n25660 = n15937 & n25659 ;
  assign n25661 = n663 & n25660 ;
  assign n25662 = ~n5339 & n16981 ;
  assign n25663 = n13043 & n25662 ;
  assign n25664 = n1054 ^ n917 ^ 1'b0 ;
  assign n25665 = n2205 | n10456 ;
  assign n25666 = n8223 ^ n3453 ^ 1'b0 ;
  assign n25667 = ~n3868 & n25666 ;
  assign n25668 = ( ~n13283 & n25665 ) | ( ~n13283 & n25667 ) | ( n25665 & n25667 ) ;
  assign n25669 = n25664 | n25668 ;
  assign n25670 = n10167 ^ n1339 ^ 1'b0 ;
  assign n25671 = ( n5144 & ~n25614 ) | ( n5144 & n25670 ) | ( ~n25614 & n25670 ) ;
  assign n25672 = n24947 ^ n3186 ^ 1'b0 ;
  assign n25673 = n11443 & n19467 ;
  assign n25674 = n25673 ^ n17629 ^ 1'b0 ;
  assign n25675 = n4134 | n25674 ;
  assign n25676 = n4460 | n17549 ;
  assign n25677 = n13776 | n25676 ;
  assign n25678 = n18137 ^ n9876 ^ 1'b0 ;
  assign n25679 = n10393 & n25678 ;
  assign n25680 = ~n7993 & n16439 ;
  assign n25681 = ~n25679 & n25680 ;
  assign n25684 = n2571 | n16426 ;
  assign n25685 = n25684 ^ n2993 ^ 1'b0 ;
  assign n25682 = n2885 & ~n8530 ;
  assign n25683 = n1081 & ~n25682 ;
  assign n25686 = n25685 ^ n25683 ^ 1'b0 ;
  assign n25687 = n8500 ^ n1723 ^ 1'b0 ;
  assign n25688 = n6184 & n25687 ;
  assign n25689 = n956 | n17765 ;
  assign n25690 = ~n1046 & n25689 ;
  assign n25691 = n3868 & n12926 ;
  assign n25692 = ~n1650 & n13372 ;
  assign n25693 = ~n4272 & n25692 ;
  assign n25694 = n8709 ^ n6452 ^ 1'b0 ;
  assign n25695 = ~x15 & n25694 ;
  assign n25696 = n23653 ^ n11851 ^ 1'b0 ;
  assign n25701 = n13171 | n18900 ;
  assign n25702 = n1646 & ~n25701 ;
  assign n25697 = n8589 | n8730 ;
  assign n25698 = n25697 ^ n9594 ^ 1'b0 ;
  assign n25699 = n25698 ^ n6542 ^ n3578 ;
  assign n25700 = n6931 & ~n25699 ;
  assign n25703 = n25702 ^ n25700 ^ 1'b0 ;
  assign n25704 = n2447 & n8374 ;
  assign n25705 = n4496 & n25704 ;
  assign n25706 = n1658 ^ n566 ^ 1'b0 ;
  assign n25707 = ~n3903 & n13431 ;
  assign n25708 = ~n11149 & n25707 ;
  assign n25709 = n25708 ^ n13886 ^ 1'b0 ;
  assign n25710 = n24050 & ~n25709 ;
  assign n25711 = n25710 ^ n22481 ^ 1'b0 ;
  assign n25712 = n872 & ~n25711 ;
  assign n25713 = n6338 & ~n11128 ;
  assign n25714 = n956 & n24459 ;
  assign n25723 = n9981 & n13909 ;
  assign n25724 = n25723 ^ n2021 ^ 1'b0 ;
  assign n25715 = n3264 | n20197 ;
  assign n25716 = n3264 & ~n25715 ;
  assign n25717 = n5287 & ~n25716 ;
  assign n25718 = ~n5287 & n25717 ;
  assign n25719 = n9137 & ~n25718 ;
  assign n25720 = n25719 ^ n5864 ^ n4972 ;
  assign n25721 = n25720 ^ n10573 ^ n6889 ;
  assign n25722 = n8503 | n25721 ;
  assign n25725 = n25724 ^ n25722 ^ 1'b0 ;
  assign n25726 = n2848 ^ n1503 ^ 1'b0 ;
  assign n25727 = n9119 | n25726 ;
  assign n25728 = n18029 ^ n1436 ^ 1'b0 ;
  assign n25729 = ~n6958 & n13708 ;
  assign n25730 = n25729 ^ n6627 ^ 1'b0 ;
  assign n25731 = n24320 & ~n25730 ;
  assign n25732 = n18464 & n25731 ;
  assign n25733 = n7290 & ~n13428 ;
  assign n25734 = n3274 | n11655 ;
  assign n25735 = n23751 | n25734 ;
  assign n25736 = ~n17344 & n20819 ;
  assign n25737 = n1928 & n8508 ;
  assign n25738 = n4709 & n25737 ;
  assign n25739 = n3687 & ~n17826 ;
  assign n25740 = n25738 & n25739 ;
  assign n25741 = ( ~n13073 & n16576 ) | ( ~n13073 & n25740 ) | ( n16576 & n25740 ) ;
  assign n25742 = n13241 ^ n8543 ^ 1'b0 ;
  assign n25743 = ( n1587 & n1637 ) | ( n1587 & ~n7359 ) | ( n1637 & ~n7359 ) ;
  assign n25744 = n25742 & ~n25743 ;
  assign n25745 = n3505 & ~n5600 ;
  assign n25746 = ~n6541 & n22975 ;
  assign n25747 = n16152 & ~n18362 ;
  assign n25748 = n384 | n4586 ;
  assign n25749 = n25748 ^ n21203 ^ n17311 ;
  assign n25750 = n8559 & n25519 ;
  assign n25751 = n23702 ^ n5896 ^ 1'b0 ;
  assign n25752 = n966 & n8049 ;
  assign n25753 = n25752 ^ n1549 ^ 1'b0 ;
  assign n25754 = n12070 ^ n9331 ^ n4314 ;
  assign n25755 = ~n923 & n23761 ;
  assign n25757 = n14122 & n17378 ;
  assign n25756 = ~n4695 & n16552 ;
  assign n25758 = n25757 ^ n25756 ^ 1'b0 ;
  assign n25759 = ~n9911 & n11848 ;
  assign n25760 = n10401 & ~n25759 ;
  assign n25761 = ~n14675 & n25760 ;
  assign n25762 = n22800 ^ n12500 ^ 1'b0 ;
  assign n25763 = n809 & n25762 ;
  assign n25764 = n6745 ^ n2486 ^ 1'b0 ;
  assign n25765 = n5672 & n25764 ;
  assign n25766 = n1410 | n12820 ;
  assign n25767 = n25209 & ~n25766 ;
  assign n25768 = n25767 ^ n12310 ^ 1'b0 ;
  assign n25769 = n25768 ^ n21739 ^ 1'b0 ;
  assign n25770 = n2550 ^ n519 ^ 1'b0 ;
  assign n25771 = n15744 & ~n25770 ;
  assign n25772 = n813 & ~n2385 ;
  assign n25773 = n5067 & ~n7367 ;
  assign n25774 = ~n13543 & n25773 ;
  assign n25775 = n4118 | n25774 ;
  assign n25776 = n25775 ^ n4689 ^ 1'b0 ;
  assign n25777 = n25776 ^ n25583 ^ n16079 ;
  assign n25778 = n25772 & ~n25777 ;
  assign n25779 = ~n10567 & n25778 ;
  assign n25780 = ~n18061 & n18679 ;
  assign n25781 = n25780 ^ n11454 ^ 1'b0 ;
  assign n25782 = n345 & n1361 ;
  assign n25783 = ~n10869 & n25782 ;
  assign n25784 = n25783 ^ n12249 ^ 1'b0 ;
  assign n25785 = n12725 | n25784 ;
  assign n25786 = n6403 & ~n25785 ;
  assign n25787 = n25786 ^ x105 ^ 1'b0 ;
  assign n25788 = n5275 & ~n8444 ;
  assign n25789 = ~n16452 & n25788 ;
  assign n25790 = n17443 | n17516 ;
  assign n25791 = n25790 ^ n16848 ^ 1'b0 ;
  assign n25792 = n18862 ^ n11226 ^ 1'b0 ;
  assign n25793 = n10164 | n12128 ;
  assign n25794 = ~n21340 & n25793 ;
  assign n25795 = n3731 & n9438 ;
  assign n25796 = n7671 ^ n1589 ^ 1'b0 ;
  assign n25797 = n24495 ^ n5418 ^ 1'b0 ;
  assign n25798 = n25797 ^ n24928 ^ 1'b0 ;
  assign n25799 = ~n8771 & n21361 ;
  assign n25800 = n25798 & n25799 ;
  assign n25801 = n8360 ^ n5610 ^ 1'b0 ;
  assign n25802 = ~n456 & n25801 ;
  assign n25803 = ~n2135 & n19235 ;
  assign n25804 = ~n25802 & n25803 ;
  assign n25805 = n1515 & ~n19098 ;
  assign n25806 = n6574 | n17695 ;
  assign n25807 = n25805 & ~n25806 ;
  assign n25808 = n22481 ^ n20621 ^ n5809 ;
  assign n25809 = n12956 & n25808 ;
  assign n25810 = n25586 ^ n2215 ^ 1'b0 ;
  assign n25811 = n2024 & ~n7227 ;
  assign n25812 = n3292 | n25811 ;
  assign n25813 = n12904 & ~n25812 ;
  assign n25814 = n1347 & n7867 ;
  assign n25815 = ~n8324 & n25814 ;
  assign n25816 = ~n14613 & n17182 ;
  assign n25817 = ( x200 & ~n11005 ) | ( x200 & n17685 ) | ( ~n11005 & n17685 ) ;
  assign n25818 = n4909 & ~n7057 ;
  assign n25819 = n25817 | n25818 ;
  assign n25820 = ~n8941 & n13022 ;
  assign n25821 = n3906 & n25820 ;
  assign n25822 = n20454 ^ n19639 ^ 1'b0 ;
  assign n25823 = ~n25821 & n25822 ;
  assign n25824 = ~n1234 & n4618 ;
  assign n25825 = ~n11851 & n21586 ;
  assign n25826 = n13475 & ~n22318 ;
  assign n25827 = ~n1901 & n17825 ;
  assign n25828 = n25363 ^ n4570 ^ 1'b0 ;
  assign n25829 = ~n14091 & n25828 ;
  assign n25830 = n9547 ^ n9035 ^ 1'b0 ;
  assign n25831 = n5316 & n25830 ;
  assign n25832 = n1517 | n8425 ;
  assign n25833 = n488 & ~n22674 ;
  assign n25834 = n4438 | n4828 ;
  assign n25835 = n1451 & ~n25834 ;
  assign n25836 = n4787 & ~n25835 ;
  assign n25837 = n15829 & n25836 ;
  assign n25838 = ( ~n18846 & n24971 ) | ( ~n18846 & n25345 ) | ( n24971 & n25345 ) ;
  assign n25839 = n12248 ^ n3387 ^ 1'b0 ;
  assign n25840 = n4630 & n14379 ;
  assign n25841 = ~n4630 & n25840 ;
  assign n25842 = n8403 | n25841 ;
  assign n25843 = x108 & n566 ;
  assign n25844 = ~x108 & n25843 ;
  assign n25845 = n4682 | n25844 ;
  assign n25846 = n1485 & ~n25845 ;
  assign n25847 = n25842 & n25846 ;
  assign n25848 = n25847 ^ n11392 ^ 1'b0 ;
  assign n25849 = ~n22676 & n25848 ;
  assign n25850 = n3501 & n5385 ;
  assign n25851 = n25850 ^ n17928 ^ 1'b0 ;
  assign n25855 = n3578 & n5801 ;
  assign n25856 = n1725 | n25855 ;
  assign n25857 = ~n1299 & n14265 ;
  assign n25858 = n15743 | n25857 ;
  assign n25859 = ~n2333 & n25858 ;
  assign n25860 = n25859 ^ n21200 ^ 1'b0 ;
  assign n25861 = n25860 ^ n7585 ^ 1'b0 ;
  assign n25862 = n25856 & ~n25861 ;
  assign n25852 = n7515 ^ n2248 ^ 1'b0 ;
  assign n25853 = n15952 & ~n25852 ;
  assign n25854 = ~n618 & n25853 ;
  assign n25863 = n25862 ^ n25854 ^ 1'b0 ;
  assign n25864 = n23125 ^ n939 ^ 1'b0 ;
  assign n25865 = n9183 | n25864 ;
  assign n25866 = n5851 | n23399 ;
  assign n25867 = n15757 ^ n6243 ^ 1'b0 ;
  assign n25871 = n1048 & n3559 ;
  assign n25872 = n25871 ^ n12527 ^ 1'b0 ;
  assign n25868 = n22063 ^ n18644 ^ 1'b0 ;
  assign n25869 = n1841 & ~n25868 ;
  assign n25870 = n3181 & n25869 ;
  assign n25873 = n25872 ^ n25870 ^ 1'b0 ;
  assign n25874 = n3292 & ~n7938 ;
  assign n25875 = n7323 | n25874 ;
  assign n25876 = n1727 ^ n292 ^ 1'b0 ;
  assign n25877 = n22803 ^ n6165 ^ 1'b0 ;
  assign n25878 = n19256 & ~n20156 ;
  assign n25879 = n25878 ^ n13912 ^ 1'b0 ;
  assign n25880 = n24409 ^ x33 ^ 1'b0 ;
  assign n25881 = n25880 ^ n5955 ^ 1'b0 ;
  assign n25882 = n17810 & n23776 ;
  assign n25883 = n5861 & n25882 ;
  assign n25884 = n1776 | n9050 ;
  assign n25885 = n25884 ^ n4291 ^ 1'b0 ;
  assign n25886 = n2463 & ~n25885 ;
  assign n25887 = n25886 ^ n17982 ^ 1'b0 ;
  assign n25888 = ~n5478 & n25887 ;
  assign n25889 = n25888 ^ n1657 ^ 1'b0 ;
  assign n25890 = ~n5445 & n25889 ;
  assign n25891 = ~n10061 & n25188 ;
  assign n25892 = n13214 & ~n20988 ;
  assign n25893 = n25892 ^ n269 ^ 1'b0 ;
  assign n25894 = n897 & n10401 ;
  assign n25895 = n25894 ^ n876 ^ 1'b0 ;
  assign n25896 = n25895 ^ n8492 ^ 1'b0 ;
  assign n25898 = n6999 ^ n2886 ^ n1683 ;
  assign n25897 = n17140 & n17560 ;
  assign n25899 = n25898 ^ n25897 ^ 1'b0 ;
  assign n25900 = n25896 | n25899 ;
  assign n25901 = n11519 | n25900 ;
  assign n25902 = ~n546 & n17588 ;
  assign n25903 = ~n6199 & n9087 ;
  assign n25904 = n4970 & n25903 ;
  assign n25905 = ~n11007 & n25904 ;
  assign n25906 = ~n631 & n17957 ;
  assign n25907 = n10584 & n25906 ;
  assign n25908 = n25907 ^ n10505 ^ 1'b0 ;
  assign n25909 = n8523 | n25908 ;
  assign n25910 = n16197 ^ n10021 ^ 1'b0 ;
  assign n25911 = ~n956 & n15737 ;
  assign n25912 = n25911 ^ n15146 ^ 1'b0 ;
  assign n25913 = n9163 & ~n10823 ;
  assign n25914 = n16448 & n25913 ;
  assign n25915 = n11486 | n22396 ;
  assign n25916 = n2861 & ~n25915 ;
  assign n25917 = n13802 & n25880 ;
  assign n25918 = n3828 & n25917 ;
  assign n25919 = n2034 ^ n1656 ^ 1'b0 ;
  assign n25920 = n14501 ^ n4178 ^ n3667 ;
  assign n25921 = n25919 & n25920 ;
  assign n25922 = n11536 & ~n21660 ;
  assign n25923 = n18289 ^ n14711 ^ 1'b0 ;
  assign n25924 = n12121 & ~n25923 ;
  assign n25925 = n25924 ^ n17801 ^ n7839 ;
  assign n25926 = n1642 | n3022 ;
  assign n25927 = n25248 ^ n23020 ^ 1'b0 ;
  assign n25928 = n15903 ^ n3229 ^ 1'b0 ;
  assign n25929 = n25927 & n25928 ;
  assign n25930 = ~n1843 & n2677 ;
  assign n25932 = ~n1859 & n3467 ;
  assign n25933 = n25932 ^ n2827 ^ 1'b0 ;
  assign n25934 = n6568 & ~n25933 ;
  assign n25931 = n4905 & ~n10150 ;
  assign n25935 = n25934 ^ n25931 ^ 1'b0 ;
  assign n25936 = n23761 ^ n3789 ^ 1'b0 ;
  assign n25937 = n2482 & n3416 ;
  assign n25938 = n6473 & n25937 ;
  assign n25939 = n4338 & ~n7674 ;
  assign n25940 = n7021 & n25939 ;
  assign n25941 = n17046 & n25940 ;
  assign n25943 = n1594 | n6081 ;
  assign n25944 = n401 & ~n25943 ;
  assign n25945 = n25944 ^ n15841 ^ 1'b0 ;
  assign n25942 = n6015 & ~n8703 ;
  assign n25946 = n25945 ^ n25942 ^ n21172 ;
  assign n25947 = n3548 ^ n2685 ^ 1'b0 ;
  assign n25948 = n3206 & ~n25947 ;
  assign n25949 = n25948 ^ n21443 ^ 1'b0 ;
  assign n25950 = x218 & ~n8770 ;
  assign n25951 = ~n10814 & n24016 ;
  assign n25952 = ~n5625 & n9061 ;
  assign n25953 = n25952 ^ n405 ^ 1'b0 ;
  assign n25954 = n5748 & n15737 ;
  assign n25956 = n11441 ^ x100 ^ 1'b0 ;
  assign n25957 = n25956 ^ n1145 ^ 1'b0 ;
  assign n25955 = n4575 | n18842 ;
  assign n25958 = n25957 ^ n25955 ^ 1'b0 ;
  assign n25959 = n3047 & n5573 ;
  assign n25960 = n25959 ^ n18174 ^ 1'b0 ;
  assign n25961 = ~n3870 & n25960 ;
  assign n25962 = n25961 ^ n7421 ^ 1'b0 ;
  assign n25963 = n1727 & n11894 ;
  assign n25964 = n25963 ^ n4366 ^ 1'b0 ;
  assign n25965 = n7978 & ~n19568 ;
  assign n25966 = n13804 ^ n871 ^ 1'b0 ;
  assign n25967 = n2175 & ~n25966 ;
  assign n25968 = n12203 & n16901 ;
  assign n25969 = n18409 & n19508 ;
  assign n25970 = n8668 ^ n1930 ^ 1'b0 ;
  assign n25971 = ~n20871 & n25970 ;
  assign n25972 = ~n1738 & n18116 ;
  assign n25973 = n6375 & n25972 ;
  assign n25974 = n25973 ^ n25857 ^ 1'b0 ;
  assign n25975 = n1429 & n11815 ;
  assign n25976 = n25975 ^ n2011 ^ 1'b0 ;
  assign n25977 = n1016 & n25976 ;
  assign n25978 = n13863 & n25977 ;
  assign n25979 = n25880 & ~n25978 ;
  assign n25980 = n13455 ^ x115 ^ 1'b0 ;
  assign n25981 = n8411 & n25980 ;
  assign n25982 = n20722 & ~n25981 ;
  assign n25983 = n8503 ^ n2264 ^ 1'b0 ;
  assign n25984 = n13596 & n25983 ;
  assign n25985 = n16580 & ~n17698 ;
  assign n25986 = n7148 & n25985 ;
  assign n25987 = n17811 | n18913 ;
  assign n25988 = n7274 | n17975 ;
  assign n25989 = n25988 ^ n11688 ^ 1'b0 ;
  assign n25990 = n22305 & n25989 ;
  assign n25991 = n22737 ^ n8386 ^ 1'b0 ;
  assign n25992 = n12157 | n17514 ;
  assign n25993 = n25992 ^ n18951 ^ 1'b0 ;
  assign n25994 = ~n7558 & n10781 ;
  assign n25995 = ~n3223 & n24108 ;
  assign n25996 = n4943 | n10785 ;
  assign n25997 = n25996 ^ n25874 ^ 1'b0 ;
  assign n25999 = n18046 ^ n6276 ^ 1'b0 ;
  assign n25998 = n470 | n21727 ;
  assign n26000 = n25999 ^ n25998 ^ 1'b0 ;
  assign n26001 = n577 | n11585 ;
  assign n26002 = x208 & ~n4333 ;
  assign n26003 = ~x54 & n26002 ;
  assign n26004 = n26003 ^ n21611 ^ n4575 ;
  assign n26005 = n26001 | n26004 ;
  assign n26006 = n11259 & ~n15622 ;
  assign n26007 = n1280 | n10229 ;
  assign n26008 = n4668 | n26007 ;
  assign n26009 = ~x50 & n1429 ;
  assign n26010 = x5 & ~n4147 ;
  assign n26011 = n19957 & n26010 ;
  assign n26012 = x95 | n16209 ;
  assign n26013 = n26011 & ~n26012 ;
  assign n26014 = n8415 ^ n1843 ^ 1'b0 ;
  assign n26015 = ~n1514 & n26014 ;
  assign n26016 = n26015 ^ n5956 ^ 1'b0 ;
  assign n26017 = n3786 & n16034 ;
  assign n26018 = ( n6704 & n26016 ) | ( n6704 & n26017 ) | ( n26016 & n26017 ) ;
  assign n26019 = n3150 & ~n18932 ;
  assign n26020 = n12988 | n19854 ;
  assign n26021 = n19542 | n26020 ;
  assign n26022 = ~n6078 & n8449 ;
  assign n26023 = n26021 & ~n26022 ;
  assign n26024 = ( n9828 & n11424 ) | ( n9828 & n21040 ) | ( n11424 & n21040 ) ;
  assign n26025 = n26024 ^ n7970 ^ 1'b0 ;
  assign n26026 = ~n14168 & n15682 ;
  assign n26027 = n9475 & n26026 ;
  assign n26028 = n4460 ^ n710 ^ 1'b0 ;
  assign n26029 = n10398 ^ n5171 ^ 1'b0 ;
  assign n26030 = n9312 & n12959 ;
  assign n26031 = n2693 & n4467 ;
  assign n26032 = n26030 & n26031 ;
  assign n26033 = n2315 ^ x127 ^ 1'b0 ;
  assign n26034 = n17580 & n26033 ;
  assign n26036 = ~n4413 & n10053 ;
  assign n26037 = n9374 | n26036 ;
  assign n26035 = ~n5563 & n8504 ;
  assign n26038 = n26037 ^ n26035 ^ 1'b0 ;
  assign n26039 = ~n4625 & n15318 ;
  assign n26040 = n2584 & n26039 ;
  assign n26041 = n754 | n26040 ;
  assign n26042 = n13821 & ~n26041 ;
  assign n26043 = n26038 & n26042 ;
  assign n26044 = n3498 & n4375 ;
  assign n26045 = n6298 | n14178 ;
  assign n26046 = n26045 ^ n13253 ^ 1'b0 ;
  assign n26047 = n5598 & ~n26046 ;
  assign n26048 = n8014 ^ n1521 ^ 1'b0 ;
  assign n26049 = n26048 ^ n917 ^ 1'b0 ;
  assign n26050 = n9760 ^ n5031 ^ 1'b0 ;
  assign n26051 = n9471 | n26050 ;
  assign n26052 = n26049 & ~n26051 ;
  assign n26053 = n26052 ^ n6162 ^ 1'b0 ;
  assign n26054 = n10756 | n26053 ;
  assign n26055 = n4784 & ~n9545 ;
  assign n26056 = ~n1713 & n26055 ;
  assign n26057 = n5607 | n26056 ;
  assign n26058 = n26057 ^ n2022 ^ 1'b0 ;
  assign n26059 = ~n19854 & n26058 ;
  assign n26060 = n4001 & n5828 ;
  assign n26061 = n26060 ^ n13585 ^ 1'b0 ;
  assign n26062 = ~n8311 & n26061 ;
  assign n26067 = n3314 & ~n3813 ;
  assign n26065 = n5471 ^ n2208 ^ 1'b0 ;
  assign n26066 = n3143 & n26065 ;
  assign n26063 = n10019 | n16346 ;
  assign n26064 = n10276 & ~n26063 ;
  assign n26068 = n26067 ^ n26066 ^ n26064 ;
  assign n26069 = n21598 | n26068 ;
  assign n26070 = n10782 ^ n9460 ^ 1'b0 ;
  assign n26071 = n7000 & n8902 ;
  assign n26072 = n26071 ^ n14241 ^ 1'b0 ;
  assign n26073 = n19439 & ~n24936 ;
  assign n26074 = n26072 | n26073 ;
  assign n26075 = n3473 & n25262 ;
  assign n26076 = n7888 & ~n20862 ;
  assign n26077 = ~n1488 & n10222 ;
  assign n26078 = n8027 ^ n3678 ^ 1'b0 ;
  assign n26079 = x246 & ~n26078 ;
  assign n26080 = n26079 ^ n4261 ^ n3754 ;
  assign n26081 = n1861 | n4532 ;
  assign n26084 = n6903 & ~n8428 ;
  assign n26082 = ~n8806 & n11370 ;
  assign n26083 = n26082 ^ n17126 ^ 1'b0 ;
  assign n26085 = n26084 ^ n26083 ^ 1'b0 ;
  assign n26086 = n10440 & ~n26085 ;
  assign n26087 = n26086 ^ n24111 ^ 1'b0 ;
  assign n26088 = n26081 & n26087 ;
  assign n26089 = n12633 ^ n5023 ^ 1'b0 ;
  assign n26090 = n7321 ^ n415 ^ 1'b0 ;
  assign n26091 = n26090 ^ n1354 ^ 1'b0 ;
  assign n26092 = n26091 ^ n18812 ^ 1'b0 ;
  assign n26093 = n12015 & ~n26092 ;
  assign n26094 = n26093 ^ n7991 ^ 1'b0 ;
  assign n26095 = n13498 & ~n22760 ;
  assign n26096 = n26095 ^ n19452 ^ 1'b0 ;
  assign n26097 = n21513 ^ n16164 ^ 1'b0 ;
  assign n26098 = n6584 & ~n7903 ;
  assign n26104 = n14388 ^ n2426 ^ 1'b0 ;
  assign n26099 = n1865 | n5136 ;
  assign n26100 = n4673 | n26099 ;
  assign n26101 = n753 | n7548 ;
  assign n26102 = n581 | n26101 ;
  assign n26103 = n26100 & n26102 ;
  assign n26105 = n26104 ^ n26103 ^ 1'b0 ;
  assign n26106 = n2602 | n6813 ;
  assign n26107 = n10564 ^ n7406 ^ 1'b0 ;
  assign n26108 = ~n5125 & n5733 ;
  assign n26111 = n5809 & n8889 ;
  assign n26112 = n26111 ^ n3754 ^ 1'b0 ;
  assign n26109 = n13547 ^ n9634 ^ 1'b0 ;
  assign n26110 = n8191 | n26109 ;
  assign n26113 = n26112 ^ n26110 ^ n2541 ;
  assign n26114 = n21669 ^ n5485 ^ n5279 ;
  assign n26115 = n979 & ~n26114 ;
  assign n26116 = n26115 ^ n9276 ^ 1'b0 ;
  assign n26117 = n11964 ^ n5196 ^ 1'b0 ;
  assign n26118 = ~n7117 & n26117 ;
  assign n26119 = n25037 ^ n3150 ^ 1'b0 ;
  assign n26120 = n23151 ^ n16037 ^ 1'b0 ;
  assign n26121 = ( n7630 & n8713 ) | ( n7630 & n18770 ) | ( n8713 & n18770 ) ;
  assign n26122 = n17755 | n26121 ;
  assign n26123 = n2179 ^ n677 ^ 1'b0 ;
  assign n26124 = ~n713 & n26123 ;
  assign n26125 = ~x84 & n26124 ;
  assign n26126 = n14908 | n26125 ;
  assign n26127 = n26126 ^ n4513 ^ 1'b0 ;
  assign n26128 = n401 & ~n16186 ;
  assign n26130 = n296 & ~n734 ;
  assign n26131 = n734 & n26130 ;
  assign n26129 = n6670 | n7046 ;
  assign n26132 = n26131 ^ n26129 ^ 1'b0 ;
  assign n26133 = n6428 & ~n26132 ;
  assign n26134 = n26132 & n26133 ;
  assign n26135 = ( ~n415 & n17375 ) | ( ~n415 & n26134 ) | ( n17375 & n26134 ) ;
  assign n26136 = n13411 & ~n15907 ;
  assign n26137 = n13723 & n15128 ;
  assign n26138 = n7884 | n11449 ;
  assign n26139 = n26138 ^ n7223 ^ 1'b0 ;
  assign n26140 = n901 | n1077 ;
  assign n26141 = n2283 & ~n11140 ;
  assign n26142 = n26141 ^ n21040 ^ 1'b0 ;
  assign n26143 = n14982 | n26142 ;
  assign n26144 = n26143 ^ n9873 ^ 1'b0 ;
  assign n26145 = n26140 & n26144 ;
  assign n26146 = ~n26139 & n26145 ;
  assign n26147 = n7548 ^ x142 ^ 1'b0 ;
  assign n26148 = n4545 | n26147 ;
  assign n26149 = n610 | n26148 ;
  assign n26150 = ( n1694 & n20657 ) | ( n1694 & n26149 ) | ( n20657 & n26149 ) ;
  assign n26151 = n2103 & n10387 ;
  assign n26152 = n26151 ^ n20491 ^ n9317 ;
  assign n26153 = n20194 ^ n13978 ^ 1'b0 ;
  assign n26154 = n2818 & ~n26153 ;
  assign n26162 = ~n3134 & n5468 ;
  assign n26158 = n3938 & n13129 ;
  assign n26159 = n2393 & n5332 ;
  assign n26160 = n26158 & n26159 ;
  assign n26155 = n5468 | n10663 ;
  assign n26156 = n26155 ^ n263 ^ 1'b0 ;
  assign n26157 = ~n4112 & n26156 ;
  assign n26161 = n26160 ^ n26157 ^ 1'b0 ;
  assign n26163 = n26162 ^ n26161 ^ 1'b0 ;
  assign n26164 = n12667 & n26163 ;
  assign n26165 = n26164 ^ n15933 ^ 1'b0 ;
  assign n26166 = n9723 & n26165 ;
  assign n26167 = n24978 ^ n10403 ^ 1'b0 ;
  assign n26168 = n17453 ^ n6437 ^ 1'b0 ;
  assign n26169 = ~n26167 & n26168 ;
  assign n26170 = ~n13609 & n26169 ;
  assign n26171 = n4367 & n20790 ;
  assign n26172 = n5490 & ~n9166 ;
  assign n26173 = n13051 & n26172 ;
  assign n26174 = n1832 & ~n11228 ;
  assign n26175 = n1758 & ~n26174 ;
  assign n26176 = ~n26173 & n26175 ;
  assign n26177 = n15249 & n18797 ;
  assign n26178 = n3302 & n12846 ;
  assign n26179 = n26178 ^ n2296 ^ 1'b0 ;
  assign n26180 = n16993 ^ n11255 ^ 1'b0 ;
  assign n26181 = n20591 & n26180 ;
  assign n26182 = ~n26179 & n26181 ;
  assign n26183 = ~n8137 & n14400 ;
  assign n26184 = n21519 & n26183 ;
  assign n26185 = n8427 & n13538 ;
  assign n26186 = ~x118 & n1106 ;
  assign n26187 = n26186 ^ n8122 ^ 1'b0 ;
  assign n26188 = ~n4340 & n5067 ;
  assign n26189 = n26187 & n26188 ;
  assign n26190 = n6014 | n24060 ;
  assign n26191 = ( n4487 & n6273 ) | ( n4487 & ~n7243 ) | ( n6273 & ~n7243 ) ;
  assign n26192 = n26191 ^ n11203 ^ 1'b0 ;
  assign n26193 = ~n3181 & n26192 ;
  assign n26194 = n25705 | n26193 ;
  assign n26195 = n4043 | n10955 ;
  assign n26196 = n26195 ^ n4521 ^ 1'b0 ;
  assign n26197 = ( ~n10767 & n14965 ) | ( ~n10767 & n26196 ) | ( n14965 & n26196 ) ;
  assign n26198 = n16978 & ~n26197 ;
  assign n26199 = n14196 ^ n11904 ^ 1'b0 ;
  assign n26200 = n11934 ^ x23 ^ 1'b0 ;
  assign n26201 = ~n3951 & n26200 ;
  assign n26202 = ( ~n2416 & n11107 ) | ( ~n2416 & n26201 ) | ( n11107 & n26201 ) ;
  assign n26203 = n1196 | n5366 ;
  assign n26204 = ~n708 & n26203 ;
  assign n26205 = n26204 ^ n4785 ^ 1'b0 ;
  assign n26206 = ~n1994 & n9584 ;
  assign n26207 = n26206 ^ n5010 ^ 1'b0 ;
  assign n26211 = ~n394 & n3239 ;
  assign n26208 = ~n1753 & n7526 ;
  assign n26209 = n26208 ^ n14248 ^ 1'b0 ;
  assign n26210 = n610 & ~n26209 ;
  assign n26212 = n26211 ^ n26210 ^ 1'b0 ;
  assign n26213 = n26207 & n26212 ;
  assign n26214 = n26213 ^ n26062 ^ 1'b0 ;
  assign n26215 = ~n533 & n26214 ;
  assign n26216 = n4982 & n22430 ;
  assign n26217 = n7126 ^ n2715 ^ 1'b0 ;
  assign n26218 = n26216 & n26217 ;
  assign n26219 = n23195 & n26218 ;
  assign n26220 = n26219 ^ n4071 ^ 1'b0 ;
  assign n26221 = n24041 ^ n2464 ^ 1'b0 ;
  assign n26222 = ~n8647 & n26221 ;
  assign n26223 = n21113 ^ n19742 ^ 1'b0 ;
  assign n26224 = n9333 & n22296 ;
  assign n26225 = ~n18427 & n26224 ;
  assign n26226 = n26225 ^ n5634 ^ 1'b0 ;
  assign n26227 = n19901 ^ n977 ^ 1'b0 ;
  assign n26228 = n16112 | n26227 ;
  assign n26229 = n3995 & ~n5468 ;
  assign n26230 = n7347 & n26229 ;
  assign n26231 = n26228 | n26230 ;
  assign n26232 = n26231 ^ n10856 ^ 1'b0 ;
  assign n26233 = ~n3256 & n7755 ;
  assign n26234 = n17779 | n26233 ;
  assign n26235 = n4811 & ~n26234 ;
  assign n26236 = n26235 ^ n6471 ^ 1'b0 ;
  assign n26237 = n15326 & n26236 ;
  assign n26238 = n648 & n3342 ;
  assign n26239 = ~n8211 & n26238 ;
  assign n26240 = n26239 ^ n18380 ^ 1'b0 ;
  assign n26241 = n18241 ^ n13738 ^ 1'b0 ;
  assign n26242 = n8187 | n26241 ;
  assign n26243 = n17738 ^ n6823 ^ 1'b0 ;
  assign n26244 = n26243 ^ n9341 ^ 1'b0 ;
  assign n26245 = n13664 & n26244 ;
  assign n26246 = n7174 & ~n26245 ;
  assign n26247 = n25135 ^ n8277 ^ 1'b0 ;
  assign n26248 = n10851 | n18695 ;
  assign n26249 = n26248 ^ n8190 ^ 1'b0 ;
  assign n26250 = n26249 ^ n2135 ^ 1'b0 ;
  assign n26251 = n22705 ^ n1793 ^ 1'b0 ;
  assign n26252 = n10108 & n26251 ;
  assign n26253 = n10686 ^ n3255 ^ 1'b0 ;
  assign n26254 = n20292 & ~n26253 ;
  assign n26255 = n26254 ^ n1104 ^ 1'b0 ;
  assign n26256 = n7560 & n19622 ;
  assign n26257 = ~n24233 & n26256 ;
  assign n26259 = n2647 & ~n14198 ;
  assign n26258 = ~n4185 & n11894 ;
  assign n26260 = n26259 ^ n26258 ^ 1'b0 ;
  assign n26261 = n2001 & n14605 ;
  assign n26262 = ~n11264 & n26261 ;
  assign n26263 = n26262 ^ n1926 ^ 1'b0 ;
  assign n26264 = n10817 & n15812 ;
  assign n26265 = n15060 & n26264 ;
  assign n26266 = n26263 & n26265 ;
  assign n26267 = n11078 & ~n21273 ;
  assign n26269 = n4173 ^ n1291 ^ 1'b0 ;
  assign n26268 = ~n2157 & n12841 ;
  assign n26270 = n26269 ^ n26268 ^ 1'b0 ;
  assign n26271 = n10631 & n16598 ;
  assign n26272 = ( n1214 & n5422 ) | ( n1214 & n9707 ) | ( n5422 & n9707 ) ;
  assign n26273 = n8731 & ~n9755 ;
  assign n26274 = ~n4541 & n13379 ;
  assign n26275 = n7133 ^ n4118 ^ 1'b0 ;
  assign n26276 = ~n7622 & n7829 ;
  assign n26277 = n26276 ^ n23538 ^ 1'b0 ;
  assign n26278 = n17948 ^ x100 ^ 1'b0 ;
  assign n26279 = ~n13000 & n19840 ;
  assign n26280 = n11685 & n26279 ;
  assign n26281 = n17907 & n26280 ;
  assign n26282 = n12359 & ~n14241 ;
  assign n26283 = ( ~n4316 & n13116 ) | ( ~n4316 & n26282 ) | ( n13116 & n26282 ) ;
  assign n26284 = ~n11974 & n25418 ;
  assign n26285 = n26284 ^ n15362 ^ 1'b0 ;
  assign n26286 = n6214 ^ n844 ^ 1'b0 ;
  assign n26287 = n13580 & n26286 ;
  assign n26288 = n1477 & ~n8424 ;
  assign n26289 = ~n4524 & n26288 ;
  assign n26290 = ~n840 & n9087 ;
  assign n26292 = n1912 & n3637 ;
  assign n26293 = n366 & n26292 ;
  assign n26291 = n4048 | n5750 ;
  assign n26294 = n26293 ^ n26291 ^ 1'b0 ;
  assign n26295 = x247 & n4316 ;
  assign n26296 = n26295 ^ n17907 ^ 1'b0 ;
  assign n26297 = n1594 | n23035 ;
  assign n26298 = n26297 ^ n9165 ^ 1'b0 ;
  assign n26299 = n10098 ^ n9908 ^ 1'b0 ;
  assign n26300 = x193 | n26299 ;
  assign n26301 = n5592 | n6255 ;
  assign n26302 = n14852 | n26301 ;
  assign n26303 = ~n15529 & n16814 ;
  assign n26304 = n21601 & n26303 ;
  assign n26305 = n26304 ^ n20391 ^ 1'b0 ;
  assign n26306 = n7020 & n8395 ;
  assign n26307 = n26306 ^ n14386 ^ n9223 ;
  assign n26308 = x122 & n343 ;
  assign n26309 = n24374 & n26308 ;
  assign n26310 = n19669 ^ n13391 ^ 1'b0 ;
  assign n26311 = n7496 | n14771 ;
  assign n26312 = n24291 & ~n26311 ;
  assign n26313 = ~n921 & n26312 ;
  assign n26314 = n26313 ^ n14201 ^ 1'b0 ;
  assign n26315 = n22207 ^ n2873 ^ n789 ;
  assign n26316 = n4169 ^ n3659 ^ 1'b0 ;
  assign n26317 = ~n3781 & n26316 ;
  assign n26318 = n5774 & n26317 ;
  assign n26319 = n7998 ^ n2287 ^ 1'b0 ;
  assign n26320 = ~n23065 & n26319 ;
  assign n26321 = ~n4063 & n7762 ;
  assign n26322 = ~n17583 & n26321 ;
  assign n26323 = n886 | n17856 ;
  assign n26324 = n14495 ^ x230 ^ 1'b0 ;
  assign n26325 = n1335 ^ n1252 ^ 1'b0 ;
  assign n26326 = n26325 ^ n4118 ^ 1'b0 ;
  assign n26327 = n26326 ^ n3419 ^ 1'b0 ;
  assign n26328 = n24241 ^ n5193 ^ 1'b0 ;
  assign n26329 = ~n26327 & n26328 ;
  assign n26330 = n8362 | n21042 ;
  assign n26331 = n6110 & n8609 ;
  assign n26332 = n11572 & n26331 ;
  assign n26333 = n8317 | n26332 ;
  assign n26334 = x170 | n15328 ;
  assign n26335 = n22174 ^ n17254 ^ 1'b0 ;
  assign n26336 = ~n17869 & n26207 ;
  assign n26337 = n2185 | n3239 ;
  assign n26338 = n11269 & ~n26337 ;
  assign n26339 = n3181 | n9773 ;
  assign n26340 = n1847 & n9285 ;
  assign n26341 = ~n13155 & n26340 ;
  assign n26342 = n24867 ^ n12051 ^ 1'b0 ;
  assign n26343 = ~n3249 & n16927 ;
  assign n26344 = n21275 & ~n26343 ;
  assign n26345 = n21209 & n26344 ;
  assign n26346 = n5116 & n12616 ;
  assign n26347 = n994 | n26346 ;
  assign n26348 = n2298 | n13585 ;
  assign n26349 = n1886 & ~n8515 ;
  assign n26350 = n21435 | n23256 ;
  assign n26351 = n6413 & ~n26350 ;
  assign n26352 = n8276 | n26351 ;
  assign n26353 = n26352 ^ n827 ^ 1'b0 ;
  assign n26354 = ~n641 & n26353 ;
  assign n26355 = n26354 ^ n21943 ^ 1'b0 ;
  assign n26356 = n2391 | n26355 ;
  assign n26357 = n3582 ^ n2159 ^ 1'b0 ;
  assign n26358 = n22927 | n26357 ;
  assign n26359 = n16552 ^ n6486 ^ 1'b0 ;
  assign n26360 = n4034 & n26359 ;
  assign n26361 = x180 & n1252 ;
  assign n26362 = n3068 | n6473 ;
  assign n26363 = n7431 ^ n5302 ^ 1'b0 ;
  assign n26364 = n3999 & n26363 ;
  assign n26365 = n26364 ^ n7454 ^ 1'b0 ;
  assign n26366 = n9651 & n26365 ;
  assign n26367 = n16330 & n26366 ;
  assign n26368 = ~n26362 & n26367 ;
  assign n26369 = ~n6193 & n9776 ;
  assign n26370 = n10189 & n26369 ;
  assign n26371 = n6100 & ~n26370 ;
  assign n26372 = n26368 | n26371 ;
  assign n26373 = n24472 ^ n20760 ^ n18136 ;
  assign n26374 = ~n4072 & n26373 ;
  assign n26375 = n6756 ^ n5675 ^ 1'b0 ;
  assign n26376 = ~n7098 & n26375 ;
  assign n26377 = ~n7565 & n26376 ;
  assign n26378 = n22635 & n26377 ;
  assign n26379 = n4258 & ~n6109 ;
  assign n26380 = n17056 ^ n2495 ^ 1'b0 ;
  assign n26381 = n19216 | n26380 ;
  assign n26382 = n4237 & n7900 ;
  assign n26383 = x116 & ~n26382 ;
  assign n26384 = n26383 ^ n6857 ^ 1'b0 ;
  assign n26385 = n8849 & ~n26384 ;
  assign n26386 = n3803 & n9386 ;
  assign n26387 = n26386 ^ n23256 ^ 1'b0 ;
  assign n26388 = n26216 ^ n16953 ^ 1'b0 ;
  assign n26389 = n26387 & ~n26388 ;
  assign n26390 = n26385 & n26389 ;
  assign n26391 = n26390 ^ x21 ^ 1'b0 ;
  assign n26392 = n2312 & n13364 ;
  assign n26393 = ~n22401 & n25036 ;
  assign n26394 = n23395 ^ n7448 ^ 1'b0 ;
  assign n26395 = n26394 ^ n11625 ^ 1'b0 ;
  assign n26396 = ~n7829 & n26395 ;
  assign n26397 = ~n26395 & n26396 ;
  assign n26398 = n25578 | n26397 ;
  assign n26399 = n26397 & ~n26398 ;
  assign n26400 = x5 & ~n2431 ;
  assign n26401 = n22846 | n26400 ;
  assign n26402 = n4520 | n7709 ;
  assign n26403 = n16792 & ~n26402 ;
  assign n26404 = ~n1099 & n3239 ;
  assign n26405 = n26404 ^ n10723 ^ 1'b0 ;
  assign n26406 = n26405 ^ n7624 ^ 1'b0 ;
  assign n26407 = ~n1195 & n22249 ;
  assign n26408 = n7500 | n15824 ;
  assign n26409 = n16846 & ~n26408 ;
  assign n26410 = n4539 & n20555 ;
  assign n26411 = n1965 & n19100 ;
  assign n26412 = ~n26410 & n26411 ;
  assign n26413 = n3323 & n26412 ;
  assign n26414 = n18591 & ~n20928 ;
  assign n26415 = n26414 ^ n12673 ^ n10002 ;
  assign n26416 = n26415 ^ n11453 ^ 1'b0 ;
  assign n26417 = n4024 | n9210 ;
  assign n26418 = n26417 ^ n3419 ^ 1'b0 ;
  assign n26419 = n10017 ^ n7554 ^ 1'b0 ;
  assign n26420 = n26419 ^ n22173 ^ 1'b0 ;
  assign n26421 = n17168 & n17285 ;
  assign n26422 = n2399 & ~n4968 ;
  assign n26423 = n26422 ^ n9489 ^ 1'b0 ;
  assign n26424 = n1917 & ~n4631 ;
  assign n26425 = n1879 | n26424 ;
  assign n26426 = n26425 ^ n11587 ^ 1'b0 ;
  assign n26427 = n26426 ^ n904 ^ 1'b0 ;
  assign n26428 = ~n24926 & n26427 ;
  assign n26429 = n5613 & n18226 ;
  assign n26430 = n633 & ~n26429 ;
  assign n26431 = n26430 ^ n3171 ^ 1'b0 ;
  assign n26432 = n723 & n13426 ;
  assign n26433 = n26432 ^ n22301 ^ 1'b0 ;
  assign n26434 = n26431 | n26433 ;
  assign n26435 = ~n6817 & n8630 ;
  assign n26436 = n26435 ^ n6407 ^ 1'b0 ;
  assign n26437 = n13115 ^ n7675 ^ 1'b0 ;
  assign n26438 = n26436 | n26437 ;
  assign n26439 = n26438 ^ n14795 ^ n2330 ;
  assign n26440 = n5155 & n21338 ;
  assign n26441 = n14593 | n26440 ;
  assign n26442 = n9815 | n26441 ;
  assign n26443 = n4447 & ~n8070 ;
  assign n26444 = n26443 ^ n16911 ^ 1'b0 ;
  assign n26445 = n15956 | n26444 ;
  assign n26446 = n10240 ^ n7392 ^ 1'b0 ;
  assign n26447 = n6225 & ~n26446 ;
  assign n26448 = ~n23691 & n26447 ;
  assign n26449 = n16813 | n19341 ;
  assign n26450 = n26449 ^ n24853 ^ 1'b0 ;
  assign n26452 = n5334 & n10527 ;
  assign n26453 = n11794 & n26452 ;
  assign n26451 = n3941 | n20179 ;
  assign n26454 = n26453 ^ n26451 ^ 1'b0 ;
  assign n26455 = n703 | n9819 ;
  assign n26456 = n3487 | n26455 ;
  assign n26457 = n26456 ^ n25839 ^ 1'b0 ;
  assign n26458 = n26048 ^ n522 ^ 1'b0 ;
  assign n26459 = n1657 & ~n26458 ;
  assign n26460 = n2637 | n12349 ;
  assign n26465 = n23026 ^ n14374 ^ 1'b0 ;
  assign n26466 = n9562 & ~n26465 ;
  assign n26467 = ~n8512 & n26466 ;
  assign n26468 = ~n6258 & n26467 ;
  assign n26461 = n8200 & n12425 ;
  assign n26462 = ~n11116 & n12963 ;
  assign n26463 = ~n26461 & n26462 ;
  assign n26464 = x247 & ~n26463 ;
  assign n26469 = n26468 ^ n26464 ^ 1'b0 ;
  assign n26471 = n5384 & n5695 ;
  assign n26472 = n26471 ^ n3556 ^ 1'b0 ;
  assign n26470 = ~n2668 & n5125 ;
  assign n26473 = n26472 ^ n26470 ^ 1'b0 ;
  assign n26474 = n5398 & n21729 ;
  assign n26475 = n23960 ^ n6085 ^ 1'b0 ;
  assign n26476 = n12423 & ~n26475 ;
  assign n26477 = n614 | n9122 ;
  assign n26478 = n26477 ^ n2903 ^ 1'b0 ;
  assign n26479 = n24181 ^ n16058 ^ 1'b0 ;
  assign n26480 = n26478 | n26479 ;
  assign n26481 = n4364 & n18448 ;
  assign n26482 = n23254 ^ n3747 ^ 1'b0 ;
  assign n26483 = n8150 | n26482 ;
  assign n26484 = n4720 | n10392 ;
  assign n26485 = n26484 ^ n22977 ^ 1'b0 ;
  assign n26486 = n3563 & ~n14995 ;
  assign n26487 = n26486 ^ n5639 ^ 1'b0 ;
  assign n26488 = n10929 & n26487 ;
  assign n26489 = ( n11268 & n21277 ) | ( n11268 & n26488 ) | ( n21277 & n26488 ) ;
  assign n26490 = ~n6005 & n26489 ;
  assign n26491 = n26490 ^ n685 ^ 1'b0 ;
  assign n26492 = n26491 ^ n13314 ^ 1'b0 ;
  assign n26493 = n3618 | n9553 ;
  assign n26494 = n18530 ^ n15867 ^ 1'b0 ;
  assign n26495 = n9900 & n15891 ;
  assign n26496 = ~n12963 & n16054 ;
  assign n26497 = n9102 & n10054 ;
  assign n26498 = ~n10054 & n26497 ;
  assign n26499 = n11886 | n26498 ;
  assign n26500 = n754 | n26499 ;
  assign n26501 = n14652 ^ n10097 ^ 1'b0 ;
  assign n26502 = n9076 & n26501 ;
  assign n26503 = ~n5498 & n20983 ;
  assign n26504 = ~n26502 & n26503 ;
  assign n26505 = ( ~n6145 & n10965 ) | ( ~n6145 & n19387 ) | ( n10965 & n19387 ) ;
  assign n26506 = n6297 & ~n21626 ;
  assign n26507 = n26506 ^ n10887 ^ 1'b0 ;
  assign n26508 = n19046 ^ n17607 ^ n2072 ;
  assign n26509 = n15135 ^ n3664 ^ 1'b0 ;
  assign n26510 = n26508 | n26509 ;
  assign n26511 = n4949 & n5976 ;
  assign n26512 = ~n526 & n944 ;
  assign n26513 = ~n6998 & n26512 ;
  assign n26514 = n9418 & ~n26513 ;
  assign n26515 = ~n6985 & n16015 ;
  assign n26516 = n19644 ^ n7991 ^ 1'b0 ;
  assign n26517 = ~n9594 & n10295 ;
  assign n26518 = n10778 & n12940 ;
  assign n26519 = n1663 | n21121 ;
  assign n26520 = n26519 ^ n16004 ^ 1'b0 ;
  assign n26521 = n26518 | n26520 ;
  assign n26522 = n3702 & ~n20931 ;
  assign n26523 = n13082 & ~n26522 ;
  assign n26524 = x63 & n4999 ;
  assign n26525 = n1159 & n26524 ;
  assign n26526 = n9092 | n26525 ;
  assign n26527 = n16667 | n26526 ;
  assign n26528 = n19319 ^ n4433 ^ 1'b0 ;
  assign n26529 = n26527 & n26528 ;
  assign n26532 = n13445 ^ n6401 ^ 1'b0 ;
  assign n26530 = n15690 ^ n11242 ^ n1514 ;
  assign n26531 = n6100 & ~n26530 ;
  assign n26533 = n26532 ^ n26531 ^ 1'b0 ;
  assign n26534 = ~n2362 & n17174 ;
  assign n26536 = n25061 ^ x91 ^ 1'b0 ;
  assign n26535 = n3283 | n13307 ;
  assign n26537 = n26536 ^ n26535 ^ 1'b0 ;
  assign n26538 = n5360 ^ n3288 ^ 1'b0 ;
  assign n26539 = n13458 | n26538 ;
  assign n26540 = n26539 ^ n15956 ^ 1'b0 ;
  assign n26541 = n17923 | n26540 ;
  assign n26542 = n7402 & ~n26541 ;
  assign n26543 = n19253 ^ n6043 ^ 1'b0 ;
  assign n26544 = ~n610 & n26543 ;
  assign n26545 = n15090 ^ n7964 ^ 1'b0 ;
  assign n26546 = n19269 & n26545 ;
  assign n26547 = n11892 ^ n3960 ^ 1'b0 ;
  assign n26548 = n21358 ^ n1850 ^ 1'b0 ;
  assign n26549 = n26547 & ~n26548 ;
  assign n26550 = x125 & n6693 ;
  assign n26551 = n3314 & n15657 ;
  assign n26552 = ( ~n5560 & n6651 ) | ( ~n5560 & n8059 ) | ( n6651 & n8059 ) ;
  assign n26553 = n17167 | n26552 ;
  assign n26554 = n26553 ^ n20177 ^ 1'b0 ;
  assign n26555 = n15088 | n15217 ;
  assign n26556 = n9211 ^ n3943 ^ n1703 ;
  assign n26557 = n26556 ^ n2247 ^ 1'b0 ;
  assign n26558 = n6381 | n8402 ;
  assign n26559 = n26558 ^ n2955 ^ 1'b0 ;
  assign n26560 = n26559 ^ n820 ^ 1'b0 ;
  assign n26562 = n15611 ^ n1605 ^ 1'b0 ;
  assign n26563 = n15316 & n26562 ;
  assign n26561 = n1173 & n2239 ;
  assign n26564 = n26563 ^ n26561 ^ 1'b0 ;
  assign n26565 = n26564 ^ n1588 ^ 1'b0 ;
  assign n26566 = ~n7064 & n21886 ;
  assign n26567 = n13795 | n16333 ;
  assign n26568 = n13892 & ~n26567 ;
  assign n26569 = n12848 & ~n26568 ;
  assign n26570 = n26569 ^ n20871 ^ 1'b0 ;
  assign n26571 = n5686 & ~n22041 ;
  assign n26572 = n16387 | n20685 ;
  assign n26573 = n3924 & ~n23280 ;
  assign n26574 = n20241 & n26573 ;
  assign n26575 = n2910 | n26574 ;
  assign n26576 = n26575 ^ n13602 ^ 1'b0 ;
  assign n26577 = n26572 & ~n26576 ;
  assign n26578 = ~n8771 & n8937 ;
  assign n26579 = n14856 & n26578 ;
  assign n26580 = n11063 ^ n10265 ^ 1'b0 ;
  assign n26581 = ~n3723 & n26580 ;
  assign n26582 = n17980 | n25774 ;
  assign n26583 = n8041 | n13899 ;
  assign n26584 = n2083 | n26583 ;
  assign n26585 = n3145 & ~n4358 ;
  assign n26586 = n4158 & n26585 ;
  assign n26587 = ~n21801 & n26586 ;
  assign n26588 = ~n26584 & n26587 ;
  assign n26589 = ~n2257 & n3171 ;
  assign n26590 = ~n4880 & n26589 ;
  assign n26591 = n26590 ^ n2469 ^ 1'b0 ;
  assign n26592 = ~n1556 & n18430 ;
  assign n26593 = n16887 & n26592 ;
  assign n26594 = x176 | n732 ;
  assign n26595 = n26594 ^ n18015 ^ 1'b0 ;
  assign n26596 = n15241 ^ n13697 ^ 1'b0 ;
  assign n26597 = n2786 | n12930 ;
  assign n26598 = n12657 ^ n10691 ^ 1'b0 ;
  assign n26599 = ~n7888 & n13271 ;
  assign n26600 = n21069 & n26599 ;
  assign n26601 = n6872 & n14601 ;
  assign n26602 = n1843 & n2039 ;
  assign n26603 = n26602 ^ n2892 ^ n2467 ;
  assign n26604 = n12667 & ~n26603 ;
  assign n26605 = n26604 ^ n7276 ^ 1'b0 ;
  assign n26606 = n5072 & ~n5996 ;
  assign n26607 = n4712 ^ n4021 ^ 1'b0 ;
  assign n26608 = n20350 ^ n19023 ^ 1'b0 ;
  assign n26609 = n26607 & n26608 ;
  assign n26610 = n5218 | n11538 ;
  assign n26611 = n21915 | n26610 ;
  assign n26612 = n9339 & ~n26611 ;
  assign n26613 = n16923 & n20398 ;
  assign n26614 = n26613 ^ n1419 ^ 1'b0 ;
  assign n26615 = n26614 ^ n13941 ^ 1'b0 ;
  assign n26616 = n6823 | n13256 ;
  assign n26617 = ~n6637 & n6999 ;
  assign n26618 = ~n26616 & n26617 ;
  assign n26619 = ~n1608 & n26618 ;
  assign n26620 = n8668 ^ n2577 ^ 1'b0 ;
  assign n26621 = ~n4622 & n26620 ;
  assign n26622 = n26621 ^ n7757 ^ 1'b0 ;
  assign n26623 = n10051 ^ n7508 ^ 1'b0 ;
  assign n26624 = ~n26622 & n26623 ;
  assign n26625 = ( n1256 & n3463 ) | ( n1256 & ~n18605 ) | ( n3463 & ~n18605 ) ;
  assign n26626 = n26625 ^ n1237 ^ 1'b0 ;
  assign n26627 = ~n3045 & n3735 ;
  assign n26628 = ~n793 & n26627 ;
  assign n26629 = n8182 | n8811 ;
  assign n26630 = ~x31 & n2887 ;
  assign n26631 = n4289 ^ n2689 ^ 1'b0 ;
  assign n26632 = n23039 & ~n26631 ;
  assign n26633 = n26632 ^ n7437 ^ 1'b0 ;
  assign n26634 = ~n26630 & n26633 ;
  assign n26635 = n14872 ^ n4675 ^ 1'b0 ;
  assign n26636 = ~n3727 & n26635 ;
  assign n26637 = ~n2228 & n26636 ;
  assign n26638 = n3062 ^ n2237 ^ 1'b0 ;
  assign n26639 = n26637 & ~n26638 ;
  assign n26640 = ~x180 & n4671 ;
  assign n26641 = n3622 & ~n15090 ;
  assign n26642 = ( n4899 & n20944 ) | ( n4899 & n26641 ) | ( n20944 & n26641 ) ;
  assign n26643 = n4470 & ~n26642 ;
  assign n26644 = n566 | n22106 ;
  assign n26645 = n10213 & ~n15098 ;
  assign n26646 = n11803 ^ n4300 ^ n816 ;
  assign n26647 = ~n1405 & n3733 ;
  assign n26648 = n15641 ^ n12694 ^ n11538 ;
  assign n26651 = n20514 ^ n10498 ^ 1'b0 ;
  assign n26649 = n15341 ^ n4334 ^ 1'b0 ;
  assign n26650 = n15913 & n26649 ;
  assign n26652 = n26651 ^ n26650 ^ 1'b0 ;
  assign n26653 = n26648 & n26652 ;
  assign n26654 = n2493 | n3274 ;
  assign n26655 = n13905 | n14632 ;
  assign n26657 = n4949 & n22658 ;
  assign n26658 = n21764 & n26657 ;
  assign n26656 = n1286 & ~n18859 ;
  assign n26659 = n26658 ^ n26656 ^ 1'b0 ;
  assign n26660 = n21093 ^ n14501 ^ 1'b0 ;
  assign n26661 = n26651 ^ n24967 ^ 1'b0 ;
  assign n26663 = ~n4540 & n6682 ;
  assign n26662 = n14197 | n18465 ;
  assign n26664 = n26663 ^ n26662 ^ 1'b0 ;
  assign n26665 = n18700 | n26664 ;
  assign n26666 = n26665 ^ n11266 ^ 1'b0 ;
  assign n26667 = n8432 & ~n23432 ;
  assign n26668 = n18755 ^ n9249 ^ 1'b0 ;
  assign n26669 = n11137 ^ n8877 ^ 1'b0 ;
  assign n26670 = n1757 & ~n13295 ;
  assign n26671 = n12389 ^ n3245 ^ 1'b0 ;
  assign n26672 = n23020 ^ n16898 ^ x123 ;
  assign n26673 = n2539 | n26672 ;
  assign n26674 = n17683 & n23739 ;
  assign n26675 = ~n11689 & n26674 ;
  assign n26676 = n2629 & ~n19540 ;
  assign n26677 = n24966 ^ n10548 ^ 1'b0 ;
  assign n26678 = ~n715 & n4971 ;
  assign n26679 = ~n26677 & n26678 ;
  assign n26680 = n2148 & ~n7448 ;
  assign n26681 = ~n1311 & n26680 ;
  assign n26682 = n833 | n3669 ;
  assign n26683 = n18305 & ~n26682 ;
  assign n26684 = n26681 & n26683 ;
  assign n26685 = n25543 ^ n4680 ^ 1'b0 ;
  assign n26686 = n9057 & ~n26685 ;
  assign n26687 = n14858 ^ n8921 ^ 1'b0 ;
  assign n26688 = n1291 | n26687 ;
  assign n26689 = n6617 | n20359 ;
  assign n26690 = n10677 | n25388 ;
  assign n26691 = n26690 ^ n3994 ^ 1'b0 ;
  assign n26692 = n5259 ^ n2858 ^ 1'b0 ;
  assign n26693 = n11242 & ~n26692 ;
  assign n26694 = ~n26691 & n26693 ;
  assign n26695 = ~n6623 & n11214 ;
  assign n26696 = n17821 & n26695 ;
  assign n26697 = n26696 ^ n2720 ^ 1'b0 ;
  assign n26698 = n26694 | n26697 ;
  assign n26699 = ~n7331 & n10843 ;
  assign n26700 = n3639 & ~n11662 ;
  assign n26701 = n11919 & n26700 ;
  assign n26703 = ~n6892 & n25066 ;
  assign n26702 = n8408 & ~n22897 ;
  assign n26704 = n26703 ^ n26702 ^ 1'b0 ;
  assign n26705 = ~n2063 & n15630 ;
  assign n26706 = n10063 | n26705 ;
  assign n26707 = n26706 ^ n11934 ^ 1'b0 ;
  assign n26708 = n987 & ~n26707 ;
  assign n26709 = n7427 ^ n5317 ^ 1'b0 ;
  assign n26711 = n26602 ^ n2892 ^ 1'b0 ;
  assign n26712 = n26711 ^ n2467 ^ 1'b0 ;
  assign n26710 = x116 & ~n4568 ;
  assign n26713 = n26712 ^ n26710 ^ 1'b0 ;
  assign n26714 = n16326 ^ n1501 ^ 1'b0 ;
  assign n26715 = n448 & n26714 ;
  assign n26716 = ( n8892 & ~n9816 ) | ( n8892 & n10604 ) | ( ~n9816 & n10604 ) ;
  assign n26717 = ~n17282 & n26716 ;
  assign n26718 = n26717 ^ n1880 ^ 1'b0 ;
  assign n26720 = n3248 & ~n13293 ;
  assign n26721 = n26720 ^ n7164 ^ 1'b0 ;
  assign n26722 = n26721 ^ n589 ^ 1'b0 ;
  assign n26719 = ~n15829 & n24644 ;
  assign n26723 = n26722 ^ n26719 ^ 1'b0 ;
  assign n26724 = n14693 & ~n26653 ;
  assign n26725 = ~n7895 & n8256 ;
  assign n26726 = ~n17005 & n26725 ;
  assign n26727 = n2966 ^ n1071 ^ 1'b0 ;
  assign n26728 = n16766 & ~n26727 ;
  assign n26729 = n26728 ^ n19474 ^ 1'b0 ;
  assign n26730 = ~n26726 & n26729 ;
  assign n26731 = n12760 ^ n6051 ^ 1'b0 ;
  assign n26732 = n10346 & ~n26731 ;
  assign n26733 = n2044 & n26732 ;
  assign n26734 = n26733 ^ n3695 ^ 1'b0 ;
  assign n26735 = ~n10690 & n18613 ;
  assign n26736 = n26735 ^ n8550 ^ 1'b0 ;
  assign n26737 = n20174 & n24261 ;
  assign n26738 = n13496 ^ n9651 ^ 1'b0 ;
  assign n26739 = n13206 ^ n5420 ^ 1'b0 ;
  assign n26740 = ~n26738 & n26739 ;
  assign n26741 = n7888 ^ n4340 ^ 1'b0 ;
  assign n26742 = n2423 & n26741 ;
  assign n26743 = ~n10223 & n26742 ;
  assign n26744 = n790 & n12962 ;
  assign n26745 = n1415 & ~n26744 ;
  assign n26746 = n26745 ^ n24364 ^ 1'b0 ;
  assign n26747 = n26746 ^ n9068 ^ 1'b0 ;
  assign n26748 = x106 & n26747 ;
  assign n26749 = n7749 & n9427 ;
  assign n26750 = n26749 ^ n4891 ^ 1'b0 ;
  assign n26751 = ~x157 & n10591 ;
  assign n26752 = n1202 & n26751 ;
  assign n26753 = n781 & ~n26752 ;
  assign n26754 = x25 & n26753 ;
  assign n26755 = n26754 ^ n25712 ^ 1'b0 ;
  assign n26756 = n16770 ^ n641 ^ 1'b0 ;
  assign n26757 = n1850 & ~n16608 ;
  assign n26758 = n26757 ^ n9413 ^ 1'b0 ;
  assign n26759 = ~n5443 & n15789 ;
  assign n26760 = ~n26758 & n26759 ;
  assign n26761 = ~x228 & n2179 ;
  assign n26762 = n26761 ^ n5903 ^ n3210 ;
  assign n26765 = n20474 ^ n6015 ^ 1'b0 ;
  assign n26766 = n11478 & ~n26765 ;
  assign n26763 = n948 | n2627 ;
  assign n26764 = n20171 & n26763 ;
  assign n26767 = n26766 ^ n26764 ^ 1'b0 ;
  assign n26768 = n15458 & ~n26767 ;
  assign n26769 = n13286 ^ n3903 ^ 1'b0 ;
  assign n26770 = n1507 | n26769 ;
  assign n26771 = n2185 | n11101 ;
  assign n26776 = n22160 ^ n13477 ^ 1'b0 ;
  assign n26772 = n25933 ^ n8333 ^ 1'b0 ;
  assign n26773 = n14285 ^ n3298 ^ 1'b0 ;
  assign n26774 = ~n26772 & n26773 ;
  assign n26775 = ~n18459 & n26774 ;
  assign n26777 = n26776 ^ n26775 ^ 1'b0 ;
  assign n26778 = ~n1481 & n22067 ;
  assign n26779 = n26778 ^ n6231 ^ 1'b0 ;
  assign n26780 = n4741 & n8279 ;
  assign n26781 = n26780 ^ n2437 ^ 1'b0 ;
  assign n26782 = n12846 & n17036 ;
  assign n26783 = n26782 ^ n24389 ^ 1'b0 ;
  assign n26784 = n17591 ^ n9910 ^ 1'b0 ;
  assign n26785 = n5883 ^ n4648 ^ 1'b0 ;
  assign n26786 = n26784 & ~n26785 ;
  assign n26787 = n26786 ^ n6757 ^ 1'b0 ;
  assign n26788 = n2615 & n26787 ;
  assign n26789 = x102 & n16460 ;
  assign n26790 = ~n26788 & n26789 ;
  assign n26791 = n26790 ^ n20751 ^ 1'b0 ;
  assign n26792 = n896 ^ n492 ^ 1'b0 ;
  assign n26793 = n8962 & n26792 ;
  assign n26794 = ~n2219 & n26793 ;
  assign n26795 = n26794 ^ n17054 ^ 1'b0 ;
  assign n26796 = ~n3059 & n6435 ;
  assign n26797 = n1475 & n26796 ;
  assign n26798 = ~n26411 & n26797 ;
  assign n26800 = n5465 & ~n7750 ;
  assign n26801 = n9331 & n26800 ;
  assign n26799 = n12136 & n18448 ;
  assign n26802 = n26801 ^ n26799 ^ 1'b0 ;
  assign n26803 = n1773 & ~n16811 ;
  assign n26804 = n20621 ^ n788 ^ 1'b0 ;
  assign n26805 = n13161 | n21570 ;
  assign n26806 = n26805 ^ n19469 ^ 1'b0 ;
  assign n26807 = n6824 | n14053 ;
  assign n26808 = n985 & ~n26807 ;
  assign n26809 = ~n3187 & n20359 ;
  assign n26810 = ~n5516 & n16007 ;
  assign n26811 = n26810 ^ n11683 ^ 1'b0 ;
  assign n26812 = n26811 ^ n16777 ^ 1'b0 ;
  assign n26813 = n10650 ^ n458 ^ 1'b0 ;
  assign n26814 = x181 & ~n26409 ;
  assign n26815 = n26814 ^ n8126 ^ 1'b0 ;
  assign n26816 = n8048 & n8242 ;
  assign n26817 = n19017 & n26816 ;
  assign n26818 = n26817 ^ n13630 ^ 1'b0 ;
  assign n26819 = n26818 ^ n2310 ^ 1'b0 ;
  assign n26820 = n6762 & ~n12151 ;
  assign n26821 = n669 | n9432 ;
  assign n26822 = n26821 ^ n23435 ^ 1'b0 ;
  assign n26823 = n26820 & n26822 ;
  assign n26824 = n15768 & ~n20809 ;
  assign n26825 = n26824 ^ n23948 ^ 1'b0 ;
  assign n26826 = n11294 & ~n22361 ;
  assign n26827 = n26826 ^ n15620 ^ 1'b0 ;
  assign n26828 = n16463 & ~n26827 ;
  assign n26829 = n26825 | n26828 ;
  assign n26830 = n2701 | n26829 ;
  assign n26832 = n12014 ^ n1765 ^ 1'b0 ;
  assign n26831 = n8692 | n15075 ;
  assign n26833 = n26832 ^ n26831 ^ 1'b0 ;
  assign n26834 = n7721 | n12911 ;
  assign n26835 = n8491 & ~n25173 ;
  assign n26836 = n10735 ^ x106 ^ 1'b0 ;
  assign n26837 = n9477 & n18684 ;
  assign n26838 = n11694 ^ n3713 ^ 1'b0 ;
  assign n26839 = n26838 ^ n2599 ^ 1'b0 ;
  assign n26840 = ~n25178 & n26839 ;
  assign n26841 = ~n14599 & n26840 ;
  assign n26842 = n18630 ^ n4217 ^ 1'b0 ;
  assign n26843 = ~n813 & n2449 ;
  assign n26844 = ~n5994 & n18576 ;
  assign n26845 = n1651 & ~n1859 ;
  assign n26846 = n4931 ^ n2790 ^ 1'b0 ;
  assign n26847 = n26846 ^ n24134 ^ 1'b0 ;
  assign n26848 = n26845 & n26847 ;
  assign n26849 = n23983 ^ n5282 ^ 1'b0 ;
  assign n26850 = ~n15860 & n26849 ;
  assign n26851 = n15803 | n26445 ;
  assign n26852 = n26851 ^ n7910 ^ 1'b0 ;
  assign n26853 = n2248 | n3465 ;
  assign n26854 = n994 | n26853 ;
  assign n26855 = n26854 ^ n16798 ^ 1'b0 ;
  assign n26856 = n11929 & ~n26855 ;
  assign n26857 = ~n950 & n5175 ;
  assign n26858 = n26857 ^ n5492 ^ 1'b0 ;
  assign n26859 = n12849 & ~n14058 ;
  assign n26860 = ~n8613 & n26859 ;
  assign n26861 = n2404 & ~n26860 ;
  assign n26862 = n9832 & n26861 ;
  assign n26863 = n21148 ^ n5838 ^ 1'b0 ;
  assign n26864 = n1228 & ~n26863 ;
  assign n26865 = n19652 ^ n12256 ^ n8874 ;
  assign n26866 = n15959 & n19054 ;
  assign n26867 = n12364 & ~n26866 ;
  assign n26868 = n5419 | n7438 ;
  assign n26869 = n6783 | n26868 ;
  assign n26870 = ~n7109 & n26869 ;
  assign n26871 = n4526 & n26870 ;
  assign n26872 = n666 & ~n1472 ;
  assign n26873 = n26872 ^ n9776 ^ 1'b0 ;
  assign n26874 = n19895 ^ n9902 ^ n5634 ;
  assign n26875 = n26874 ^ x20 ^ 1'b0 ;
  assign n26876 = ~n26873 & n26875 ;
  assign n26877 = n15423 & ~n20579 ;
  assign n26878 = n26877 ^ n23617 ^ 1'b0 ;
  assign n26879 = n1739 | n26878 ;
  assign n26880 = ~n1195 & n12164 ;
  assign n26881 = ~n13570 & n26880 ;
  assign n26882 = n15183 & ~n17068 ;
  assign n26883 = n5326 | n5597 ;
  assign n26884 = n26883 ^ n1368 ^ 1'b0 ;
  assign n26885 = n10300 ^ n3153 ^ 1'b0 ;
  assign n26886 = n4789 & ~n24645 ;
  assign n26887 = n23294 ^ n2610 ^ 1'b0 ;
  assign n26888 = n26886 & ~n26887 ;
  assign n26889 = n5390 ^ n2587 ^ 1'b0 ;
  assign n26890 = n1658 | n26889 ;
  assign n26891 = n818 | n26890 ;
  assign n26892 = ~n18048 & n26891 ;
  assign n26893 = ~n25465 & n26892 ;
  assign n26894 = n19851 ^ n10886 ^ 1'b0 ;
  assign n26895 = ~n19534 & n24321 ;
  assign n26896 = n19341 & n26895 ;
  assign n26897 = ~n1644 & n10630 ;
  assign n26898 = ~n20517 & n26897 ;
  assign n26899 = n26898 ^ n14817 ^ 1'b0 ;
  assign n26900 = ( ~n4122 & n11217 ) | ( ~n4122 & n15533 ) | ( n11217 & n15533 ) ;
  assign n26901 = n10418 & ~n26900 ;
  assign n26902 = n936 & ~n8586 ;
  assign n26903 = n26902 ^ n14195 ^ 1'b0 ;
  assign n26904 = n8090 ^ n6468 ^ 1'b0 ;
  assign n26905 = n14495 & ~n26904 ;
  assign n26906 = n2001 | n3902 ;
  assign n26907 = ~n2210 & n26906 ;
  assign n26913 = ~n2157 & n21995 ;
  assign n26914 = ~n6747 & n26913 ;
  assign n26908 = n936 & n14852 ;
  assign n26909 = n832 & n26908 ;
  assign n26910 = n13046 & n26909 ;
  assign n26911 = n7425 & ~n26910 ;
  assign n26912 = n26911 ^ n10530 ^ 1'b0 ;
  assign n26915 = n26914 ^ n26912 ^ 1'b0 ;
  assign n26916 = n26915 ^ n17269 ^ 1'b0 ;
  assign n26917 = ~n1535 & n5799 ;
  assign n26918 = ~n4928 & n26917 ;
  assign n26919 = ( n4705 & n13876 ) | ( n4705 & n26918 ) | ( n13876 & n26918 ) ;
  assign n26920 = n15471 & n22789 ;
  assign n26921 = n9183 & n26920 ;
  assign n26922 = ~n8520 & n10904 ;
  assign n26923 = n26921 & n26922 ;
  assign n26924 = n6849 & n8442 ;
  assign n26925 = n26924 ^ n17521 ^ 1'b0 ;
  assign n26926 = ~n5285 & n26925 ;
  assign n26927 = n14399 ^ n5250 ^ 1'b0 ;
  assign n26928 = n10567 | n13763 ;
  assign n26929 = ~n3197 & n7448 ;
  assign n26930 = ~n11855 & n22705 ;
  assign n26931 = ~n6351 & n26930 ;
  assign n26932 = n26931 ^ n16694 ^ 1'b0 ;
  assign n26933 = n9682 & n17193 ;
  assign n26934 = ~n15161 & n26933 ;
  assign n26935 = n8992 & n9300 ;
  assign n26936 = n18762 | n25631 ;
  assign n26937 = n26935 | n26936 ;
  assign n26938 = ~n18629 & n26937 ;
  assign n26939 = n26938 ^ n14798 ^ 1'b0 ;
  assign n26940 = n10771 & n17061 ;
  assign n26941 = n26940 ^ n2860 ^ 1'b0 ;
  assign n26942 = n6141 ^ n6052 ^ 1'b0 ;
  assign n26943 = n2292 & n26942 ;
  assign n26944 = n13673 ^ n690 ^ 1'b0 ;
  assign n26945 = n26944 ^ n631 ^ 1'b0 ;
  assign n26946 = n26943 & n26945 ;
  assign n26947 = ~n16209 & n17520 ;
  assign n26948 = n10500 & n26947 ;
  assign n26949 = n3624 & n8209 ;
  assign n26950 = n4910 | n23512 ;
  assign n26951 = n7017 & n9040 ;
  assign n26952 = n21764 & n26951 ;
  assign n26953 = n26357 ^ n13901 ^ 1'b0 ;
  assign n26954 = n19275 ^ n13235 ^ 1'b0 ;
  assign n26955 = n26953 & n26954 ;
  assign n26956 = n19716 ^ n5157 ^ 1'b0 ;
  assign n26957 = n20584 | n26956 ;
  assign n26958 = ~n2003 & n16802 ;
  assign n26959 = ~n16802 & n26958 ;
  assign n26960 = n8616 | n26959 ;
  assign n26961 = n9636 & ~n17599 ;
  assign n26962 = n17599 & n26961 ;
  assign n26963 = n26960 | n26962 ;
  assign n26964 = ( n5207 & ~n9778 ) | ( n5207 & n26963 ) | ( ~n9778 & n26963 ) ;
  assign n26965 = ~n17514 & n17611 ;
  assign n26966 = n6343 & n26965 ;
  assign n26967 = n7905 & n15535 ;
  assign n26968 = n26967 ^ n9086 ^ 1'b0 ;
  assign n26969 = n23149 | n25311 ;
  assign n26970 = n20408 | n26969 ;
  assign n26971 = n2480 & ~n7185 ;
  assign n26972 = n26971 ^ n9857 ^ 1'b0 ;
  assign n26973 = ~n3703 & n26972 ;
  assign n26974 = n21807 ^ n15233 ^ 1'b0 ;
  assign n26975 = n1819 & n26974 ;
  assign n26976 = n16028 & ~n18572 ;
  assign n26977 = n21328 ^ n17748 ^ 1'b0 ;
  assign n26978 = ~n18471 & n26977 ;
  assign n26979 = ~n8054 & n17741 ;
  assign n26980 = n26979 ^ n5457 ^ 1'b0 ;
  assign n26981 = n3988 & n17061 ;
  assign n26982 = n26981 ^ n1826 ^ 1'b0 ;
  assign n26983 = ~n2495 & n14951 ;
  assign n26984 = n13426 ^ n12154 ^ n1877 ;
  assign n26985 = n5608 & ~n26984 ;
  assign n26986 = n26985 ^ n14105 ^ 1'b0 ;
  assign n26987 = n5201 & ~n14417 ;
  assign n26988 = n26987 ^ n13919 ^ 1'b0 ;
  assign n26989 = n5140 | n26988 ;
  assign n26990 = n22616 ^ n16109 ^ 1'b0 ;
  assign n26991 = n2063 & n3661 ;
  assign n26992 = ~n526 & n3124 ;
  assign n26993 = n26992 ^ n17931 ^ 1'b0 ;
  assign n26994 = n26991 | n26993 ;
  assign n26995 = n17111 ^ n937 ^ 1'b0 ;
  assign n26996 = n2153 & n22096 ;
  assign n26997 = n2768 & n23245 ;
  assign n26998 = n2976 ^ n1014 ^ 1'b0 ;
  assign n26999 = n1368 & n26998 ;
  assign n27000 = n7689 | n8841 ;
  assign n27001 = n26999 | n27000 ;
  assign n27002 = ~n4681 & n5712 ;
  assign n27003 = n27002 ^ n11526 ^ 1'b0 ;
  assign n27004 = n6432 | n9352 ;
  assign n27005 = x50 & ~n3759 ;
  assign n27007 = n2761 & ~n9076 ;
  assign n27008 = n8555 ^ n4714 ^ 1'b0 ;
  assign n27009 = n27007 & ~n27008 ;
  assign n27006 = n1117 | n11655 ;
  assign n27010 = n27009 ^ n27006 ^ 1'b0 ;
  assign n27011 = n27010 ^ n6333 ^ 1'b0 ;
  assign n27012 = n27005 & ~n27011 ;
  assign n27013 = n4681 ^ n4291 ^ 1'b0 ;
  assign n27016 = n1668 & n14937 ;
  assign n27017 = n27016 ^ n2854 ^ 1'b0 ;
  assign n27018 = ~n9223 & n27017 ;
  assign n27014 = n11740 ^ x170 ^ 1'b0 ;
  assign n27015 = n2653 & n27014 ;
  assign n27019 = n27018 ^ n27015 ^ n4644 ;
  assign n27020 = ( n4804 & n6838 ) | ( n4804 & n7345 ) | ( n6838 & n7345 ) ;
  assign n27021 = ~n8202 & n27020 ;
  assign n27022 = n26017 | n27021 ;
  assign n27023 = n27022 ^ n20345 ^ 1'b0 ;
  assign n27024 = n20627 & ~n27023 ;
  assign n27025 = ~n3882 & n12402 ;
  assign n27026 = n27025 ^ n4409 ^ 1'b0 ;
  assign n27027 = n1554 & n27026 ;
  assign n27028 = ~n901 & n18119 ;
  assign n27029 = n27028 ^ n9707 ^ 1'b0 ;
  assign n27030 = n27027 | n27029 ;
  assign n27031 = n27030 ^ n7199 ^ 1'b0 ;
  assign n27032 = n21495 ^ n978 ^ 1'b0 ;
  assign n27033 = n1383 & n2006 ;
  assign n27034 = n10221 ^ n2068 ^ 1'b0 ;
  assign n27035 = n27033 & ~n27034 ;
  assign n27036 = n21499 & ~n23325 ;
  assign n27037 = ~n26811 & n27036 ;
  assign n27038 = n20186 & ~n27037 ;
  assign n27039 = n27038 ^ n6192 ^ 1'b0 ;
  assign n27042 = n12020 ^ n11387 ^ 1'b0 ;
  assign n27043 = ~n13072 & n27042 ;
  assign n27040 = n14563 ^ n7736 ^ 1'b0 ;
  assign n27041 = ~n19602 & n27040 ;
  assign n27044 = n27043 ^ n27041 ^ 1'b0 ;
  assign n27045 = n16931 & n27044 ;
  assign n27046 = n8348 ^ n3255 ^ 1'b0 ;
  assign n27047 = ~n13630 & n27046 ;
  assign n27048 = ( ~n6152 & n10154 ) | ( ~n6152 & n27047 ) | ( n10154 & n27047 ) ;
  assign n27049 = n1680 | n10330 ;
  assign n27050 = n18806 ^ n8029 ^ n1758 ;
  assign n27051 = ~n22886 & n26211 ;
  assign n27052 = n27051 ^ n10757 ^ 1'b0 ;
  assign n27053 = n6191 | n6560 ;
  assign n27054 = n27053 ^ n1835 ^ 1'b0 ;
  assign n27055 = n18723 ^ n12410 ^ 1'b0 ;
  assign n27056 = n7258 & n27055 ;
  assign n27057 = n1404 | n25442 ;
  assign n27058 = ~n1093 & n4788 ;
  assign n27059 = n27058 ^ n10583 ^ 1'b0 ;
  assign n27060 = n13255 | n27059 ;
  assign n27061 = n27060 ^ n12911 ^ 1'b0 ;
  assign n27062 = n16028 | n19086 ;
  assign n27063 = n13707 | n27062 ;
  assign n27064 = n27061 | n27063 ;
  assign n27065 = n27064 ^ n1126 ^ 1'b0 ;
  assign n27066 = n7727 | n27065 ;
  assign n27067 = n7826 & n26326 ;
  assign n27068 = n14058 ^ n4400 ^ 1'b0 ;
  assign n27069 = n5522 & ~n27068 ;
  assign n27070 = ~n5887 & n27069 ;
  assign n27071 = n17307 & n27070 ;
  assign n27072 = n19137 ^ n8278 ^ 1'b0 ;
  assign n27073 = n19359 ^ n5974 ^ 1'b0 ;
  assign n27074 = n26293 ^ n6146 ^ 1'b0 ;
  assign n27076 = n20677 ^ n1604 ^ 1'b0 ;
  assign n27075 = n10451 & ~n14043 ;
  assign n27077 = n27076 ^ n27075 ^ 1'b0 ;
  assign n27078 = ~n25796 & n27077 ;
  assign n27079 = n27078 ^ n19229 ^ 1'b0 ;
  assign n27080 = n5903 & ~n6523 ;
  assign n27081 = ~n5903 & n27080 ;
  assign n27082 = n7942 | n27081 ;
  assign n27083 = n27081 & ~n27082 ;
  assign n27084 = ~n909 & n25774 ;
  assign n27085 = n450 | n6712 ;
  assign n27086 = n17384 ^ n16454 ^ 1'b0 ;
  assign n27087 = n923 & ~n1269 ;
  assign n27088 = n20790 & n27087 ;
  assign n27089 = n1175 | n26632 ;
  assign n27090 = n17958 ^ n3340 ^ 1'b0 ;
  assign n27091 = n23023 ^ n21122 ^ 1'b0 ;
  assign n27092 = n24808 ^ n22558 ^ 1'b0 ;
  assign n27093 = n5203 | n14404 ;
  assign n27094 = n6616 ^ n5024 ^ 1'b0 ;
  assign n27095 = n2046 & n7583 ;
  assign n27096 = ~n2351 & n27095 ;
  assign n27097 = n27096 ^ n14447 ^ 1'b0 ;
  assign n27098 = n27094 | n27097 ;
  assign n27099 = n25712 & ~n27098 ;
  assign n27100 = n14508 & ~n17084 ;
  assign n27101 = n27100 ^ n11656 ^ 1'b0 ;
  assign n27102 = n841 & ~n12154 ;
  assign n27103 = n27102 ^ n2358 ^ 1'b0 ;
  assign n27104 = n11743 | n27103 ;
  assign n27105 = n6516 & ~n27104 ;
  assign n27106 = n27105 ^ n1510 ^ 1'b0 ;
  assign n27107 = n3281 & ~n12142 ;
  assign n27108 = n26385 ^ n20263 ^ 1'b0 ;
  assign n27109 = n20144 ^ n13241 ^ n5761 ;
  assign n27110 = n4395 & ~n8667 ;
  assign n27111 = ~x21 & n27110 ;
  assign n27112 = n6517 & n15083 ;
  assign n27113 = n27111 & n27112 ;
  assign n27114 = n6375 ^ n5529 ^ 1'b0 ;
  assign n27115 = n27113 | n27114 ;
  assign n27116 = ~n2392 & n10813 ;
  assign n27117 = ~x77 & n27116 ;
  assign n27118 = ~n3385 & n13268 ;
  assign n27119 = n16658 | n27118 ;
  assign n27120 = n10678 | n27119 ;
  assign n27121 = n3386 | n8509 ;
  assign n27122 = n1914 & n10507 ;
  assign n27123 = n3546 | n14637 ;
  assign n27125 = n10714 ^ n5222 ^ 1'b0 ;
  assign n27126 = n9320 & n27125 ;
  assign n27124 = n11885 | n20263 ;
  assign n27127 = n27126 ^ n27124 ^ 1'b0 ;
  assign n27128 = n2470 | n13833 ;
  assign n27129 = n3060 | n27128 ;
  assign n27130 = n4749 & n27129 ;
  assign n27131 = n27130 ^ n2089 ^ 1'b0 ;
  assign n27132 = n2744 & n5519 ;
  assign n27133 = n2264 | n3565 ;
  assign n27134 = n27133 ^ n1964 ^ 1'b0 ;
  assign n27135 = n5740 & ~n27134 ;
  assign n27136 = n27135 ^ n14238 ^ 1'b0 ;
  assign n27137 = n5192 & n15379 ;
  assign n27138 = n27137 ^ n9083 ^ 1'b0 ;
  assign n27139 = n11758 & n27138 ;
  assign n27140 = ~n3127 & n27139 ;
  assign n27141 = n27140 ^ n13428 ^ 1'b0 ;
  assign n27142 = n15531 & n27141 ;
  assign n27143 = n4267 | n14639 ;
  assign n27144 = n27143 ^ n16645 ^ 1'b0 ;
  assign n27145 = n19621 | n27144 ;
  assign n27146 = n4723 & n17499 ;
  assign n27147 = n14550 ^ n6496 ^ 1'b0 ;
  assign n27148 = n6396 & ~n23868 ;
  assign n27149 = ~n2305 & n26463 ;
  assign n27150 = n4888 | n21365 ;
  assign n27151 = n27150 ^ n24947 ^ 1'b0 ;
  assign n27152 = n13752 ^ n4321 ^ 1'b0 ;
  assign n27153 = n22825 & ~n27152 ;
  assign n27154 = n1557 ^ n292 ^ 1'b0 ;
  assign n27155 = n880 & ~n27154 ;
  assign n27156 = n27155 ^ n17038 ^ 1'b0 ;
  assign n27157 = n7704 ^ n630 ^ 1'b0 ;
  assign n27158 = n7884 | n27157 ;
  assign n27159 = n11166 | n27158 ;
  assign n27160 = n27156 | n27159 ;
  assign n27161 = n1299 & ~n11814 ;
  assign n27162 = n729 & ~n2826 ;
  assign n27163 = ~n12502 & n27162 ;
  assign n27164 = n4705 & ~n9550 ;
  assign n27165 = n27164 ^ n15475 ^ 1'b0 ;
  assign n27167 = n12543 & ~n14937 ;
  assign n27166 = n2629 & ~n2722 ;
  assign n27168 = n27167 ^ n27166 ^ 1'b0 ;
  assign n27169 = n17546 ^ n12379 ^ 1'b0 ;
  assign n27170 = n2143 | n26630 ;
  assign n27171 = n27169 & n27170 ;
  assign n27172 = n8284 & n27171 ;
  assign n27173 = x212 & ~n27172 ;
  assign n27174 = ~n27168 & n27173 ;
  assign n27175 = n5711 & ~n24936 ;
  assign n27176 = n14645 & n27175 ;
  assign n27177 = n27176 ^ n18452 ^ 1'b0 ;
  assign n27178 = n5052 | n20844 ;
  assign n27179 = n6861 | n27178 ;
  assign n27180 = ~n9074 & n27179 ;
  assign n27181 = n27180 ^ n4703 ^ 1'b0 ;
  assign n27182 = n7529 & n24336 ;
  assign n27183 = ~n4840 & n25829 ;
  assign n27184 = n27183 ^ n4185 ^ 1'b0 ;
  assign n27185 = n10458 ^ n8611 ^ 1'b0 ;
  assign n27186 = n5560 | n11219 ;
  assign n27187 = n27186 ^ n5021 ^ 1'b0 ;
  assign n27188 = n5903 | n27187 ;
  assign n27189 = n27188 ^ n3966 ^ 1'b0 ;
  assign n27190 = n7350 & ~n27189 ;
  assign n27191 = n11335 & n16244 ;
  assign n27192 = ~n5265 & n27191 ;
  assign n27193 = n21445 ^ n14803 ^ 1'b0 ;
  assign n27194 = n7582 | n27193 ;
  assign n27195 = n27194 ^ n22410 ^ 1'b0 ;
  assign n27196 = ~n10757 & n17004 ;
  assign n27197 = ~n11983 & n27196 ;
  assign n27198 = n1990 & ~n27197 ;
  assign n27199 = n3321 & n4701 ;
  assign n27200 = n27198 & n27199 ;
  assign n27201 = n24198 & n27200 ;
  assign n27202 = n27201 ^ n8679 ^ 1'b0 ;
  assign n27203 = n4700 & n9869 ;
  assign n27204 = n27203 ^ n1622 ^ 1'b0 ;
  assign n27205 = n19313 ^ n3703 ^ 1'b0 ;
  assign n27206 = ~n22356 & n27205 ;
  assign n27207 = n2652 ^ n476 ^ 1'b0 ;
  assign n27208 = ( n1650 & n6461 ) | ( n1650 & n27207 ) | ( n6461 & n27207 ) ;
  assign n27209 = n2837 & n27208 ;
  assign n27210 = n27209 ^ n15847 ^ 1'b0 ;
  assign n27211 = n16994 ^ n7287 ^ 1'b0 ;
  assign n27212 = n2274 & n2561 ;
  assign n27213 = n27211 | n27212 ;
  assign n27214 = n11543 | n12991 ;
  assign n27215 = n27214 ^ n946 ^ 1'b0 ;
  assign n27216 = n2243 & ~n27215 ;
  assign n27217 = n4824 ^ n2955 ^ 1'b0 ;
  assign n27218 = n2947 & ~n27217 ;
  assign n27219 = n8065 & n27218 ;
  assign n27220 = ~x43 & n15396 ;
  assign n27221 = n27220 ^ n15048 ^ 1'b0 ;
  assign n27222 = ~n3119 & n4723 ;
  assign n27223 = n27222 ^ n8087 ^ 1'b0 ;
  assign n27224 = n8935 | n27223 ;
  assign n27225 = n1488 & n13776 ;
  assign n27226 = ~n20657 & n27225 ;
  assign n27227 = x61 | n14589 ;
  assign n27228 = n2539 | n27227 ;
  assign n27229 = n528 ^ x25 ^ 1'b0 ;
  assign n27230 = n22396 ^ n16465 ^ 1'b0 ;
  assign n27231 = n10199 ^ n10010 ^ 1'b0 ;
  assign n27232 = n14508 & ~n27231 ;
  assign n27233 = n14541 | n21421 ;
  assign n27242 = n17050 ^ n9801 ^ 1'b0 ;
  assign n27234 = n22424 ^ n16744 ^ 1'b0 ;
  assign n27236 = n1775 & ~n12087 ;
  assign n27235 = n7608 & n14805 ;
  assign n27237 = n27236 ^ n27235 ^ 1'b0 ;
  assign n27238 = ( ~n5110 & n27234 ) | ( ~n5110 & n27237 ) | ( n27234 & n27237 ) ;
  assign n27239 = n13269 ^ n4827 ^ 1'b0 ;
  assign n27240 = n1361 & n27239 ;
  assign n27241 = n27238 | n27240 ;
  assign n27243 = n27242 ^ n27241 ^ n22177 ;
  assign n27244 = n2411 & n7133 ;
  assign n27245 = n22562 & ~n27244 ;
  assign n27246 = n2837 & ~n7446 ;
  assign n27247 = n16645 | n27246 ;
  assign n27248 = ~n414 & n25193 ;
  assign n27249 = n21026 & n27248 ;
  assign n27250 = n27249 ^ n6001 ^ 1'b0 ;
  assign n27251 = ~n13322 & n27250 ;
  assign n27252 = n27212 ^ n1618 ^ 1'b0 ;
  assign n27253 = n14803 & n27252 ;
  assign n27254 = n6343 & n27253 ;
  assign n27255 = n5176 & n10333 ;
  assign n27256 = n15930 ^ n4575 ^ 1'b0 ;
  assign n27257 = n13787 & n27256 ;
  assign n27258 = n22794 & n27257 ;
  assign n27259 = n27255 & n27258 ;
  assign n27260 = n8456 ^ n4473 ^ 1'b0 ;
  assign n27261 = n7175 & ~n27260 ;
  assign n27262 = n2589 & n11574 ;
  assign n27263 = n27261 & n27262 ;
  assign n27264 = n2487 & n27263 ;
  assign n27265 = ~n6075 & n17590 ;
  assign n27266 = n18737 & n27265 ;
  assign n27267 = n417 | n3125 ;
  assign n27268 = n5991 ^ n2463 ^ 1'b0 ;
  assign n27269 = n6008 & ~n14825 ;
  assign n27270 = n2219 & ~n14891 ;
  assign n27271 = n532 | n27270 ;
  assign n27272 = x72 & ~n27271 ;
  assign n27273 = ~n16579 & n27272 ;
  assign n27274 = n2145 | n20882 ;
  assign n27275 = n6805 | n8837 ;
  assign n27276 = n27275 ^ n4834 ^ 1'b0 ;
  assign n27277 = n7683 ^ n5571 ^ 1'b0 ;
  assign n27278 = n9731 & n27277 ;
  assign n27279 = n27278 ^ n2153 ^ 1'b0 ;
  assign n27280 = n12230 & n27279 ;
  assign n27281 = ~n4417 & n4521 ;
  assign n27282 = n6950 & ~n27281 ;
  assign n27283 = n6229 & n6342 ;
  assign n27284 = n27283 ^ x130 ^ 1'b0 ;
  assign n27285 = n27282 & ~n27284 ;
  assign n27286 = n13000 ^ n1137 ^ 1'b0 ;
  assign n27287 = n27286 ^ n13515 ^ 1'b0 ;
  assign n27288 = n6635 & ~n13892 ;
  assign n27289 = n472 | n20770 ;
  assign n27290 = n27288 & n27289 ;
  assign n27291 = n13054 & ~n22825 ;
  assign n27295 = n3950 & n12798 ;
  assign n27296 = n6662 | n27295 ;
  assign n27297 = n27296 ^ n21074 ^ n10138 ;
  assign n27292 = n17586 ^ n11272 ^ 1'b0 ;
  assign n27293 = n19024 & ~n27292 ;
  assign n27294 = ~n1449 & n27293 ;
  assign n27298 = n27297 ^ n27294 ^ 1'b0 ;
  assign n27299 = x14 & n22793 ;
  assign n27300 = n8493 & n8968 ;
  assign n27301 = n27300 ^ n7984 ^ 1'b0 ;
  assign n27302 = n6278 | n27301 ;
  assign n27303 = n20869 & ~n21191 ;
  assign n27304 = ( n6207 & n13541 ) | ( n6207 & ~n17192 ) | ( n13541 & ~n17192 ) ;
  assign n27305 = n747 & n8072 ;
  assign n27306 = n27305 ^ n8028 ^ 1'b0 ;
  assign n27307 = n14294 & ~n27306 ;
  assign n27308 = n399 & n5730 ;
  assign n27309 = n27308 ^ n22801 ^ 1'b0 ;
  assign n27310 = n27309 ^ n7737 ^ n6149 ;
  assign n27311 = ~n4408 & n27310 ;
  assign n27314 = ~n1234 & n2319 ;
  assign n27315 = n27314 ^ n22746 ^ 1'b0 ;
  assign n27316 = n27315 ^ n17519 ^ n7416 ;
  assign n27317 = n27316 ^ n532 ^ 1'b0 ;
  assign n27312 = n5242 & ~n17741 ;
  assign n27313 = n19181 & ~n27312 ;
  assign n27318 = n27317 ^ n27313 ^ 1'b0 ;
  assign n27319 = ~n11866 & n23125 ;
  assign n27320 = n27319 ^ n11159 ^ 1'b0 ;
  assign n27321 = n27320 ^ n6721 ^ 1'b0 ;
  assign n27322 = n25296 & n27321 ;
  assign n27323 = ~n13027 & n27322 ;
  assign n27326 = n12419 & n17690 ;
  assign n27324 = n17384 ^ n13938 ^ 1'b0 ;
  assign n27325 = n3032 & n27324 ;
  assign n27327 = n27326 ^ n27325 ^ 1'b0 ;
  assign n27328 = n16731 & ~n25135 ;
  assign n27329 = n23333 ^ n2006 ^ 1'b0 ;
  assign n27330 = n24722 | n27329 ;
  assign n27331 = n2644 & ~n13980 ;
  assign n27332 = n2120 | n17232 ;
  assign n27333 = ~n2689 & n27332 ;
  assign n27334 = ~n27331 & n27333 ;
  assign n27335 = ~n2011 & n16719 ;
  assign n27336 = n27335 ^ n11105 ^ 1'b0 ;
  assign n27337 = n1356 | n27336 ;
  assign n27338 = n5136 | n9121 ;
  assign n27339 = n2306 & ~n27338 ;
  assign n27340 = n27339 ^ n19771 ^ n4024 ;
  assign n27341 = n27340 ^ n1648 ^ 1'b0 ;
  assign n27342 = ~x203 & n26943 ;
  assign n27343 = n27342 ^ n15388 ^ 1'b0 ;
  assign n27344 = n27341 & n27343 ;
  assign n27345 = n2314 & n6089 ;
  assign n27346 = n25139 & n27345 ;
  assign n27347 = n13965 ^ n4122 ^ 1'b0 ;
  assign n27348 = n7890 & n18232 ;
  assign n27349 = n2277 & ~n7640 ;
  assign n27350 = n20437 & n27349 ;
  assign n27351 = n6341 ^ n4641 ^ 1'b0 ;
  assign n27352 = n27351 ^ n12046 ^ 1'b0 ;
  assign n27353 = n27350 & ~n27352 ;
  assign n27354 = n17188 ^ n5897 ^ 1'b0 ;
  assign n27355 = n21302 & ~n27354 ;
  assign n27356 = ~n824 & n4643 ;
  assign n27357 = n27356 ^ n436 ^ 1'b0 ;
  assign n27358 = n5965 & ~n14226 ;
  assign n27359 = n27357 & ~n27358 ;
  assign n27360 = x97 & n2891 ;
  assign n27361 = n7124 | n18900 ;
  assign n27362 = n27361 ^ n13932 ^ 1'b0 ;
  assign n27363 = n474 | n749 ;
  assign n27364 = n27362 | n27363 ;
  assign n27365 = n11747 & n27364 ;
  assign n27366 = n9807 ^ n4099 ^ 1'b0 ;
  assign n27367 = n3630 & n27366 ;
  assign n27368 = n27367 ^ n12656 ^ 1'b0 ;
  assign n27369 = n1212 | n1769 ;
  assign n27370 = n543 & ~n27369 ;
  assign n27371 = n12971 & ~n27370 ;
  assign n27372 = ~n7667 & n27371 ;
  assign n27373 = n7824 ^ n2929 ^ 1'b0 ;
  assign n27374 = n926 & ~n27373 ;
  assign n27375 = n27374 ^ n24413 ^ 1'b0 ;
  assign n27376 = n20437 ^ n2728 ^ 1'b0 ;
  assign n27377 = n21447 & n27376 ;
  assign n27378 = ~n8048 & n8854 ;
  assign n27379 = ~n2180 & n27378 ;
  assign n27380 = n1038 & n27379 ;
  assign n27381 = n1514 & ~n4813 ;
  assign n27382 = ~n6250 & n27381 ;
  assign n27383 = n15752 & ~n27382 ;
  assign n27384 = ~n26362 & n27383 ;
  assign n27385 = n27384 ^ n8326 ^ 1'b0 ;
  assign n27386 = ~n4709 & n27385 ;
  assign n27387 = n9114 ^ n3229 ^ 1'b0 ;
  assign n27388 = n577 | n27387 ;
  assign n27389 = n27388 ^ n14173 ^ 1'b0 ;
  assign n27390 = n25919 ^ n7880 ^ 1'b0 ;
  assign n27391 = ~n3924 & n14981 ;
  assign n27392 = n20723 & n27391 ;
  assign n27393 = n23385 & n27392 ;
  assign n27394 = ~n9585 & n27393 ;
  assign n27395 = n27394 ^ n14696 ^ 1'b0 ;
  assign n27396 = ~n5857 & n6045 ;
  assign n27397 = n27396 ^ n6500 ^ 1'b0 ;
  assign n27398 = ~x54 & n5047 ;
  assign n27399 = n27398 ^ n15853 ^ 1'b0 ;
  assign n27400 = n19727 ^ n9193 ^ 1'b0 ;
  assign n27401 = n3872 | n15225 ;
  assign n27402 = n20715 ^ n6297 ^ 1'b0 ;
  assign n27403 = n13036 & n25265 ;
  assign n27404 = n27403 ^ n12527 ^ 1'b0 ;
  assign n27405 = n7140 & ~n9062 ;
  assign n27406 = n5056 ^ n2242 ^ 1'b0 ;
  assign n27407 = n298 | n411 ;
  assign n27408 = n27407 ^ n22094 ^ 1'b0 ;
  assign n27409 = n2478 & n27408 ;
  assign n27411 = n2827 & ~n4720 ;
  assign n27410 = n7252 & ~n8214 ;
  assign n27412 = n27411 ^ n27410 ^ 1'b0 ;
  assign n27413 = n13580 | n27412 ;
  assign n27414 = n642 & ~n9530 ;
  assign n27415 = n27414 ^ n15440 ^ 1'b0 ;
  assign n27416 = n1605 | n27415 ;
  assign n27417 = n12250 ^ n11439 ^ 1'b0 ;
  assign n27418 = ~n468 & n9205 ;
  assign n27419 = n27418 ^ n10019 ^ 1'b0 ;
  assign n27420 = n4788 & n11572 ;
  assign n27421 = ~n27419 & n27420 ;
  assign n27422 = ~n3568 & n5192 ;
  assign n27423 = ~n23853 & n27422 ;
  assign n27424 = n25933 ^ n23335 ^ n5535 ;
  assign n27425 = n1651 & n21974 ;
  assign n27426 = ~n1810 & n27425 ;
  assign n27427 = x200 & n27426 ;
  assign n27428 = n10829 & n27427 ;
  assign n27429 = n17007 & n26023 ;
  assign n27430 = ~n8223 & n27429 ;
  assign n27431 = n1969 & n12753 ;
  assign n27432 = n27431 ^ n4631 ^ 1'b0 ;
  assign n27433 = n13215 & ~n27432 ;
  assign n27434 = n23627 | n27433 ;
  assign n27435 = n27434 ^ n1784 ^ 1'b0 ;
  assign n27436 = n14700 ^ n8202 ^ 1'b0 ;
  assign n27437 = ~n27435 & n27436 ;
  assign n27438 = ~n2575 & n17580 ;
  assign n27439 = n27438 ^ n320 ^ 1'b0 ;
  assign n27440 = n16472 ^ n8352 ^ 1'b0 ;
  assign n27441 = n27290 ^ x218 ^ 1'b0 ;
  assign n27442 = n27440 | n27441 ;
  assign n27443 = n10272 & ~n13121 ;
  assign n27444 = n10750 & n27443 ;
  assign n27445 = n27444 ^ n11157 ^ 1'b0 ;
  assign n27446 = ~n3505 & n27445 ;
  assign n27447 = n9954 & n27446 ;
  assign n27448 = n27447 ^ n7461 ^ 1'b0 ;
  assign n27449 = n18271 ^ n13633 ^ n1521 ;
  assign n27450 = ~n3676 & n27449 ;
  assign n27451 = n21121 & n27450 ;
  assign n27452 = n1126 & ~n15678 ;
  assign n27453 = n26286 ^ n22700 ^ n11736 ;
  assign n27454 = n14765 ^ n1217 ^ 1'b0 ;
  assign n27455 = n26084 & ~n27454 ;
  assign n27456 = n8628 | n23254 ;
  assign n27457 = n12894 | n27456 ;
  assign n27458 = n10643 & ~n13978 ;
  assign n27459 = n5372 & n27458 ;
  assign n27461 = ~n2914 & n11891 ;
  assign n27462 = ~n4246 & n27461 ;
  assign n27460 = n1596 | n5809 ;
  assign n27463 = n27462 ^ n27460 ^ 1'b0 ;
  assign n27464 = n27463 ^ n17112 ^ 1'b0 ;
  assign n27465 = n9022 | n18540 ;
  assign n27466 = ~n24348 & n25828 ;
  assign n27467 = n3817 & n15206 ;
  assign n27470 = n9400 ^ n1646 ^ 1'b0 ;
  assign n27468 = n7768 | n9923 ;
  assign n27469 = n27468 ^ n5447 ^ 1'b0 ;
  assign n27471 = n27470 ^ n27469 ^ 1'b0 ;
  assign n27472 = x232 & n3073 ;
  assign n27473 = n27472 ^ n18671 ^ 1'b0 ;
  assign n27474 = n10800 & n14061 ;
  assign n27475 = n10097 ^ n7708 ^ 1'b0 ;
  assign n27476 = n11481 & ~n27475 ;
  assign n27477 = ~n1704 & n27476 ;
  assign n27478 = n26376 ^ n14349 ^ 1'b0 ;
  assign n27479 = n19455 ^ n8646 ^ 1'b0 ;
  assign n27480 = n12515 ^ n1328 ^ 1'b0 ;
  assign n27481 = n17526 | n25431 ;
  assign n27482 = n25617 | n27481 ;
  assign n27483 = n3376 & n6893 ;
  assign n27484 = n27483 ^ n23273 ^ n13502 ;
  assign n27485 = n6762 ^ n4124 ^ 1'b0 ;
  assign n27486 = n12625 | n22099 ;
  assign n27487 = n1696 & ~n27486 ;
  assign n27488 = n16083 ^ n5861 ^ 1'b0 ;
  assign n27489 = ~n4617 & n11235 ;
  assign n27490 = n4119 ^ n566 ^ 1'b0 ;
  assign n27491 = ~n27489 & n27490 ;
  assign n27492 = x110 & n15019 ;
  assign n27493 = ~n4664 & n9177 ;
  assign n27494 = n13369 & ~n20165 ;
  assign n27495 = ~n8912 & n16234 ;
  assign n27496 = n27495 ^ n6891 ^ 1'b0 ;
  assign n27497 = n23254 ^ n8479 ^ 1'b0 ;
  assign n27498 = n5269 & ~n6572 ;
  assign n27499 = n7690 ^ n1085 ^ 1'b0 ;
  assign n27500 = n3635 & ~n17812 ;
  assign n27501 = n2180 | n18388 ;
  assign n27502 = n7415 & ~n18590 ;
  assign n27503 = n19696 | n27502 ;
  assign n27504 = ~n2750 & n27503 ;
  assign n27505 = n19349 ^ n7743 ^ n2279 ;
  assign n27506 = n11231 & n15019 ;
  assign n27507 = n4005 | n6531 ;
  assign n27508 = n10935 & ~n27507 ;
  assign n27509 = n4848 ^ n4484 ^ 1'b0 ;
  assign n27510 = n27509 ^ n24122 ^ 1'b0 ;
  assign n27511 = n27510 ^ n8111 ^ 1'b0 ;
  assign n27512 = n5105 | n18833 ;
  assign n27513 = ~n4747 & n23252 ;
  assign n27514 = n11705 ^ n11578 ^ n1286 ;
  assign n27515 = n4026 & ~n6895 ;
  assign n27516 = n2961 & ~n27515 ;
  assign n27517 = n27516 ^ n19622 ^ 1'b0 ;
  assign n27518 = ~n2038 & n21328 ;
  assign n27519 = n26722 & n27518 ;
  assign n27520 = n9340 & n12543 ;
  assign n27521 = ~n10051 & n27520 ;
  assign n27522 = x234 & n27521 ;
  assign n27523 = n27522 ^ n22766 ^ 1'b0 ;
  assign n27524 = n14654 ^ n8095 ^ 1'b0 ;
  assign n27525 = n966 & n23207 ;
  assign n27526 = n27524 & n27525 ;
  assign n27527 = n14895 & n22092 ;
  assign n27528 = n9606 & ~n11224 ;
  assign n27529 = n27528 ^ n1751 ^ 1'b0 ;
  assign n27530 = n7132 & ~n21435 ;
  assign n27531 = n24342 | n27530 ;
  assign n27532 = ~n9092 & n13780 ;
  assign n27533 = ~n3676 & n12425 ;
  assign n27534 = n1661 & n25837 ;
  assign n27535 = ~n13725 & n27497 ;
  assign n27536 = ~n14981 & n27535 ;
  assign n27537 = n3257 & n9495 ;
  assign n27538 = n27537 ^ n9923 ^ 1'b0 ;
  assign n27539 = n8893 & n27538 ;
  assign n27540 = n27539 ^ n11711 ^ 1'b0 ;
  assign n27541 = n5300 | n11565 ;
  assign n27542 = n27541 ^ n24666 ^ 1'b0 ;
  assign n27543 = n27542 ^ n6571 ^ 1'b0 ;
  assign n27544 = n2421 & ~n27543 ;
  assign n27545 = n19821 ^ n15350 ^ 1'b0 ;
  assign n27546 = ~n24778 & n25223 ;
  assign n27547 = ~n25998 & n26334 ;
  assign n27548 = ( n9598 & n14323 ) | ( n9598 & ~n17126 ) | ( n14323 & ~n17126 ) ;
  assign n27549 = ~n6009 & n27548 ;
  assign n27550 = n15131 ^ n841 ^ 1'b0 ;
  assign n27551 = n27549 & n27550 ;
  assign n27552 = ~n3796 & n5806 ;
  assign n27553 = n27552 ^ n17757 ^ 1'b0 ;
  assign n27554 = n22713 ^ x160 ^ 1'b0 ;
  assign n27555 = n25404 & ~n27554 ;
  assign n27556 = ~n13553 & n19304 ;
  assign n27557 = n1485 & n17380 ;
  assign n27558 = ~n17286 & n27557 ;
  assign n27559 = n26091 ^ n19753 ^ 1'b0 ;
  assign n27560 = ~n7083 & n26871 ;
  assign n27561 = n1514 & n3745 ;
  assign n27562 = n19682 & ~n27561 ;
  assign n27563 = n21595 ^ n10996 ^ 1'b0 ;
  assign n27564 = n3501 | n27563 ;
  assign n27565 = n1926 | n27564 ;
  assign n27566 = n2685 | n27565 ;
  assign n27567 = n4769 & n18443 ;
  assign n27568 = ~n27566 & n27567 ;
  assign n27569 = n22268 ^ n19719 ^ 1'b0 ;
  assign n27570 = n4385 | n15106 ;
  assign n27571 = ~n7720 & n27570 ;
  assign n27572 = n7017 & n24523 ;
  assign n27573 = ~n16734 & n27572 ;
  assign n27574 = n1352 | n27573 ;
  assign n27575 = n27574 ^ n12182 ^ 1'b0 ;
  assign n27576 = n12789 ^ n3657 ^ 1'b0 ;
  assign n27577 = ( ~n9985 & n14335 ) | ( ~n9985 & n27576 ) | ( n14335 & n27576 ) ;
  assign n27578 = n2712 & n7440 ;
  assign n27579 = n388 ^ n298 ^ 1'b0 ;
  assign n27580 = ~n12242 & n27579 ;
  assign n27581 = n3392 | n5597 ;
  assign n27582 = ~n10438 & n27581 ;
  assign n27583 = ( ~n3819 & n22450 ) | ( ~n3819 & n27582 ) | ( n22450 & n27582 ) ;
  assign n27584 = ~n11982 & n27583 ;
  assign n27585 = n27207 ^ n288 ^ 1'b0 ;
  assign n27586 = n23132 & n27585 ;
  assign n27587 = n3532 | n14507 ;
  assign n27588 = n3089 | n27587 ;
  assign n27589 = n13155 & n17743 ;
  assign n27590 = n27175 & ~n27589 ;
  assign n27591 = n16322 ^ n12882 ^ 1'b0 ;
  assign n27592 = n12020 | n27591 ;
  assign n27593 = n13514 | n27592 ;
  assign n27594 = n3926 | n9972 ;
  assign n27595 = n23729 | n24470 ;
  assign n27596 = n13740 ^ n1742 ^ 1'b0 ;
  assign n27597 = ~n5485 & n27596 ;
  assign n27598 = ~x47 & n27597 ;
  assign n27599 = n19176 ^ n979 ^ 1'b0 ;
  assign n27600 = ~n15215 & n27599 ;
  assign n27601 = n4789 & ~n27600 ;
  assign n27602 = n18717 ^ n10986 ^ n2271 ;
  assign n27603 = x248 & ~n12235 ;
  assign n27604 = n4499 | n27603 ;
  assign n27605 = x60 & ~n27604 ;
  assign n27606 = n27605 ^ n2582 ^ 1'b0 ;
  assign n27607 = n3798 ^ n1507 ^ 1'b0 ;
  assign n27608 = ~n3379 & n16493 ;
  assign n27609 = n7120 & n24322 ;
  assign n27610 = n26809 & n27609 ;
  assign n27611 = n1379 & n4545 ;
  assign n27612 = n19017 & n25316 ;
  assign n27613 = n2432 | n24173 ;
  assign n27614 = n3745 | n27613 ;
  assign n27615 = x44 & n6031 ;
  assign n27616 = n9428 & ~n27615 ;
  assign n27617 = n27616 ^ n3006 ^ 1'b0 ;
  assign n27618 = n11574 & n13400 ;
  assign n27619 = n27618 ^ n18066 ^ 1'b0 ;
  assign n27620 = n27617 & n27619 ;
  assign n27621 = ~n27614 & n27620 ;
  assign n27622 = n18268 ^ n2770 ^ 1'b0 ;
  assign n27623 = ~n27621 & n27622 ;
  assign n27624 = n14694 ^ n14605 ^ 1'b0 ;
  assign n27625 = n1035 & n27624 ;
  assign n27626 = n21221 & n27625 ;
  assign n27627 = n13927 & n15248 ;
  assign n27628 = ~n780 & n2885 ;
  assign n27629 = n27628 ^ x231 ^ 1'b0 ;
  assign n27630 = n27627 & n27629 ;
  assign n27631 = n4027 & ~n14451 ;
  assign n27632 = n27631 ^ n8733 ^ 1'b0 ;
  assign n27633 = n19821 | n27632 ;
  assign n27634 = ~n6205 & n18400 ;
  assign n27635 = n2555 | n15142 ;
  assign n27636 = n23737 & ~n27635 ;
  assign n27637 = n14045 & n27636 ;
  assign n27640 = ~n798 & n4170 ;
  assign n27638 = n10815 ^ n4720 ^ 1'b0 ;
  assign n27639 = n9834 & n27638 ;
  assign n27641 = n27640 ^ n27639 ^ 1'b0 ;
  assign n27642 = n19334 ^ n17523 ^ n5394 ;
  assign n27643 = n20319 ^ n18505 ^ 1'b0 ;
  assign n27644 = n27643 ^ n8261 ^ 1'b0 ;
  assign n27645 = ~n15469 & n27644 ;
  assign n27646 = ~n2232 & n27645 ;
  assign n27647 = n27646 ^ n21297 ^ 1'b0 ;
  assign n27648 = n9589 ^ n2671 ^ 1'b0 ;
  assign n27649 = ~n9416 & n27648 ;
  assign n27650 = ~n14506 & n25712 ;
  assign n27651 = n1423 & n16269 ;
  assign n27652 = n23802 & n27651 ;
  assign n27653 = n5525 & ~n27652 ;
  assign n27654 = n465 & ~n2909 ;
  assign n27655 = n27654 ^ n7151 ^ 1'b0 ;
  assign n27656 = ~n4804 & n27655 ;
  assign n27657 = n13671 ^ n8480 ^ 1'b0 ;
  assign n27658 = n3481 & ~n4857 ;
  assign n27659 = n9690 | n27658 ;
  assign n27660 = n27659 ^ n22292 ^ 1'b0 ;
  assign n27661 = n27660 ^ n3373 ^ 1'b0 ;
  assign n27662 = n2543 & n17841 ;
  assign n27663 = n13073 & ~n27662 ;
  assign n27664 = n17214 ^ n1365 ^ 1'b0 ;
  assign n27665 = n14937 ^ n3940 ^ 1'b0 ;
  assign n27666 = n27665 ^ n12848 ^ 1'b0 ;
  assign n27667 = n1192 | n13206 ;
  assign n27668 = ~n9493 & n9503 ;
  assign n27669 = ~n27667 & n27668 ;
  assign n27670 = ~n27666 & n27669 ;
  assign n27671 = n1045 & ~n11509 ;
  assign n27672 = n27671 ^ n16481 ^ 1'b0 ;
  assign n27673 = n1692 & n2766 ;
  assign n27674 = n2586 ^ n1195 ^ 1'b0 ;
  assign n27675 = n5176 & n27674 ;
  assign n27676 = ~n27673 & n27675 ;
  assign n27677 = ~n283 & n3850 ;
  assign n27678 = n27677 ^ n6169 ^ 1'b0 ;
  assign n27679 = n21063 ^ n1188 ^ 1'b0 ;
  assign n27680 = n15556 ^ n7777 ^ 1'b0 ;
  assign n27681 = n7507 | n27680 ;
  assign n27682 = n27681 ^ n14803 ^ 1'b0 ;
  assign n27683 = x122 ^ x11 ^ 1'b0 ;
  assign n27684 = n4540 ^ n3578 ^ 1'b0 ;
  assign n27685 = ~n27683 & n27684 ;
  assign n27686 = n298 & n3397 ;
  assign n27687 = n3559 & ~n4948 ;
  assign n27688 = n6553 & n27687 ;
  assign n27689 = n13922 & n15201 ;
  assign n27690 = ~n21483 & n27544 ;
  assign n27691 = n3146 & n27690 ;
  assign n27692 = ~n4128 & n17030 ;
  assign n27693 = ~n19101 & n27692 ;
  assign n27694 = n26306 ^ n14386 ^ 1'b0 ;
  assign n27695 = n27694 ^ n13267 ^ 1'b0 ;
  assign n27696 = ~n8719 & n27695 ;
  assign n27697 = n10540 ^ n414 ^ 1'b0 ;
  assign n27698 = n15587 | n27697 ;
  assign n27699 = n27698 ^ n23914 ^ 1'b0 ;
  assign n27700 = n1651 | n14993 ;
  assign n27701 = n866 & n4258 ;
  assign n27702 = n27701 ^ n5907 ^ 1'b0 ;
  assign n27703 = n9598 & ~n12862 ;
  assign n27704 = n27703 ^ n1112 ^ 1'b0 ;
  assign n27705 = ~n1366 & n6273 ;
  assign n27706 = n27705 ^ n16015 ^ 1'b0 ;
  assign n27707 = n21495 | n27706 ;
  assign n27708 = n18846 | n19172 ;
  assign n27709 = n27708 ^ n14501 ^ 1'b0 ;
  assign n27710 = n7695 ^ n7463 ^ 1'b0 ;
  assign n27711 = n27710 ^ n23335 ^ n8725 ;
  assign n27712 = ~n3230 & n6931 ;
  assign n27713 = n11803 ^ n3637 ^ 1'b0 ;
  assign n27714 = n6060 & ~n27713 ;
  assign n27715 = n27714 ^ n7902 ^ 1'b0 ;
  assign n27716 = n4225 | n27715 ;
  assign n27717 = n18355 ^ n16015 ^ 1'b0 ;
  assign n27718 = n27717 ^ n17774 ^ 1'b0 ;
  assign n27719 = n24374 ^ n22220 ^ 1'b0 ;
  assign n27720 = n2042 & ~n27719 ;
  assign n27721 = n26361 ^ n1273 ^ 1'b0 ;
  assign n27722 = n11810 & n27721 ;
  assign n27723 = n11136 ^ n2393 ^ 1'b0 ;
  assign n27724 = n10689 ^ n4819 ^ 1'b0 ;
  assign n27725 = n4040 & ~n27724 ;
  assign n27726 = n1787 & ~n10292 ;
  assign n27727 = n10205 ^ n2883 ^ 1'b0 ;
  assign n27729 = n5500 ^ n4605 ^ 1'b0 ;
  assign n27728 = ~n12616 & n21064 ;
  assign n27730 = n27729 ^ n27728 ^ 1'b0 ;
  assign n27731 = n19800 & ~n20275 ;
  assign n27732 = n27731 ^ n6110 ^ 1'b0 ;
  assign n27733 = n7684 | n10507 ;
  assign n27734 = n4940 ^ n1177 ^ 1'b0 ;
  assign n27735 = n2179 | n27734 ;
  assign n27736 = n809 & ~n21715 ;
  assign n27737 = n2221 & ~n6950 ;
  assign n27738 = n27737 ^ n16879 ^ 1'b0 ;
  assign n27739 = n19021 & n22380 ;
  assign n27740 = ~n18067 & n27739 ;
  assign n27741 = n3687 | n27740 ;
  assign n27742 = n14349 | n17464 ;
  assign n27743 = n27742 ^ n15949 ^ 1'b0 ;
  assign n27744 = n5587 | n10785 ;
  assign n27745 = n3316 ^ n445 ^ 1'b0 ;
  assign n27746 = n27744 & n27745 ;
  assign n27747 = n1573 & ~n3213 ;
  assign n27748 = n15477 | n18932 ;
  assign n27749 = n1397 & ~n26293 ;
  assign n27750 = ~n22035 & n27749 ;
  assign n27751 = n23040 ^ n16000 ^ n11209 ;
  assign n27752 = n19370 ^ n5034 ^ 1'b0 ;
  assign n27753 = n27751 & ~n27752 ;
  assign n27754 = n16439 ^ n7144 ^ 1'b0 ;
  assign n27755 = n9087 & ~n13077 ;
  assign n27756 = n27755 ^ n2853 ^ 1'b0 ;
  assign n27757 = ( ~n13054 & n27754 ) | ( ~n13054 & n27756 ) | ( n27754 & n27756 ) ;
  assign n27758 = ( n1653 & n6010 ) | ( n1653 & n8960 ) | ( n6010 & n8960 ) ;
  assign n27763 = n2055 | n2441 ;
  assign n27764 = n27763 ^ n10306 ^ 1'b0 ;
  assign n27765 = ~n17785 & n27764 ;
  assign n27766 = ~x83 & n27765 ;
  assign n27759 = n5207 | n6012 ;
  assign n27760 = n27759 ^ n5682 ^ 1'b0 ;
  assign n27761 = n24694 & ~n27760 ;
  assign n27762 = n5476 | n27761 ;
  assign n27767 = n27766 ^ n27762 ^ 1'b0 ;
  assign n27768 = n5507 ^ n605 ^ 1'b0 ;
  assign n27769 = n12432 & n27768 ;
  assign n27770 = n7687 | n9717 ;
  assign n27771 = n27770 ^ n19176 ^ 1'b0 ;
  assign n27772 = ~n7019 & n16156 ;
  assign n27773 = n5328 | n9092 ;
  assign n27774 = n27773 ^ n275 ^ 1'b0 ;
  assign n27775 = n15531 | n27774 ;
  assign n27776 = n3961 | n7474 ;
  assign n27777 = n2239 & n27776 ;
  assign n27778 = n27777 ^ n15681 ^ 1'b0 ;
  assign n27779 = n502 & n19592 ;
  assign n27780 = n15168 & n23457 ;
  assign n27781 = n27780 ^ n17851 ^ 1'b0 ;
  assign n27782 = n8531 & ~n18016 ;
  assign n27783 = n5136 ^ n608 ^ 1'b0 ;
  assign n27784 = ~n18504 & n27783 ;
  assign n27785 = ~n8686 & n27784 ;
  assign n27786 = n10241 & ~n24208 ;
  assign n27787 = n10458 & n27786 ;
  assign n27788 = n12304 ^ n9880 ^ 1'b0 ;
  assign n27789 = ~n1991 & n27788 ;
  assign n27790 = n27789 ^ n7408 ^ 1'b0 ;
  assign n27791 = n12686 ^ n6008 ^ 1'b0 ;
  assign n27792 = n9323 & n27791 ;
  assign n27793 = n27792 ^ n12898 ^ 1'b0 ;
  assign n27794 = n27793 ^ n15681 ^ 1'b0 ;
  assign n27795 = n26778 ^ n23249 ^ 1'b0 ;
  assign n27798 = n5273 ^ n401 ^ 1'b0 ;
  assign n27799 = n1059 | n27798 ;
  assign n27796 = ~n9717 & n13570 ;
  assign n27797 = n27796 ^ n20515 ^ 1'b0 ;
  assign n27800 = n27799 ^ n27797 ^ n17383 ;
  assign n27802 = x136 & n2035 ;
  assign n27801 = n6326 & ~n8503 ;
  assign n27803 = n27802 ^ n27801 ^ 1'b0 ;
  assign n27804 = n15409 & n27803 ;
  assign n27805 = ~n20162 & n27804 ;
  assign n27806 = n2159 & n8384 ;
  assign n27807 = ~n6550 & n11672 ;
  assign n27808 = n27806 & n27807 ;
  assign n27809 = n6288 & n23975 ;
  assign n27810 = x42 | n14133 ;
  assign n27811 = n20121 ^ n2420 ^ 1'b0 ;
  assign n27812 = n7512 ^ n2316 ^ 1'b0 ;
  assign n27814 = n1154 & ~n1740 ;
  assign n27813 = n25578 | n27342 ;
  assign n27815 = n27814 ^ n27813 ^ 1'b0 ;
  assign n27816 = n11607 & n27815 ;
  assign n27817 = n3377 & ~n27816 ;
  assign n27818 = n5293 | n8281 ;
  assign n27819 = n27818 ^ n6766 ^ 1'b0 ;
  assign n27820 = ~n2725 & n19474 ;
  assign n27821 = n1580 | n2124 ;
  assign n27822 = n18377 ^ n18039 ^ 1'b0 ;
  assign n27823 = ~n10509 & n27822 ;
  assign n27824 = n744 & n3862 ;
  assign n27825 = n27824 ^ n3165 ^ 1'b0 ;
  assign n27826 = n27825 ^ n6986 ^ 1'b0 ;
  assign n27827 = n655 & ~n10608 ;
  assign n27828 = n22753 ^ n8686 ^ 1'b0 ;
  assign n27829 = n9081 & n19241 ;
  assign n27830 = n13619 & n27829 ;
  assign n27831 = n5525 | n26413 ;
  assign n27832 = ~n3473 & n14403 ;
  assign n27833 = n11771 & n27832 ;
  assign n27834 = n23767 & ~n27833 ;
  assign n27835 = n27834 ^ n9811 ^ 1'b0 ;
  assign n27836 = n1709 & n27835 ;
  assign n27837 = n9607 ^ n1772 ^ 1'b0 ;
  assign n27838 = n11131 & ~n27837 ;
  assign n27839 = n12438 & n27838 ;
  assign n27840 = n27839 ^ n6846 ^ 1'b0 ;
  assign n27841 = n7881 & ~n19325 ;
  assign n27842 = n23977 ^ n23933 ^ n9239 ;
  assign n27843 = n6054 & n21989 ;
  assign n27844 = ~n12185 & n27843 ;
  assign n27845 = ~n4459 & n16876 ;
  assign n27846 = n9484 | n27845 ;
  assign n27847 = n27812 ^ n25543 ^ 1'b0 ;
  assign n27848 = n4857 & n27847 ;
  assign n27849 = n4838 ^ n3855 ^ 1'b0 ;
  assign n27850 = n4688 & ~n27849 ;
  assign n27851 = n27850 ^ n26081 ^ n16697 ;
  assign n27852 = ~n3754 & n16798 ;
  assign n27853 = n18180 ^ n7671 ^ 1'b0 ;
  assign n27854 = ~n2785 & n27853 ;
  assign n27855 = n8146 & ~n12070 ;
  assign n27876 = n1841 & ~n15027 ;
  assign n27877 = n15027 & n27876 ;
  assign n27878 = x115 | n5956 ;
  assign n27879 = n27877 | n27878 ;
  assign n27880 = n14527 & ~n27879 ;
  assign n27881 = n9723 & n17658 ;
  assign n27882 = n14066 & n27881 ;
  assign n27883 = n8942 | n27882 ;
  assign n27884 = n27882 & ~n27883 ;
  assign n27885 = n27880 | n27884 ;
  assign n27886 = n27880 & ~n27885 ;
  assign n27869 = n10557 & ~n12496 ;
  assign n27856 = ~n1223 & n22443 ;
  assign n27857 = x50 & n27856 ;
  assign n27858 = n891 & n3123 ;
  assign n27859 = ~n891 & n27858 ;
  assign n27860 = n27857 & n27859 ;
  assign n27861 = x31 & ~n548 ;
  assign n27862 = n548 & n27861 ;
  assign n27863 = n1689 | n1753 ;
  assign n27864 = n27862 & ~n27863 ;
  assign n27865 = n5619 | n27864 ;
  assign n27866 = n27865 ^ n9503 ^ 1'b0 ;
  assign n27867 = n27860 & n27866 ;
  assign n27868 = n6401 & n27867 ;
  assign n27870 = n27869 ^ n27868 ^ 1'b0 ;
  assign n27871 = ~n8866 & n9547 ;
  assign n27872 = ~n27870 & n27871 ;
  assign n27873 = n16224 | n27872 ;
  assign n27874 = n27872 & ~n27873 ;
  assign n27875 = n18362 & ~n27874 ;
  assign n27887 = n27886 ^ n27875 ^ 1'b0 ;
  assign n27888 = ~n3298 & n21096 ;
  assign n27889 = n27888 ^ n3760 ^ 1'b0 ;
  assign n27890 = n7864 & n27889 ;
  assign n27891 = ~n20788 & n27890 ;
  assign n27892 = n16454 ^ n2406 ^ 1'b0 ;
  assign n27893 = ~n983 & n1048 ;
  assign n27894 = n10744 & n27893 ;
  assign n27895 = n27892 & ~n27894 ;
  assign n27896 = n10988 ^ n7508 ^ n6646 ;
  assign n27897 = ~n3509 & n27896 ;
  assign n27898 = n26152 ^ n21128 ^ 1'b0 ;
  assign n27899 = n10382 ^ n4151 ^ 1'b0 ;
  assign n27900 = n17276 | n18723 ;
  assign n27901 = ~n8212 & n12095 ;
  assign n27902 = n27901 ^ n7878 ^ 1'b0 ;
  assign n27904 = n8706 & ~n14830 ;
  assign n27903 = n9310 & ~n20419 ;
  assign n27905 = n27904 ^ n27903 ^ 1'b0 ;
  assign n27906 = ~n14767 & n27905 ;
  assign n27907 = n27902 & n27906 ;
  assign n27908 = n19531 ^ n788 ^ 1'b0 ;
  assign n27909 = ( n1139 & n15711 ) | ( n1139 & n27596 ) | ( n15711 & n27596 ) ;
  assign n27910 = n5233 & n12238 ;
  assign n27911 = n7968 & n9040 ;
  assign n27912 = n27911 ^ n6307 ^ 1'b0 ;
  assign n27913 = n17309 & ~n27912 ;
  assign n27914 = ~n17848 & n21751 ;
  assign n27915 = n13231 & ~n22460 ;
  assign n27916 = n18969 & n27915 ;
  assign n27917 = ~n18907 & n25449 ;
  assign n27918 = n3678 | n9819 ;
  assign n27919 = n27918 ^ n401 ^ 1'b0 ;
  assign n27920 = n13330 ^ n9327 ^ 1'b0 ;
  assign n27921 = n3503 | n6191 ;
  assign n27922 = n18565 & ~n27921 ;
  assign n27923 = ~n1562 & n14508 ;
  assign n27924 = n27923 ^ n22813 ^ 1'b0 ;
  assign n27925 = n18074 ^ n4785 ^ 1'b0 ;
  assign n27926 = ~n15674 & n27925 ;
  assign n27927 = n18341 ^ n7630 ^ 1'b0 ;
  assign n27928 = ~n18768 & n20621 ;
  assign n27929 = n11758 & ~n12713 ;
  assign n27930 = n27929 ^ n892 ^ 1'b0 ;
  assign n27931 = n16681 & n24079 ;
  assign n27932 = n3799 & n27931 ;
  assign n27933 = n14589 ^ n10160 ^ 1'b0 ;
  assign n27934 = n18241 & n27933 ;
  assign n27937 = n7567 ^ n6945 ^ 1'b0 ;
  assign n27935 = n4459 & ~n5717 ;
  assign n27936 = n7194 | n27935 ;
  assign n27938 = n27937 ^ n27936 ^ 1'b0 ;
  assign n27939 = n2747 & n21938 ;
  assign n27940 = ~n3678 & n8509 ;
  assign n27941 = n14859 & n27940 ;
  assign n27942 = n27941 ^ n16676 ^ 1'b0 ;
  assign n27943 = n12238 & n27942 ;
  assign n27944 = n16808 & n25514 ;
  assign n27945 = n6028 & ~n15057 ;
  assign n27946 = n13520 ^ n5552 ^ 1'b0 ;
  assign n27947 = n8448 & ~n27946 ;
  assign n27948 = ~n27945 & n27947 ;
  assign n27949 = n23610 ^ n345 ^ 1'b0 ;
  assign n27950 = ~n13619 & n27949 ;
  assign n27951 = ~n25433 & n27950 ;
  assign n27952 = n21801 & n27951 ;
  assign n27953 = n6617 ^ n5067 ^ 1'b0 ;
  assign n27954 = ~n6084 & n27953 ;
  assign n27955 = n19560 ^ n7601 ^ 1'b0 ;
  assign n27956 = ~n405 & n27955 ;
  assign n27957 = ( ~n11699 & n16520 ) | ( ~n11699 & n27956 ) | ( n16520 & n27956 ) ;
  assign n27958 = n10813 ^ n8165 ^ x61 ;
  assign n27959 = n27957 & ~n27958 ;
  assign n27960 = n4253 ^ n3162 ^ n2475 ;
  assign n27961 = n1152 & n8058 ;
  assign n27962 = n27961 ^ n6566 ^ 1'b0 ;
  assign n27963 = n27960 | n27962 ;
  assign n27964 = n27963 ^ n1696 ^ 1'b0 ;
  assign n27965 = n24471 & ~n27964 ;
  assign n27966 = n9898 | n15260 ;
  assign n27967 = n602 | n27966 ;
  assign n27968 = n805 | n5325 ;
  assign n27969 = n7190 | n27968 ;
  assign n27970 = ~n11327 & n25619 ;
  assign n27971 = ~n27969 & n27970 ;
  assign n27972 = n10813 ^ n5443 ^ 1'b0 ;
  assign n27973 = ~n3112 & n27972 ;
  assign n27974 = n1297 | n23855 ;
  assign n27975 = n602 & n13511 ;
  assign n27976 = n2629 & n27975 ;
  assign n27977 = ~n27974 & n27976 ;
  assign n27978 = n24472 ^ n18835 ^ n16712 ;
  assign n27979 = n6751 ^ n2047 ^ 1'b0 ;
  assign n27980 = n15363 & ~n27979 ;
  assign n27981 = n5411 & ~n24877 ;
  assign n27982 = ~n3929 & n27981 ;
  assign n27983 = n11857 ^ n631 ^ 1'b0 ;
  assign n27984 = n7833 & ~n27983 ;
  assign n27985 = x220 | n13763 ;
  assign n27986 = n4592 & n13603 ;
  assign n27987 = n3184 | n27986 ;
  assign n27988 = n27987 ^ n2660 ^ 1'b0 ;
  assign n27989 = n498 & n27988 ;
  assign n27990 = n9358 ^ n7132 ^ 1'b0 ;
  assign n27991 = n1738 & n18770 ;
  assign n27992 = n856 & n11864 ;
  assign n27993 = n5328 ^ n3694 ^ n3625 ;
  assign n27994 = n3796 & n14403 ;
  assign n27995 = n7671 | n27994 ;
  assign n27996 = n27995 ^ n24895 ^ 1'b0 ;
  assign n27997 = n8959 ^ n8890 ^ 1'b0 ;
  assign n27998 = n27997 ^ n8829 ^ 1'b0 ;
  assign n27999 = ~n3971 & n5343 ;
  assign n28000 = ~n17634 & n27999 ;
  assign n28001 = ~n6193 & n18904 ;
  assign n28002 = n7917 ^ n2744 ^ 1'b0 ;
  assign n28003 = ~n21188 & n28002 ;
  assign n28004 = n25456 ^ n9158 ^ 1'b0 ;
  assign n28005 = ~n13026 & n28004 ;
  assign n28006 = ( n1668 & n6967 ) | ( n1668 & ~n28005 ) | ( n6967 & ~n28005 ) ;
  assign n28008 = n1443 ^ x178 ^ 1'b0 ;
  assign n28009 = n28008 ^ n12521 ^ 1'b0 ;
  assign n28007 = ~n7384 & n27410 ;
  assign n28010 = n28009 ^ n28007 ^ 1'b0 ;
  assign n28011 = n1596 | n7510 ;
  assign n28012 = n28011 ^ n7997 ^ 1'b0 ;
  assign n28013 = ~n1339 & n8625 ;
  assign n28014 = n6191 & n28013 ;
  assign n28015 = ~n2402 & n9690 ;
  assign n28016 = ~n7813 & n12141 ;
  assign n28017 = n28016 ^ n12351 ^ 1'b0 ;
  assign n28018 = n1890 | n25814 ;
  assign n28019 = n10668 | n25034 ;
  assign n28020 = n22968 ^ n985 ^ 1'b0 ;
  assign n28021 = n28019 & n28020 ;
  assign n28022 = n15136 ^ n9495 ^ 1'b0 ;
  assign n28023 = ~n11612 & n28022 ;
  assign n28024 = ~n6489 & n28023 ;
  assign n28026 = n12765 ^ n7692 ^ 1'b0 ;
  assign n28025 = n5706 & ~n15783 ;
  assign n28027 = n28026 ^ n28025 ^ 1'b0 ;
  assign n28028 = ~n7175 & n17825 ;
  assign n28029 = n618 ^ x253 ^ 1'b0 ;
  assign n28030 = n3968 & ~n28029 ;
  assign n28031 = n283 | n27604 ;
  assign n28032 = n28030 | n28031 ;
  assign n28033 = n24088 ^ n19564 ^ 1'b0 ;
  assign n28034 = ~n9051 & n28033 ;
  assign n28035 = n320 & n28034 ;
  assign n28036 = ~n19533 & n20133 ;
  assign n28037 = n7133 & ~n28036 ;
  assign n28038 = n28037 ^ n5670 ^ 1'b0 ;
  assign n28039 = n16558 ^ n11892 ^ 1'b0 ;
  assign n28040 = n3239 & ~n28039 ;
  assign n28041 = n27444 & ~n28040 ;
  assign n28042 = n5929 | n13817 ;
  assign n28043 = n7718 | n28042 ;
  assign n28044 = ( ~n4271 & n14843 ) | ( ~n4271 & n28043 ) | ( n14843 & n28043 ) ;
  assign n28045 = n2611 | n3993 ;
  assign n28046 = n8132 ^ n1896 ^ 1'b0 ;
  assign n28047 = ~n17749 & n28046 ;
  assign n28048 = n18829 & n24337 ;
  assign n28049 = n1286 & n28048 ;
  assign n28050 = n486 | n3874 ;
  assign n28051 = n1613 & ~n28050 ;
  assign n28052 = ( n821 & ~n23074 ) | ( n821 & n28051 ) | ( ~n23074 & n28051 ) ;
  assign n28053 = x206 | n4133 ;
  assign n28054 = n28053 ^ n26150 ^ 1'b0 ;
  assign n28055 = n8137 ^ n3054 ^ 1'b0 ;
  assign n28056 = ~n11743 & n28055 ;
  assign n28057 = ~n2389 & n11472 ;
  assign n28058 = n28057 ^ n3578 ^ 1'b0 ;
  assign n28059 = n28056 & n28058 ;
  assign n28060 = n8258 ^ n6685 ^ 1'b0 ;
  assign n28061 = n18262 | n20569 ;
  assign n28062 = n28061 ^ n19722 ^ 1'b0 ;
  assign n28063 = n20158 ^ n3212 ^ 1'b0 ;
  assign n28064 = n26332 & n28063 ;
  assign n28065 = ~n2161 & n28064 ;
  assign n28066 = n13439 ^ n7192 ^ 1'b0 ;
  assign n28067 = n13064 & n21116 ;
  assign n28068 = n19864 ^ n3343 ^ 1'b0 ;
  assign n28069 = n3280 & n25343 ;
  assign n28070 = n4244 ^ n3630 ^ 1'b0 ;
  assign n28071 = n28070 ^ n14309 ^ 1'b0 ;
  assign n28072 = ~n12069 & n26179 ;
  assign n28073 = n28072 ^ n2938 ^ 1'b0 ;
  assign n28074 = n11456 & n28073 ;
  assign n28075 = n27643 ^ n17508 ^ 1'b0 ;
  assign n28076 = n3434 | n4147 ;
  assign n28077 = n18120 | n28076 ;
  assign n28078 = n4092 & n15630 ;
  assign n28079 = n4197 & n28078 ;
  assign n28080 = n1977 | n28079 ;
  assign n28081 = n28080 ^ n20900 ^ 1'b0 ;
  assign n28082 = x11 & x111 ;
  assign n28083 = n1429 & n28082 ;
  assign n28084 = n28083 ^ n15230 ^ 1'b0 ;
  assign n28085 = n9073 & n28084 ;
  assign n28086 = n22774 ^ n2336 ^ 1'b0 ;
  assign n28087 = n13164 ^ n3953 ^ 1'b0 ;
  assign n28088 = n18954 ^ n6413 ^ 1'b0 ;
  assign n28089 = n28087 & ~n28088 ;
  assign n28090 = n2486 & n28089 ;
  assign n28091 = n16422 & n28090 ;
  assign n28092 = n26456 ^ n6026 ^ 1'b0 ;
  assign n28093 = n6226 | n13245 ;
  assign n28094 = n6226 & ~n28093 ;
  assign n28095 = x133 & ~n2087 ;
  assign n28096 = n18173 & n19073 ;
  assign n28097 = ~n28095 & n28096 ;
  assign n28098 = n9438 & ~n28097 ;
  assign n28099 = n28094 & n28098 ;
  assign n28100 = n24949 | n28099 ;
  assign n28101 = n28099 & ~n28100 ;
  assign n28102 = x240 & n1301 ;
  assign n28103 = ~x240 & n28102 ;
  assign n28104 = n4903 & n28103 ;
  assign n28105 = n24094 & n28104 ;
  assign n28106 = ~n24094 & n28105 ;
  assign n28107 = n28106 ^ n8860 ^ 1'b0 ;
  assign n28108 = ~n28101 & n28107 ;
  assign n28109 = n18322 ^ n4068 ^ 1'b0 ;
  assign n28110 = n19044 & ~n26630 ;
  assign n28111 = n28110 ^ n10434 ^ 1'b0 ;
  assign n28112 = ~n2928 & n5574 ;
  assign n28113 = n3332 | n13842 ;
  assign n28114 = n28112 & ~n28113 ;
  assign n28115 = n12862 & n15910 ;
  assign n28116 = n11687 ^ n4108 ^ 1'b0 ;
  assign n28118 = n4208 | n13761 ;
  assign n28119 = n2495 & n5006 ;
  assign n28120 = n28119 ^ n8733 ^ 1'b0 ;
  assign n28121 = n28118 & n28120 ;
  assign n28122 = ~n13213 & n28121 ;
  assign n28123 = n28122 ^ n13043 ^ 1'b0 ;
  assign n28117 = n5205 & n6542 ;
  assign n28124 = n28123 ^ n28117 ^ 1'b0 ;
  assign n28125 = n10485 & n21999 ;
  assign n28126 = n3124 & ~n6640 ;
  assign n28127 = ~n6317 & n28126 ;
  assign n28128 = n4399 | n28127 ;
  assign n28130 = n7278 | n14919 ;
  assign n28129 = x61 | n7575 ;
  assign n28131 = n28130 ^ n28129 ^ n14986 ;
  assign n28132 = n2164 & n28131 ;
  assign n28133 = n10540 ^ n3812 ^ 1'b0 ;
  assign n28134 = n8905 ^ n7218 ^ x36 ;
  assign n28135 = n15976 & n28134 ;
  assign n28136 = n5762 & ~n28135 ;
  assign n28137 = ~n5256 & n5494 ;
  assign n28138 = ~n11191 & n28137 ;
  assign n28139 = n5725 ^ n3574 ^ 1'b0 ;
  assign n28140 = n28139 ^ n27435 ^ 1'b0 ;
  assign n28141 = x206 & ~n8352 ;
  assign n28142 = n8352 & n28141 ;
  assign n28143 = n564 & ~n2455 ;
  assign n28144 = n2455 & n28143 ;
  assign n28145 = n8481 & ~n28144 ;
  assign n28146 = ~n8481 & n28145 ;
  assign n28147 = ~n5937 & n28146 ;
  assign n28148 = n9385 | n28147 ;
  assign n28149 = n28142 | n28148 ;
  assign n28150 = n28142 & ~n28149 ;
  assign n28151 = n25295 ^ n2464 ^ 1'b0 ;
  assign n28152 = ~n577 & n28151 ;
  assign n28153 = ~n11293 & n12352 ;
  assign n28154 = n18251 & n28153 ;
  assign n28155 = n21297 ^ n12977 ^ 1'b0 ;
  assign n28157 = ~n1559 & n11050 ;
  assign n28158 = n28157 ^ n9251 ^ 1'b0 ;
  assign n28156 = n9191 & n19508 ;
  assign n28159 = n28158 ^ n28156 ^ 1'b0 ;
  assign n28160 = n23308 ^ n4536 ^ 1'b0 ;
  assign n28161 = n22618 | n24614 ;
  assign n28162 = n6647 & n26245 ;
  assign n28163 = ~n14685 & n28162 ;
  assign n28164 = x82 & ~n16252 ;
  assign n28165 = ~x82 & n28164 ;
  assign n28166 = n8160 | n28165 ;
  assign n28167 = n5525 & ~n28166 ;
  assign n28168 = n27109 | n28167 ;
  assign n28169 = n28168 ^ n21121 ^ 1'b0 ;
  assign n28170 = n22369 ^ n903 ^ 1'b0 ;
  assign n28171 = ~n4931 & n28170 ;
  assign n28172 = ~n15351 & n27533 ;
  assign n28173 = n15927 ^ n8416 ^ 1'b0 ;
  assign n28174 = n28172 | n28173 ;
  assign n28175 = x228 & ~n4580 ;
  assign n28176 = n1409 & ~n1423 ;
  assign n28177 = n28175 | n28176 ;
  assign n28182 = n3212 ^ n436 ^ 1'b0 ;
  assign n28183 = n4758 | n28182 ;
  assign n28178 = n445 & ~n5347 ;
  assign n28179 = ~n25573 & n28178 ;
  assign n28180 = n27671 ^ n5579 ^ 1'b0 ;
  assign n28181 = n28179 | n28180 ;
  assign n28184 = n28183 ^ n28181 ^ 1'b0 ;
  assign n28185 = n1740 & n8240 ;
  assign n28186 = n28185 ^ n3137 ^ 1'b0 ;
  assign n28187 = n10913 & ~n28186 ;
  assign n28188 = n1560 | n26873 ;
  assign n28189 = ~n1145 & n4834 ;
  assign n28190 = ~n4834 & n28189 ;
  assign n28191 = n16648 | n28190 ;
  assign n28192 = n8980 | n28191 ;
  assign n28193 = n8980 & ~n28192 ;
  assign n28194 = ~n23628 & n25548 ;
  assign n28195 = n28193 & n28194 ;
  assign n28197 = n15362 ^ n11523 ^ 1'b0 ;
  assign n28196 = ~n7265 & n12353 ;
  assign n28198 = n28197 ^ n28196 ^ 1'b0 ;
  assign n28199 = n4673 & ~n28198 ;
  assign n28200 = n28199 ^ n19770 ^ 1'b0 ;
  assign n28201 = ~n3575 & n28200 ;
  assign n28202 = n16855 & n28201 ;
  assign n28203 = n22782 ^ n14484 ^ 1'b0 ;
  assign n28204 = n8392 ^ n4002 ^ n1637 ;
  assign n28205 = n1549 & n28204 ;
  assign n28206 = n28205 ^ n5956 ^ 1'b0 ;
  assign n28207 = n4857 & ~n28206 ;
  assign n28208 = n7748 | n11934 ;
  assign n28209 = n28207 & ~n28208 ;
  assign n28210 = n2098 & ~n21671 ;
  assign n28211 = n28210 ^ n2385 ^ 1'b0 ;
  assign n28212 = n8378 ^ n5076 ^ n568 ;
  assign n28213 = n1192 | n17867 ;
  assign n28214 = n12777 | n28213 ;
  assign n28215 = n28214 ^ n23403 ^ 1'b0 ;
  assign n28216 = n11868 & n28215 ;
  assign n28217 = n9389 | n20181 ;
  assign n28218 = n28217 ^ n19925 ^ 1'b0 ;
  assign n28219 = n3774 & ~n28218 ;
  assign n28221 = ~n8427 & n14903 ;
  assign n28222 = n28221 ^ n3462 ^ 1'b0 ;
  assign n28220 = n8756 & n18276 ;
  assign n28223 = n28222 ^ n28220 ^ 1'b0 ;
  assign n28224 = n28223 ^ n27944 ^ 1'b0 ;
  assign n28225 = n11279 & ~n28224 ;
  assign n28233 = x64 & n27362 ;
  assign n28234 = ~n4283 & n28233 ;
  assign n28228 = n8948 ^ n5843 ^ 1'b0 ;
  assign n28229 = n25182 & ~n28228 ;
  assign n28226 = n994 ^ n756 ^ 1'b0 ;
  assign n28227 = ~n5417 & n28226 ;
  assign n28230 = n28229 ^ n28227 ^ 1'b0 ;
  assign n28231 = n10259 & n28230 ;
  assign n28232 = n28231 ^ n1512 ^ 1'b0 ;
  assign n28235 = n28234 ^ n28232 ^ 1'b0 ;
  assign n28236 = n11541 & n28235 ;
  assign n28237 = ~n2311 & n3419 ;
  assign n28238 = ~x204 & n28237 ;
  assign n28240 = n7809 & n11504 ;
  assign n28239 = n3772 & ~n14681 ;
  assign n28241 = n28240 ^ n28239 ^ n6271 ;
  assign n28242 = ~n10318 & n28241 ;
  assign n28243 = n26162 ^ n17736 ^ 1'b0 ;
  assign n28244 = n14392 ^ n8184 ^ 1'b0 ;
  assign n28245 = n28244 ^ n3872 ^ 1'b0 ;
  assign n28246 = n18128 ^ x73 ^ 1'b0 ;
  assign n28247 = n4843 & ~n9095 ;
  assign n28248 = n28247 ^ n18641 ^ 1'b0 ;
  assign n28249 = n2572 & ~n22950 ;
  assign n28250 = ~x35 & n10762 ;
  assign n28252 = n3297 & n5268 ;
  assign n28251 = n5256 & n16287 ;
  assign n28253 = n28252 ^ n28251 ^ 1'b0 ;
  assign n28254 = n28253 ^ n10222 ^ 1'b0 ;
  assign n28255 = n1642 ^ x33 ^ 1'b0 ;
  assign n28256 = n2939 & n28255 ;
  assign n28257 = ~n2668 & n10401 ;
  assign n28258 = n9655 ^ n2868 ^ 1'b0 ;
  assign n28259 = n28257 & ~n28258 ;
  assign n28260 = n2272 & n28259 ;
  assign n28261 = n2184 | n7578 ;
  assign n28262 = n28261 ^ n15652 ^ 1'b0 ;
  assign n28263 = n23991 ^ n13036 ^ 1'b0 ;
  assign n28264 = n8752 | n28263 ;
  assign n28265 = n28264 ^ n1096 ^ 1'b0 ;
  assign n28266 = n27814 ^ n841 ^ 1'b0 ;
  assign n28267 = n16784 & n17375 ;
  assign n28268 = n15081 ^ n3334 ^ 1'b0 ;
  assign n28269 = n12080 & n28268 ;
  assign n28270 = n11847 | n28269 ;
  assign n28271 = n23140 ^ n5021 ^ 1'b0 ;
  assign n28272 = n2577 & n16865 ;
  assign n28273 = n28272 ^ x50 ^ 1'b0 ;
  assign n28274 = n13794 & ~n28273 ;
  assign n28275 = n2627 & ~n28274 ;
  assign n28276 = ~n1042 & n28275 ;
  assign n28277 = n20450 ^ n9857 ^ 1'b0 ;
  assign n28278 = n5615 & ~n28277 ;
  assign n28279 = n6085 & n6857 ;
  assign n28280 = n9142 ^ n1441 ^ 1'b0 ;
  assign n28281 = n11274 & n28280 ;
  assign n28282 = ~n4333 & n6109 ;
  assign n28283 = n28282 ^ n9879 ^ 1'b0 ;
  assign n28284 = n28281 & n28283 ;
  assign n28285 = n12536 ^ n2437 ^ 1'b0 ;
  assign n28286 = n3298 | n28285 ;
  assign n28288 = n2765 | n8256 ;
  assign n28287 = n10914 ^ n9592 ^ 1'b0 ;
  assign n28289 = n28288 ^ n28287 ^ 1'b0 ;
  assign n28290 = ~n23305 & n28289 ;
  assign n28291 = ~n4020 & n28290 ;
  assign n28292 = n6359 & n11479 ;
  assign n28293 = n28292 ^ n7697 ^ 1'b0 ;
  assign n28294 = ~n1608 & n10760 ;
  assign n28295 = n28294 ^ n14353 ^ 1'b0 ;
  assign n28296 = n27959 & ~n28295 ;
  assign n28297 = n2068 | n16332 ;
  assign n28298 = ~n3581 & n28297 ;
  assign n28299 = n1638 | n12395 ;
  assign n28300 = ~n4382 & n28299 ;
  assign n28301 = n28300 ^ n13133 ^ 1'b0 ;
  assign n28302 = ~n10325 & n18030 ;
  assign n28303 = n28302 ^ n4615 ^ 1'b0 ;
  assign n28304 = n22387 ^ n2618 ^ 1'b0 ;
  assign n28305 = n1833 | n28304 ;
  assign n28306 = n15724 ^ n407 ^ 1'b0 ;
  assign n28307 = n15161 & n28306 ;
  assign n28308 = n5844 | n7074 ;
  assign n28309 = n14352 & ~n26364 ;
  assign n28312 = n26585 ^ n15829 ^ 1'b0 ;
  assign n28310 = n15309 & ~n22658 ;
  assign n28311 = n8604 & n28310 ;
  assign n28313 = n28312 ^ n28311 ^ 1'b0 ;
  assign n28314 = ~n611 & n12148 ;
  assign n28315 = n28314 ^ n15609 ^ 1'b0 ;
  assign n28316 = n26090 & ~n28315 ;
  assign n28317 = n808 & n2925 ;
  assign n28318 = n3983 ^ n2740 ^ 1'b0 ;
  assign n28319 = n20149 ^ n10222 ^ 1'b0 ;
  assign n28320 = n7325 & ~n28319 ;
  assign n28321 = n8259 | n28320 ;
  assign n28322 = n14197 ^ n9982 ^ 1'b0 ;
  assign n28323 = n4048 | n28322 ;
  assign n28324 = n28321 | n28323 ;
  assign n28325 = n4652 | n28324 ;
  assign n28326 = n28325 ^ n20164 ^ x102 ;
  assign n28327 = n28318 & ~n28326 ;
  assign n28328 = n9084 & ~n10744 ;
  assign n28329 = n28328 ^ n27825 ^ 1'b0 ;
  assign n28330 = n2518 & ~n28329 ;
  assign n28331 = n17588 ^ n1233 ^ 1'b0 ;
  assign n28332 = n16102 & n28331 ;
  assign n28333 = n28332 ^ n19699 ^ 1'b0 ;
  assign n28334 = n9075 & n28333 ;
  assign n28335 = n28334 ^ n27937 ^ 1'b0 ;
  assign n28336 = n361 & n5493 ;
  assign n28337 = n28336 ^ n6944 ^ n6884 ;
  assign n28338 = n10325 | n28337 ;
  assign n28339 = n22049 | n28338 ;
  assign n28340 = n14193 | n28339 ;
  assign n28341 = n28340 ^ n10204 ^ 1'b0 ;
  assign n28343 = n5945 ^ n2739 ^ x51 ;
  assign n28342 = n4819 & n10375 ;
  assign n28344 = n28343 ^ n28342 ^ 1'b0 ;
  assign n28345 = ~n2949 & n4429 ;
  assign n28347 = n8602 | n17361 ;
  assign n28348 = n4622 & ~n28347 ;
  assign n28346 = n1285 & ~n3426 ;
  assign n28349 = n28348 ^ n28346 ^ 1'b0 ;
  assign n28350 = n24459 ^ n5004 ^ 1'b0 ;
  assign n28351 = n10718 & n28350 ;
  assign n28352 = n4424 & ~n27581 ;
  assign n28353 = n28352 ^ n394 ^ 1'b0 ;
  assign n28354 = n17362 & ~n25747 ;
  assign n28355 = n4260 | n14859 ;
  assign n28356 = n28355 ^ n20519 ^ 1'b0 ;
  assign n28357 = n28356 ^ n6842 ^ 1'b0 ;
  assign n28358 = n10678 ^ n5070 ^ 1'b0 ;
  assign n28359 = ~n1837 & n28358 ;
  assign n28360 = n12065 & n28359 ;
  assign n28361 = ~n12201 & n28360 ;
  assign n28362 = n12378 | n28361 ;
  assign n28363 = ~n5327 & n11156 ;
  assign n28364 = n6261 ^ n4714 ^ 1'b0 ;
  assign n28365 = n11005 & n28364 ;
  assign n28366 = n28365 ^ n13675 ^ 1'b0 ;
  assign n28367 = n18417 & ~n28366 ;
  assign n28368 = n800 & n7737 ;
  assign n28369 = ~n10813 & n28368 ;
  assign n28370 = n10572 & ~n13704 ;
  assign n28371 = n1866 & ~n28370 ;
  assign n28372 = n28371 ^ n14324 ^ 1'b0 ;
  assign n28373 = n13172 | n28372 ;
  assign n28374 = n28369 | n28373 ;
  assign n28376 = ~n20975 & n21024 ;
  assign n28375 = n17611 & n28297 ;
  assign n28377 = n28376 ^ n28375 ^ 1'b0 ;
  assign n28378 = n5427 ^ n1112 ^ 1'b0 ;
  assign n28379 = n13029 & ~n28378 ;
  assign n28380 = ~n1378 & n28379 ;
  assign n28381 = n28380 ^ n21714 ^ 1'b0 ;
  assign n28382 = ~n263 & n9177 ;
  assign n28383 = n8142 & ~n13226 ;
  assign n28384 = ~n28382 & n28383 ;
  assign n28385 = n8201 & ~n13979 ;
  assign n28386 = n10236 ^ n7421 ^ 1'b0 ;
  assign n28387 = n20007 | n28386 ;
  assign n28388 = n11152 & ~n14546 ;
  assign n28389 = n28388 ^ n5525 ^ 1'b0 ;
  assign n28390 = n20405 & ~n28389 ;
  assign n28391 = n13945 ^ n7685 ^ 1'b0 ;
  assign n28392 = n28390 & ~n28391 ;
  assign n28393 = n8847 & ~n12686 ;
  assign n28394 = ~n5631 & n28393 ;
  assign n28395 = n3744 | n3929 ;
  assign n28396 = n1764 & n6655 ;
  assign n28397 = ~n14861 & n28396 ;
  assign n28398 = ~n28395 & n28397 ;
  assign n28399 = n12182 ^ n4154 ^ 1'b0 ;
  assign n28400 = n15225 | n28399 ;
  assign n28401 = n20538 ^ n1681 ^ 1'b0 ;
  assign n28402 = n2914 | n28401 ;
  assign n28403 = n2731 | n28402 ;
  assign n28404 = n28403 ^ n12002 ^ 1'b0 ;
  assign n28405 = n28404 ^ n16617 ^ 1'b0 ;
  assign n28406 = n909 | n9249 ;
  assign n28407 = n8919 & ~n28406 ;
  assign n28408 = n12040 | n28407 ;
  assign n28409 = n28408 ^ n7466 ^ 1'b0 ;
  assign n28410 = ( n5838 & ~n18629 ) | ( n5838 & n28409 ) | ( ~n18629 & n28409 ) ;
  assign n28411 = n13804 ^ n5880 ^ 1'b0 ;
  assign n28412 = n20506 | n28411 ;
  assign n28413 = n10389 ^ n6407 ^ 1'b0 ;
  assign n28414 = n3518 ^ n1690 ^ 1'b0 ;
  assign n28415 = n5915 & ~n7624 ;
  assign n28416 = ~n5151 & n28415 ;
  assign n28417 = ~n28229 & n28416 ;
  assign n28418 = n1081 & n7325 ;
  assign n28419 = n2508 & n28418 ;
  assign n28420 = n28419 ^ n7858 ^ 1'b0 ;
  assign n28421 = ~n28417 & n28420 ;
  assign n28422 = n5105 & ~n16236 ;
  assign n28423 = ~n5563 & n16895 ;
  assign n28424 = n3601 & ~n22697 ;
  assign n28425 = n28423 & n28424 ;
  assign n28426 = n15675 ^ n8657 ^ n3673 ;
  assign n28427 = n28426 ^ n4627 ^ 1'b0 ;
  assign n28428 = n5427 & n28427 ;
  assign n28429 = n28428 ^ n7940 ^ 1'b0 ;
  assign n28430 = n2839 | n4301 ;
  assign n28431 = ~n7538 & n18961 ;
  assign n28432 = ~n28430 & n28431 ;
  assign n28433 = n7175 | n28432 ;
  assign n28434 = n17537 & ~n19095 ;
  assign n28435 = n5381 & n21960 ;
  assign n28436 = n28435 ^ n19075 ^ 1'b0 ;
  assign n28437 = n9239 ^ n516 ^ 1'b0 ;
  assign n28438 = x211 | n28437 ;
  assign n28439 = n10701 & ~n24058 ;
  assign n28440 = n5418 & ~n26518 ;
  assign n28441 = n10619 ^ n3872 ^ 1'b0 ;
  assign n28442 = n13887 ^ n12522 ^ 1'b0 ;
  assign n28443 = n24414 & ~n28442 ;
  assign n28444 = n3421 & n28443 ;
  assign n28445 = n28444 ^ n10309 ^ 1'b0 ;
  assign n28446 = n5969 & n26215 ;
  assign n28447 = n27312 ^ x21 ^ 1'b0 ;
  assign n28448 = x232 & ~n895 ;
  assign n28449 = ~n2518 & n28448 ;
  assign n28450 = n2187 | n4734 ;
  assign n28451 = n718 & ~n28450 ;
  assign n28452 = n28451 ^ n2487 ^ 1'b0 ;
  assign n28453 = n28452 ^ n1190 ^ 1'b0 ;
  assign n28454 = n14871 ^ n14664 ^ 1'b0 ;
  assign n28455 = ~n21277 & n28454 ;
  assign n28456 = n21524 | n28455 ;
  assign n28460 = n12200 ^ n923 ^ 1'b0 ;
  assign n28461 = n9942 & n28460 ;
  assign n28457 = n7490 & n7721 ;
  assign n28458 = n3938 & ~n28457 ;
  assign n28459 = n9232 & n28458 ;
  assign n28462 = n28461 ^ n28459 ^ 1'b0 ;
  assign n28463 = ~n9307 & n27362 ;
  assign n28467 = n4024 & n6376 ;
  assign n28468 = ~n4024 & n28467 ;
  assign n28464 = n5918 | n6362 ;
  assign n28465 = n6362 & ~n28464 ;
  assign n28466 = n8919 | n28465 ;
  assign n28469 = n28468 ^ n28466 ^ 1'b0 ;
  assign n28470 = n28469 ^ n5893 ^ 1'b0 ;
  assign n28471 = n14647 | n28470 ;
  assign n28472 = n28471 ^ n13993 ^ 1'b0 ;
  assign n28473 = n6990 & ~n19387 ;
  assign n28474 = ~n6990 & n28473 ;
  assign n28475 = n28472 & ~n28474 ;
  assign n28476 = ~n28472 & n28475 ;
  assign n28477 = ( n5562 & n6014 ) | ( n5562 & n15483 ) | ( n6014 & n15483 ) ;
  assign n28478 = n5144 & ~n16487 ;
  assign n28479 = n3485 & n10122 ;
  assign n28480 = n28478 & n28479 ;
  assign n28482 = n23456 ^ n13788 ^ 1'b0 ;
  assign n28481 = n2704 & n5852 ;
  assign n28483 = n28482 ^ n28481 ^ 1'b0 ;
  assign n28484 = ( n4104 & ~n17488 ) | ( n4104 & n18313 ) | ( ~n17488 & n18313 ) ;
  assign n28485 = ~n7074 & n10988 ;
  assign n28487 = n12419 ^ n4854 ^ 1'b0 ;
  assign n28488 = n6861 & ~n28487 ;
  assign n28489 = n20868 & n28488 ;
  assign n28490 = n15435 & n28489 ;
  assign n28486 = n2186 | n5980 ;
  assign n28491 = n28490 ^ n28486 ^ n3888 ;
  assign n28492 = n14468 | n28026 ;
  assign n28493 = n28492 ^ n2252 ^ 1'b0 ;
  assign n28494 = n28493 ^ n23697 ^ 1'b0 ;
  assign n28495 = ~n8175 & n28494 ;
  assign n28496 = n2387 & n28495 ;
  assign n28497 = n9716 & ~n28496 ;
  assign n28498 = n28497 ^ n3107 ^ 1'b0 ;
  assign n28500 = n3357 & n4395 ;
  assign n28501 = n7970 & n28500 ;
  assign n28499 = n637 | n16862 ;
  assign n28502 = n28501 ^ n28499 ^ 1'b0 ;
  assign n28503 = x111 & ~n28502 ;
  assign n28504 = n12820 | n15748 ;
  assign n28505 = n3827 | n28504 ;
  assign n28506 = n7584 & n28505 ;
  assign n28509 = ~n2982 & n4769 ;
  assign n28510 = ~n5382 & n6557 ;
  assign n28511 = ~n28509 & n28510 ;
  assign n28512 = n28511 ^ n7736 ^ 1'b0 ;
  assign n28507 = n4310 & n8547 ;
  assign n28508 = n6053 & ~n28507 ;
  assign n28513 = n28512 ^ n28508 ^ 1'b0 ;
  assign n28514 = n7701 ^ n4284 ^ 1'b0 ;
  assign n28515 = n7077 & n7535 ;
  assign n28516 = n14876 ^ n8244 ^ 1'b0 ;
  assign n28517 = ~n23928 & n28516 ;
  assign n28518 = ~n8602 & n27652 ;
  assign n28519 = n8748 ^ n4602 ^ 1'b0 ;
  assign n28520 = ~n1675 & n28519 ;
  assign n28521 = ~n13759 & n14351 ;
  assign n28522 = n8582 & n28521 ;
  assign n28523 = n4092 | n28522 ;
  assign n28524 = ~n3566 & n8228 ;
  assign n28525 = n28524 ^ n19084 ^ 1'b0 ;
  assign n28526 = n8018 | n17874 ;
  assign n28527 = x16 & ~n28526 ;
  assign n28529 = n4730 & n23371 ;
  assign n28530 = n28529 ^ n3964 ^ 1'b0 ;
  assign n28528 = n5812 ^ n1969 ^ 1'b0 ;
  assign n28531 = n28530 ^ n28528 ^ 1'b0 ;
  assign n28532 = n2524 | n26908 ;
  assign n28533 = ~n2873 & n18180 ;
  assign n28534 = n12200 ^ n311 ^ 1'b0 ;
  assign n28535 = n11237 | n28534 ;
  assign n28536 = n17797 ^ n1572 ^ 1'b0 ;
  assign n28537 = n12414 & n28536 ;
  assign n28538 = n14501 ^ n2846 ^ 1'b0 ;
  assign n28539 = ~n13291 & n28538 ;
  assign n28540 = ~n22820 & n28539 ;
  assign n28541 = n5422 & n28540 ;
  assign n28542 = n6434 & n26079 ;
  assign n28543 = ~n12531 & n16939 ;
  assign n28545 = n23353 ^ n17254 ^ 1'b0 ;
  assign n28544 = n12601 | n18972 ;
  assign n28546 = n28545 ^ n28544 ^ 1'b0 ;
  assign n28547 = n1368 & ~n11003 ;
  assign n28548 = ~n3109 & n28547 ;
  assign n28551 = n2752 & n24060 ;
  assign n28552 = ~n10733 & n28551 ;
  assign n28553 = ~n6712 & n28552 ;
  assign n28549 = n20583 ^ n4502 ^ 1'b0 ;
  assign n28550 = n2382 & n28549 ;
  assign n28554 = n28553 ^ n28550 ^ 1'b0 ;
  assign n28555 = n12465 & n23138 ;
  assign n28556 = ~n18661 & n28555 ;
  assign n28557 = n4671 & n28556 ;
  assign n28558 = n28557 ^ n16711 ^ 1'b0 ;
  assign n28562 = n5835 ^ n3583 ^ 1'b0 ;
  assign n28563 = n9657 & ~n28562 ;
  assign n28559 = ~n901 & n16908 ;
  assign n28560 = ~n7522 & n28559 ;
  assign n28561 = n28560 ^ n19507 ^ x26 ;
  assign n28564 = n28563 ^ n28561 ^ 1'b0 ;
  assign n28565 = n9523 ^ n2846 ^ 1'b0 ;
  assign n28566 = ~n23703 & n28565 ;
  assign n28567 = n25554 & ~n28566 ;
  assign n28568 = ~n23558 & n28567 ;
  assign n28569 = ~n10663 & n14887 ;
  assign n28570 = n5168 & ~n7613 ;
  assign n28571 = ~n5168 & n28570 ;
  assign n28572 = n610 & n11094 ;
  assign n28573 = ~n11094 & n28572 ;
  assign n28574 = n11115 & n28573 ;
  assign n28575 = n28571 | n28574 ;
  assign n28576 = n26970 | n28575 ;
  assign n28577 = n6009 & ~n28576 ;
  assign n28578 = n13838 ^ n644 ^ 1'b0 ;
  assign n28579 = n21767 | n28578 ;
  assign n28580 = n1684 & ~n24949 ;
  assign n28581 = n28579 & n28580 ;
  assign n28582 = n15135 & ~n16457 ;
  assign n28583 = n6268 | n26900 ;
  assign n28584 = n15065 ^ n9051 ^ 1'b0 ;
  assign n28585 = x36 & ~n28584 ;
  assign n28586 = n11185 & n17769 ;
  assign n28587 = n3707 & n3760 ;
  assign n28588 = ~n14568 & n28587 ;
  assign n28589 = n28588 ^ n12220 ^ n1499 ;
  assign n28590 = ~n10603 & n28589 ;
  assign n28591 = n3676 & n28590 ;
  assign n28592 = n4537 ^ n3899 ^ 1'b0 ;
  assign n28593 = n7666 | n28592 ;
  assign n28594 = n21532 ^ n2975 ^ 1'b0 ;
  assign n28595 = n19542 & ~n28594 ;
  assign n28596 = n28595 ^ n17076 ^ 1'b0 ;
  assign n28597 = n2083 & n28596 ;
  assign n28598 = ~n2292 & n3611 ;
  assign n28599 = n9749 & ~n17298 ;
  assign n28600 = n15956 ^ n4537 ^ x208 ;
  assign n28601 = n14634 ^ n5392 ^ 1'b0 ;
  assign n28602 = n28601 ^ x62 ^ 1'b0 ;
  assign n28603 = n6357 & ~n22956 ;
  assign n28604 = ~n880 & n16186 ;
  assign n28605 = n2075 & ~n14476 ;
  assign n28606 = n28604 & n28605 ;
  assign n28607 = n4877 | n8074 ;
  assign n28608 = n28607 ^ n19088 ^ 1'b0 ;
  assign n28609 = x115 | n28608 ;
  assign n28610 = ~n19317 & n25293 ;
  assign n28611 = n28610 ^ n18883 ^ 1'b0 ;
  assign n28612 = n2482 & ~n3429 ;
  assign n28613 = n24823 & n28612 ;
  assign n28614 = n3700 & ~n11128 ;
  assign n28615 = n21620 ^ n19325 ^ 1'b0 ;
  assign n28616 = n8132 ^ n2006 ^ 1'b0 ;
  assign n28617 = n1684 | n28616 ;
  assign n28618 = n7108 | n10908 ;
  assign n28619 = n19088 | n28618 ;
  assign n28620 = n21755 ^ n10018 ^ n9051 ;
  assign n28621 = ~n9896 & n18498 ;
  assign n28622 = n4271 & n28621 ;
  assign n28623 = n12777 ^ n9449 ^ n6851 ;
  assign n28624 = ~n4796 & n17831 ;
  assign n28625 = n28624 ^ n12140 ^ 1'b0 ;
  assign n28626 = n2283 & ~n18270 ;
  assign n28627 = n28626 ^ x177 ^ 1'b0 ;
  assign n28628 = n27275 | n28627 ;
  assign n28629 = ~n7550 & n27315 ;
  assign n28630 = n19774 & ~n28629 ;
  assign n28631 = n2420 & n28630 ;
  assign n28632 = n16902 & ~n28631 ;
  assign n28633 = ~n28628 & n28632 ;
  assign n28634 = n9412 ^ n4827 ^ 1'b0 ;
  assign n28635 = n26139 & n28634 ;
  assign n28636 = n12152 & n28635 ;
  assign n28637 = n5750 & n28636 ;
  assign n28638 = n7333 ^ n5916 ^ 1'b0 ;
  assign n28639 = n3071 & n28638 ;
  assign n28640 = n10694 & n28639 ;
  assign n28641 = ~n14080 & n24087 ;
  assign n28642 = x159 & ~n1299 ;
  assign n28643 = ~n27695 & n28642 ;
  assign n28644 = n7732 ^ n6592 ^ 1'b0 ;
  assign n28645 = n16502 | n28644 ;
  assign n28646 = n6525 ^ n5509 ^ 1'b0 ;
  assign n28647 = n10637 | n28646 ;
  assign n28648 = n28647 ^ n21221 ^ 1'b0 ;
  assign n28649 = ~n6133 & n28648 ;
  assign n28650 = n18678 | n28649 ;
  assign n28651 = ~n13710 & n17770 ;
  assign n28652 = n1696 & ~n27053 ;
  assign n28653 = n28652 ^ n15720 ^ 1'b0 ;
  assign n28656 = n1159 & ~n11979 ;
  assign n28654 = n8123 ^ n8043 ^ 1'b0 ;
  assign n28655 = n5768 | n28654 ;
  assign n28657 = n28656 ^ n28655 ^ 1'b0 ;
  assign n28658 = ~n16208 & n24108 ;
  assign n28659 = n20087 ^ n12709 ^ 1'b0 ;
  assign n28660 = n10286 & n28659 ;
  assign n28661 = n6986 | n10221 ;
  assign n28662 = n13517 | n28661 ;
  assign n28663 = n1639 & n28662 ;
  assign n28664 = n28663 ^ n2668 ^ 1'b0 ;
  assign n28665 = n13788 | n28664 ;
  assign n28666 = n2510 | n7032 ;
  assign n28667 = n387 & ~n28666 ;
  assign n28668 = n4149 & n11443 ;
  assign n28670 = n12816 ^ n6022 ^ 1'b0 ;
  assign n28671 = n1459 & ~n28670 ;
  assign n28672 = n28671 ^ n3017 ^ 1'b0 ;
  assign n28669 = n6038 & ~n6585 ;
  assign n28673 = n28672 ^ n28669 ^ 1'b0 ;
  assign n28674 = n17971 ^ n12927 ^ 1'b0 ;
  assign n28675 = n2487 & ~n4979 ;
  assign n28676 = n4993 & n28675 ;
  assign n28677 = n28676 ^ n1646 ^ 1'b0 ;
  assign n28678 = ~n1697 & n2517 ;
  assign n28679 = n4529 & ~n28314 ;
  assign n28680 = n28679 ^ n818 ^ 1'b0 ;
  assign n28681 = n28564 ^ n17189 ^ 1'b0 ;
  assign n28682 = n21699 ^ n20113 ^ 1'b0 ;
  assign n28683 = n788 & n9186 ;
  assign n28684 = n28683 ^ n20769 ^ 1'b0 ;
  assign n28685 = n28684 ^ n7421 ^ 1'b0 ;
  assign n28686 = n3319 & ~n14365 ;
  assign n28687 = n972 & n3163 ;
  assign n28688 = n17070 & n20774 ;
  assign n28689 = n28688 ^ n5026 ^ 1'b0 ;
  assign n28690 = ( n6950 & n28687 ) | ( n6950 & n28689 ) | ( n28687 & n28689 ) ;
  assign n28691 = n1580 | n18766 ;
  assign n28692 = n28691 ^ n9518 ^ 1'b0 ;
  assign n28693 = ~n4333 & n28692 ;
  assign n28694 = ~n7594 & n14397 ;
  assign n28695 = n7666 & n28694 ;
  assign n28696 = ~n5956 & n5990 ;
  assign n28697 = ~n519 & n28696 ;
  assign n28698 = n2213 & n13385 ;
  assign n28699 = n12451 & ~n25158 ;
  assign n28700 = ~n3548 & n28699 ;
  assign n28701 = ~n352 & n2900 ;
  assign n28702 = ~n8349 & n28701 ;
  assign n28703 = n22769 ^ n6241 ^ 1'b0 ;
  assign n28704 = ~n28702 & n28703 ;
  assign n28705 = n5198 & n28532 ;
  assign n28706 = n28705 ^ n23658 ^ 1'b0 ;
  assign n28707 = n6995 ^ n5138 ^ 1'b0 ;
  assign n28708 = n26351 ^ n5121 ^ n4496 ;
  assign n28709 = n26325 ^ n24728 ^ 1'b0 ;
  assign n28710 = n28709 ^ n18971 ^ 1'b0 ;
  assign n28711 = ~n6174 & n28710 ;
  assign n28712 = n825 | n27281 ;
  assign n28713 = n11483 | n27342 ;
  assign n28714 = ( ~n9768 & n10697 ) | ( ~n9768 & n28713 ) | ( n10697 & n28713 ) ;
  assign n28715 = n21704 | n21965 ;
  assign n28716 = n2909 | n8731 ;
  assign n28717 = n21669 | n28716 ;
  assign n28718 = n28717 ^ n21299 ^ 1'b0 ;
  assign n28719 = ~n7951 & n10126 ;
  assign n28720 = ~n387 & n28719 ;
  assign n28721 = n5887 | n25667 ;
  assign n28722 = n7531 & ~n21767 ;
  assign n28723 = n12149 & ~n28722 ;
  assign n28724 = n4587 ^ n3984 ^ 1'b0 ;
  assign n28725 = ~n533 & n28724 ;
  assign n28726 = n22721 & n28725 ;
  assign n28727 = n28726 ^ n5706 ^ 1'b0 ;
  assign n28728 = n23744 & ~n28727 ;
  assign n28729 = n1100 & ~n25314 ;
  assign n28730 = n8175 & n28729 ;
  assign n28731 = n956 ^ n298 ^ 1'b0 ;
  assign n28732 = n10077 & n28731 ;
  assign n28733 = n28732 ^ n23266 ^ 1'b0 ;
  assign n28734 = n24713 & ~n28733 ;
  assign n28735 = n3888 & n28734 ;
  assign n28736 = n10287 ^ n7135 ^ n5371 ;
  assign n28738 = n6401 | n21660 ;
  assign n28737 = n2899 & ~n27001 ;
  assign n28739 = n28738 ^ n28737 ^ 1'b0 ;
  assign n28740 = n8095 ^ n4455 ^ 1'b0 ;
  assign n28741 = n28740 ^ n27526 ^ 1'b0 ;
  assign n28742 = ~n12233 & n28741 ;
  assign n28743 = n3960 | n17499 ;
  assign n28744 = ~n2715 & n13651 ;
  assign n28745 = n28744 ^ n15189 ^ 1'b0 ;
  assign n28746 = ~n25493 & n26315 ;
  assign n28747 = ~n3078 & n9128 ;
  assign n28748 = n9907 & ~n20855 ;
  assign n28749 = n1666 & n22376 ;
  assign n28750 = n9177 & n14000 ;
  assign n28751 = n23763 & n28750 ;
  assign n28752 = n4636 | n18822 ;
  assign n28753 = n20860 ^ n17601 ^ 1'b0 ;
  assign n28754 = n4980 ^ n1354 ^ 1'b0 ;
  assign n28755 = n7907 & n28754 ;
  assign n28756 = n12035 ^ n6089 ^ 1'b0 ;
  assign n28757 = n28755 & ~n28756 ;
  assign n28758 = n8621 ^ n7359 ^ 1'b0 ;
  assign n28759 = n5843 | n28758 ;
  assign n28760 = ~n747 & n4074 ;
  assign n28761 = n28760 ^ n5991 ^ 1'b0 ;
  assign n28762 = n13056 ^ n5877 ^ 1'b0 ;
  assign n28763 = n19697 & n28762 ;
  assign n28764 = n4238 ^ n2356 ^ 1'b0 ;
  assign n28765 = n6468 & n28764 ;
  assign n28766 = n5600 & n28765 ;
  assign n28767 = n3798 | n28766 ;
  assign n28768 = n17512 ^ n470 ^ 1'b0 ;
  assign n28769 = n3672 | n4423 ;
  assign n28770 = ~n5124 & n28769 ;
  assign n28771 = n21487 ^ n19533 ^ 1'b0 ;
  assign n28772 = n28770 & ~n28771 ;
  assign n28773 = x71 & n10778 ;
  assign n28774 = n4545 & ~n10847 ;
  assign n28775 = n10672 & n23294 ;
  assign n28776 = n11359 ^ n9688 ^ 1'b0 ;
  assign n28777 = n10354 & ~n28776 ;
  assign n28778 = n7076 & ~n15455 ;
  assign n28779 = ~n28777 & n28778 ;
  assign n28780 = n6681 | n23601 ;
  assign n28781 = n7528 & ~n28780 ;
  assign n28782 = ~n1249 & n21335 ;
  assign n28783 = n14675 ^ n13727 ^ 1'b0 ;
  assign n28784 = n20225 ^ n5484 ^ 1'b0 ;
  assign n28785 = n6727 ^ n3280 ^ 1'b0 ;
  assign n28786 = ~n26438 & n27320 ;
  assign n28787 = n10403 ^ n3487 ^ 1'b0 ;
  assign n28788 = ~n6710 & n28787 ;
  assign n28789 = n3888 | n6290 ;
  assign n28790 = n28789 ^ n22737 ^ 1'b0 ;
  assign n28791 = n28297 ^ n8735 ^ 1'b0 ;
  assign n28792 = n28790 & ~n28791 ;
  assign n28795 = n7113 ^ n5744 ^ n1596 ;
  assign n28793 = n6073 ^ n1299 ^ 1'b0 ;
  assign n28794 = n28793 ^ n4094 ^ 1'b0 ;
  assign n28796 = n28795 ^ n28794 ^ 1'b0 ;
  assign n28797 = n4939 & ~n28796 ;
  assign n28798 = n2275 & n28797 ;
  assign n28799 = n8290 | n8947 ;
  assign n28800 = n9340 & ~n28799 ;
  assign n28801 = n6702 | n28800 ;
  assign n28802 = n10861 ^ n5500 ^ 1'b0 ;
  assign n28803 = x64 & ~n28802 ;
  assign n28804 = n10633 & n11688 ;
  assign n28805 = x20 & n28804 ;
  assign n28806 = n28805 ^ n4590 ^ 1'b0 ;
  assign n28807 = n27731 | n28806 ;
  assign n28808 = n4500 & n10276 ;
  assign n28809 = n7580 & ~n22290 ;
  assign n28810 = n28808 & n28809 ;
  assign n28814 = n15077 ^ n7539 ^ n2725 ;
  assign n28811 = n5877 & ~n27244 ;
  assign n28812 = n28811 ^ n16067 ^ 1'b0 ;
  assign n28813 = ~n5798 & n28812 ;
  assign n28815 = n28814 ^ n28813 ^ n12220 ;
  assign n28816 = ~n3013 & n9380 ;
  assign n28817 = ~n7214 & n15999 ;
  assign n28818 = n3022 | n11269 ;
  assign n28819 = n28818 ^ n19754 ^ 1'b0 ;
  assign n28821 = ~n2523 & n23199 ;
  assign n28822 = n28821 ^ n9755 ^ 1'b0 ;
  assign n28820 = n5308 ^ n4290 ^ 1'b0 ;
  assign n28823 = n28822 ^ n28820 ^ 1'b0 ;
  assign n28824 = n13029 | n28823 ;
  assign n28825 = n18725 ^ n14029 ^ 1'b0 ;
  assign n28826 = n25640 ^ x130 ^ 1'b0 ;
  assign n28827 = n20752 & ~n21415 ;
  assign n28828 = n28827 ^ n7132 ^ 1'b0 ;
  assign n28829 = x59 | n1791 ;
  assign n28830 = n28461 & ~n28829 ;
  assign n28831 = n28830 ^ n4241 ^ 1'b0 ;
  assign n28832 = n16610 | n25520 ;
  assign n28833 = n2911 ^ n1847 ^ 1'b0 ;
  assign n28834 = n28833 ^ n22018 ^ 1'b0 ;
  assign n28835 = n11048 | n11096 ;
  assign n28836 = ( n832 & n21551 ) | ( n832 & n28835 ) | ( n21551 & n28835 ) ;
  assign n28837 = n1449 ^ x193 ^ 1'b0 ;
  assign n28838 = n21545 ^ n1470 ^ 1'b0 ;
  assign n28839 = n28837 & ~n28838 ;
  assign n28840 = n20922 ^ n12202 ^ 1'b0 ;
  assign n28841 = n17777 ^ n1212 ^ 1'b0 ;
  assign n28842 = n13585 ^ n10721 ^ 1'b0 ;
  assign n28843 = ~n4888 & n23926 ;
  assign n28844 = n21024 & n26915 ;
  assign n28846 = n5686 & n7192 ;
  assign n28847 = ~n1808 & n28846 ;
  assign n28848 = n11065 & ~n28847 ;
  assign n28845 = n8334 & n24531 ;
  assign n28849 = n28848 ^ n28845 ^ 1'b0 ;
  assign n28850 = n1160 & n6998 ;
  assign n28851 = ~n1264 & n3533 ;
  assign n28852 = n28851 ^ n5107 ^ 1'b0 ;
  assign n28853 = n20515 & n28852 ;
  assign n28854 = ~n3920 & n15842 ;
  assign n28855 = n28854 ^ n3803 ^ 1'b0 ;
  assign n28856 = n2066 & n5073 ;
  assign n28857 = n18333 ^ n1446 ^ 1'b0 ;
  assign n28858 = n4382 | n10035 ;
  assign n28859 = n25379 & ~n28858 ;
  assign n28860 = ~n2665 & n11504 ;
  assign n28861 = n891 & ~n14395 ;
  assign n28862 = ~n1100 & n24778 ;
  assign n28863 = ~n6030 & n13656 ;
  assign n28864 = ~n2129 & n2648 ;
  assign n28865 = n6712 ^ n6583 ^ 1'b0 ;
  assign n28866 = ~n27320 & n28865 ;
  assign n28867 = n27512 ^ n25458 ^ 1'b0 ;
  assign n28868 = ~n19800 & n28867 ;
  assign n28871 = ~n2021 & n13598 ;
  assign n28872 = ~x161 & n28871 ;
  assign n28870 = ~n18723 & n23048 ;
  assign n28873 = n28872 ^ n28870 ^ 1'b0 ;
  assign n28869 = n9471 | n9911 ;
  assign n28874 = n28873 ^ n28869 ^ 1'b0 ;
  assign n28875 = n12581 & ~n28874 ;
  assign n28876 = n23035 ^ n12329 ^ 1'b0 ;
  assign n28877 = n27833 & ~n28163 ;
  assign n28878 = n10367 ^ n5050 ^ 1'b0 ;
  assign n28879 = n20720 ^ n858 ^ 1'b0 ;
  assign n28880 = ~n12180 & n28879 ;
  assign n28881 = n27667 ^ n3558 ^ 1'b0 ;
  assign n28882 = n28880 | n28881 ;
  assign n28883 = n880 & ~n19533 ;
  assign n28884 = n8944 & n28883 ;
  assign n28885 = n4132 & n27497 ;
  assign n28886 = n5358 & ~n27911 ;
  assign n28887 = n1731 & ~n6969 ;
  assign n28888 = n28887 ^ n12758 ^ 1'b0 ;
  assign n28889 = ~n28886 & n28888 ;
  assign n28890 = n9771 & ~n28889 ;
  assign n28891 = n28890 ^ n25428 ^ 1'b0 ;
  assign n28893 = n17936 ^ n3095 ^ 1'b0 ;
  assign n28892 = n5095 & ~n26426 ;
  assign n28894 = n28893 ^ n28892 ^ 1'b0 ;
  assign n28895 = ~n8944 & n28894 ;
  assign n28896 = n28895 ^ n8534 ^ 1'b0 ;
  assign n28897 = n1164 & ~n26900 ;
  assign n28898 = n25673 ^ n22073 ^ n21216 ;
  assign n28899 = n28795 & n28898 ;
  assign n28900 = n2230 | n8294 ;
  assign n28901 = n21563 ^ n13279 ^ 1'b0 ;
  assign n28902 = n23212 & ~n28901 ;
  assign n28903 = n1016 & n28902 ;
  assign n28904 = ( ~n4289 & n27077 ) | ( ~n4289 & n28903 ) | ( n27077 & n28903 ) ;
  assign n28905 = n2074 ^ n1066 ^ 1'b0 ;
  assign n28906 = n1786 & ~n28905 ;
  assign n28907 = ~n4076 & n28906 ;
  assign n28908 = n14818 ^ n7710 ^ 1'b0 ;
  assign n28909 = n16497 & ~n28908 ;
  assign n28910 = n5275 ^ n4154 ^ 1'b0 ;
  assign n28911 = ~n22290 & n28910 ;
  assign n28912 = ~n5424 & n14057 ;
  assign n28913 = n1646 | n2503 ;
  assign n28914 = n17628 ^ n1007 ^ 1'b0 ;
  assign n28915 = n17681 & ~n18519 ;
  assign n28916 = n28915 ^ n8033 ^ 1'b0 ;
  assign n28917 = n18828 ^ n16574 ^ 1'b0 ;
  assign n28918 = n21786 & n24262 ;
  assign n28919 = n19966 ^ n3611 ^ n2955 ;
  assign n28921 = n16222 ^ n5911 ^ 1'b0 ;
  assign n28922 = n6552 & n28921 ;
  assign n28920 = ~n4815 & n9097 ;
  assign n28923 = n28922 ^ n28920 ^ 1'b0 ;
  assign n28924 = n5457 & ~n10711 ;
  assign n28925 = n28924 ^ n18557 ^ 1'b0 ;
  assign n28926 = ~n2140 & n7259 ;
  assign n28927 = n28925 & n28926 ;
  assign n28929 = n5223 & n20156 ;
  assign n28928 = x157 & ~n2022 ;
  assign n28930 = n28929 ^ n28928 ^ 1'b0 ;
  assign n28931 = n24825 ^ n4178 ^ 1'b0 ;
  assign n28932 = ~n23512 & n28931 ;
  assign n28933 = n6777 & ~n23803 ;
  assign n28934 = n644 & n7193 ;
  assign n28935 = n13481 & ~n28934 ;
  assign n28936 = ~n3593 & n16722 ;
  assign n28937 = n5648 ^ n3703 ^ 1'b0 ;
  assign n28938 = n28936 & n28937 ;
  assign n28939 = ~n11859 & n14993 ;
  assign n28940 = n11599 | n28939 ;
  assign n28941 = n24431 ^ n2451 ^ 1'b0 ;
  assign n28942 = n6812 | n28941 ;
  assign n28943 = n6263 & n11093 ;
  assign n28944 = n1424 & n20072 ;
  assign n28946 = n2527 & n22886 ;
  assign n28945 = n776 & n14275 ;
  assign n28947 = n28946 ^ n28945 ^ 1'b0 ;
  assign n28948 = ~n4955 & n8198 ;
  assign n28949 = ~n11364 & n13428 ;
  assign n28950 = n28949 ^ n2083 ^ 1'b0 ;
  assign n28951 = ~n28948 & n28950 ;
  assign n28952 = n23977 ^ n16789 ^ 1'b0 ;
  assign n28954 = n387 & ~n12744 ;
  assign n28953 = ~n12707 & n16868 ;
  assign n28955 = n28954 ^ n28953 ^ 1'b0 ;
  assign n28956 = n11918 & ~n21154 ;
  assign n28957 = n28956 ^ n5343 ^ 1'b0 ;
  assign n28958 = n20908 | n28957 ;
  assign n28959 = n1978 & ~n10689 ;
  assign n28960 = n14685 & n28959 ;
  assign n28961 = n11651 & n28960 ;
  assign n28962 = n313 & n15061 ;
  assign n28963 = ~n22284 & n28962 ;
  assign n28964 = n409 & n28963 ;
  assign n28965 = n28964 ^ n7768 ^ 1'b0 ;
  assign n28966 = n1239 & n2893 ;
  assign n28967 = n28966 ^ n18527 ^ 1'b0 ;
  assign n28968 = n10002 & ~n26910 ;
  assign n28979 = n1042 & ~n1882 ;
  assign n28980 = ~n1042 & n28979 ;
  assign n28981 = ~n4358 & n28980 ;
  assign n28982 = ~n1337 & n28981 ;
  assign n28970 = ~n2826 & n11029 ;
  assign n28971 = n8395 & n28970 ;
  assign n28972 = n2909 & ~n4840 ;
  assign n28973 = n4840 & n28972 ;
  assign n28974 = n28973 ^ n5185 ^ 1'b0 ;
  assign n28975 = n28971 & n28974 ;
  assign n28976 = n17656 & n21554 ;
  assign n28977 = n28976 ^ n7275 ^ 1'b0 ;
  assign n28978 = n28975 & ~n28977 ;
  assign n28983 = n28982 ^ n28978 ^ 1'b0 ;
  assign n28969 = n3006 | n19460 ;
  assign n28984 = n28983 ^ n28969 ^ 1'b0 ;
  assign n28985 = n15543 & n23046 ;
  assign n28986 = n2633 & ~n28985 ;
  assign n28987 = n28986 ^ n15842 ^ 1'b0 ;
  assign n28988 = n7680 & n13970 ;
  assign n28989 = ~n24778 & n28988 ;
  assign n28990 = ~n14593 & n28509 ;
  assign n28991 = n28990 ^ n18541 ^ 1'b0 ;
  assign n28992 = n5521 | n28991 ;
  assign n28996 = n10094 ^ n9012 ^ 1'b0 ;
  assign n28997 = n3413 | n28996 ;
  assign n28993 = n6557 ^ n2429 ^ 1'b0 ;
  assign n28994 = n4103 & n28993 ;
  assign n28995 = n4179 & n28994 ;
  assign n28998 = n28997 ^ n28995 ^ 1'b0 ;
  assign n28999 = n22995 ^ n2074 ^ 1'b0 ;
  assign n29000 = n2466 ^ n948 ^ 1'b0 ;
  assign n29001 = n28999 & ~n29000 ;
  assign n29002 = n2959 & n26337 ;
  assign n29003 = x95 & n29002 ;
  assign n29004 = n29003 ^ n14869 ^ 1'b0 ;
  assign n29005 = n29004 ^ n16709 ^ n4598 ;
  assign n29006 = n21172 & ~n26098 ;
  assign n29007 = ~n4711 & n29006 ;
  assign n29008 = n9103 ^ n8251 ^ 1'b0 ;
  assign n29009 = n23385 & n28217 ;
  assign n29010 = n17139 ^ n10652 ^ n8414 ;
  assign n29011 = n10305 & ~n29010 ;
  assign n29012 = n27410 ^ n25173 ^ n17669 ;
  assign n29013 = n29012 ^ n17332 ^ 1'b0 ;
  assign n29014 = ( n929 & n12302 ) | ( n929 & n29013 ) | ( n12302 & n29013 ) ;
  assign n29015 = ~n2637 & n29014 ;
  assign n29017 = ~n788 & n18588 ;
  assign n29016 = n4316 & n22621 ;
  assign n29018 = n29017 ^ n29016 ^ 1'b0 ;
  assign n29019 = n22836 ^ n8283 ^ 1'b0 ;
  assign n29020 = ~n2040 & n26418 ;
  assign n29021 = n11668 & n29020 ;
  assign n29022 = n3739 & ~n15060 ;
  assign n29023 = ~n21260 & n29022 ;
  assign n29024 = n23680 & n29023 ;
  assign n29025 = n17752 ^ n8388 ^ 1'b0 ;
  assign n29026 = n12529 & ~n29025 ;
  assign n29027 = n6287 & n8912 ;
  assign n29028 = ~n19727 & n29027 ;
  assign n29029 = n12988 ^ n6589 ^ 1'b0 ;
  assign n29030 = n29028 | n29029 ;
  assign n29031 = n4103 & ~n9239 ;
  assign n29032 = n5129 & n29031 ;
  assign n29033 = n26491 | n29032 ;
  assign n29034 = n17731 & ~n23305 ;
  assign n29035 = ~n29033 & n29034 ;
  assign n29036 = ~n3329 & n18696 ;
  assign n29037 = ( x152 & n298 ) | ( x152 & ~n15312 ) | ( n298 & ~n15312 ) ;
  assign n29038 = ~n15566 & n29037 ;
  assign n29039 = ~x186 & n29038 ;
  assign n29040 = n29039 ^ n1353 ^ 1'b0 ;
  assign n29041 = n24645 ^ n14871 ^ n7785 ;
  assign n29045 = n7007 & n13115 ;
  assign n29042 = n10027 | n17226 ;
  assign n29043 = n22842 | n29042 ;
  assign n29044 = ~n7421 & n29043 ;
  assign n29046 = n29045 ^ n29044 ^ 1'b0 ;
  assign n29047 = n21034 ^ n815 ^ 1'b0 ;
  assign n29048 = n27437 & n29047 ;
  assign n29049 = ~n1575 & n18585 ;
  assign n29050 = ( ~n13106 & n21182 ) | ( ~n13106 & n28962 ) | ( n21182 & n28962 ) ;
  assign n29051 = n11259 ^ n5231 ^ 1'b0 ;
  assign n29052 = n8332 & ~n29051 ;
  assign n29053 = n1260 & ~n3939 ;
  assign n29054 = n23021 ^ n12172 ^ 1'b0 ;
  assign n29055 = n8094 | n29054 ;
  assign n29056 = n2185 & n18134 ;
  assign n29057 = n29056 ^ n4582 ^ 1'b0 ;
  assign n29058 = n21158 ^ n10330 ^ 1'b0 ;
  assign n29059 = n8562 ^ n2115 ^ 1'b0 ;
  assign n29060 = ~n4526 & n5968 ;
  assign n29061 = ~n24263 & n26385 ;
  assign n29062 = n29061 ^ n10590 ^ 1'b0 ;
  assign n29063 = n1337 | n1472 ;
  assign n29064 = n29063 ^ n11520 ^ 1'b0 ;
  assign n29065 = n26510 | n29064 ;
  assign n29066 = n29062 | n29065 ;
  assign n29067 = n8750 & ~n22771 ;
  assign n29068 = ~n29066 & n29067 ;
  assign n29069 = ( n9273 & ~n13468 ) | ( n9273 & n18660 ) | ( ~n13468 & n18660 ) ;
  assign n29070 = n23293 ^ n8251 ^ 1'b0 ;
  assign n29071 = n17804 & n29070 ;
  assign n29072 = ~n9178 & n25647 ;
  assign n29073 = n10397 ^ n4157 ^ 1'b0 ;
  assign n29074 = ~n10018 & n21281 ;
  assign n29077 = ~n6473 & n14069 ;
  assign n29078 = n29077 ^ n3368 ^ 1'b0 ;
  assign n29075 = ~x76 & n3905 ;
  assign n29076 = n3933 & n29075 ;
  assign n29079 = n29078 ^ n29076 ^ 1'b0 ;
  assign n29080 = n29079 ^ n22819 ^ 1'b0 ;
  assign n29081 = n2477 ^ n1337 ^ 1'b0 ;
  assign n29082 = n29081 ^ n21601 ^ 1'b0 ;
  assign n29083 = n15927 ^ n14308 ^ 1'b0 ;
  assign n29086 = ~n4827 & n7220 ;
  assign n29087 = n14820 ^ n6412 ^ 1'b0 ;
  assign n29088 = n29086 & ~n29087 ;
  assign n29085 = ( ~n871 & n9721 ) | ( ~n871 & n12026 ) | ( n9721 & n12026 ) ;
  assign n29084 = n4562 & ~n5692 ;
  assign n29089 = n29088 ^ n29085 ^ n29084 ;
  assign n29090 = n11979 ^ n5495 ^ 1'b0 ;
  assign n29091 = n1920 | n29090 ;
  assign n29092 = n3292 ^ n2561 ^ 1'b0 ;
  assign n29093 = n3093 & n21995 ;
  assign n29094 = ~n3619 & n29093 ;
  assign n29095 = n22354 ^ n5719 ^ 1'b0 ;
  assign n29096 = n9803 & n29095 ;
  assign n29097 = n9005 | n29096 ;
  assign n29100 = n1076 & ~n2019 ;
  assign n29098 = n14071 | n18986 ;
  assign n29099 = n22756 & ~n29098 ;
  assign n29101 = n29100 ^ n29099 ^ n22110 ;
  assign n29102 = n1028 & n19174 ;
  assign n29103 = n9716 ^ n2119 ^ 1'b0 ;
  assign n29104 = n29102 | n29103 ;
  assign n29105 = n6031 | n6550 ;
  assign n29106 = n16371 ^ n2503 ^ 1'b0 ;
  assign n29107 = n15260 ^ n987 ^ 1'b0 ;
  assign n29108 = n2809 & ~n29107 ;
  assign n29109 = n29108 ^ n9307 ^ 1'b0 ;
  assign n29111 = n9535 ^ n907 ^ 1'b0 ;
  assign n29110 = n5702 & ~n26530 ;
  assign n29112 = n29111 ^ n29110 ^ n18478 ;
  assign n29113 = n14335 | n29112 ;
  assign n29114 = n6208 ^ n1266 ^ 1'b0 ;
  assign n29115 = n29114 ^ n18366 ^ 1'b0 ;
  assign n29116 = n7146 ^ n1264 ^ n635 ;
  assign n29117 = n9232 & ~n29116 ;
  assign n29118 = n29117 ^ n2131 ^ 1'b0 ;
  assign n29119 = n15898 ^ n8343 ^ 1'b0 ;
  assign n29120 = n1725 ^ n734 ^ 1'b0 ;
  assign n29121 = n29120 ^ n13243 ^ 1'b0 ;
  assign n29122 = ~n20690 & n29121 ;
  assign n29123 = n26017 ^ n14192 ^ 1'b0 ;
  assign n29124 = n16284 ^ n2279 ^ 1'b0 ;
  assign n29125 = n5334 & n29124 ;
  assign n29126 = n29125 ^ n603 ^ 1'b0 ;
  assign n29127 = n6372 & ~n29126 ;
  assign n29128 = n29123 | n29127 ;
  assign n29129 = n7117 & ~n14231 ;
  assign n29130 = n27406 & n28509 ;
  assign n29131 = ~n4118 & n29130 ;
  assign n29132 = n18454 & ~n26921 ;
  assign n29133 = n25178 ^ n2845 ^ 1'b0 ;
  assign n29134 = ~n29132 & n29133 ;
  assign n29135 = n21112 ^ n11061 ^ 1'b0 ;
  assign n29136 = ~n20000 & n29135 ;
  assign n29137 = n9340 & n29136 ;
  assign n29138 = n930 & n4698 ;
  assign n29139 = n28005 ^ n14032 ^ n12543 ;
  assign n29140 = n3583 & ~n10856 ;
  assign n29141 = n4677 & n17562 ;
  assign n29142 = n29141 ^ n21377 ^ 1'b0 ;
  assign n29144 = x5 & n15933 ;
  assign n29145 = n11240 & ~n29144 ;
  assign n29143 = n3068 & n8641 ;
  assign n29146 = n29145 ^ n29143 ^ 1'b0 ;
  assign n29147 = n10090 ^ n3754 ^ 1'b0 ;
  assign n29148 = n3903 & ~n29147 ;
  assign n29149 = n2798 ^ n1608 ^ 1'b0 ;
  assign n29150 = n7017 & n29149 ;
  assign n29151 = n15169 ^ n2681 ^ 1'b0 ;
  assign n29152 = n29150 & n29151 ;
  assign n29153 = n10888 | n15565 ;
  assign n29154 = ~n2749 & n4627 ;
  assign n29155 = n4536 & ~n6670 ;
  assign n29156 = n4400 & ~n29155 ;
  assign n29157 = n29154 & n29156 ;
  assign n29158 = n25518 & ~n29157 ;
  assign n29159 = n29158 ^ n5601 ^ 1'b0 ;
  assign n29160 = n29153 | n29159 ;
  assign n29161 = n16584 ^ n11203 ^ 1'b0 ;
  assign n29162 = n23463 & ~n29161 ;
  assign n29163 = n29162 ^ n3245 ^ 1'b0 ;
  assign n29164 = n1684 & n29163 ;
  assign n29165 = n2768 & ~n29164 ;
  assign n29166 = n637 & n1249 ;
  assign n29167 = ~n1249 & n29166 ;
  assign n29168 = n29167 ^ n13125 ^ 1'b0 ;
  assign n29169 = n807 & n2079 ;
  assign n29170 = ~n2079 & n29169 ;
  assign n29171 = ~n3505 & n9410 ;
  assign n29172 = n3505 & n29171 ;
  assign n29173 = n12334 & n29172 ;
  assign n29174 = n29170 | n29173 ;
  assign n29175 = n29168 & ~n29174 ;
  assign n29176 = n11518 | n20232 ;
  assign n29177 = n9076 | n29176 ;
  assign n29178 = n14192 ^ n1195 ^ n797 ;
  assign n29179 = n12783 & n29178 ;
  assign n29180 = n29177 & n29179 ;
  assign n29181 = n1693 & n29180 ;
  assign n29182 = n315 | n3984 ;
  assign n29183 = n29182 ^ n7539 ^ 1'b0 ;
  assign n29184 = n3762 | n3764 ;
  assign n29185 = n6749 & ~n29184 ;
  assign n29186 = ~n10623 & n16329 ;
  assign n29187 = n25391 ^ n3137 ^ 1'b0 ;
  assign n29188 = n29186 & ~n29187 ;
  assign n29189 = ~x47 & n2440 ;
  assign n29190 = n29189 ^ n13551 ^ n11451 ;
  assign n29191 = n841 & ~n15675 ;
  assign n29192 = ~n19517 & n29191 ;
  assign n29193 = n5134 | n29192 ;
  assign n29194 = n13854 & ~n29193 ;
  assign n29195 = n25631 & n28954 ;
  assign n29196 = ~n15587 & n19212 ;
  assign n29197 = n29196 ^ n2863 ^ 1'b0 ;
  assign n29198 = n4238 & n29197 ;
  assign n29199 = ~n18821 & n29198 ;
  assign n29200 = n29199 ^ n28438 ^ 1'b0 ;
  assign n29201 = ( n19940 & n28204 ) | ( n19940 & n28564 ) | ( n28204 & n28564 ) ;
  assign n29202 = n2097 | n13127 ;
  assign n29203 = n1766 & ~n6437 ;
  assign n29204 = n29203 ^ n10900 ^ 1'b0 ;
  assign n29205 = n25030 ^ n9012 ^ 1'b0 ;
  assign n29206 = n29204 | n29205 ;
  assign n29207 = n2463 | n6112 ;
  assign n29208 = n29207 ^ n5076 ^ 1'b0 ;
  assign n29209 = ~n23329 & n29208 ;
  assign n29210 = n1320 & n29209 ;
  assign n29211 = n4933 | n29210 ;
  assign n29212 = ~n2311 & n3813 ;
  assign n29213 = n29212 ^ n5504 ^ 1'b0 ;
  assign n29214 = n5579 & n29213 ;
  assign n29215 = n29214 ^ n9966 ^ 1'b0 ;
  assign n29216 = n13027 & ~n29215 ;
  assign n29217 = n4428 ^ n807 ^ 1'b0 ;
  assign n29218 = n29186 & n29217 ;
  assign n29219 = n10605 ^ n7148 ^ 1'b0 ;
  assign n29220 = n7695 & n29219 ;
  assign n29221 = n4215 | n6342 ;
  assign n29222 = n1977 & n6712 ;
  assign n29223 = ~n5398 & n29222 ;
  assign n29224 = n17376 | n29223 ;
  assign n29225 = n6358 & n29224 ;
  assign n29226 = n15812 & n21684 ;
  assign n29227 = n29226 ^ n7308 ^ 1'b0 ;
  assign n29228 = n8725 | n11445 ;
  assign n29229 = n29228 ^ n5006 ^ 1'b0 ;
  assign n29230 = ~n21493 & n29229 ;
  assign n29231 = n5074 & ~n12000 ;
  assign n29233 = ~n8111 & n8541 ;
  assign n29232 = n9998 ^ n8160 ^ n4680 ;
  assign n29234 = n29233 ^ n29232 ^ 1'b0 ;
  assign n29235 = n15884 ^ n13857 ^ 1'b0 ;
  assign n29236 = n26456 & ~n29235 ;
  assign n29237 = n3217 ^ x167 ^ 1'b0 ;
  assign n29238 = n29237 ^ n12956 ^ 1'b0 ;
  assign n29239 = ~n23158 & n29238 ;
  assign n29240 = n22025 ^ n1062 ^ 1'b0 ;
  assign n29241 = ( ~n13279 & n18236 ) | ( ~n13279 & n29240 ) | ( n18236 & n29240 ) ;
  assign n29242 = n4720 & n6945 ;
  assign n29243 = n29242 ^ n2491 ^ 1'b0 ;
  assign n29244 = n16204 ^ n11207 ^ 1'b0 ;
  assign n29245 = n29243 & ~n29244 ;
  assign n29246 = n8116 ^ n3893 ^ 1'b0 ;
  assign n29247 = n11572 & ~n29246 ;
  assign n29248 = n29247 ^ n2472 ^ 1'b0 ;
  assign n29249 = ~n1451 & n29248 ;
  assign n29250 = n7281 ^ n1021 ^ 1'b0 ;
  assign n29251 = n5965 & ~n29250 ;
  assign n29252 = n1969 & n6744 ;
  assign n29253 = x145 & ~n29252 ;
  assign n29254 = ~n29251 & n29253 ;
  assign n29255 = n9881 & ~n11486 ;
  assign n29256 = n29255 ^ n9097 ^ 1'b0 ;
  assign n29257 = n5922 | n8944 ;
  assign n29258 = n20864 & ~n29257 ;
  assign n29259 = n27997 ^ n21525 ^ 1'b0 ;
  assign n29260 = n15815 & n29259 ;
  assign n29261 = n24878 ^ n1361 ^ 1'b0 ;
  assign n29262 = n20302 ^ n15126 ^ 1'b0 ;
  assign n29263 = ~n718 & n29262 ;
  assign n29264 = n14192 & n29263 ;
  assign n29265 = n29264 ^ n21480 ^ 1'b0 ;
  assign n29266 = n5627 | n14839 ;
  assign n29267 = n29266 ^ n548 ^ 1'b0 ;
  assign n29268 = n9361 & ~n13813 ;
  assign n29269 = n5518 & n29268 ;
  assign n29270 = n8602 | n29099 ;
  assign n29271 = n23658 | n29270 ;
  assign n29272 = n15737 ^ n3426 ^ 1'b0 ;
  assign n29273 = n10867 & n29272 ;
  assign n29274 = x160 & n29273 ;
  assign n29275 = ~n7043 & n29274 ;
  assign n29276 = n538 & ~n27297 ;
  assign n29277 = ~n19418 & n29276 ;
  assign n29278 = ~n5337 & n27758 ;
  assign n29279 = n4220 & n29278 ;
  assign n29280 = n2047 ^ n1571 ^ 1'b0 ;
  assign n29281 = n2402 | n29280 ;
  assign n29282 = n29281 ^ n17563 ^ n13044 ;
  assign n29283 = n5492 & ~n15515 ;
  assign n29284 = n11956 & ~n27806 ;
  assign n29285 = n27411 ^ n4573 ^ 1'b0 ;
  assign n29286 = n22684 | n29285 ;
  assign n29287 = ~n6605 & n13054 ;
  assign n29288 = ~n7508 & n29287 ;
  assign n29289 = n354 & n1249 ;
  assign n29290 = n29288 & n29289 ;
  assign n29291 = ( n12720 & n28769 ) | ( n12720 & ~n29290 ) | ( n28769 & ~n29290 ) ;
  assign n29293 = n4676 & n9214 ;
  assign n29292 = n14327 & n18361 ;
  assign n29294 = n29293 ^ n29292 ^ 1'b0 ;
  assign n29295 = n8811 ^ n722 ^ 1'b0 ;
  assign n29296 = n571 & n29295 ;
  assign n29297 = n29296 ^ n29024 ^ 1'b0 ;
  assign n29298 = n5413 & n14022 ;
  assign n29299 = ~n2633 & n29298 ;
  assign n29300 = n5287 & ~n22051 ;
  assign n29301 = n10186 & n29300 ;
  assign n29302 = n12980 | n15975 ;
  assign n29303 = n12940 & ~n29302 ;
  assign n29304 = n3487 & n3727 ;
  assign n29305 = ~n5821 & n7451 ;
  assign n29306 = ~n1544 & n9181 ;
  assign n29307 = ( n27941 & n29305 ) | ( n27941 & n29306 ) | ( n29305 & n29306 ) ;
  assign n29308 = n1658 & ~n6443 ;
  assign n29310 = n5384 ^ n2615 ^ 1'b0 ;
  assign n29309 = ~x22 & n22073 ;
  assign n29311 = n29310 ^ n29309 ^ 1'b0 ;
  assign n29312 = n14678 | n29311 ;
  assign n29313 = n6019 ^ n2744 ^ 1'b0 ;
  assign n29314 = n12060 & ~n29313 ;
  assign n29315 = n15891 ^ n1724 ^ 1'b0 ;
  assign n29316 = n1920 ^ n498 ^ 1'b0 ;
  assign n29317 = n6480 ^ n3217 ^ 1'b0 ;
  assign n29318 = n9874 & n29317 ;
  assign n29319 = ~n10519 & n29318 ;
  assign n29320 = n12997 ^ n4203 ^ 1'b0 ;
  assign n29321 = n4571 & n25648 ;
  assign n29322 = n13879 | n29321 ;
  assign n29323 = n13213 ^ n12331 ^ 1'b0 ;
  assign n29324 = n22771 ^ n6963 ^ 1'b0 ;
  assign n29325 = ( n4122 & ~n19052 ) | ( n4122 & n21008 ) | ( ~n19052 & n21008 ) ;
  assign n29326 = n29325 ^ n8888 ^ 1'b0 ;
  assign n29327 = n29324 & n29326 ;
  assign n29328 = n14994 | n20883 ;
  assign n29329 = n12242 & n18141 ;
  assign n29330 = n10547 ^ n6816 ^ 1'b0 ;
  assign n29331 = n11854 & ~n29330 ;
  assign n29332 = ~n3069 & n7559 ;
  assign n29333 = ~n29331 & n29332 ;
  assign n29334 = n5756 | n19775 ;
  assign n29335 = n3713 & ~n4544 ;
  assign n29336 = ~n4464 & n6005 ;
  assign n29337 = n4217 & ~n29336 ;
  assign n29338 = ~n7888 & n20993 ;
  assign n29339 = n3223 | n18041 ;
  assign n29340 = n29208 & n29339 ;
  assign n29341 = n1663 & ~n23327 ;
  assign n29345 = n4398 & ~n5828 ;
  assign n29344 = ~n10808 & n21932 ;
  assign n29342 = ~n12766 & n28373 ;
  assign n29343 = n29342 ^ n28797 ^ 1'b0 ;
  assign n29346 = n29345 ^ n29344 ^ n29343 ;
  assign n29347 = ( ~n11987 & n17535 ) | ( ~n11987 & n29346 ) | ( n17535 & n29346 ) ;
  assign n29348 = n8809 & ~n11816 ;
  assign n29349 = ~n25231 & n25838 ;
  assign n29350 = n27089 ^ n2505 ^ 1'b0 ;
  assign n29351 = ~n1130 & n18916 ;
  assign n29352 = n29351 ^ n27628 ^ 1'b0 ;
  assign n29353 = n24717 | n29352 ;
  assign n29354 = ~n4228 & n8551 ;
  assign n29355 = n9759 ^ n5105 ^ 1'b0 ;
  assign n29356 = n3527 & n7557 ;
  assign n29357 = n29356 ^ x231 ^ 1'b0 ;
  assign n29358 = n10767 & ~n29357 ;
  assign n29359 = ~n24284 & n29358 ;
  assign n29360 = n18067 & n26598 ;
  assign n29361 = n11927 & n29360 ;
  assign n29362 = ~n3657 & n26037 ;
  assign n29363 = n29362 ^ n16217 ^ 1'b0 ;
  assign n29364 = n21008 ^ n10437 ^ 1'b0 ;
  assign n29365 = n14338 & ~n29364 ;
  assign n29366 = n5755 ^ n3123 ^ 1'b0 ;
  assign n29367 = ~n20138 & n29366 ;
  assign n29368 = ~n15061 & n29367 ;
  assign n29369 = n24927 ^ n11720 ^ 1'b0 ;
  assign n29370 = n28639 | n29369 ;
  assign n29371 = n19279 ^ n13644 ^ n3064 ;
  assign n29372 = n16164 ^ n5637 ^ 1'b0 ;
  assign n29373 = n17597 ^ n17364 ^ 1'b0 ;
  assign n29374 = n1099 ^ x182 ^ 1'b0 ;
  assign n29375 = ~n17361 & n29374 ;
  assign n29376 = n1974 & n9483 ;
  assign n29377 = ~n1805 & n29376 ;
  assign n29378 = ~n14103 & n17409 ;
  assign n29379 = n29378 ^ n12894 ^ 1'b0 ;
  assign n29380 = n25596 ^ n8927 ^ 1'b0 ;
  assign n29381 = n8225 & ~n12241 ;
  assign n29382 = n24052 & ~n26376 ;
  assign n29383 = n4493 ^ n1324 ^ 1'b0 ;
  assign n29384 = n3392 | n8257 ;
  assign n29385 = n29383 | n29384 ;
  assign n29386 = n6464 ^ n4753 ^ 1'b0 ;
  assign n29387 = n23132 & n29386 ;
  assign n29388 = n29387 ^ n14866 ^ 1'b0 ;
  assign n29389 = n11242 & n27591 ;
  assign n29390 = ~n573 & n13109 ;
  assign n29391 = n29390 ^ n13203 ^ 1'b0 ;
  assign n29392 = n16221 & n29391 ;
  assign n29393 = ~n12407 & n29392 ;
  assign n29394 = n9542 & n24880 ;
  assign n29395 = n977 & n29394 ;
  assign n29396 = n4278 & ~n5865 ;
  assign n29397 = n5821 & n29396 ;
  assign n29398 = n3324 ^ n1925 ^ 1'b0 ;
  assign n29399 = ~n3308 & n29398 ;
  assign n29400 = n29397 & n29399 ;
  assign n29401 = n29400 ^ n9578 ^ 1'b0 ;
  assign n29402 = n1459 | n29401 ;
  assign n29403 = n8045 & n19078 ;
  assign n29404 = n29403 ^ n20228 ^ 1'b0 ;
  assign n29405 = ~n6995 & n29404 ;
  assign n29406 = n2115 & ~n8548 ;
  assign n29407 = ~n29405 & n29406 ;
  assign n29409 = ~n2853 & n5261 ;
  assign n29408 = ~n3768 & n15139 ;
  assign n29410 = n29409 ^ n29408 ^ 1'b0 ;
  assign n29411 = ~n5277 & n5846 ;
  assign n29412 = n29411 ^ n1424 ^ 1'b0 ;
  assign n29413 = n23136 | n29412 ;
  assign n29414 = n20198 ^ x160 ^ 1'b0 ;
  assign n29415 = n9877 | n29414 ;
  assign n29416 = n8564 | n29415 ;
  assign n29417 = n6858 ^ n3024 ^ 1'b0 ;
  assign n29418 = n22567 & n29417 ;
  assign n29419 = n29418 ^ n21096 ^ 1'b0 ;
  assign n29420 = n21018 | n23722 ;
  assign n29423 = n16206 ^ n10753 ^ 1'b0 ;
  assign n29421 = n6834 | n15302 ;
  assign n29422 = n10316 | n29421 ;
  assign n29424 = n29423 ^ n29422 ^ n7281 ;
  assign n29425 = n4398 & ~n24499 ;
  assign n29426 = n29425 ^ n7043 ^ 1'b0 ;
  assign n29427 = n5141 & ~n14818 ;
  assign n29428 = n29427 ^ n7659 ^ 1'b0 ;
  assign n29429 = n6296 | n29428 ;
  assign n29430 = n13523 & ~n23005 ;
  assign n29431 = n29430 ^ n14941 ^ 1'b0 ;
  assign n29432 = n28528 & n29431 ;
  assign n29433 = n4122 ^ n2015 ^ 1'b0 ;
  assign n29434 = n1661 & ~n29433 ;
  assign n29435 = n7415 ^ n3480 ^ 1'b0 ;
  assign n29436 = ~n11856 & n29435 ;
  assign n29437 = n11803 ^ x93 ^ 1'b0 ;
  assign n29438 = n13916 & n29437 ;
  assign n29439 = n15463 & n29438 ;
  assign n29440 = n21174 & ~n28912 ;
  assign n29441 = x155 & n18189 ;
  assign n29442 = ~n12613 & n16074 ;
  assign n29443 = n12754 & n29442 ;
  assign n29444 = n6484 | n29441 ;
  assign n29445 = n23075 & ~n28884 ;
  assign n29446 = n15856 ^ n2451 ^ 1'b0 ;
  assign n29447 = ~n22313 & n29446 ;
  assign n29448 = x166 | n1557 ;
  assign n29449 = n3348 | n5702 ;
  assign n29450 = n29449 ^ n29208 ^ 1'b0 ;
  assign n29451 = n4261 & ~n8518 ;
  assign n29452 = ( ~n1007 & n2436 ) | ( ~n1007 & n29451 ) | ( n2436 & n29451 ) ;
  assign n29453 = ~n12867 & n24852 ;
  assign n29454 = n19089 ^ n12824 ^ 1'b0 ;
  assign n29455 = n1656 & n29454 ;
  assign n29456 = ~n17302 & n29455 ;
  assign n29457 = ~n12980 & n14643 ;
  assign n29458 = ~n2604 & n13998 ;
  assign n29459 = ~n14355 & n29458 ;
  assign n29460 = n29459 ^ n6740 ^ 1'b0 ;
  assign n29461 = n17218 | n23979 ;
  assign n29462 = n7314 ^ n6621 ^ 1'b0 ;
  assign n29463 = n10240 & ~n29462 ;
  assign n29464 = n20627 ^ n13248 ^ 1'b0 ;
  assign n29465 = n18342 & ~n18402 ;
  assign n29466 = n10809 | n12329 ;
  assign n29467 = n9941 & ~n29466 ;
  assign n29468 = n18236 & n29467 ;
  assign n29469 = n4160 | n15667 ;
  assign n29470 = n2273 & ~n24152 ;
  assign n29471 = ~n15990 & n29470 ;
  assign n29472 = n3184 | n13756 ;
  assign n29473 = n5575 & ~n29472 ;
  assign n29474 = n4364 & ~n29473 ;
  assign n29475 = n8333 ^ n8068 ^ 1'b0 ;
  assign n29476 = n2990 & n3198 ;
  assign n29477 = ~n3433 & n6014 ;
  assign n29478 = ~n2521 & n29477 ;
  assign n29479 = n12898 & ~n29478 ;
  assign n29480 = n16233 ^ n4803 ^ 1'b0 ;
  assign n29481 = n25311 ^ n1808 ^ 1'b0 ;
  assign n29482 = n7501 & n29481 ;
  assign n29483 = n29482 ^ n10284 ^ 1'b0 ;
  assign n29484 = n16420 | n23547 ;
  assign n29485 = n29484 ^ n17499 ^ 1'b0 ;
  assign n29486 = n2624 & n24996 ;
  assign n29487 = n11924 ^ n7251 ^ 1'b0 ;
  assign n29488 = n8733 & n18892 ;
  assign n29489 = n18229 | n24301 ;
  assign n29490 = n4822 & ~n14374 ;
  assign n29491 = n1152 & n24551 ;
  assign n29492 = n1268 & ~n5750 ;
  assign n29493 = ~n11778 & n29492 ;
  assign n29494 = ~n944 & n7202 ;
  assign n29495 = n6817 | n17390 ;
  assign n29496 = n1457 & ~n2491 ;
  assign n29497 = ~n2185 & n29496 ;
  assign n29501 = n8635 & ~n12781 ;
  assign n29500 = n1657 | n13659 ;
  assign n29502 = n29501 ^ n29500 ^ 1'b0 ;
  assign n29498 = x150 & n7266 ;
  assign n29499 = n694 | n29498 ;
  assign n29503 = n29502 ^ n29499 ^ 1'b0 ;
  assign n29504 = n28082 ^ n1983 ^ 1'b0 ;
  assign n29505 = ~n24298 & n29504 ;
  assign n29506 = n15297 & n19130 ;
  assign n29507 = ( n1440 & n8430 ) | ( n1440 & ~n29506 ) | ( n8430 & ~n29506 ) ;
  assign n29508 = n20081 & ~n29507 ;
  assign n29509 = n10988 ^ n827 ^ 1'b0 ;
  assign n29510 = n2175 & n29509 ;
  assign n29511 = n12306 & ~n13656 ;
  assign n29512 = n4917 | n29511 ;
  assign n29513 = n4358 | n8399 ;
  assign n29514 = n29513 ^ n16708 ^ 1'b0 ;
  assign n29515 = ~n7314 & n29514 ;
  assign n29516 = ~n2486 & n29515 ;
  assign n29517 = n29516 ^ n19822 ^ 1'b0 ;
  assign n29518 = n29517 ^ n17554 ^ 1'b0 ;
  assign n29519 = n17952 & n29518 ;
  assign n29520 = n29519 ^ n1199 ^ 1'b0 ;
  assign n29521 = n2315 ^ n1344 ^ 1'b0 ;
  assign n29522 = n13850 & ~n29521 ;
  assign n29523 = ~n10969 & n29177 ;
  assign n29524 = n6158 & n29523 ;
  assign n29525 = ~n12841 & n18619 ;
  assign n29526 = n15960 | n29525 ;
  assign n29527 = n29526 ^ n13255 ^ 1'b0 ;
  assign n29528 = n27624 ^ n13613 ^ 1'b0 ;
  assign n29529 = ~n26718 & n29528 ;
  assign n29530 = ( n7060 & n26508 ) | ( n7060 & n28977 ) | ( n26508 & n28977 ) ;
  assign n29531 = n23353 ^ n22229 ^ 1'b0 ;
  assign n29532 = ~n9001 & n11689 ;
  assign n29533 = n5592 & ~n29532 ;
  assign n29535 = n24643 ^ n4814 ^ 1'b0 ;
  assign n29534 = n4896 | n5870 ;
  assign n29536 = n29535 ^ n29534 ^ 1'b0 ;
  assign n29537 = n10450 | n14933 ;
  assign n29538 = n11388 & ~n24735 ;
  assign n29539 = n5922 & n11431 ;
  assign n29540 = n5695 & n24673 ;
  assign n29541 = n20916 ^ n6498 ^ 1'b0 ;
  assign n29542 = n20705 ^ n3933 ^ 1'b0 ;
  assign n29544 = n698 ^ x6 ^ 1'b0 ;
  assign n29543 = ~n10441 & n20607 ;
  assign n29545 = n29544 ^ n29543 ^ 1'b0 ;
  assign n29546 = ( n10908 & ~n29542 ) | ( n10908 & n29545 ) | ( ~n29542 & n29545 ) ;
  assign n29547 = n7836 & n28530 ;
  assign n29548 = n15748 | n16608 ;
  assign n29549 = n29548 ^ n1646 ^ 1'b0 ;
  assign n29550 = ( n2054 & n5768 ) | ( n2054 & n10898 ) | ( n5768 & n10898 ) ;
  assign n29551 = ( n21064 & n29549 ) | ( n21064 & n29550 ) | ( n29549 & n29550 ) ;
  assign n29552 = n8665 | n14572 ;
  assign n29553 = n8915 ^ n2546 ^ n1978 ;
  assign n29554 = n25419 ^ n4385 ^ 1'b0 ;
  assign n29555 = n6056 & n8513 ;
  assign n29556 = n29555 ^ n5354 ^ 1'b0 ;
  assign n29557 = n3343 | n29556 ;
  assign n29558 = n29556 & ~n29557 ;
  assign n29559 = ~n5964 & n6663 ;
  assign n29561 = ~n7296 & n15687 ;
  assign n29560 = n7867 & ~n23504 ;
  assign n29562 = n29561 ^ n29560 ^ 1'b0 ;
  assign n29563 = n5086 & ~n29562 ;
  assign n29564 = n29563 ^ n11299 ^ 1'b0 ;
  assign n29565 = n7650 & n10058 ;
  assign n29566 = x21 & n12386 ;
  assign n29567 = n29566 ^ n8200 ^ 1'b0 ;
  assign n29568 = n5707 | n21224 ;
  assign n29569 = n1354 | n7449 ;
  assign n29570 = n29569 ^ n22330 ^ 1'b0 ;
  assign n29571 = n9815 ^ n4402 ^ 1'b0 ;
  assign n29572 = ~n3340 & n29571 ;
  assign n29573 = ~n1149 & n7918 ;
  assign n29574 = ~n29572 & n29573 ;
  assign n29575 = n3392 | n14977 ;
  assign n29576 = ( ~n6712 & n27341 ) | ( ~n6712 & n29575 ) | ( n27341 & n29575 ) ;
  assign n29577 = n809 & n6111 ;
  assign n29578 = n923 & n29577 ;
  assign n29579 = ~n7098 & n14554 ;
  assign n29580 = n9027 & n29579 ;
  assign n29581 = n29580 ^ n28770 ^ 1'b0 ;
  assign n29582 = n26695 ^ n4553 ^ 1'b0 ;
  assign n29583 = n29582 ^ x196 ^ 1'b0 ;
  assign n29584 = n29583 ^ n24009 ^ 1'b0 ;
  assign n29585 = x130 | n29584 ;
  assign n29586 = n12037 & ~n29585 ;
  assign n29587 = n3181 & ~n12028 ;
  assign n29588 = n3710 & n28797 ;
  assign n29589 = n29588 ^ n3349 ^ 1'b0 ;
  assign n29590 = n15872 ^ n5217 ^ 1'b0 ;
  assign n29591 = n12033 & ~n29590 ;
  assign n29592 = n781 | n6152 ;
  assign n29593 = n29591 & n29592 ;
  assign n29594 = n29593 ^ n9734 ^ 1'b0 ;
  assign n29595 = n23810 | n29594 ;
  assign n29596 = n5577 | n6742 ;
  assign n29597 = n29596 ^ n24391 ^ 1'b0 ;
  assign n29598 = n25293 ^ n20622 ^ 1'b0 ;
  assign n29599 = ~n7700 & n29598 ;
  assign n29600 = n22312 ^ n18423 ^ 1'b0 ;
  assign n29601 = ~n5426 & n13388 ;
  assign n29602 = n2022 & n29601 ;
  assign n29603 = n8578 ^ n1575 ^ 1'b0 ;
  assign n29604 = n26500 | n29603 ;
  assign n29605 = n17024 & n18164 ;
  assign n29606 = n13129 & n29605 ;
  assign n29607 = n12071 & ~n13527 ;
  assign n29608 = n3636 & ~n7115 ;
  assign n29609 = n12087 ^ n8408 ^ 1'b0 ;
  assign n29610 = n5316 & ~n29609 ;
  assign n29611 = n29610 ^ n9454 ^ 1'b0 ;
  assign n29612 = ~n29608 & n29611 ;
  assign n29613 = n11584 ^ n7133 ^ 1'b0 ;
  assign n29614 = n9132 ^ n6478 ^ 1'b0 ;
  assign n29615 = n29613 | n29614 ;
  assign n29616 = n29615 ^ n15568 ^ 1'b0 ;
  assign n29617 = ( x73 & ~n2492 ) | ( x73 & n6557 ) | ( ~n2492 & n6557 ) ;
  assign n29618 = n8002 & n29617 ;
  assign n29619 = n29618 ^ n5958 ^ 1'b0 ;
  assign n29620 = n29619 ^ n8229 ^ 1'b0 ;
  assign n29621 = n29616 | n29620 ;
  assign n29622 = ~x60 & n7945 ;
  assign n29623 = n29622 ^ n7769 ^ 1'b0 ;
  assign n29624 = n29623 ^ n5615 ^ n4258 ;
  assign n29625 = n9032 & ~n14298 ;
  assign n29626 = ~n8685 & n9624 ;
  assign n29627 = n29625 | n29626 ;
  assign n29628 = n5837 & ~n10318 ;
  assign n29629 = n29628 ^ n3622 ^ 1'b0 ;
  assign n29630 = ( n2846 & n20868 ) | ( n2846 & ~n29629 ) | ( n20868 & ~n29629 ) ;
  assign n29631 = x115 & ~n9461 ;
  assign n29632 = n9269 & n29631 ;
  assign n29633 = n2058 & n16889 ;
  assign n29634 = n29633 ^ n5635 ^ 1'b0 ;
  assign n29635 = n9964 & ~n11655 ;
  assign n29636 = ~n29634 & n29635 ;
  assign n29637 = n10194 | n14274 ;
  assign n29638 = n14661 ^ n2426 ^ 1'b0 ;
  assign n29639 = n29638 ^ n15564 ^ 1'b0 ;
  assign n29640 = n26309 & ~n29639 ;
  assign n29644 = n1623 & n7407 ;
  assign n29645 = n2071 & n29644 ;
  assign n29643 = n19386 & n29563 ;
  assign n29646 = n29645 ^ n29643 ^ 1'b0 ;
  assign n29641 = n13194 ^ n8821 ^ 1'b0 ;
  assign n29642 = n12456 | n29641 ;
  assign n29647 = n29646 ^ n29642 ^ 1'b0 ;
  assign n29650 = ( n3606 & ~n13160 ) | ( n3606 & n13262 ) | ( ~n13160 & n13262 ) ;
  assign n29648 = n12919 ^ n7079 ^ 1'b0 ;
  assign n29649 = n2340 | n29648 ;
  assign n29651 = n29650 ^ n29649 ^ 1'b0 ;
  assign n29652 = n1751 | n19586 ;
  assign n29653 = n5984 & ~n29652 ;
  assign n29654 = n29653 ^ n994 ^ 1'b0 ;
  assign n29655 = n29124 & ~n29654 ;
  assign n29656 = n8458 & ~n21184 ;
  assign n29657 = ~n25579 & n29656 ;
  assign n29658 = n12089 ^ n2486 ^ 1'b0 ;
  assign n29659 = n14602 ^ n1240 ^ 1'b0 ;
  assign n29660 = ~n14759 & n29659 ;
  assign n29661 = n29660 ^ x139 ^ 1'b0 ;
  assign n29662 = n12686 ^ n730 ^ 1'b0 ;
  assign n29663 = n13084 ^ n421 ^ 1'b0 ;
  assign n29664 = n10465 & n29663 ;
  assign n29665 = ~n29662 & n29664 ;
  assign n29666 = n8954 & n10997 ;
  assign n29667 = ~n8954 & n29666 ;
  assign n29668 = n29667 ^ n10044 ^ n4002 ;
  assign n29669 = n9565 & ~n24926 ;
  assign n29670 = n29668 & n29669 ;
  assign n29671 = n1646 & n18315 ;
  assign n29672 = n1470 | n1575 ;
  assign n29673 = n29672 ^ n29208 ^ n4092 ;
  assign n29674 = n3781 & ~n29673 ;
  assign n29675 = n29674 ^ n4112 ^ 1'b0 ;
  assign n29677 = ~n6067 & n8145 ;
  assign n29678 = n2670 & n29677 ;
  assign n29679 = n29678 ^ n6682 ^ 1'b0 ;
  assign n29680 = n5411 & n17588 ;
  assign n29681 = n29679 & n29680 ;
  assign n29676 = n5490 | n10681 ;
  assign n29682 = n29681 ^ n29676 ^ 1'b0 ;
  assign n29683 = n9144 | n12753 ;
  assign n29684 = n20662 & ~n29683 ;
  assign n29685 = ~n1651 & n9681 ;
  assign n29686 = n13142 ^ n4031 ^ 1'b0 ;
  assign n29687 = ~n29685 & n29686 ;
  assign n29688 = n28589 ^ n13207 ^ n6570 ;
  assign n29689 = n8679 & n11255 ;
  assign n29690 = n5945 | n17466 ;
  assign n29691 = n10379 ^ n4217 ^ 1'b0 ;
  assign n29692 = n1890 & n29691 ;
  assign n29695 = n3905 & ~n20321 ;
  assign n29696 = n29695 ^ n8760 ^ 1'b0 ;
  assign n29693 = n19469 ^ n4813 ^ 1'b0 ;
  assign n29694 = n11165 & n29693 ;
  assign n29697 = n29696 ^ n29694 ^ 1'b0 ;
  assign n29698 = x238 & ~n918 ;
  assign n29699 = ~n11796 & n29698 ;
  assign n29700 = n28901 & n29699 ;
  assign n29701 = n29700 ^ n11829 ^ 1'b0 ;
  assign n29702 = n20672 ^ n18766 ^ 1'b0 ;
  assign n29703 = n2029 ^ n1920 ^ 1'b0 ;
  assign n29704 = n628 | n29703 ;
  assign n29705 = n9646 & n29704 ;
  assign n29706 = n29705 ^ n20145 ^ 1'b0 ;
  assign n29707 = n13671 & ~n29706 ;
  assign n29708 = n4048 & ~n14859 ;
  assign n29709 = n5473 ^ n3981 ^ 1'b0 ;
  assign n29710 = n29709 ^ n15216 ^ 1'b0 ;
  assign n29711 = n29708 & ~n29710 ;
  assign n29712 = n11851 | n29711 ;
  assign n29713 = n4115 | n9869 ;
  assign n29714 = n9027 ^ n1299 ^ 1'b0 ;
  assign n29715 = n29714 ^ n4103 ^ 1'b0 ;
  assign n29716 = n22182 ^ n3488 ^ 1'b0 ;
  assign n29717 = n15575 ^ n14913 ^ 1'b0 ;
  assign n29718 = n18661 & n29717 ;
  assign n29719 = ~n13785 & n29718 ;
  assign n29720 = ~n18479 & n19464 ;
  assign n29721 = n29720 ^ n15824 ^ n988 ;
  assign n29731 = n15866 ^ n11914 ^ 1'b0 ;
  assign n29722 = n1597 | n2806 ;
  assign n29723 = n2806 & ~n29722 ;
  assign n29724 = n29723 ^ n12257 ^ 1'b0 ;
  assign n29725 = n22925 ^ n15927 ^ 1'b0 ;
  assign n29726 = n29724 & ~n29725 ;
  assign n29727 = ~n1694 & n10580 ;
  assign n29728 = ~n10580 & n29727 ;
  assign n29729 = n29728 ^ n6471 ^ 1'b0 ;
  assign n29730 = n29726 & ~n29729 ;
  assign n29732 = n29731 ^ n29730 ^ 1'b0 ;
  assign n29733 = n772 & n5645 ;
  assign n29734 = ~n5645 & n29733 ;
  assign n29735 = n6267 | n29734 ;
  assign n29736 = n2822 & ~n7154 ;
  assign n29737 = ~n10108 & n29736 ;
  assign n29738 = ~n29736 & n29737 ;
  assign n29739 = n29735 | n29738 ;
  assign n29740 = n29739 ^ n17790 ^ 1'b0 ;
  assign n29741 = n6421 | n16776 ;
  assign n29742 = n832 & ~n1589 ;
  assign n29743 = n29742 ^ n11758 ^ 1'b0 ;
  assign n29744 = n15515 ^ n4265 ^ 1'b0 ;
  assign n29745 = n4576 ^ n500 ^ 1'b0 ;
  assign n29746 = n5796 & ~n10619 ;
  assign n29747 = n29746 ^ n28265 ^ n2072 ;
  assign n29748 = n472 & ~n6194 ;
  assign n29749 = n29748 ^ n17135 ^ 1'b0 ;
  assign n29750 = n22526 & ~n29749 ;
  assign n29751 = n7628 & ~n14580 ;
  assign n29752 = n5942 ^ n3793 ^ 1'b0 ;
  assign n29753 = ~n9461 & n29752 ;
  assign n29754 = n29753 ^ n26547 ^ n4094 ;
  assign n29755 = n3195 ^ n2870 ^ 1'b0 ;
  assign n29756 = ~n2087 & n14938 ;
  assign n29757 = ~n16144 & n21995 ;
  assign n29758 = n11910 ^ n5398 ^ 1'b0 ;
  assign n29759 = n12703 | n29758 ;
  assign n29760 = n1978 & n8234 ;
  assign n29761 = n29760 ^ n3855 ^ 1'b0 ;
  assign n29762 = n29761 ^ n11657 ^ 1'b0 ;
  assign n29763 = n5108 | n23159 ;
  assign n29764 = n4469 ^ n2855 ^ 1'b0 ;
  assign n29765 = ~n12389 & n29764 ;
  assign n29766 = n994 | n29765 ;
  assign n29767 = n27372 | n29766 ;
  assign n29768 = n20963 | n29767 ;
  assign n29769 = n16608 ^ n7266 ^ 1'b0 ;
  assign n29770 = n1724 & ~n29769 ;
  assign n29771 = ~n2254 & n3800 ;
  assign n29772 = n17981 ^ n1305 ^ 1'b0 ;
  assign n29773 = n29771 & ~n29772 ;
  assign n29774 = n14030 ^ n10764 ^ 1'b0 ;
  assign n29775 = n3611 & ~n13724 ;
  assign n29776 = n29775 ^ n18477 ^ 1'b0 ;
  assign n29777 = n3339 ^ x165 ^ 1'b0 ;
  assign n29778 = n29776 | n29777 ;
  assign n29779 = ~n21442 & n24370 ;
  assign n29780 = n29779 ^ n12703 ^ 1'b0 ;
  assign n29781 = n20514 ^ n12841 ^ 1'b0 ;
  assign n29782 = n3277 & ~n29781 ;
  assign n29783 = n2973 & n29782 ;
  assign n29784 = n29783 ^ n3251 ^ 1'b0 ;
  assign n29785 = ~n16876 & n19364 ;
  assign n29786 = n8259 | n29785 ;
  assign n29787 = ~n13854 & n22938 ;
  assign n29788 = n11491 ^ n990 ^ 1'b0 ;
  assign n29789 = n5607 & n5776 ;
  assign n29790 = n29789 ^ n11806 ^ n7667 ;
  assign n29791 = x9 & ~n1831 ;
  assign n29792 = n16580 ^ n12807 ^ 1'b0 ;
  assign n29793 = n29792 ^ n12298 ^ 1'b0 ;
  assign n29794 = n29791 & ~n29793 ;
  assign n29795 = n1152 | n4257 ;
  assign n29796 = n29795 ^ n9612 ^ 1'b0 ;
  assign n29797 = n919 | n2283 ;
  assign n29798 = n1910 & ~n29797 ;
  assign n29799 = n19613 | n29798 ;
  assign n29800 = ~n1988 & n19728 ;
  assign n29801 = n1724 & ~n29800 ;
  assign n29802 = ~n12473 & n29801 ;
  assign n29803 = n8095 & n29802 ;
  assign n29804 = n10728 & ~n11301 ;
  assign n29805 = n27780 | n29804 ;
  assign n29806 = n29803 & ~n29805 ;
  assign n29807 = n11612 & n24792 ;
  assign n29808 = n17195 | n19867 ;
  assign n29809 = ~n13676 & n23230 ;
  assign n29810 = ~n2553 & n12772 ;
  assign n29811 = n29809 & n29810 ;
  assign n29812 = n12247 ^ n7449 ^ 1'b0 ;
  assign n29813 = n2392 & ~n11217 ;
  assign n29814 = n10290 | n29813 ;
  assign n29815 = n3370 & ~n7478 ;
  assign n29816 = n29815 ^ n6189 ^ 1'b0 ;
  assign n29817 = n3577 & n29816 ;
  assign n29818 = n4172 & n8203 ;
  assign n29819 = n14461 | n20676 ;
  assign n29820 = n29819 ^ n25777 ^ 1'b0 ;
  assign n29821 = n1578 ^ x25 ^ 1'b0 ;
  assign n29822 = n19521 & ~n29821 ;
  assign n29823 = ~n28601 & n29822 ;
  assign n29824 = n29823 ^ n12136 ^ 1'b0 ;
  assign n29825 = n3794 | n3926 ;
  assign n29826 = n2476 | n10437 ;
  assign n29827 = n4580 & ~n29826 ;
  assign n29828 = n29827 ^ n8507 ^ n8237 ;
  assign n29829 = n4267 & n29828 ;
  assign n29832 = ~n8390 & n20841 ;
  assign n29830 = n6522 & n12581 ;
  assign n29831 = n29830 ^ n5308 ^ 1'b0 ;
  assign n29833 = n29832 ^ n29831 ^ n3624 ;
  assign n29834 = n4827 & n23038 ;
  assign n29835 = n10604 & n29834 ;
  assign n29836 = n4059 ^ n1094 ^ 1'b0 ;
  assign n29837 = n19592 & n29836 ;
  assign n29838 = n29837 ^ n24831 ^ 1'b0 ;
  assign n29839 = n11272 ^ n4656 ^ 1'b0 ;
  assign n29840 = ~n12452 & n17322 ;
  assign n29841 = n3877 & ~n6149 ;
  assign n29842 = n9249 ^ n7800 ^ 1'b0 ;
  assign n29843 = n13052 ^ n7668 ^ 1'b0 ;
  assign n29844 = n16351 & ~n23228 ;
  assign n29845 = n29844 ^ n3355 ^ 1'b0 ;
  assign n29846 = n2076 & n26642 ;
  assign n29847 = n29846 ^ n19744 ^ 1'b0 ;
  assign n29848 = n430 & n3721 ;
  assign n29849 = n9910 ^ n8619 ^ 1'b0 ;
  assign n29851 = n7769 ^ n1818 ^ 1'b0 ;
  assign n29850 = x74 & n28917 ;
  assign n29852 = n29851 ^ n29850 ^ 1'b0 ;
  assign n29853 = n5861 ^ n1490 ^ 1'b0 ;
  assign n29854 = ~n13038 & n29853 ;
  assign n29855 = n4727 | n8944 ;
  assign n29856 = n17143 | n29855 ;
  assign n29857 = n6431 & n29856 ;
  assign n29858 = n1170 & ~n1172 ;
  assign n29859 = n29858 ^ n9364 ^ n2350 ;
  assign n29868 = n964 & ~n1391 ;
  assign n29869 = ~n964 & n29868 ;
  assign n29870 = n3694 & ~n29869 ;
  assign n29861 = ~n4661 & n6271 ;
  assign n29862 = n4661 & n29861 ;
  assign n29863 = n8525 | n29862 ;
  assign n29864 = n8525 & ~n29863 ;
  assign n29865 = n29864 ^ n15003 ^ 1'b0 ;
  assign n29866 = n14449 & ~n29865 ;
  assign n29867 = ~n14449 & n29866 ;
  assign n29871 = n29870 ^ n29867 ^ 1'b0 ;
  assign n29860 = n25782 ^ n8879 ^ 1'b0 ;
  assign n29872 = n29871 ^ n29860 ^ 1'b0 ;
  assign n29873 = ~n2071 & n29872 ;
  assign n29874 = n5146 & n29873 ;
  assign n29875 = n7590 & ~n14829 ;
  assign n29876 = ~n19977 & n28765 ;
  assign n29877 = ~n2807 & n29876 ;
  assign n29878 = n12854 | n13180 ;
  assign n29879 = n5450 & ~n29878 ;
  assign n29880 = ~n2179 & n9264 ;
  assign n29881 = ~n15280 & n29880 ;
  assign n29882 = n1832 & n28543 ;
  assign n29883 = ~n20048 & n29882 ;
  assign n29884 = n15380 & ~n21930 ;
  assign n29885 = n8728 & ~n20907 ;
  assign n29886 = n29885 ^ x178 ^ 1'b0 ;
  assign n29887 = n13053 & ~n26172 ;
  assign n29888 = ~n9123 & n16731 ;
  assign n29889 = n5116 & n9380 ;
  assign n29890 = n14477 | n23129 ;
  assign n29892 = n3463 | n21691 ;
  assign n29891 = n2333 | n2743 ;
  assign n29893 = n29892 ^ n29891 ^ 1'b0 ;
  assign n29894 = n2330 | n21761 ;
  assign n29895 = n29894 ^ n3540 ^ 1'b0 ;
  assign n29896 = n9696 | n15579 ;
  assign n29897 = n24003 | n29896 ;
  assign n29898 = n19508 ^ n7358 ^ n5728 ;
  assign n29899 = n16333 ^ n2445 ^ 1'b0 ;
  assign n29900 = n29898 & n29899 ;
  assign n29901 = n7692 & ~n9794 ;
  assign n29902 = n16012 & ~n28926 ;
  assign n29903 = n29902 ^ n28940 ^ 1'b0 ;
  assign n29904 = n3751 | n15019 ;
  assign n29905 = n16327 | n29904 ;
  assign n29906 = n14608 ^ n12667 ^ 1'b0 ;
  assign n29907 = n18558 & ~n29906 ;
  assign n29908 = ~n29905 & n29907 ;
  assign n29909 = n428 ^ x199 ^ 1'b0 ;
  assign n29910 = n19282 | n29909 ;
  assign n29911 = ~n1782 & n3988 ;
  assign n29912 = n8305 & n29911 ;
  assign n29913 = ~n14481 & n29912 ;
  assign n29914 = n18862 ^ n14981 ^ 1'b0 ;
  assign n29915 = n29914 ^ n8138 ^ 1'b0 ;
  assign n29916 = ~n23721 & n29915 ;
  assign n29917 = ~n1216 & n24874 ;
  assign n29918 = ~n28325 & n29917 ;
  assign n29919 = n7667 ^ x72 ^ 1'b0 ;
  assign n29920 = n2576 & ~n8821 ;
  assign n29921 = n8808 & ~n26626 ;
  assign n29922 = ( n11402 & ~n15090 ) | ( n11402 & n19387 ) | ( ~n15090 & n19387 ) ;
  assign n29923 = ~n19871 & n29922 ;
  assign n29924 = n1546 & ~n6786 ;
  assign n29925 = n15952 | n20460 ;
  assign n29926 = ~n7357 & n12273 ;
  assign n29927 = n29926 ^ n3272 ^ 1'b0 ;
  assign n29928 = n27295 | n29927 ;
  assign n29929 = n1474 & n10214 ;
  assign n29930 = n12971 ^ n6100 ^ 1'b0 ;
  assign n29931 = n21636 & n29930 ;
  assign n29932 = n6049 & n29931 ;
  assign n29933 = n21404 ^ n5988 ^ 1'b0 ;
  assign n29934 = n25130 & n29933 ;
  assign n29935 = n9941 | n13483 ;
  assign n29936 = n8734 ^ n827 ^ 1'b0 ;
  assign n29937 = n29936 ^ n17882 ^ 1'b0 ;
  assign n29938 = x94 & ~n29937 ;
  assign n29939 = n29938 ^ n14967 ^ 1'b0 ;
  assign n29940 = ~n29935 & n29939 ;
  assign n29941 = n3953 | n7755 ;
  assign n29942 = n1290 & n17094 ;
  assign n29945 = x130 & ~n15007 ;
  assign n29943 = n26271 ^ n8317 ^ x192 ;
  assign n29944 = n9415 & ~n29943 ;
  assign n29946 = n29945 ^ n29944 ^ 1'b0 ;
  assign n29947 = ~n11987 & n12694 ;
  assign n29948 = ( ~n10328 & n28437 ) | ( ~n10328 & n29947 ) | ( n28437 & n29947 ) ;
  assign n29949 = n21693 & ~n28132 ;
  assign n29950 = n1305 & n21230 ;
  assign n29951 = ~n5752 & n8135 ;
  assign n29952 = n6084 & n29951 ;
  assign n29953 = n29952 ^ n10587 ^ 1'b0 ;
  assign n29954 = ~n11427 & n21472 ;
  assign n29955 = n29954 ^ n1160 ^ 1'b0 ;
  assign n29956 = n24628 & ~n26472 ;
  assign n29957 = n994 & n7089 ;
  assign n29958 = n5242 & n29957 ;
  assign n29959 = n7531 & n29958 ;
  assign n29960 = ~n7531 & n29959 ;
  assign n29961 = n14742 ^ n732 ^ 1'b0 ;
  assign n29962 = n29957 & ~n29961 ;
  assign n29963 = n29962 ^ n3678 ^ 1'b0 ;
  assign n29964 = ~n11553 & n29963 ;
  assign n29965 = ~n29960 & n29964 ;
  assign n29966 = n29960 & n29965 ;
  assign n29967 = x208 | n9598 ;
  assign n29968 = n10283 & ~n29967 ;
  assign n29971 = n13492 ^ n11187 ^ n8122 ;
  assign n29969 = n22392 & ~n22993 ;
  assign n29970 = ~n13585 & n29969 ;
  assign n29972 = n29971 ^ n29970 ^ 1'b0 ;
  assign n29973 = n9855 & ~n20082 ;
  assign n29974 = n12026 ^ n4689 ^ 1'b0 ;
  assign n29975 = n29973 & ~n29974 ;
  assign n29976 = ~n1857 & n17820 ;
  assign n29977 = ~n29975 & n29976 ;
  assign n29978 = n29977 ^ n9880 ^ 1'b0 ;
  assign n29979 = n9290 & n17586 ;
  assign n29980 = n29979 ^ n14415 ^ 1'b0 ;
  assign n29981 = n715 & n29980 ;
  assign n29982 = n19533 ^ n16724 ^ 1'b0 ;
  assign n29983 = ~n10652 & n12340 ;
  assign n29984 = n6423 & n29983 ;
  assign n29985 = n10721 & ~n29984 ;
  assign n29986 = n7364 & n29985 ;
  assign n29987 = n22440 | n29986 ;
  assign n29988 = n2343 ^ x109 ^ 1'b0 ;
  assign n29990 = n11433 & n17214 ;
  assign n29989 = x174 & n5139 ;
  assign n29991 = n29990 ^ n29989 ^ 1'b0 ;
  assign n29992 = n10360 | n29991 ;
  assign n29993 = n8010 ^ n3565 ^ 1'b0 ;
  assign n29994 = n11725 & n20680 ;
  assign n29995 = ( n2403 & n3812 ) | ( n2403 & n8969 ) | ( n3812 & n8969 ) ;
  assign n29996 = n9128 ^ n4967 ^ 1'b0 ;
  assign n29997 = n17167 | n29996 ;
  assign n29998 = ~n7373 & n29997 ;
  assign n29999 = n1382 | n11280 ;
  assign n30000 = n4913 & ~n29999 ;
  assign n30001 = n5364 & ~n6400 ;
  assign n30002 = n30001 ^ n25828 ^ 1'b0 ;
  assign n30003 = n23234 & ~n26326 ;
  assign n30004 = ~n4306 & n8110 ;
  assign n30005 = n30004 ^ n5312 ^ 1'b0 ;
  assign n30006 = n4191 & n24343 ;
  assign n30007 = n3181 & ~n6938 ;
  assign n30008 = n4930 & ~n30007 ;
  assign n30009 = ~n24284 & n30008 ;
  assign n30010 = n1832 ^ n1232 ^ 1'b0 ;
  assign n30011 = n3314 & ~n30010 ;
  assign n30014 = n11988 ^ n8559 ^ 1'b0 ;
  assign n30015 = n11130 & ~n30014 ;
  assign n30012 = n7293 | n11392 ;
  assign n30013 = n5571 & ~n30012 ;
  assign n30016 = n30015 ^ n30013 ^ n20824 ;
  assign n30017 = n30011 & n30016 ;
  assign n30018 = x191 | n1017 ;
  assign n30019 = ~n685 & n1661 ;
  assign n30020 = n30019 ^ n16580 ^ 1'b0 ;
  assign n30021 = n29595 | n30020 ;
  assign n30022 = n30021 ^ n17893 ^ 1'b0 ;
  assign n30023 = n13708 & n17554 ;
  assign n30024 = n30023 ^ n6561 ^ 1'b0 ;
  assign n30025 = n3774 & n20312 ;
  assign n30026 = n30025 ^ n18695 ^ 1'b0 ;
  assign n30027 = n1195 & n11983 ;
  assign n30028 = n7933 & n30027 ;
  assign n30029 = ~n11817 & n29096 ;
  assign n30030 = n9550 ^ n8928 ^ 1'b0 ;
  assign n30031 = n24052 & ~n29660 ;
  assign n30032 = n19300 ^ n1402 ^ 1'b0 ;
  assign n30033 = n23473 | n30032 ;
  assign n30034 = n1397 & ~n10955 ;
  assign n30035 = n30034 ^ n23840 ^ 1'b0 ;
  assign n30036 = n18464 ^ n11400 ^ 1'b0 ;
  assign n30037 = n2172 | n30036 ;
  assign n30038 = n450 | n30037 ;
  assign n30039 = ~n6338 & n18461 ;
  assign n30040 = n5012 & n30039 ;
  assign n30041 = n9143 & ~n11649 ;
  assign n30042 = n30041 ^ n15578 ^ 1'b0 ;
  assign n30043 = n4172 & ~n30042 ;
  assign n30044 = n12887 ^ n12726 ^ 1'b0 ;
  assign n30045 = x14 & n30044 ;
  assign n30046 = n3071 & n30045 ;
  assign n30047 = n12302 & ~n24292 ;
  assign n30048 = n1173 | n30047 ;
  assign n30049 = n26882 ^ n2995 ^ 1'b0 ;
  assign n30050 = n12546 | n30049 ;
  assign n30051 = n13804 & ~n26431 ;
  assign n30052 = n30051 ^ n4859 ^ 1'b0 ;
  assign n30053 = n15524 | n24373 ;
  assign n30054 = n6045 | n8902 ;
  assign n30055 = n24976 & n30054 ;
  assign n30056 = n14770 ^ n9451 ^ 1'b0 ;
  assign n30058 = n9253 & n16654 ;
  assign n30059 = ~n5540 & n30058 ;
  assign n30057 = n6676 & n8290 ;
  assign n30060 = n30059 ^ n30057 ^ 1'b0 ;
  assign n30061 = ~n621 & n8390 ;
  assign n30062 = n21482 ^ n19917 ^ 1'b0 ;
  assign n30063 = ~n12805 & n23729 ;
  assign n30064 = n30063 ^ n17156 ^ 1'b0 ;
  assign n30065 = n21820 ^ n15172 ^ 1'b0 ;
  assign n30066 = n593 & n30065 ;
  assign n30067 = n24868 ^ n8111 ^ 1'b0 ;
  assign n30068 = ~n7545 & n30067 ;
  assign n30069 = n13789 ^ n10382 ^ 1'b0 ;
  assign n30070 = n17238 ^ n11927 ^ 1'b0 ;
  assign n30071 = n14788 ^ n2472 ^ 1'b0 ;
  assign n30072 = n924 & ~n30071 ;
  assign n30073 = n8612 & n30072 ;
  assign n30074 = n10915 | n12950 ;
  assign n30075 = n28280 ^ n5290 ^ 1'b0 ;
  assign n30077 = n8041 ^ n2188 ^ 1'b0 ;
  assign n30078 = x236 & ~n30077 ;
  assign n30076 = n11903 & n12596 ;
  assign n30079 = n30078 ^ n30076 ^ 1'b0 ;
  assign n30080 = ~n13426 & n30079 ;
  assign n30081 = n10555 & n17214 ;
  assign n30082 = ( n3364 & n13586 ) | ( n3364 & ~n26771 ) | ( n13586 & ~n26771 ) ;
  assign n30083 = n14414 & ~n28198 ;
  assign n30084 = n30083 ^ n19911 ^ 1'b0 ;
  assign n30085 = ~n6346 & n30084 ;
  assign n30086 = n15101 | n20827 ;
  assign n30087 = n3316 & ~n30086 ;
  assign n30088 = n15031 | n19311 ;
  assign n30089 = n17819 ^ n12563 ^ 1'b0 ;
  assign n30090 = n3179 & n25345 ;
  assign n30091 = ~n11920 & n30090 ;
  assign n30092 = n30091 ^ n4586 ^ 1'b0 ;
  assign n30093 = x27 & ~n4115 ;
  assign n30094 = n10556 | n15362 ;
  assign n30095 = n1818 | n30094 ;
  assign n30096 = n542 & ~n5781 ;
  assign n30097 = n3731 & n30096 ;
  assign n30098 = n30097 ^ n13580 ^ 1'b0 ;
  assign n30099 = n30095 & ~n30098 ;
  assign n30100 = n7810 ^ n2727 ^ x93 ;
  assign n30101 = n13133 | n30100 ;
  assign n30102 = n7446 | n30101 ;
  assign n30103 = n13567 & n30102 ;
  assign n30104 = n7232 & n21435 ;
  assign n30105 = n11965 | n30104 ;
  assign n30106 = ~n6566 & n12245 ;
  assign n30107 = ~n19442 & n30106 ;
  assign n30109 = n7769 ^ n1684 ^ 1'b0 ;
  assign n30108 = n20623 & n27288 ;
  assign n30110 = n30109 ^ n30108 ^ 1'b0 ;
  assign n30111 = n1806 | n2014 ;
  assign n30112 = n2561 & n30111 ;
  assign n30113 = n6874 & ~n10458 ;
  assign n30114 = n30113 ^ n29086 ^ 1'b0 ;
  assign n30115 = n7230 & ~n30114 ;
  assign n30116 = ~n7862 & n28229 ;
  assign n30117 = n3021 | n6050 ;
  assign n30118 = n30117 ^ n17632 ^ n12762 ;
  assign n30119 = x76 & n13297 ;
  assign n30124 = n16880 ^ n13949 ^ 1'b0 ;
  assign n30125 = n11281 ^ n8761 ^ 1'b0 ;
  assign n30126 = ~n30124 & n30125 ;
  assign n30120 = n5052 ^ x178 ^ 1'b0 ;
  assign n30121 = n4118 & n30120 ;
  assign n30122 = ~n9239 & n30121 ;
  assign n30123 = ~n3461 & n30122 ;
  assign n30127 = n30126 ^ n30123 ^ 1'b0 ;
  assign n30128 = n5989 & ~n28204 ;
  assign n30129 = n24917 ^ n24022 ^ 1'b0 ;
  assign n30130 = n17004 ^ n14492 ^ n1521 ;
  assign n30134 = n8836 & ~n20715 ;
  assign n30131 = n14103 ^ n9001 ^ 1'b0 ;
  assign n30132 = n19058 | n30131 ;
  assign n30133 = n7536 | n30132 ;
  assign n30135 = n30134 ^ n30133 ^ 1'b0 ;
  assign n30136 = n16508 & ~n21321 ;
  assign n30137 = ~n4238 & n16506 ;
  assign n30138 = n23549 & n30137 ;
  assign n30139 = n4220 ^ n2460 ^ 1'b0 ;
  assign n30140 = n11427 ^ n6362 ^ 1'b0 ;
  assign n30141 = n345 | n3890 ;
  assign n30142 = n3890 & ~n30141 ;
  assign n30143 = ~n3488 & n30142 ;
  assign n30144 = x33 & ~n481 ;
  assign n30145 = ~x33 & n30144 ;
  assign n30146 = n30143 | n30145 ;
  assign n30147 = n30143 & ~n30146 ;
  assign n30148 = ~n4801 & n30147 ;
  assign n30149 = ~n2944 & n30148 ;
  assign n30150 = ~n4483 & n30149 ;
  assign n30151 = n29705 | n30150 ;
  assign n30152 = n30150 & ~n30151 ;
  assign n30153 = n549 & ~n30152 ;
  assign n30154 = n30152 & n30153 ;
  assign n30155 = n30140 | n30154 ;
  assign n30156 = n30139 & ~n30155 ;
  assign n30157 = n3472 | n17219 ;
  assign n30158 = n1857 | n30157 ;
  assign n30159 = n13590 & ~n30158 ;
  assign n30160 = n18790 ^ n10797 ^ 1'b0 ;
  assign n30161 = n1593 & ~n30160 ;
  assign n30162 = n30159 & n30161 ;
  assign n30163 = n5804 ^ x195 ^ 1'b0 ;
  assign n30164 = n25601 | n30163 ;
  assign n30165 = n5372 & n17897 ;
  assign n30166 = n10178 & n30165 ;
  assign n30167 = ( n1080 & n1499 ) | ( n1080 & n5898 ) | ( n1499 & n5898 ) ;
  assign n30168 = n29832 ^ n4143 ^ 1'b0 ;
  assign n30169 = n17677 & ~n30168 ;
  assign n30170 = n3189 & n19511 ;
  assign n30171 = n27950 ^ n20140 ^ 1'b0 ;
  assign n30172 = n30170 & ~n30171 ;
  assign n30173 = ~n7697 & n30172 ;
  assign n30174 = n30173 ^ n21365 ^ 1'b0 ;
  assign n30175 = n19936 ^ n17754 ^ 1'b0 ;
  assign n30176 = n24736 ^ n1773 ^ 1'b0 ;
  assign n30177 = n8454 & n30176 ;
  assign n30178 = n26666 ^ n13301 ^ 1'b0 ;
  assign n30179 = n2374 | n30178 ;
  assign n30180 = n15626 & n25907 ;
  assign n30181 = ~n7367 & n20627 ;
  assign n30182 = n3298 | n12116 ;
  assign n30183 = n30182 ^ n4385 ^ 1'b0 ;
  assign n30184 = ~n15161 & n30183 ;
  assign n30185 = n5305 & n18468 ;
  assign n30186 = n9788 | n14786 ;
  assign n30187 = n30185 | n30186 ;
  assign n30188 = n20328 & n21444 ;
  assign n30189 = n18491 ^ n2143 ^ x223 ;
  assign n30190 = n30189 ^ n15039 ^ 1'b0 ;
  assign n30191 = n6432 | n30190 ;
  assign n30192 = ~n10795 & n13391 ;
  assign n30193 = x81 & n14171 ;
  assign n30194 = ~n18310 & n24139 ;
  assign n30196 = n5482 & n22997 ;
  assign n30197 = n30196 ^ n17586 ^ 1'b0 ;
  assign n30195 = n20948 & n22249 ;
  assign n30198 = n30197 ^ n30195 ^ 1'b0 ;
  assign n30199 = n11273 ^ n1269 ^ 1'b0 ;
  assign n30200 = x7 & ~n30199 ;
  assign n30201 = n22961 & n30200 ;
  assign n30202 = ( n452 & n2093 ) | ( n452 & ~n10171 ) | ( n2093 & ~n10171 ) ;
  assign n30203 = n30202 ^ n21965 ^ 1'b0 ;
  assign n30204 = n28457 & n30203 ;
  assign n30205 = n2287 ^ n327 ^ 1'b0 ;
  assign n30206 = n28797 ^ n5977 ^ 1'b0 ;
  assign n30207 = n16326 & n30206 ;
  assign n30208 = n29294 ^ n17067 ^ 1'b0 ;
  assign n30209 = n1709 ^ x202 ^ 1'b0 ;
  assign n30210 = n9160 & n18954 ;
  assign n30211 = n11810 & ~n24899 ;
  assign n30212 = n21388 & n30211 ;
  assign n30213 = ~n15091 & n17859 ;
  assign n30214 = n19101 & n30213 ;
  assign n30215 = n30214 ^ n25828 ^ 1'b0 ;
  assign n30216 = n6954 | n14241 ;
  assign n30217 = n2877 | n30216 ;
  assign n30218 = n30217 ^ n25044 ^ n18131 ;
  assign n30219 = ~n13568 & n30218 ;
  assign n30220 = n1271 | n19958 ;
  assign n30221 = n9632 & ~n30220 ;
  assign n30222 = n30221 ^ n1977 ^ 1'b0 ;
  assign n30223 = n11778 ^ n3381 ^ 1'b0 ;
  assign n30224 = n30222 | n30223 ;
  assign n30225 = ~n1672 & n11037 ;
  assign n30226 = n2431 & n13647 ;
  assign n30227 = n3083 & ~n30226 ;
  assign n30228 = ~n12725 & n30227 ;
  assign n30229 = n30228 ^ n1337 ^ 1'b0 ;
  assign n30230 = n18221 | n23559 ;
  assign n30231 = ~n17803 & n19801 ;
  assign n30232 = n30231 ^ n3984 ^ 1'b0 ;
  assign n30233 = n3735 & n5898 ;
  assign n30234 = ~n5512 & n30233 ;
  assign n30235 = n3647 | n30234 ;
  assign n30236 = n8685 | n30235 ;
  assign n30237 = n19577 ^ n4302 ^ 1'b0 ;
  assign n30238 = n1697 & n6661 ;
  assign n30239 = n18228 & ~n30238 ;
  assign n30240 = n30239 ^ n7512 ^ 1'b0 ;
  assign n30241 = n5422 | n13521 ;
  assign n30242 = n5439 | n13269 ;
  assign n30243 = n25916 ^ n12458 ^ 1'b0 ;
  assign n30244 = n11458 & n30243 ;
  assign n30245 = n13226 ^ n10354 ^ 1'b0 ;
  assign n30246 = ~n11237 & n30245 ;
  assign n30247 = ~n13761 & n30246 ;
  assign n30248 = n24113 & n30247 ;
  assign n30257 = n5332 & ~n17717 ;
  assign n30258 = n30257 ^ n5495 ^ 1'b0 ;
  assign n30249 = n2701 & n6740 ;
  assign n30250 = ~n2701 & n30249 ;
  assign n30251 = n9765 | n30250 ;
  assign n30252 = n1366 | n1419 ;
  assign n30253 = n1366 & ~n30252 ;
  assign n30254 = ~n3329 & n30253 ;
  assign n30255 = n12205 | n30254 ;
  assign n30256 = n30251 | n30255 ;
  assign n30259 = n30258 ^ n30256 ^ 1'b0 ;
  assign n30260 = n2877 & n22603 ;
  assign n30261 = n12645 ^ n11354 ^ n2534 ;
  assign n30262 = n313 | n25353 ;
  assign n30263 = n30262 ^ n5675 ^ 1'b0 ;
  assign n30264 = n22385 ^ n7942 ^ 1'b0 ;
  assign n30265 = n3308 | n30264 ;
  assign n30266 = n1688 & ~n12845 ;
  assign n30267 = ~n26840 & n30266 ;
  assign n30268 = ~n2207 & n11989 ;
  assign n30269 = n30268 ^ n7279 ^ 1'b0 ;
  assign n30270 = n30269 ^ n11720 ^ 1'b0 ;
  assign n30271 = n7680 | n10416 ;
  assign n30272 = n30271 ^ n2055 ^ 1'b0 ;
  assign n30273 = n1174 | n10116 ;
  assign n30274 = n7662 ^ n3814 ^ 1'b0 ;
  assign n30275 = n16792 & ~n27905 ;
  assign n30276 = n1939 ^ n1313 ^ 1'b0 ;
  assign n30277 = x212 & ~n30276 ;
  assign n30278 = n30277 ^ n21146 ^ 1'b0 ;
  assign n30279 = n6989 ^ n5176 ^ 1'b0 ;
  assign n30280 = n29295 & n30279 ;
  assign n30281 = n9759 | n30179 ;
  assign n30283 = n16012 ^ n5592 ^ n2264 ;
  assign n30284 = n12213 & ~n30283 ;
  assign n30282 = n1672 | n13159 ;
  assign n30285 = n30284 ^ n30282 ^ 1'b0 ;
  assign n30286 = n7766 & n19830 ;
  assign n30287 = n30286 ^ n2668 ^ 1'b0 ;
  assign n30288 = n9436 & n23213 ;
  assign n30289 = n16161 & ~n20164 ;
  assign n30290 = n30289 ^ n7031 ^ 1'b0 ;
  assign n30291 = n30234 | n30290 ;
  assign n30292 = n1108 | n25428 ;
  assign n30293 = n30292 ^ n18069 ^ 1'b0 ;
  assign n30294 = ~n9384 & n30293 ;
  assign n30295 = ~n17518 & n30294 ;
  assign n30296 = n2761 | n5670 ;
  assign n30297 = n30296 ^ n13647 ^ 1'b0 ;
  assign n30298 = n25556 | n30297 ;
  assign n30299 = n2516 ^ n797 ^ 1'b0 ;
  assign n30300 = n7659 ^ n645 ^ 1'b0 ;
  assign n30301 = n30299 & n30300 ;
  assign n30302 = n30301 ^ n6479 ^ 1'b0 ;
  assign n30303 = n1886 | n22146 ;
  assign n30304 = n30303 ^ n3520 ^ 1'b0 ;
  assign n30305 = n7902 | n30304 ;
  assign n30306 = n30302 & ~n30305 ;
  assign n30307 = n20587 ^ n17570 ^ n9886 ;
  assign n30308 = n3848 ^ n3219 ^ 1'b0 ;
  assign n30309 = ~n26721 & n30308 ;
  assign n30311 = n6381 | n12636 ;
  assign n30312 = n30311 ^ n5201 ^ 1'b0 ;
  assign n30310 = n21352 | n22782 ;
  assign n30313 = n30312 ^ n30310 ^ 1'b0 ;
  assign n30314 = x200 & ~n15250 ;
  assign n30315 = ~n22294 & n30314 ;
  assign n30316 = n30315 ^ n4696 ^ x17 ;
  assign n30317 = n25914 ^ n13886 ^ 1'b0 ;
  assign n30318 = n30316 & n30317 ;
  assign n30319 = n21660 ^ n5176 ^ 1'b0 ;
  assign n30320 = n14428 ^ n1139 ^ 1'b0 ;
  assign n30321 = n3714 & ~n30320 ;
  assign n30322 = n3226 & n6405 ;
  assign n30323 = n30322 ^ n3588 ^ 1'b0 ;
  assign n30324 = n23141 ^ n1638 ^ 1'b0 ;
  assign n30325 = n2809 | n8559 ;
  assign n30326 = n30325 ^ n19309 ^ 1'b0 ;
  assign n30327 = ( ~n7536 & n23978 ) | ( ~n7536 & n30326 ) | ( n23978 & n30326 ) ;
  assign n30328 = n2610 & n30327 ;
  assign n30329 = n30328 ^ n15584 ^ 1'b0 ;
  assign n30330 = ~n13899 & n27563 ;
  assign n30331 = n30330 ^ n10488 ^ 1'b0 ;
  assign n30332 = n8145 & ~n26957 ;
  assign n30333 = ~n30331 & n30332 ;
  assign n30337 = n2487 ^ x155 ^ 1'b0 ;
  assign n30338 = n4190 & ~n30337 ;
  assign n30334 = ~n18677 & n26648 ;
  assign n30335 = n30334 ^ n4810 ^ 1'b0 ;
  assign n30336 = n14448 & ~n30335 ;
  assign n30339 = n30338 ^ n30336 ^ 1'b0 ;
  assign n30340 = x248 & ~n6262 ;
  assign n30341 = n30339 | n30340 ;
  assign n30342 = ( n4600 & n5182 ) | ( n4600 & ~n28378 ) | ( n5182 & ~n28378 ) ;
  assign n30343 = n6001 & ~n10516 ;
  assign n30344 = n30342 & n30343 ;
  assign n30345 = n18806 & n24348 ;
  assign n30346 = ~n15298 & n30345 ;
  assign n30347 = n19756 ^ n9965 ^ 1'b0 ;
  assign n30348 = n14981 ^ n13823 ^ 1'b0 ;
  assign n30349 = n13742 ^ n7408 ^ 1'b0 ;
  assign n30350 = n9951 & n30349 ;
  assign n30351 = n3003 & ~n27992 ;
  assign n30352 = n17762 & n30351 ;
  assign n30353 = n28869 ^ n3499 ^ 1'b0 ;
  assign n30354 = n8969 | n14652 ;
  assign n30355 = n420 & ~n30354 ;
  assign n30356 = n26616 ^ n4406 ^ 1'b0 ;
  assign n30357 = n28622 ^ n4988 ^ n1978 ;
  assign n30358 = n20741 ^ n12309 ^ 1'b0 ;
  assign n30359 = n2250 & n7179 ;
  assign n30360 = n30359 ^ n15175 ^ 1'b0 ;
  assign n30361 = ~n2296 & n30360 ;
  assign n30362 = n30361 ^ n14632 ^ 1'b0 ;
  assign n30363 = n7897 & n30362 ;
  assign n30372 = n13500 ^ n5043 ^ 1'b0 ;
  assign n30371 = ~n1018 & n8226 ;
  assign n30373 = n30372 ^ n30371 ^ 1'b0 ;
  assign n30370 = n7630 & ~n23109 ;
  assign n30374 = n30373 ^ n30370 ^ 1'b0 ;
  assign n30364 = ~n1597 & n4726 ;
  assign n30365 = ~n4726 & n30364 ;
  assign n30366 = ~n2141 & n30365 ;
  assign n30367 = n1196 | n30366 ;
  assign n30368 = n1196 & ~n30367 ;
  assign n30369 = n6031 | n30368 ;
  assign n30375 = n30374 ^ n30369 ^ 1'b0 ;
  assign n30376 = n24103 ^ n1360 ^ 1'b0 ;
  assign n30377 = n2143 & n9013 ;
  assign n30378 = n30377 ^ n17260 ^ 1'b0 ;
  assign n30379 = n7217 & n16485 ;
  assign n30380 = n17955 ^ n12024 ^ 1'b0 ;
  assign n30381 = n30379 & n30380 ;
  assign n30382 = n1521 & n30381 ;
  assign n30383 = n30382 ^ n16898 ^ 1'b0 ;
  assign n30384 = n17460 & ~n30383 ;
  assign n30385 = n30384 ^ n12033 ^ 1'b0 ;
  assign n30386 = n10384 & n19433 ;
  assign n30387 = n30386 ^ n21387 ^ 1'b0 ;
  assign n30391 = n9643 & n15225 ;
  assign n30388 = n18387 ^ n14498 ^ n5619 ;
  assign n30389 = n30388 ^ n1058 ^ 1'b0 ;
  assign n30390 = n7241 & ~n30389 ;
  assign n30392 = n30391 ^ n30390 ^ 1'b0 ;
  assign n30393 = n20499 ^ n15291 ^ 1'b0 ;
  assign n30394 = n11055 ^ n9626 ^ 1'b0 ;
  assign n30395 = ~n2629 & n30394 ;
  assign n30396 = n30395 ^ n18402 ^ 1'b0 ;
  assign n30397 = n5887 & n15447 ;
  assign n30398 = n30397 ^ n4562 ^ 1'b0 ;
  assign n30399 = n10038 & ~n24479 ;
  assign n30400 = n17026 ^ n9539 ^ 1'b0 ;
  assign n30401 = n14053 ^ n9043 ^ 1'b0 ;
  assign n30402 = n12997 & ~n30401 ;
  assign n30403 = n17652 ^ x235 ^ 1'b0 ;
  assign n30404 = n15135 ^ n11976 ^ 1'b0 ;
  assign n30405 = n29766 | n30404 ;
  assign n30406 = n18131 | n19639 ;
  assign n30407 = n8626 ^ n3165 ^ 1'b0 ;
  assign n30408 = n30407 ^ n22114 ^ 1'b0 ;
  assign n30409 = n19445 ^ n12006 ^ 1'b0 ;
  assign n30410 = n2476 & ~n27187 ;
  assign n30411 = n2626 & ~n30410 ;
  assign n30412 = n25445 & n30411 ;
  assign n30413 = n20791 ^ n8532 ^ 1'b0 ;
  assign n30414 = n1378 & n19670 ;
  assign n30415 = n13613 & ~n15168 ;
  assign n30416 = ~n10106 & n30415 ;
  assign n30417 = n19181 ^ n14871 ^ 1'b0 ;
  assign n30418 = n28372 ^ n7898 ^ 1'b0 ;
  assign n30419 = n18215 & ~n28579 ;
  assign n30420 = n3748 & n30419 ;
  assign n30421 = n1518 | n10150 ;
  assign n30422 = n30421 ^ n29509 ^ 1'b0 ;
  assign n30423 = ~n30420 & n30422 ;
  assign n30424 = ~n30418 & n30423 ;
  assign n30425 = ~n2542 & n29852 ;
  assign n30426 = n19363 ^ n6375 ^ 1'b0 ;
  assign n30427 = n4442 | n23855 ;
  assign n30428 = n465 & n30427 ;
  assign n30429 = n30428 ^ n23972 ^ 1'b0 ;
  assign n30430 = n7291 & n8309 ;
  assign n30431 = n22383 | n30430 ;
  assign n30432 = n30431 ^ n3803 ^ 1'b0 ;
  assign n30433 = n13775 & n30432 ;
  assign n30434 = x33 | n6558 ;
  assign n30435 = n16988 | n30434 ;
  assign n30436 = n30435 ^ n26836 ^ 1'b0 ;
  assign n30440 = x87 & n1310 ;
  assign n30441 = ~n1310 & n30440 ;
  assign n30442 = n1670 & n30441 ;
  assign n30443 = ~n320 & n30442 ;
  assign n30444 = n887 & n3441 ;
  assign n30445 = ~n887 & n30444 ;
  assign n30446 = n30443 & ~n30445 ;
  assign n30447 = ~n30443 & n30446 ;
  assign n30437 = n25576 ^ n21288 ^ 1'b0 ;
  assign n30438 = n30437 ^ n10912 ^ 1'b0 ;
  assign n30439 = n16125 & ~n30438 ;
  assign n30448 = n30447 ^ n30439 ^ n24881 ;
  assign n30449 = n10422 | n12621 ;
  assign n30450 = n30449 ^ n26461 ^ 1'b0 ;
  assign n30451 = n996 & ~n9576 ;
  assign n30452 = n9335 & n30451 ;
  assign n30453 = ~n11918 & n30452 ;
  assign n30454 = n30453 ^ n2061 ^ 1'b0 ;
  assign n30455 = ~n3581 & n30454 ;
  assign n30456 = n30455 ^ n28030 ^ 1'b0 ;
  assign n30457 = n22133 ^ n9177 ^ 1'b0 ;
  assign n30458 = n7295 | n30457 ;
  assign n30459 = n1239 & ~n6308 ;
  assign n30460 = ~n4961 & n23734 ;
  assign n30461 = n26409 & n30460 ;
  assign n30462 = ( n5950 & n7291 ) | ( n5950 & n8137 ) | ( n7291 & n8137 ) ;
  assign n30463 = n6586 & ~n27350 ;
  assign n30464 = n16401 & n27959 ;
  assign n30465 = n30464 ^ n26233 ^ 1'b0 ;
  assign n30466 = n20414 ^ n1573 ^ 1'b0 ;
  assign n30467 = n27450 ^ n12177 ^ 1'b0 ;
  assign n30468 = n14598 ^ n12230 ^ 1'b0 ;
  assign n30469 = n15151 & n30468 ;
  assign n30470 = n1402 & ~n30469 ;
  assign n30471 = n10048 & n10864 ;
  assign n30472 = n30471 ^ n26070 ^ 1'b0 ;
  assign n30473 = n13225 & n27164 ;
  assign n30474 = n30473 ^ n5512 ^ 1'b0 ;
  assign n30475 = n5470 | n10985 ;
  assign n30476 = n21551 & ~n23688 ;
  assign n30477 = n30476 ^ n4549 ^ 1'b0 ;
  assign n30478 = n399 & n3793 ;
  assign n30479 = n20669 & ~n30478 ;
  assign n30480 = n22989 | n30479 ;
  assign n30481 = x65 & n1345 ;
  assign n30482 = n30481 ^ n11042 ^ 1'b0 ;
  assign n30483 = ~n30121 & n30482 ;
  assign n30484 = x208 & n3608 ;
  assign n30485 = ~x181 & n30484 ;
  assign n30486 = n12256 & ~n30485 ;
  assign n30487 = n30486 ^ n24234 ^ 1'b0 ;
  assign n30488 = n10685 ^ n5729 ^ 1'b0 ;
  assign n30489 = ~n20617 & n29925 ;
  assign n30490 = n30489 ^ n16028 ^ 1'b0 ;
  assign n30491 = n17201 ^ n7124 ^ 1'b0 ;
  assign n30492 = n5076 ^ n747 ^ 1'b0 ;
  assign n30493 = n7796 & ~n30492 ;
  assign n30494 = ~n3445 & n15498 ;
  assign n30495 = n21509 & ~n30494 ;
  assign n30496 = n21995 | n24041 ;
  assign n30497 = n22919 ^ n2404 ^ 1'b0 ;
  assign n30498 = n18777 | n30497 ;
  assign n30500 = n5692 & n8416 ;
  assign n30501 = n30500 ^ n2057 ^ 1'b0 ;
  assign n30499 = ~n1689 & n24103 ;
  assign n30502 = n30501 ^ n30499 ^ 1'b0 ;
  assign n30503 = ~n8314 & n30502 ;
  assign n30504 = n30498 & n30503 ;
  assign n30505 = ( x226 & n4024 ) | ( x226 & n25348 ) | ( n4024 & n25348 ) ;
  assign n30506 = n20458 | n28213 ;
  assign n30507 = n17777 ^ n9789 ^ 1'b0 ;
  assign n30508 = n22711 ^ n7269 ^ 1'b0 ;
  assign n30509 = n12991 & n26701 ;
  assign n30510 = n7022 ^ n4293 ^ 1'b0 ;
  assign n30511 = ~n5077 & n30510 ;
  assign n30512 = n30511 ^ n20772 ^ 1'b0 ;
  assign n30513 = n8445 & n22786 ;
  assign n30514 = n8049 | n15739 ;
  assign n30515 = n13943 ^ n1339 ^ 1'b0 ;
  assign n30516 = n29085 & n30515 ;
  assign n30517 = n30516 ^ n5818 ^ 1'b0 ;
  assign n30518 = n6427 & n8738 ;
  assign n30519 = n22886 ^ n3416 ^ 1'b0 ;
  assign n30520 = n18045 ^ n7431 ^ 1'b0 ;
  assign n30521 = ~n30519 & n30520 ;
  assign n30522 = ( n8654 & ~n30518 ) | ( n8654 & n30521 ) | ( ~n30518 & n30521 ) ;
  assign n30523 = n24877 ^ n2133 ^ 1'b0 ;
  assign n30524 = n27106 & ~n30523 ;
  assign n30525 = n30524 ^ n16170 ^ 1'b0 ;
  assign n30526 = n21878 | n30525 ;
  assign n30527 = n15239 ^ n5982 ^ 1'b0 ;
  assign n30528 = ~n6134 & n30527 ;
  assign n30530 = n21358 & n21388 ;
  assign n30529 = ~n6879 & n21230 ;
  assign n30531 = n30530 ^ n30529 ^ 1'b0 ;
  assign n30532 = n3661 | n12032 ;
  assign n30533 = n21573 & ~n30532 ;
  assign n30534 = n10327 | n19211 ;
  assign n30535 = n27301 ^ n2909 ^ 1'b0 ;
  assign n30536 = n9879 & n10217 ;
  assign n30537 = n30536 ^ n21911 ^ 1'b0 ;
  assign n30538 = n5634 | n8753 ;
  assign n30539 = n17632 | n22150 ;
  assign n30540 = ~n17817 & n28452 ;
  assign n30541 = ~n3540 & n3868 ;
  assign n30542 = n30540 & n30541 ;
  assign n30543 = n17752 ^ n16291 ^ 1'b0 ;
  assign n30544 = n30543 ^ n19407 ^ 1'b0 ;
  assign n30545 = n29831 | n30544 ;
  assign n30546 = n11616 ^ n1311 ^ 1'b0 ;
  assign n30547 = n11851 & ~n30546 ;
  assign n30548 = n9765 ^ x237 ^ 1'b0 ;
  assign n30549 = n30547 & ~n30548 ;
  assign n30550 = ~n13420 & n17103 ;
  assign n30551 = n20511 ^ n12619 ^ 1'b0 ;
  assign n30552 = n30550 & n30551 ;
  assign n30553 = n6990 ^ n1997 ^ 1'b0 ;
  assign n30554 = n4260 & n30553 ;
  assign n30555 = n30554 ^ n9985 ^ 1'b0 ;
  assign n30556 = n21253 ^ n7500 ^ 1'b0 ;
  assign n30557 = n30555 & ~n30556 ;
  assign n30558 = n30557 ^ n22607 ^ 1'b0 ;
  assign n30559 = n12546 & ~n18268 ;
  assign n30560 = n30559 ^ n18849 ^ n9285 ;
  assign n30561 = n3385 | n22292 ;
  assign n30562 = n23070 | n30561 ;
  assign n30563 = n3265 | n12590 ;
  assign n30564 = n12710 ^ n956 ^ 1'b0 ;
  assign n30565 = n30563 | n30564 ;
  assign n30566 = n15694 ^ x209 ^ 1'b0 ;
  assign n30567 = n3154 & ~n22669 ;
  assign n30568 = n30567 ^ n18536 ^ 1'b0 ;
  assign n30569 = n1035 | n16077 ;
  assign n30570 = n15636 ^ n1608 ^ 1'b0 ;
  assign n30571 = n21297 ^ n7907 ^ 1'b0 ;
  assign n30572 = ~n25030 & n30571 ;
  assign n30573 = n30572 ^ n4301 ^ 1'b0 ;
  assign n30574 = n30570 | n30573 ;
  assign n30575 = n16157 & n16364 ;
  assign n30576 = n3417 & n30575 ;
  assign n30577 = n30576 ^ n13036 ^ 1'b0 ;
  assign n30578 = ~n1045 & n7177 ;
  assign n30579 = ( n4449 & n10631 ) | ( n4449 & ~n30578 ) | ( n10631 & ~n30578 ) ;
  assign n30580 = n10888 ^ n2959 ^ 1'b0 ;
  assign n30581 = n4727 | n30580 ;
  assign n30582 = ~n8054 & n18171 ;
  assign n30583 = n30581 & n30582 ;
  assign n30584 = n760 & ~n3107 ;
  assign n30585 = n7683 ^ n7559 ^ 1'b0 ;
  assign n30586 = n10714 & ~n30585 ;
  assign n30587 = n30586 ^ n23069 ^ 1'b0 ;
  assign n30588 = n16213 & ~n26233 ;
  assign n30591 = n13593 ^ n2165 ^ 1'b0 ;
  assign n30592 = n6226 | n30591 ;
  assign n30589 = n15469 & n20965 ;
  assign n30590 = n30589 ^ n1328 ^ 1'b0 ;
  assign n30593 = n30592 ^ n30590 ^ n11387 ;
  assign n30594 = n19796 & n25538 ;
  assign n30595 = n20094 ^ n2420 ^ 1'b0 ;
  assign n30596 = n5120 & ~n28197 ;
  assign n30597 = n10027 & ~n10803 ;
  assign n30598 = n11345 & ~n30597 ;
  assign n30599 = n9445 & ~n30598 ;
  assign n30600 = n30599 ^ n17007 ^ 1'b0 ;
  assign n30601 = n15543 ^ x67 ^ 1'b0 ;
  assign n30602 = n2693 & ~n30601 ;
  assign n30603 = ~n11040 & n15158 ;
  assign n30604 = n30603 ^ n17825 ^ 1'b0 ;
  assign n30605 = n12934 & n28947 ;
  assign n30606 = n4159 | n5238 ;
  assign n30607 = n30606 ^ n23349 ^ 1'b0 ;
  assign n30608 = n22756 & ~n30607 ;
  assign n30609 = n22728 ^ n15171 ^ 1'b0 ;
  assign n30610 = n21099 ^ n11441 ^ 1'b0 ;
  assign n30611 = n18380 & ~n18444 ;
  assign n30612 = n20161 & ~n30611 ;
  assign n30613 = n1618 & ~n13033 ;
  assign n30614 = n2423 & n30613 ;
  assign n30615 = n11928 | n13800 ;
  assign n30616 = ~n30493 & n30615 ;
  assign n30617 = n19758 & ~n30616 ;
  assign n30618 = ~n3143 & n30617 ;
  assign n30619 = n3476 & ~n30618 ;
  assign n30620 = n30614 & n30619 ;
  assign n30621 = n27163 ^ n12380 ^ 1'b0 ;
  assign n30622 = n5392 & n8758 ;
  assign n30623 = n3740 & n30622 ;
  assign n30624 = n8329 & n27249 ;
  assign n30625 = n7015 & ~n7469 ;
  assign n30626 = n15728 & n26825 ;
  assign n30627 = n30626 ^ n7395 ^ 1'b0 ;
  assign n30628 = n2887 & n18967 ;
  assign n30629 = ~x243 & n29418 ;
  assign n30630 = n5124 & n30629 ;
  assign n30631 = n11586 & n30630 ;
  assign n30632 = ~n8112 & n14199 ;
  assign n30633 = ~n16131 & n30632 ;
  assign n30634 = n13705 & ~n20001 ;
  assign n30635 = ~n30633 & n30634 ;
  assign n30636 = ~n2664 & n30635 ;
  assign n30637 = ~n2310 & n5938 ;
  assign n30638 = ~n9309 & n30637 ;
  assign n30639 = n7442 | n18881 ;
  assign n30640 = ~n10996 & n23353 ;
  assign n30641 = n1038 & n6416 ;
  assign n30642 = n5458 & ~n21736 ;
  assign n30643 = n19935 ^ n15531 ^ 1'b0 ;
  assign n30644 = ~n16952 & n30643 ;
  assign n30645 = n30597 ^ n22616 ^ x221 ;
  assign n30646 = n5379 ^ n1621 ^ 1'b0 ;
  assign n30647 = ~n23522 & n30646 ;
  assign n30648 = ~n9786 & n16993 ;
  assign n30649 = n923 | n30648 ;
  assign n30650 = x79 & n722 ;
  assign n30651 = n4424 & ~n7036 ;
  assign n30652 = n30651 ^ n20579 ^ 1'b0 ;
  assign n30653 = n20741 ^ n9032 ^ 1'b0 ;
  assign n30654 = n24234 | n26120 ;
  assign n30655 = n30654 ^ n6278 ^ 1'b0 ;
  assign n30656 = n12707 ^ n257 ^ 1'b0 ;
  assign n30657 = n15739 & ~n30656 ;
  assign n30658 = n30657 ^ n26705 ^ 1'b0 ;
  assign n30659 = n23871 | n28387 ;
  assign n30660 = n30659 ^ n7679 ^ 1'b0 ;
  assign n30661 = n16399 ^ n8630 ^ 1'b0 ;
  assign n30662 = ~n17067 & n30661 ;
  assign n30663 = n8389 ^ n4236 ^ 1'b0 ;
  assign n30664 = ~n3673 & n17020 ;
  assign n30665 = n26692 & n30664 ;
  assign n30666 = x240 & ~n7605 ;
  assign n30667 = n30666 ^ n13559 ^ 1'b0 ;
  assign n30668 = ~n476 & n3616 ;
  assign n30669 = n30668 ^ n14068 ^ 1'b0 ;
  assign n30670 = ~n11465 & n20871 ;
  assign n30671 = n26307 ^ n13026 ^ 1'b0 ;
  assign n30672 = ~n2480 & n30671 ;
  assign n30673 = n1961 | n11651 ;
  assign n30674 = n9076 ^ x81 ^ 1'b0 ;
  assign n30675 = n30673 & n30674 ;
  assign n30676 = ~n2186 & n15033 ;
  assign n30677 = n30676 ^ n15399 ^ 1'b0 ;
  assign n30678 = ( n4325 & n14871 ) | ( n4325 & ~n28045 ) | ( n14871 & ~n28045 ) ;
  assign n30679 = n22603 & ~n30678 ;
  assign n30680 = ( ~n3325 & n7217 ) | ( ~n3325 & n9229 ) | ( n7217 & n9229 ) ;
  assign n30681 = n20011 | n22740 ;
  assign n30682 = n15312 ^ n2916 ^ 1'b0 ;
  assign n30683 = n2057 & n3040 ;
  assign n30684 = n30683 ^ n2720 ^ 1'b0 ;
  assign n30685 = ~n10147 & n30684 ;
  assign n30686 = n17393 | n30685 ;
  assign n30687 = n30682 & ~n30686 ;
  assign n30688 = n6583 & n15063 ;
  assign n30689 = n9614 & n23918 ;
  assign n30690 = n30090 ^ n12574 ^ 1'b0 ;
  assign n30691 = n5229 & n30690 ;
  assign n30692 = n20474 ^ n5703 ^ 1'b0 ;
  assign n30693 = n4536 | n17280 ;
  assign n30694 = n4333 | n30693 ;
  assign n30695 = ~n1000 & n5419 ;
  assign n30696 = n5875 | n30695 ;
  assign n30697 = n30696 ^ n28356 ^ 1'b0 ;
  assign n30698 = n2962 & n11302 ;
  assign n30699 = n13135 ^ n6220 ^ 1'b0 ;
  assign n30700 = ~n17874 & n24050 ;
  assign n30701 = n17971 ^ n13125 ^ 1'b0 ;
  assign n30702 = n15185 ^ n2470 ^ 1'b0 ;
  assign n30703 = n4267 | n13329 ;
  assign n30704 = n29383 | n30703 ;
  assign n30706 = n9565 & n13232 ;
  assign n30705 = n403 & n4549 ;
  assign n30707 = n30706 ^ n30705 ^ n13603 ;
  assign n30708 = ~n959 & n5110 ;
  assign n30709 = n30708 ^ n7123 ^ 1'b0 ;
  assign n30710 = n5312 | n26871 ;
  assign n30711 = n28698 ^ n9789 ^ 1'b0 ;
  assign n30715 = n20515 & ~n21483 ;
  assign n30716 = ~n12334 & n30715 ;
  assign n30712 = n4430 ^ n3507 ^ 1'b0 ;
  assign n30713 = n21221 | n30712 ;
  assign n30714 = n23818 & ~n30713 ;
  assign n30717 = n30716 ^ n30714 ^ 1'b0 ;
  assign n30718 = n16939 | n21864 ;
  assign n30719 = n30718 ^ n7232 ^ 1'b0 ;
  assign n30721 = n9203 & n27945 ;
  assign n30722 = ~n6106 & n30721 ;
  assign n30720 = n5610 & n23566 ;
  assign n30723 = n30722 ^ n30720 ^ 1'b0 ;
  assign n30724 = n12225 ^ n5971 ^ 1'b0 ;
  assign n30725 = n14057 & ~n30724 ;
  assign n30726 = n10160 ^ n8133 ^ 1'b0 ;
  assign n30727 = ~n4813 & n30726 ;
  assign n30728 = n30727 ^ n3964 ^ 1'b0 ;
  assign n30729 = n24150 ^ n8387 ^ 1'b0 ;
  assign n30730 = n13447 & ~n17012 ;
  assign n30731 = n30729 & n30730 ;
  assign n30732 = n13763 ^ n1459 ^ 1'b0 ;
  assign n30733 = n3090 & ~n9174 ;
  assign n30734 = ~n27240 & n30733 ;
  assign n30735 = n15081 ^ n10792 ^ 1'b0 ;
  assign n30736 = n13925 | n26148 ;
  assign n30737 = n30736 ^ n9336 ^ 1'b0 ;
  assign n30738 = n4671 & n7585 ;
  assign n30739 = n5419 & n30738 ;
  assign n30740 = n29638 ^ n9305 ^ 1'b0 ;
  assign n30741 = ~n7210 & n13770 ;
  assign n30742 = n30741 ^ n15743 ^ 1'b0 ;
  assign n30743 = ( ~n15067 & n16463 ) | ( ~n15067 & n30742 ) | ( n16463 & n30742 ) ;
  assign n30744 = ~n2257 & n2809 ;
  assign n30745 = n12862 ^ n3604 ^ 1'b0 ;
  assign n30746 = ~n3153 & n4617 ;
  assign n30747 = n1622 | n19296 ;
  assign n30748 = n2169 & ~n25538 ;
  assign n30749 = n24877 ^ n24821 ^ 1'b0 ;
  assign n30750 = n10140 & n10387 ;
  assign n30751 = n30749 & n30750 ;
  assign n30752 = n17110 ^ n4350 ^ 1'b0 ;
  assign n30753 = ~n4913 & n11242 ;
  assign n30754 = n10452 ^ x226 ^ 1'b0 ;
  assign n30755 = ~n4384 & n5025 ;
  assign n30756 = n17788 & ~n24023 ;
  assign n30757 = n30756 ^ n18496 ^ 1'b0 ;
  assign n30758 = ~n9466 & n11439 ;
  assign n30759 = n30758 ^ n6651 ^ 1'b0 ;
  assign n30760 = n17810 ^ n366 ^ x171 ;
  assign n30761 = x115 & n3530 ;
  assign n30762 = n24055 & n30761 ;
  assign n30763 = x221 & n1103 ;
  assign n30764 = n10630 & n30763 ;
  assign n30765 = n5382 & n30764 ;
  assign n30766 = n30762 | n30765 ;
  assign n30767 = n3319 | n3625 ;
  assign n30768 = n9389 & ~n30767 ;
  assign n30769 = ~n1623 & n16797 ;
  assign n30770 = n13537 & n18080 ;
  assign n30771 = n771 & n3395 ;
  assign n30773 = ~n21706 & n24408 ;
  assign n30774 = ~n1738 & n30773 ;
  assign n30772 = n8563 & ~n12573 ;
  assign n30775 = n30774 ^ n30772 ^ 1'b0 ;
  assign n30776 = n15463 ^ n1373 ^ 1'b0 ;
  assign n30777 = n729 | n30776 ;
  assign n30778 = n14065 | n30777 ;
  assign n30779 = n30778 ^ n23813 ^ 1'b0 ;
  assign n30780 = n10345 ^ n9653 ^ 1'b0 ;
  assign n30781 = ~n2872 & n30780 ;
  assign n30782 = ~n9295 & n30781 ;
  assign n30783 = ~n28378 & n28886 ;
  assign n30784 = n6781 & ~n30783 ;
  assign n30785 = n30784 ^ n23985 ^ 1'b0 ;
  assign n30787 = n14807 ^ n4111 ^ 1'b0 ;
  assign n30786 = n2977 & n10822 ;
  assign n30788 = n30787 ^ n30786 ^ n2505 ;
  assign n30789 = n1014 & n4010 ;
  assign n30790 = n1563 & n10758 ;
  assign n30791 = n30789 & n30790 ;
  assign n30792 = ~n13252 & n13445 ;
  assign n30793 = n10258 ^ n8921 ^ 1'b0 ;
  assign n30794 = n30407 & ~n30793 ;
  assign n30795 = ( n3563 & n30792 ) | ( n3563 & n30794 ) | ( n30792 & n30794 ) ;
  assign n30796 = n13217 & n14641 ;
  assign n30797 = n13555 ^ n296 ^ 1'b0 ;
  assign n30798 = n30796 | n30797 ;
  assign n30799 = n1939 ^ n1808 ^ 1'b0 ;
  assign n30800 = n30799 ^ n18679 ^ 1'b0 ;
  assign n30801 = n9786 & ~n30800 ;
  assign n30802 = n17499 ^ n3796 ^ 1'b0 ;
  assign n30803 = ~n5566 & n25921 ;
  assign n30804 = n30803 ^ n12185 ^ 1'b0 ;
  assign n30805 = n29132 | n30804 ;
  assign n30806 = n18686 & ~n28112 ;
  assign n30807 = n30806 ^ n3376 ^ 1'b0 ;
  assign n30808 = n8792 ^ n5000 ^ 1'b0 ;
  assign n30809 = n5931 & n30808 ;
  assign n30810 = ~n11611 & n18932 ;
  assign n30811 = ~n8797 & n30810 ;
  assign n30812 = n3884 | n18432 ;
  assign n30813 = ~n4169 & n24996 ;
  assign n30814 = n30813 ^ n24188 ^ n23430 ;
  assign n30815 = ~n10604 & n12552 ;
  assign n30816 = n25350 & n30815 ;
  assign n30817 = n8897 | n19494 ;
  assign n30818 = n30817 ^ n3272 ^ 1'b0 ;
  assign n30819 = n22173 & ~n30818 ;
  assign n30820 = ~n7744 & n30819 ;
  assign n30821 = n3978 & n9589 ;
  assign n30823 = ~n12785 & n14329 ;
  assign n30822 = n4899 & ~n7477 ;
  assign n30824 = n30823 ^ n30822 ^ 1'b0 ;
  assign n30825 = n964 & ~n13222 ;
  assign n30826 = n21040 ^ n16954 ^ 1'b0 ;
  assign n30827 = n30825 | n30826 ;
  assign n30828 = n1693 & n5604 ;
  assign n30829 = n21673 ^ x27 ^ 1'b0 ;
  assign n30830 = n5761 & ~n11486 ;
  assign n30831 = n14103 ^ n7701 ^ 1'b0 ;
  assign n30832 = n26368 | n30831 ;
  assign n30833 = n14175 ^ n12728 ^ n11171 ;
  assign n30834 = n538 & ~n15682 ;
  assign n30835 = ~n30833 & n30834 ;
  assign n30836 = n9745 & ~n12448 ;
  assign n30837 = n16523 & n23748 ;
  assign n30838 = ~n4400 & n30837 ;
  assign n30839 = n30838 ^ n7015 ^ 1'b0 ;
  assign n30840 = n3189 & ~n10855 ;
  assign n30841 = n27388 & n30840 ;
  assign n30842 = n2459 & ~n16612 ;
  assign n30843 = n8771 & ~n14246 ;
  assign n30844 = n30843 ^ n4658 ^ 1'b0 ;
  assign n30845 = n9266 ^ n7050 ^ 1'b0 ;
  assign n30846 = ~n5384 & n30845 ;
  assign n30847 = n710 & ~n25515 ;
  assign n30848 = n30847 ^ n30084 ^ 1'b0 ;
  assign n30849 = ( ~n9967 & n27756 ) | ( ~n9967 & n28265 ) | ( n27756 & n28265 ) ;
  assign n30850 = ~n5124 & n8287 ;
  assign n30851 = n20844 & n30850 ;
  assign n30852 = n25426 ^ n6977 ^ 1'b0 ;
  assign n30853 = ~n2716 & n8645 ;
  assign n30854 = n30853 ^ n5128 ^ 1'b0 ;
  assign n30855 = n1795 & n30854 ;
  assign n30856 = n4213 & n13235 ;
  assign n30857 = n30856 ^ n22748 ^ 1'b0 ;
  assign n30860 = n18672 | n28323 ;
  assign n30861 = n30860 ^ n3127 ^ 1'b0 ;
  assign n30858 = n1038 & n7467 ;
  assign n30859 = n13703 | n30858 ;
  assign n30862 = n30861 ^ n30859 ^ 1'b0 ;
  assign n30863 = n25493 ^ n15509 ^ 1'b0 ;
  assign n30864 = n20320 & n30863 ;
  assign n30865 = n5591 | n18928 ;
  assign n30866 = n29228 & ~n30865 ;
  assign n30867 = n18371 ^ n12860 ^ 1'b0 ;
  assign n30868 = n1431 & ~n30867 ;
  assign n30869 = n10953 & n30868 ;
  assign n30870 = n30869 ^ n978 ^ 1'b0 ;
  assign n30871 = n2523 & ~n10240 ;
  assign n30872 = ~n1801 & n30871 ;
  assign n30873 = n5396 & n10617 ;
  assign n30874 = n7900 & n12852 ;
  assign n30875 = ~n3265 & n30874 ;
  assign n30876 = n1703 | n17760 ;
  assign n30877 = x123 | n30876 ;
  assign n30878 = n3869 & n14677 ;
  assign n30879 = n30878 ^ n5778 ^ 1'b0 ;
  assign n30880 = n7193 | n30879 ;
  assign n30881 = n7618 | n13303 ;
  assign n30882 = n30881 ^ n3295 ^ 1'b0 ;
  assign n30883 = ~n9785 & n30882 ;
  assign n30884 = ~n4396 & n20941 ;
  assign n30885 = n30884 ^ n1733 ^ 1'b0 ;
  assign n30886 = n3342 & ~n18604 ;
  assign n30887 = n26312 & n30886 ;
  assign n30888 = n7173 & ~n16784 ;
  assign n30889 = n30888 ^ n4333 ^ 1'b0 ;
  assign n30890 = ~n1146 & n22014 ;
  assign n30891 = n30890 ^ n7618 ^ 1'b0 ;
  assign n30892 = n26277 ^ n1480 ^ 1'b0 ;
  assign n30893 = n12265 | n20820 ;
  assign n30894 = n24731 | n30893 ;
  assign n30895 = n3685 ^ n1264 ^ n649 ;
  assign n30896 = n30895 ^ n7993 ^ 1'b0 ;
  assign n30897 = ~n4300 & n30896 ;
  assign n30898 = n4857 & n30897 ;
  assign n30899 = n30898 ^ n1905 ^ 1'b0 ;
  assign n30900 = n24382 ^ n22787 ^ 1'b0 ;
  assign n30901 = n13833 ^ n4039 ^ 1'b0 ;
  assign n30904 = n2324 & n11815 ;
  assign n30902 = n10750 ^ n1594 ^ 1'b0 ;
  assign n30903 = ~n23677 & n30902 ;
  assign n30905 = n30904 ^ n30903 ^ 1'b0 ;
  assign n30906 = n891 & n25944 ;
  assign n30907 = n2875 & ~n8010 ;
  assign n30908 = ~n963 & n30907 ;
  assign n30910 = n4166 ^ n1787 ^ 1'b0 ;
  assign n30911 = n14998 | n30910 ;
  assign n30912 = ~n16074 & n30911 ;
  assign n30909 = n2731 | n11383 ;
  assign n30913 = n30912 ^ n30909 ^ 1'b0 ;
  assign n30914 = n5624 & ~n30913 ;
  assign n30915 = ~n1950 & n30914 ;
  assign n30916 = x163 & n11258 ;
  assign n30917 = ( x241 & n1048 ) | ( x241 & n25770 ) | ( n1048 & n25770 ) ;
  assign n30918 = n30917 ^ n10377 ^ 1'b0 ;
  assign n30919 = n7907 | n30918 ;
  assign n30920 = n30919 ^ n412 ^ 1'b0 ;
  assign n30921 = n3823 & ~n27524 ;
  assign n30922 = n6817 | n25591 ;
  assign n30923 = n15142 & ~n30922 ;
  assign n30924 = ~n4763 & n29512 ;
  assign n30925 = ~n18234 & n30924 ;
  assign n30926 = n1429 & n15141 ;
  assign n30927 = n5750 & n12733 ;
  assign n30928 = n5192 & n22246 ;
  assign n30929 = n30927 & n30928 ;
  assign n30930 = n9558 & ~n10185 ;
  assign n30931 = ~n15673 & n30930 ;
  assign n30932 = n30931 ^ n7967 ^ 1'b0 ;
  assign n30933 = n24722 ^ n15011 ^ n14891 ;
  assign n30934 = n1505 | n30933 ;
  assign n30935 = ( n1290 & ~n4223 ) | ( n1290 & n26928 ) | ( ~n4223 & n26928 ) ;
  assign n30936 = n14545 & ~n18888 ;
  assign n30937 = ~n1810 & n30936 ;
  assign n30938 = n30937 ^ n8059 ^ 1'b0 ;
  assign n30939 = ~n24010 & n30938 ;
  assign n30940 = n11501 ^ n6009 ^ 1'b0 ;
  assign n30941 = n6554 & n10089 ;
  assign n30942 = n30941 ^ n9217 ^ 1'b0 ;
  assign n30943 = n20560 ^ n807 ^ 1'b0 ;
  assign n30944 = n29544 | n30943 ;
  assign n30945 = n4205 | n4632 ;
  assign n30946 = n23125 & ~n30945 ;
  assign n30947 = n10631 & n15429 ;
  assign n30948 = ~n1537 & n30947 ;
  assign n30949 = ~n2698 & n30948 ;
  assign n30950 = n19552 ^ n9171 ^ n5125 ;
  assign n30951 = ~n2566 & n6034 ;
  assign n30952 = ~n3940 & n30951 ;
  assign n30953 = n9551 ^ n3227 ^ 1'b0 ;
  assign n30954 = n30953 ^ n15180 ^ 1'b0 ;
  assign n30955 = n16750 | n30954 ;
  assign n30956 = n30955 ^ n4179 ^ 1'b0 ;
  assign n30957 = n3281 & ~n30956 ;
  assign n30958 = n6207 & n30957 ;
  assign n30959 = n4396 | n11716 ;
  assign n30960 = n3714 & n30959 ;
  assign n30961 = n15689 ^ n12287 ^ 1'b0 ;
  assign n30962 = ~n13759 & n30961 ;
  assign n30963 = n30962 ^ n5916 ^ 1'b0 ;
  assign n30964 = n444 & n9487 ;
  assign n30965 = n7557 & n16099 ;
  assign n30966 = n12208 | n14757 ;
  assign n30967 = n30965 & n30966 ;
  assign n30968 = n13382 | n25442 ;
  assign n30969 = n23293 & ~n24426 ;
  assign n30970 = n20626 ^ n3326 ^ 1'b0 ;
  assign n30971 = n5384 | n14375 ;
  assign n30972 = n25520 | n30971 ;
  assign n30973 = n623 & n9321 ;
  assign n30974 = n30973 ^ n1007 ^ 1'b0 ;
  assign n30975 = n12961 & ~n27658 ;
  assign n30976 = n30975 ^ n7655 ^ 1'b0 ;
  assign n30977 = ~n6254 & n10900 ;
  assign n30978 = ~n3575 & n10149 ;
  assign n30979 = n30978 ^ n7406 ^ 1'b0 ;
  assign n30980 = n27563 ^ n2091 ^ 1'b0 ;
  assign n30981 = n24364 & n30980 ;
  assign n30982 = ~n5268 & n14960 ;
  assign n30983 = n21693 ^ n8712 ^ 1'b0 ;
  assign n30984 = n7666 | n30983 ;
  assign n30985 = n30982 | n30984 ;
  assign n30986 = ~n26542 & n30985 ;
  assign n30987 = n11900 ^ n5091 ^ n729 ;
  assign n30988 = n7659 & ~n10108 ;
  assign n30989 = ~n4660 & n10935 ;
  assign n30990 = n8759 & ~n29556 ;
  assign n30991 = n13945 ^ n1277 ^ 1'b0 ;
  assign n30992 = n8291 ^ n1023 ^ 1'b0 ;
  assign n30993 = n30991 & n30992 ;
  assign n30994 = n305 & ~n14436 ;
  assign n30995 = n1240 & ~n17282 ;
  assign n30996 = x201 & ~n14942 ;
  assign n30997 = n30996 ^ n3239 ^ 1'b0 ;
  assign n30998 = n9323 ^ n2212 ^ 1'b0 ;
  assign n30999 = ~n5419 & n30998 ;
  assign n31000 = ~n25934 & n30999 ;
  assign n31001 = n16426 ^ n10653 ^ 1'b0 ;
  assign n31002 = n10426 | n31001 ;
  assign n31003 = n24464 ^ n10491 ^ 1'b0 ;
  assign n31004 = n10602 & ~n10843 ;
  assign n31005 = n31004 ^ n27283 ^ 1'b0 ;
  assign n31006 = n14228 ^ n13155 ^ 1'b0 ;
  assign n31007 = n26527 & ~n27698 ;
  assign n31008 = n31007 ^ n23516 ^ 1'b0 ;
  assign n31009 = n7214 | n14757 ;
  assign n31010 = n23431 & ~n23548 ;
  assign n31011 = ~n17996 & n31010 ;
  assign n31012 = n3324 & n25256 ;
  assign n31013 = n22729 ^ n13426 ^ 1'b0 ;
  assign n31014 = ( n21864 & n29514 ) | ( n21864 & n31013 ) | ( n29514 & n31013 ) ;
  assign n31015 = ~n9194 & n25270 ;
  assign n31016 = n30947 ^ n21704 ^ 1'b0 ;
  assign n31017 = ~n669 & n31016 ;
  assign n31018 = ~n31015 & n31017 ;
  assign n31019 = n2426 | n2885 ;
  assign n31022 = ~n729 & n4289 ;
  assign n31023 = ~n2469 & n31022 ;
  assign n31020 = n6505 & n18588 ;
  assign n31021 = ~n7241 & n31020 ;
  assign n31024 = n31023 ^ n31021 ^ 1'b0 ;
  assign n31025 = n14385 ^ n3872 ^ 1'b0 ;
  assign n31026 = n3647 | n17453 ;
  assign n31027 = n31026 ^ n27704 ^ 1'b0 ;
  assign n31028 = n11893 ^ n9951 ^ 1'b0 ;
  assign n31029 = n13926 | n25540 ;
  assign n31030 = n4502 | n7261 ;
  assign n31031 = n12295 | n31030 ;
  assign n31032 = n3979 & n4376 ;
  assign n31033 = ~n15906 & n22512 ;
  assign n31034 = n26968 ^ n16954 ^ 1'b0 ;
  assign n31035 = n20177 & n31034 ;
  assign n31036 = n7333 ^ x230 ^ 1'b0 ;
  assign n31037 = n2660 & ~n20662 ;
  assign n31038 = ~n31036 & n31037 ;
  assign n31039 = n18504 | n31038 ;
  assign n31040 = ( n3833 & n13844 ) | ( n3833 & ~n17936 ) | ( n13844 & ~n17936 ) ;
  assign n31041 = n28427 & ~n31040 ;
  assign n31042 = n31041 ^ n19544 ^ 1'b0 ;
  assign n31043 = n10867 & ~n14800 ;
  assign n31044 = n17706 & n31043 ;
  assign n31045 = n988 | n17236 ;
  assign n31046 = n13264 | n31045 ;
  assign n31047 = n14848 & n28597 ;
  assign n31053 = n6220 ^ n1675 ^ 1'b0 ;
  assign n31054 = n5748 ^ n5239 ^ x223 ;
  assign n31055 = n31053 | n31054 ;
  assign n31049 = n1523 & ~n2555 ;
  assign n31050 = ~n1523 & n31049 ;
  assign n31048 = ~n4429 & n18392 ;
  assign n31051 = n31050 ^ n31048 ^ 1'b0 ;
  assign n31052 = n14377 & n31051 ;
  assign n31056 = n31055 ^ n31052 ^ 1'b0 ;
  assign n31058 = n4067 & ~n6231 ;
  assign n31059 = n21886 & n31058 ;
  assign n31057 = n648 & ~n19906 ;
  assign n31060 = n31059 ^ n31057 ^ 1'b0 ;
  assign n31061 = ~n27533 & n31060 ;
  assign n31062 = n4568 | n14965 ;
  assign n31063 = n31061 & ~n31062 ;
  assign n31064 = ~n6025 & n9381 ;
  assign n31065 = n31064 ^ n12251 ^ 1'b0 ;
  assign n31066 = n15644 | n31065 ;
  assign n31067 = n7111 | n8406 ;
  assign n31068 = n29079 ^ n16688 ^ 1'b0 ;
  assign n31069 = n1501 & n31068 ;
  assign n31070 = n24821 & n31069 ;
  assign n31071 = ~n1186 & n31070 ;
  assign n31072 = n641 | n7407 ;
  assign n31073 = n1610 & ~n1920 ;
  assign n31074 = n27106 ^ n18673 ^ 1'b0 ;
  assign n31075 = n27267 ^ n17136 ^ 1'b0 ;
  assign n31076 = n3240 & ~n31075 ;
  assign n31077 = n23189 ^ n16608 ^ n498 ;
  assign n31078 = ~n1027 & n11423 ;
  assign n31079 = ~n20714 & n31078 ;
  assign n31080 = n4295 & ~n5094 ;
  assign n31081 = n8033 | n12619 ;
  assign n31082 = n31080 & ~n31081 ;
  assign n31083 = n7469 | n11682 ;
  assign n31084 = n31083 ^ n14459 ^ 1'b0 ;
  assign n31085 = n13727 ^ n7833 ^ 1'b0 ;
  assign n31086 = n22699 & ~n31085 ;
  assign n31087 = n31086 ^ n1160 ^ 1'b0 ;
  assign n31088 = n13804 & ~n31087 ;
  assign n31089 = n4313 & ~n10551 ;
  assign n31090 = ( ~n3618 & n29606 ) | ( ~n3618 & n31089 ) | ( n29606 & n31089 ) ;
  assign n31091 = n4128 | n15677 ;
  assign n31092 = n13089 | n31091 ;
  assign n31093 = n17681 & ~n22678 ;
  assign n31094 = n31093 ^ n18945 ^ 1'b0 ;
  assign n31095 = ~n1118 & n31094 ;
  assign n31096 = ~n31092 & n31095 ;
  assign n31097 = ~n1854 & n15139 ;
  assign n31098 = n1725 & n31097 ;
  assign n31099 = x140 & ~n12585 ;
  assign n31100 = n11454 & ~n31099 ;
  assign n31101 = n19178 & ~n27049 ;
  assign n31102 = ~n3585 & n10605 ;
  assign n31103 = n6070 ^ n2753 ^ 1'b0 ;
  assign n31104 = n25618 ^ n10188 ^ n9256 ;
  assign n31105 = n13665 ^ n5167 ^ 1'b0 ;
  assign n31106 = ~n31104 & n31105 ;
  assign n31107 = n31106 ^ n17382 ^ 1'b0 ;
  assign n31108 = n13517 & ~n31107 ;
  assign n31109 = n2667 | n4360 ;
  assign n31110 = ~n3448 & n19650 ;
  assign n31111 = n7627 & n18530 ;
  assign n31112 = ~n10039 & n31111 ;
  assign n31113 = n3906 ^ n1867 ^ 1'b0 ;
  assign n31114 = n17112 ^ n790 ^ 1'b0 ;
  assign n31115 = n2283 & n9393 ;
  assign n31116 = n31115 ^ n8331 ^ 1'b0 ;
  assign n31117 = n8324 | n30290 ;
  assign n31118 = n20257 & ~n20946 ;
  assign n31119 = n31118 ^ n20749 ^ 1'b0 ;
  assign n31120 = ~n12067 & n12515 ;
  assign n31121 = n31120 ^ n20629 ^ 1'b0 ;
  assign n31122 = n12228 ^ n3331 ^ 1'b0 ;
  assign n31124 = n3593 | n22626 ;
  assign n31125 = n3656 & ~n31124 ;
  assign n31126 = n31125 ^ n756 ^ 1'b0 ;
  assign n31123 = n1693 | n15582 ;
  assign n31127 = n31126 ^ n31123 ^ 1'b0 ;
  assign n31128 = ~n6410 & n17172 ;
  assign n31129 = ~n17172 & n31128 ;
  assign n31130 = ( n3304 & n30648 ) | ( n3304 & ~n31129 ) | ( n30648 & ~n31129 ) ;
  assign n31131 = n28525 & ~n31130 ;
  assign n31132 = n18171 & ~n31131 ;
  assign n31133 = n31132 ^ n5021 ^ 1'b0 ;
  assign n31134 = ~n10797 & n11291 ;
  assign n31135 = n3082 & n31134 ;
  assign n31136 = n19350 & n31135 ;
  assign n31137 = n21307 & ~n26245 ;
  assign n31138 = n7595 ^ n6195 ^ 1'b0 ;
  assign n31139 = n30410 | n31138 ;
  assign n31140 = n1083 & n20375 ;
  assign n31141 = n31140 ^ n9089 ^ 1'b0 ;
  assign n31142 = n6966 & n16102 ;
  assign n31143 = n20587 & n31142 ;
  assign n31144 = n5290 & ~n12215 ;
  assign n31145 = n27400 | n31144 ;
  assign n31146 = n1859 ^ x120 ^ 1'b0 ;
  assign n31147 = n4203 | n31146 ;
  assign n31148 = n548 & n21307 ;
  assign n31149 = ~n9063 & n20430 ;
  assign n31150 = n31149 ^ n24635 ^ 1'b0 ;
  assign n31151 = n3426 | n24256 ;
  assign n31152 = n17467 ^ n2037 ^ 1'b0 ;
  assign n31153 = n31152 ^ n5368 ^ 1'b0 ;
  assign n31154 = n9102 & ~n10201 ;
  assign n31155 = n1365 & n31154 ;
  assign n31156 = x220 & ~n9377 ;
  assign n31157 = n31156 ^ n13515 ^ 1'b0 ;
  assign n31158 = n897 & n31157 ;
  assign n31159 = n12680 | n16218 ;
  assign n31160 = n31159 ^ n472 ^ 1'b0 ;
  assign n31161 = n17340 & n31160 ;
  assign n31162 = ~n5414 & n6389 ;
  assign n31163 = n7478 | n11110 ;
  assign n31164 = n31163 ^ n8276 ^ 1'b0 ;
  assign n31165 = n31164 ^ n20882 ^ 1'b0 ;
  assign n31166 = n14866 ^ n1208 ^ 1'b0 ;
  assign n31167 = n17806 & n31166 ;
  assign n31168 = ~n12471 & n30435 ;
  assign n31169 = n3181 ^ n1511 ^ 1'b0 ;
  assign n31170 = n2693 & ~n31169 ;
  assign n31171 = n18313 & n31170 ;
  assign n31172 = n7633 ^ n796 ^ 1'b0 ;
  assign n31173 = n31171 & n31172 ;
  assign n31174 = n320 & n10645 ;
  assign n31175 = n19220 | n31174 ;
  assign n31176 = ~n4347 & n8512 ;
  assign n31177 = n25512 & n31176 ;
  assign n31178 = ~n23499 & n31177 ;
  assign n31179 = n23802 ^ n17866 ^ 1'b0 ;
  assign n31180 = n6049 & n31179 ;
  assign n31181 = n31180 ^ n1402 ^ 1'b0 ;
  assign n31182 = ( ~n5286 & n14076 ) | ( ~n5286 & n19756 ) | ( n14076 & n19756 ) ;
  assign n31183 = n19444 ^ n9399 ^ 1'b0 ;
  assign n31184 = n3645 | n26282 ;
  assign n31185 = n14412 ^ n1477 ^ 1'b0 ;
  assign n31186 = ~n31184 & n31185 ;
  assign n31187 = n22889 | n26790 ;
  assign n31189 = n3604 & n8692 ;
  assign n31188 = n13764 | n13987 ;
  assign n31190 = n31189 ^ n31188 ^ 1'b0 ;
  assign n31191 = n1707 & n9277 ;
  assign n31192 = ~x145 & n31191 ;
  assign n31193 = n10818 | n28654 ;
  assign n31194 = n31193 ^ n6480 ^ 1'b0 ;
  assign n31195 = n6152 & n13585 ;
  assign n31196 = n31195 ^ n7011 ^ 1'b0 ;
  assign n31197 = n10044 ^ n1909 ^ 1'b0 ;
  assign n31198 = n7644 | n31197 ;
  assign n31199 = n8990 ^ n8532 ^ 1'b0 ;
  assign n31200 = ~n22556 & n24516 ;
  assign n31201 = n869 | n22180 ;
  assign n31202 = ( n10689 & n12448 ) | ( n10689 & n12737 ) | ( n12448 & n12737 ) ;
  assign n31203 = n9433 & n25928 ;
  assign n31204 = n21427 ^ n3076 ^ 1'b0 ;
  assign n31205 = n3088 & ~n9267 ;
  assign n31206 = ~n10046 & n31205 ;
  assign n31207 = n31204 & n31206 ;
  assign n31208 = n11417 ^ n8128 ^ 1'b0 ;
  assign n31209 = n13934 & ~n17106 ;
  assign n31210 = n31209 ^ n18216 ^ 1'b0 ;
  assign n31211 = n8378 ^ n7010 ^ 1'b0 ;
  assign n31212 = n18275 & n22986 ;
  assign n31213 = n6811 | n31212 ;
  assign n31214 = n1906 ^ n808 ^ 1'b0 ;
  assign n31217 = ~n2306 & n21767 ;
  assign n31215 = n5346 ^ n405 ^ 1'b0 ;
  assign n31216 = n23740 & n31215 ;
  assign n31218 = n31217 ^ n31216 ^ 1'b0 ;
  assign n31219 = ~n7960 & n31218 ;
  assign n31220 = n8654 ^ n8083 ^ 1'b0 ;
  assign n31221 = n2561 & ~n31220 ;
  assign n31222 = ~n2644 & n31221 ;
  assign n31223 = ~n31221 & n31222 ;
  assign n31224 = n29698 ^ n10498 ^ 1'b0 ;
  assign n31225 = n29550 | n31224 ;
  assign n31226 = n5974 ^ n4991 ^ n784 ;
  assign n31227 = n12190 ^ n7986 ^ 1'b0 ;
  assign n31228 = n1025 & n4959 ;
  assign n31229 = n31228 ^ n11519 ^ 1'b0 ;
  assign n31230 = n2307 & n3533 ;
  assign n31231 = ~n11680 & n31230 ;
  assign n31232 = n1025 & ~n31231 ;
  assign n31233 = ~x123 & n11197 ;
  assign n31234 = n25721 ^ n18849 ^ 1'b0 ;
  assign n31240 = ~n11354 & n17092 ;
  assign n31241 = n31240 ^ n20480 ^ 1'b0 ;
  assign n31242 = n14240 & ~n31241 ;
  assign n31243 = n10652 ^ n8010 ^ 1'b0 ;
  assign n31244 = n31243 ^ n5021 ^ 1'b0 ;
  assign n31245 = n31242 & n31244 ;
  assign n31246 = n17573 & ~n31245 ;
  assign n31237 = n9799 ^ x152 ^ 1'b0 ;
  assign n31235 = n19629 ^ n2320 ^ 1'b0 ;
  assign n31236 = ~n26703 & n31235 ;
  assign n31238 = n31237 ^ n31236 ^ n28994 ;
  assign n31239 = ~n21685 & n31238 ;
  assign n31247 = n31246 ^ n31239 ^ 1'b0 ;
  assign n31248 = n25570 ^ n7810 ^ 1'b0 ;
  assign n31249 = ~n10967 & n31248 ;
  assign n31250 = n1446 & n20031 ;
  assign n31251 = n31250 ^ n9959 ^ 1'b0 ;
  assign n31252 = n2185 | n14508 ;
  assign n31253 = n9916 & ~n31252 ;
  assign n31254 = n19984 | n31253 ;
  assign n31255 = n1608 & ~n31254 ;
  assign n31256 = n13578 & ~n31255 ;
  assign n31257 = n31256 ^ n621 ^ 1'b0 ;
  assign n31258 = n4336 ^ x84 ^ 1'b0 ;
  assign n31259 = ~n24884 & n31258 ;
  assign n31260 = n6558 & n31259 ;
  assign n31261 = ~n4351 & n21979 ;
  assign n31262 = n31261 ^ n29084 ^ 1'b0 ;
  assign n31263 = n9104 & ~n15711 ;
  assign n31264 = n22509 & n31263 ;
  assign n31265 = n12154 ^ n10854 ^ 1'b0 ;
  assign n31266 = n16898 & n31265 ;
  assign n31267 = ~n14980 & n31266 ;
  assign n31268 = n31264 & n31267 ;
  assign n31269 = n11219 & n15245 ;
  assign n31270 = n5591 | n31269 ;
  assign n31271 = n15783 & n31270 ;
  assign n31272 = n3409 & n31271 ;
  assign n31273 = n11302 ^ n7726 ^ 1'b0 ;
  assign n31274 = ~n19945 & n31273 ;
  assign n31275 = n31272 & n31274 ;
  assign n31276 = n6507 ^ n5162 ^ 1'b0 ;
  assign n31277 = n5296 & n31276 ;
  assign n31278 = n6676 & n9217 ;
  assign n31279 = n31278 ^ n1814 ^ 1'b0 ;
  assign n31280 = n9681 | n31279 ;
  assign n31281 = n18885 ^ n6355 ^ 1'b0 ;
  assign n31287 = n11176 ^ n1663 ^ 1'b0 ;
  assign n31288 = ~n8935 & n31287 ;
  assign n31282 = x208 & n1217 ;
  assign n31283 = ~x208 & n31282 ;
  assign n31284 = n31283 ^ n18022 ^ 1'b0 ;
  assign n31285 = n25209 | n31284 ;
  assign n31286 = n29498 | n31285 ;
  assign n31289 = n31288 ^ n31286 ^ 1'b0 ;
  assign n31290 = ~n1046 & n31289 ;
  assign n31291 = n18241 ^ n15425 ^ 1'b0 ;
  assign n31292 = n17895 & ~n31291 ;
  assign n31293 = n4412 & n31292 ;
  assign n31294 = ~n9087 & n31293 ;
  assign n31295 = ~n4089 & n15537 ;
  assign n31296 = n24626 ^ n7729 ^ n4502 ;
  assign n31297 = n4260 & n11274 ;
  assign n31298 = n1016 & ~n18393 ;
  assign n31299 = n31298 ^ n7912 ^ 1'b0 ;
  assign n31300 = x76 | n31299 ;
  assign n31301 = n3529 & ~n31300 ;
  assign n31302 = n18136 ^ n5244 ^ 1'b0 ;
  assign n31303 = n13564 | n31302 ;
  assign n31304 = n17489 ^ n8437 ^ 1'b0 ;
  assign n31305 = n31304 ^ n16908 ^ n15737 ;
  assign n31306 = n6431 & n7890 ;
  assign n31307 = n2362 & n31306 ;
  assign n31308 = n3484 & n13763 ;
  assign n31309 = n27238 ^ n10039 ^ 1'b0 ;
  assign n31310 = n16688 & n31309 ;
  assign n31311 = n31310 ^ n13256 ^ 1'b0 ;
  assign n31314 = ~n1348 & n5369 ;
  assign n31312 = n5700 & n6876 ;
  assign n31313 = n27702 | n31312 ;
  assign n31315 = n31314 ^ n31313 ^ 1'b0 ;
  assign n31316 = ~n7411 & n12592 ;
  assign n31317 = n4560 & n18226 ;
  assign n31318 = n31317 ^ n28287 ^ 1'b0 ;
  assign n31319 = n12245 ^ n10413 ^ 1'b0 ;
  assign n31320 = n21964 & ~n31319 ;
  assign n31321 = n10780 ^ n1628 ^ 1'b0 ;
  assign n31322 = n3055 & ~n31321 ;
  assign n31323 = n31322 ^ n3143 ^ 1'b0 ;
  assign n31324 = n8892 & ~n31323 ;
  assign n31325 = n4951 & ~n8495 ;
  assign n31326 = n15021 & ~n31325 ;
  assign n31327 = n20243 ^ n17466 ^ 1'b0 ;
  assign n31328 = ~n16981 & n31327 ;
  assign n31329 = n8268 | n13306 ;
  assign n31330 = n15494 & ~n31329 ;
  assign n31331 = ( n4092 & n10363 ) | ( n4092 & n11233 ) | ( n10363 & n11233 ) ;
  assign n31332 = n14969 ^ n9402 ^ 1'b0 ;
  assign n31333 = n29658 | n31332 ;
  assign n31334 = n2373 & n11059 ;
  assign n31335 = ~n1111 & n18030 ;
  assign n31336 = n31335 ^ n23803 ^ 1'b0 ;
  assign n31337 = ( ~n7888 & n15456 ) | ( ~n7888 & n30084 ) | ( n15456 & n30084 ) ;
  assign n31338 = n7241 & ~n8846 ;
  assign n31339 = n1376 & ~n1661 ;
  assign n31340 = ~n9149 & n31339 ;
  assign n31341 = ( n13590 & ~n26693 ) | ( n13590 & n31340 ) | ( ~n26693 & n31340 ) ;
  assign n31342 = n1307 & ~n8059 ;
  assign n31343 = n18046 & n31342 ;
  assign n31344 = n2136 & ~n30395 ;
  assign n31345 = n31343 & n31344 ;
  assign n31346 = n31345 ^ n1267 ^ 1'b0 ;
  assign n31347 = n31341 | n31346 ;
  assign n31348 = n7151 ^ n1959 ^ n553 ;
  assign n31349 = n24151 ^ n12004 ^ 1'b0 ;
  assign n31350 = ~n2731 & n31349 ;
  assign n31351 = n20820 ^ n19088 ^ 1'b0 ;
  assign n31352 = ~n1732 & n3152 ;
  assign n31354 = ~n590 & n782 ;
  assign n31353 = n5808 & n6097 ;
  assign n31355 = n31354 ^ n31353 ^ 1'b0 ;
  assign n31356 = n20687 ^ n11205 ^ 1'b0 ;
  assign n31357 = n23856 ^ n1511 ^ 1'b0 ;
  assign n31358 = n25579 & n31357 ;
  assign n31359 = n14807 | n28925 ;
  assign n31360 = n20374 ^ n19992 ^ 1'b0 ;
  assign n31361 = ~x25 & n31360 ;
  assign n31362 = ~n24150 & n31361 ;
  assign n31363 = n9254 & ~n29311 ;
  assign n31364 = n31363 ^ n19019 ^ 1'b0 ;
  assign n31365 = n31364 ^ n17907 ^ n9606 ;
  assign n31366 = ~n4323 & n15391 ;
  assign n31367 = x180 & ~n25460 ;
  assign n31368 = n6881 & n19332 ;
  assign n31369 = n12400 ^ n2668 ^ 1'b0 ;
  assign n31370 = ~n31368 & n31369 ;
  assign n31371 = ~n21671 & n31370 ;
  assign n31372 = n31367 & n31371 ;
  assign n31373 = ~n22424 & n23910 ;
  assign n31374 = n28282 ^ n13567 ^ 1'b0 ;
  assign n31375 = n31374 ^ n17095 ^ 1'b0 ;
  assign n31376 = n1896 & n2507 ;
  assign n31377 = ~n5354 & n31376 ;
  assign n31378 = n11524 | n31377 ;
  assign n31379 = n31375 | n31378 ;
  assign n31380 = n21342 ^ n2230 ^ 1'b0 ;
  assign n31381 = n31379 & n31380 ;
  assign n31382 = n24373 & ~n24663 ;
  assign n31383 = n22057 ^ n12379 ^ 1'b0 ;
  assign n31384 = ~n4655 & n7454 ;
  assign n31385 = ~n3566 & n5064 ;
  assign n31386 = ~n10391 & n31385 ;
  assign n31387 = n31386 ^ n17958 ^ 1'b0 ;
  assign n31388 = n31384 & n31387 ;
  assign n31389 = n16130 ^ n10516 ^ 1'b0 ;
  assign n31390 = n20968 ^ n7081 ^ 1'b0 ;
  assign n31391 = n11128 ^ n3316 ^ n2017 ;
  assign n31392 = n17817 | n31391 ;
  assign n31393 = n14299 & n31392 ;
  assign n31394 = n30823 ^ n3458 ^ 1'b0 ;
  assign n31395 = ~n7749 & n18432 ;
  assign n31396 = n30420 ^ n15854 ^ 1'b0 ;
  assign n31397 = n21246 & n26277 ;
  assign n31398 = n3097 & n31397 ;
  assign n31399 = n9542 & n19942 ;
  assign n31400 = n31399 ^ n7337 ^ n5160 ;
  assign n31401 = x208 & n31400 ;
  assign n31402 = n31401 ^ n7878 ^ 1'b0 ;
  assign n31403 = n3487 & n22071 ;
  assign n31404 = n29685 & n31403 ;
  assign n31405 = n12380 & ~n18355 ;
  assign n31406 = n31405 ^ n13261 ^ 1'b0 ;
  assign n31407 = n11196 & n31406 ;
  assign n31408 = n13213 & n31407 ;
  assign n31409 = n6972 ^ n3597 ^ 1'b0 ;
  assign n31410 = n30047 & n31409 ;
  assign n31411 = n29099 ^ n26129 ^ 1'b0 ;
  assign n31412 = ~n4647 & n13398 ;
  assign n31413 = n31412 ^ n22012 ^ 1'b0 ;
  assign n31414 = n31411 & ~n31413 ;
  assign n31415 = n19257 ^ n1900 ^ 1'b0 ;
  assign n31416 = n13053 & ~n27199 ;
  assign n31417 = ~n31292 & n31416 ;
  assign n31418 = n19297 ^ n6868 ^ 1'b0 ;
  assign n31419 = ~n8617 & n30134 ;
  assign n31420 = n6899 | n18097 ;
  assign n31421 = n31420 ^ x98 ^ 1'b0 ;
  assign n31423 = n1345 & n19635 ;
  assign n31422 = n1580 | n15930 ;
  assign n31424 = n31423 ^ n31422 ^ 1'b0 ;
  assign n31425 = n5458 & n9597 ;
  assign n31426 = n4694 & n31425 ;
  assign n31427 = n5122 ^ n1183 ^ 1'b0 ;
  assign n31428 = n14848 & ~n31427 ;
  assign n31429 = n1436 & ~n20556 ;
  assign n31430 = n20996 & n31429 ;
  assign n31431 = n30485 ^ n19682 ^ 1'b0 ;
  assign n31432 = ( n1104 & n10213 ) | ( n1104 & n31431 ) | ( n10213 & n31431 ) ;
  assign n31433 = ~n7228 & n18174 ;
  assign n31434 = n3387 | n24980 ;
  assign n31435 = n30651 ^ n2261 ^ 1'b0 ;
  assign n31436 = n14639 ^ n7077 ^ n4613 ;
  assign n31437 = n1038 & ~n6679 ;
  assign n31438 = n31437 ^ n21395 ^ 1'b0 ;
  assign n31439 = n15393 & n31438 ;
  assign n31440 = n14837 ^ n12184 ^ n10400 ;
  assign n31441 = n24545 & n31440 ;
  assign n31442 = ~n12163 & n21036 ;
  assign n31443 = n13543 ^ n4289 ^ 1'b0 ;
  assign n31444 = n8295 & ~n31443 ;
  assign n31445 = ~n5751 & n31444 ;
  assign n31446 = ~n8236 & n19059 ;
  assign n31447 = ~n18059 & n31446 ;
  assign n31448 = n29383 ^ n13099 ^ 1'b0 ;
  assign n31449 = x24 & n7049 ;
  assign n31450 = n18867 ^ n1133 ^ 1'b0 ;
  assign n31451 = n31450 ^ n9095 ^ 1'b0 ;
  assign n31452 = ~n26294 & n31451 ;
  assign n31453 = ~n13127 & n16135 ;
  assign n31454 = n6171 | n11083 ;
  assign n31455 = n18895 ^ n3524 ^ 1'b0 ;
  assign n31456 = n1992 & n31455 ;
  assign n31457 = n31456 ^ n27542 ^ n27341 ;
  assign n31458 = n18145 | n28123 ;
  assign n31459 = n18192 ^ n6382 ^ 1'b0 ;
  assign n31460 = n6250 ^ n4540 ^ 1'b0 ;
  assign n31461 = n22318 ^ n13001 ^ n9446 ;
  assign n31462 = ~n17124 & n18657 ;
  assign n31463 = ~n24881 & n31462 ;
  assign n31464 = n30463 | n31463 ;
  assign n31466 = n1195 & n23279 ;
  assign n31467 = ~n7515 & n31466 ;
  assign n31465 = ~n6989 & n13057 ;
  assign n31468 = n31467 ^ n31465 ^ 1'b0 ;
  assign n31469 = n27505 ^ n10175 ^ 1'b0 ;
  assign n31470 = ~n8742 & n29229 ;
  assign n31471 = n31470 ^ n7020 ^ 1'b0 ;
  assign n31472 = n9125 | n31471 ;
  assign n31473 = n1334 & ~n21865 ;
  assign n31474 = n12738 ^ n5125 ^ n1453 ;
  assign n31475 = n14360 | n31474 ;
  assign n31476 = n31475 ^ n9518 ^ n1814 ;
  assign n31478 = n11944 ^ n10098 ^ 1'b0 ;
  assign n31479 = n1029 & n31478 ;
  assign n31477 = ~n2286 & n9254 ;
  assign n31480 = n31479 ^ n31477 ^ 1'b0 ;
  assign n31481 = n2063 & n28415 ;
  assign n31482 = n31481 ^ n6104 ^ 1'b0 ;
  assign n31483 = n1234 | n31482 ;
  assign n31484 = n17247 ^ n1308 ^ 1'b0 ;
  assign n31485 = ~n919 & n15851 ;
  assign n31486 = n31485 ^ n17497 ^ 1'b0 ;
  assign n31487 = n11240 & n27242 ;
  assign n31488 = n5018 ^ x2 ^ 1'b0 ;
  assign n31489 = n15650 ^ n13745 ^ n3249 ;
  assign n31490 = n6271 & n7613 ;
  assign n31491 = ~n6715 & n16752 ;
  assign n31492 = n16512 & n19985 ;
  assign n31493 = ~n2730 & n31492 ;
  assign n31494 = n3687 & n4233 ;
  assign n31495 = n31494 ^ n9427 ^ 1'b0 ;
  assign n31496 = ~n23457 & n31495 ;
  assign n31497 = n3343 & n12494 ;
  assign n31498 = n1457 & n31497 ;
  assign n31499 = ~n7457 & n31498 ;
  assign n31500 = n7277 & n28646 ;
  assign n31501 = n31500 ^ n14288 ^ 1'b0 ;
  assign n31502 = n31501 ^ n9326 ^ 1'b0 ;
  assign n31503 = n8102 & ~n31502 ;
  assign n31504 = x92 & ~n20397 ;
  assign n31505 = n5021 ^ n1376 ^ 1'b0 ;
  assign n31506 = n18829 ^ n14045 ^ 1'b0 ;
  assign n31507 = n6498 ^ n1363 ^ 1'b0 ;
  assign n31508 = ~n21450 & n31507 ;
  assign n31509 = n9966 ^ n3039 ^ 1'b0 ;
  assign n31510 = n3852 & n31509 ;
  assign n31511 = n31508 & ~n31510 ;
  assign n31512 = ~n2303 & n15341 ;
  assign n31513 = ~n8659 & n31512 ;
  assign n31514 = n8851 ^ n4345 ^ 1'b0 ;
  assign n31515 = n31514 ^ n7047 ^ 1'b0 ;
  assign n31516 = n27208 & n31515 ;
  assign n31517 = n18951 ^ n12601 ^ 1'b0 ;
  assign n31518 = ~n28419 & n31517 ;
  assign n31519 = n26682 ^ n17591 ^ 1'b0 ;
  assign n31520 = n8118 & ~n9025 ;
  assign n31521 = n6809 ^ n2615 ^ 1'b0 ;
  assign n31522 = n31521 ^ n2826 ^ 1'b0 ;
  assign n31523 = n31522 ^ n14767 ^ 1'b0 ;
  assign n31524 = n4214 & n31523 ;
  assign n31525 = n6112 | n10684 ;
  assign n31526 = n31524 | n31525 ;
  assign n31527 = n5943 ^ n1727 ^ 1'b0 ;
  assign n31528 = n5862 & n18134 ;
  assign n31529 = ~n31527 & n31528 ;
  assign n31530 = n7652 | n15814 ;
  assign n31531 = n31530 ^ n16206 ^ 1'b0 ;
  assign n31532 = n21805 & ~n31531 ;
  assign n31533 = ~n5217 & n9741 ;
  assign n31534 = n31533 ^ n26552 ^ 1'b0 ;
  assign n31535 = n30304 ^ n1825 ^ 1'b0 ;
  assign n31536 = n23353 | n31535 ;
  assign n31537 = n29418 ^ n12443 ^ n4048 ;
  assign n31538 = n24941 ^ n5112 ^ 1'b0 ;
  assign n31539 = n1474 & n31538 ;
  assign n31540 = n6402 & ~n10186 ;
  assign n31541 = ~n6402 & n31540 ;
  assign n31543 = ~x193 & n7583 ;
  assign n31544 = x193 & n31543 ;
  assign n31542 = n15189 ^ n13661 ^ 1'b0 ;
  assign n31545 = n31544 ^ n31542 ^ 1'b0 ;
  assign n31546 = n31541 | n31545 ;
  assign n31547 = n21058 & n28463 ;
  assign n31548 = n5139 & n31547 ;
  assign n31549 = n368 | n17307 ;
  assign n31550 = x160 & ~n20553 ;
  assign n31551 = ~n14652 & n31550 ;
  assign n31552 = n2613 | n22266 ;
  assign n31553 = n31552 ^ n25853 ^ 1'b0 ;
  assign n31554 = ~n4699 & n7856 ;
  assign n31555 = n15918 ^ n7701 ^ 1'b0 ;
  assign n31556 = n31554 & ~n31555 ;
  assign n31557 = n27175 ^ n6532 ^ 1'b0 ;
  assign n31558 = n568 & n2257 ;
  assign n31559 = n31069 ^ n18370 ^ 1'b0 ;
  assign n31560 = n3468 & n4300 ;
  assign n31561 = ~n3468 & n31560 ;
  assign n31562 = n19924 | n31561 ;
  assign n31563 = n18466 ^ n17886 ^ 1'b0 ;
  assign n31564 = n31562 & n31563 ;
  assign n31565 = n31564 ^ n10603 ^ 1'b0 ;
  assign n31566 = n2371 | n16314 ;
  assign n31567 = n21261 ^ n4094 ^ 1'b0 ;
  assign n31568 = n18196 & ~n22338 ;
  assign n31569 = n4404 ^ n2263 ^ 1'b0 ;
  assign n31570 = n1111 & n31569 ;
  assign n31571 = ~n16855 & n31570 ;
  assign n31572 = n2018 & n31571 ;
  assign n31573 = n17465 | n31572 ;
  assign n31574 = n31573 ^ n1996 ^ 1'b0 ;
  assign n31575 = n4896 | n5704 ;
  assign n31576 = n13034 & ~n31575 ;
  assign n31577 = n12514 ^ n3695 ^ 1'b0 ;
  assign n31578 = n15509 | n31577 ;
  assign n31579 = ~n10674 & n25015 ;
  assign n31580 = n15046 ^ n2739 ^ 1'b0 ;
  assign n31581 = ~n13890 & n31580 ;
  assign n31582 = n6104 ^ n1926 ^ 1'b0 ;
  assign n31583 = ~n19254 & n25640 ;
  assign n31584 = n15548 & n17341 ;
  assign n31585 = n8065 | n31584 ;
  assign n31586 = n31585 ^ n15352 ^ 1'b0 ;
  assign n31589 = ~n436 & n540 ;
  assign n31590 = n436 & n31589 ;
  assign n31591 = n1177 & ~n31590 ;
  assign n31592 = ~n1177 & n31591 ;
  assign n31593 = ~n2550 & n31592 ;
  assign n31587 = ~n6617 & n8728 ;
  assign n31588 = ~n8728 & n31587 ;
  assign n31594 = n31593 ^ n31588 ^ 1'b0 ;
  assign n31595 = x34 & x219 ;
  assign n31596 = ~x219 & n31595 ;
  assign n31597 = n994 & ~n31596 ;
  assign n31598 = x105 & x199 ;
  assign n31599 = ~x105 & n31598 ;
  assign n31600 = n454 & ~n31599 ;
  assign n31601 = n31599 & n31600 ;
  assign n31602 = n1271 | n31601 ;
  assign n31603 = n31601 & ~n31602 ;
  assign n31604 = n31597 & n31603 ;
  assign n31605 = n2892 | n31604 ;
  assign n31606 = n31604 & ~n31605 ;
  assign n31607 = n26999 & ~n31606 ;
  assign n31608 = ~n26999 & n31607 ;
  assign n31609 = n3337 | n31608 ;
  assign n31610 = n31594 & ~n31609 ;
  assign n31611 = n3378 & n12966 ;
  assign n31612 = n31611 ^ n22544 ^ 1'b0 ;
  assign n31614 = n6162 | n19254 ;
  assign n31613 = n6091 & n10709 ;
  assign n31615 = n31614 ^ n31613 ^ 1'b0 ;
  assign n31616 = n21307 & ~n21714 ;
  assign n31617 = n31616 ^ n15337 ^ 1'b0 ;
  assign n31618 = ( n6655 & n10714 ) | ( n6655 & ~n10827 ) | ( n10714 & ~n10827 ) ;
  assign n31619 = n14133 ^ n1353 ^ 1'b0 ;
  assign n31620 = ~n944 & n21447 ;
  assign n31621 = n8764 | n21242 ;
  assign n31622 = n31621 ^ n8663 ^ 1'b0 ;
  assign n31623 = n3399 & ~n8651 ;
  assign n31624 = n22557 & n31623 ;
  assign n31625 = n17579 & ~n31624 ;
  assign n31626 = n24033 & n31625 ;
  assign n31627 = n20568 & ~n31174 ;
  assign n31628 = n31627 ^ n2127 ^ 1'b0 ;
  assign n31629 = x175 | n14428 ;
  assign n31630 = n31629 ^ n18349 ^ 1'b0 ;
  assign n31631 = n1566 & n27198 ;
  assign n31632 = ~n11001 & n11963 ;
  assign n31633 = n5759 | n31632 ;
  assign n31634 = n31633 ^ n23764 ^ 1'b0 ;
  assign n31635 = n13285 ^ n5848 ^ 1'b0 ;
  assign n31637 = n4186 & ~n9889 ;
  assign n31638 = n2939 & n31637 ;
  assign n31639 = n31638 ^ n15519 ^ 1'b0 ;
  assign n31636 = ~n1146 & n27120 ;
  assign n31640 = n31639 ^ n31636 ^ 1'b0 ;
  assign n31641 = n9438 ^ n1243 ^ 1'b0 ;
  assign n31642 = n1762 & n31641 ;
  assign n31643 = ~n4059 & n27443 ;
  assign n31645 = x165 & ~n1788 ;
  assign n31646 = n2887 | n20555 ;
  assign n31647 = n31646 ^ n3561 ^ 1'b0 ;
  assign n31648 = ~n31645 & n31647 ;
  assign n31644 = n29096 & n31586 ;
  assign n31649 = n31648 ^ n31644 ^ 1'b0 ;
  assign n31651 = ~n20928 & n24709 ;
  assign n31652 = n31651 ^ n11963 ^ 1'b0 ;
  assign n31650 = n10747 | n13222 ;
  assign n31653 = n31652 ^ n31650 ^ 1'b0 ;
  assign n31654 = n18344 ^ n7508 ^ 1'b0 ;
  assign n31655 = n9376 & ~n31654 ;
  assign n31656 = n1291 | n20447 ;
  assign n31657 = n967 | n31656 ;
  assign n31658 = n13021 ^ n562 ^ 1'b0 ;
  assign n31659 = n2368 & n20457 ;
  assign n31660 = n13115 & ~n18412 ;
  assign n31661 = n31660 ^ n13778 ^ 1'b0 ;
  assign n31662 = n1302 & n31661 ;
  assign n31663 = n7459 ^ n3071 ^ 1'b0 ;
  assign n31664 = n6928 | n9069 ;
  assign n31665 = n17256 ^ n17182 ^ 1'b0 ;
  assign n31666 = n5686 & n31665 ;
  assign n31667 = n31666 ^ n6127 ^ 1'b0 ;
  assign n31668 = n31664 & ~n31667 ;
  assign n31669 = n2315 | n11742 ;
  assign n31670 = n7135 & n14324 ;
  assign n31671 = n18304 ^ n11449 ^ 1'b0 ;
  assign n31672 = n6979 & ~n31671 ;
  assign n31673 = n11201 | n22288 ;
  assign n31674 = n7126 & ~n23273 ;
  assign n31675 = n10608 ^ n505 ^ 1'b0 ;
  assign n31676 = n31674 | n31675 ;
  assign n31677 = n11775 | n19568 ;
  assign n31678 = n3905 & ~n5384 ;
  assign n31679 = n31678 ^ n8281 ^ 1'b0 ;
  assign n31680 = n1507 | n31679 ;
  assign n31681 = n17471 | n20480 ;
  assign n31682 = n4881 & n27890 ;
  assign n31683 = n31682 ^ n29357 ^ 1'b0 ;
  assign n31684 = n590 & n1070 ;
  assign n31685 = n2561 & n6288 ;
  assign n31686 = x179 & n31685 ;
  assign n31687 = ~n19366 & n31686 ;
  assign n31688 = n17188 ^ n8240 ^ 1'b0 ;
  assign n31689 = ( n16610 & n20345 ) | ( n16610 & ~n31688 ) | ( n20345 & ~n31688 ) ;
  assign n31690 = n22164 ^ n10623 ^ 1'b0 ;
  assign n31691 = ~n13040 & n31690 ;
  assign n31692 = n23497 ^ n9517 ^ 1'b0 ;
  assign n31693 = n10829 & n31692 ;
  assign n31694 = ~n16418 & n31693 ;
  assign n31695 = ~n18749 & n20685 ;
  assign n31696 = n11933 & n31695 ;
  assign n31697 = n15248 & ~n28812 ;
  assign n31698 = ~n15434 & n31697 ;
  assign n31699 = n26218 & ~n31698 ;
  assign n31700 = ~n14805 & n31699 ;
  assign n31701 = n7338 & ~n8378 ;
  assign n31702 = ~x130 & n31701 ;
  assign n31703 = n11914 ^ n5186 ^ 1'b0 ;
  assign n31704 = x73 & ~n2470 ;
  assign n31705 = n2470 & n31704 ;
  assign n31706 = n31705 ^ n415 ^ 1'b0 ;
  assign n31707 = ~n16054 & n31706 ;
  assign n31708 = n12952 | n31707 ;
  assign n31709 = n23712 ^ n4785 ^ 1'b0 ;
  assign n31710 = n16678 & n18508 ;
  assign n31711 = n936 & n6325 ;
  assign n31712 = ~n6325 & n31711 ;
  assign n31713 = n2615 | n31712 ;
  assign n31714 = n8613 ^ n8242 ^ 1'b0 ;
  assign n31715 = n3386 ^ n1792 ^ 1'b0 ;
  assign n31716 = ~n26516 & n31715 ;
  assign n31717 = n31716 ^ n651 ^ 1'b0 ;
  assign n31718 = ~n1411 & n26376 ;
  assign n31719 = n19478 ^ n7102 ^ n3187 ;
  assign n31720 = ~n3331 & n27370 ;
  assign n31721 = ~n2895 & n23524 ;
  assign n31722 = ~n452 & n29045 ;
  assign n31723 = n3376 | n8056 ;
  assign n31724 = n30824 ^ n13388 ^ 1'b0 ;
  assign n31725 = n22576 & n31724 ;
  assign n31726 = n31725 ^ n9617 ^ 1'b0 ;
  assign n31727 = n313 & n30167 ;
  assign n31728 = ~n3255 & n4867 ;
  assign n31729 = ~n2292 & n31728 ;
  assign n31730 = n1681 | n3468 ;
  assign n31731 = n27286 ^ n859 ^ 1'b0 ;
  assign n31732 = ( n6483 & n12858 ) | ( n6483 & n30238 ) | ( n12858 & n30238 ) ;
  assign n31733 = ~n1879 & n6956 ;
  assign n31734 = ~n20941 & n31733 ;
  assign n31735 = n14335 ^ n1644 ^ 1'b0 ;
  assign n31736 = ~n10100 & n18270 ;
  assign n31737 = n6900 ^ n6001 ^ 1'b0 ;
  assign n31738 = ~n23740 & n31737 ;
  assign n31739 = ~n11694 & n16986 ;
  assign n31740 = n31739 ^ n573 ^ 1'b0 ;
  assign n31743 = ~n6205 & n12233 ;
  assign n31741 = n4321 & ~n13992 ;
  assign n31742 = n20773 & n31741 ;
  assign n31744 = n31743 ^ n31742 ^ 1'b0 ;
  assign n31745 = n31740 & ~n31744 ;
  assign n31746 = ~n7944 & n14717 ;
  assign n31748 = ( ~n1806 & n3920 ) | ( ~n1806 & n24222 ) | ( n3920 & n24222 ) ;
  assign n31747 = n1952 | n3263 ;
  assign n31749 = n31748 ^ n31747 ^ 1'b0 ;
  assign n31750 = n10237 & ~n31749 ;
  assign n31751 = n20621 ^ n2951 ^ 1'b0 ;
  assign n31752 = ~n2814 & n3187 ;
  assign n31753 = ( n9590 & ~n12470 ) | ( n9590 & n28808 ) | ( ~n12470 & n28808 ) ;
  assign n31754 = ( n31751 & n31752 ) | ( n31751 & ~n31753 ) | ( n31752 & ~n31753 ) ;
  assign n31755 = n20464 & n20608 ;
  assign n31756 = n31755 ^ n29919 ^ 1'b0 ;
  assign n31757 = ( n1518 & ~n20001 ) | ( n1518 & n28566 ) | ( ~n20001 & n28566 ) ;
  assign n31758 = n4289 & n7459 ;
  assign n31759 = n31757 & n31758 ;
  assign n31760 = n31514 ^ n2546 ^ 1'b0 ;
  assign n31761 = ~n730 & n8903 ;
  assign n31762 = n28216 & n31761 ;
  assign n31763 = n14601 ^ n8500 ^ 1'b0 ;
  assign n31764 = n7526 & ~n31763 ;
  assign n31765 = n25140 ^ n292 ^ 1'b0 ;
  assign n31766 = n31764 & n31765 ;
  assign n31767 = n11108 & ~n24971 ;
  assign n31771 = n21805 ^ n1766 ^ 1'b0 ;
  assign n31768 = n2761 & ~n21666 ;
  assign n31769 = ~n2134 & n31768 ;
  assign n31770 = n29995 | n31769 ;
  assign n31772 = n31771 ^ n31770 ^ 1'b0 ;
  assign n31773 = n7496 | n10715 ;
  assign n31774 = n31773 ^ n5991 ^ 1'b0 ;
  assign n31775 = ~n6328 & n31774 ;
  assign n31776 = ~n13515 & n31775 ;
  assign n31777 = n31776 ^ n1588 ^ 1'b0 ;
  assign n31778 = ~n6370 & n21521 ;
  assign n31779 = n13166 & n31778 ;
  assign n31780 = n4480 ^ n1522 ^ 1'b0 ;
  assign n31781 = n31780 ^ n22772 ^ 1'b0 ;
  assign n31782 = ~n31779 & n31781 ;
  assign n31783 = n20442 & ~n21395 ;
  assign n31786 = n1507 & n3171 ;
  assign n31787 = ~n1507 & n31786 ;
  assign n31784 = n22046 ^ n21944 ^ 1'b0 ;
  assign n31785 = n23508 | n31784 ;
  assign n31788 = n31787 ^ n31785 ^ 1'b0 ;
  assign n31789 = ~n19527 & n31788 ;
  assign n31790 = n2273 & ~n19730 ;
  assign n31791 = n31790 ^ n22249 ^ 1'b0 ;
  assign n31792 = n10893 & ~n29629 ;
  assign n31793 = ~n7434 & n15231 ;
  assign n31794 = n2194 | n31793 ;
  assign n31800 = n2503 & ~n7228 ;
  assign n31801 = n6373 | n31800 ;
  assign n31795 = ~n4176 & n29273 ;
  assign n31796 = n31795 ^ n14007 ^ 1'b0 ;
  assign n31797 = n31796 ^ n14845 ^ 1'b0 ;
  assign n31798 = ~n9105 & n31797 ;
  assign n31799 = n14960 & n31798 ;
  assign n31802 = n31801 ^ n31799 ^ 1'b0 ;
  assign n31803 = ~n3274 & n31802 ;
  assign n31804 = n31803 ^ n27257 ^ 1'b0 ;
  assign n31805 = n29306 ^ n17495 ^ 1'b0 ;
  assign n31806 = n21038 & n30079 ;
  assign n31807 = n15543 ^ n10754 ^ 1'b0 ;
  assign n31808 = n31806 | n31807 ;
  assign n31809 = ~n709 & n19261 ;
  assign n31810 = n31809 ^ n21278 ^ n5097 ;
  assign n31815 = n10263 | n18916 ;
  assign n31811 = ~n15294 & n16033 ;
  assign n31812 = n31811 ^ x46 ^ 1'b0 ;
  assign n31813 = n1894 & ~n31812 ;
  assign n31814 = n24480 & n31813 ;
  assign n31816 = n31815 ^ n31814 ^ 1'b0 ;
  assign n31817 = n4265 & ~n31816 ;
  assign n31818 = n4647 ^ n927 ^ 1'b0 ;
  assign n31819 = n874 & ~n21650 ;
  assign n31820 = ~n31818 & n31819 ;
  assign n31821 = ~n10859 & n13027 ;
  assign n31822 = n4225 | n8059 ;
  assign n31823 = ~n7115 & n31822 ;
  assign n31824 = ~n20901 & n28303 ;
  assign n31825 = n5928 & n31824 ;
  assign n31826 = n20708 ^ n12458 ^ 1'b0 ;
  assign n31827 = n12750 & n31826 ;
  assign n31828 = n4911 & n15694 ;
  assign n31829 = n17811 & n31828 ;
  assign n31830 = n1473 & n31829 ;
  assign n31831 = n21568 & ~n27339 ;
  assign n31832 = ~n31830 & n31831 ;
  assign n31833 = n1407 | n4595 ;
  assign n31834 = n2723 | n31833 ;
  assign n31835 = n31834 ^ n3456 ^ 1'b0 ;
  assign n31836 = n2827 & ~n30395 ;
  assign n31837 = n31836 ^ n8142 ^ 1'b0 ;
  assign n31838 = n8560 & ~n31837 ;
  assign n31839 = n6735 & ~n13810 ;
  assign n31840 = n5116 | n31839 ;
  assign n31841 = n31840 ^ n2008 ^ 1'b0 ;
  assign n31842 = ~n4620 & n12912 ;
  assign n31843 = ~n7421 & n31842 ;
  assign n31844 = n31843 ^ n978 ^ 1'b0 ;
  assign n31846 = n24975 ^ n3822 ^ 1'b0 ;
  assign n31845 = n5470 & n29531 ;
  assign n31847 = n31846 ^ n31845 ^ 1'b0 ;
  assign n31849 = n7821 | n20708 ;
  assign n31850 = n28455 | n31849 ;
  assign n31848 = n1268 | n26653 ;
  assign n31851 = n31850 ^ n31848 ^ 1'b0 ;
  assign n31852 = n5709 ^ n1071 ^ 1'b0 ;
  assign n31853 = n21415 & ~n31852 ;
  assign n31854 = n14338 ^ n13307 ^ 1'b0 ;
  assign n31855 = n10954 ^ n9751 ^ 1'b0 ;
  assign n31856 = n9497 & n27585 ;
  assign n31857 = n6427 & ~n31080 ;
  assign n31858 = x131 & n31857 ;
  assign n31860 = ~n2172 & n27658 ;
  assign n31859 = ~n4009 & n14386 ;
  assign n31861 = n31860 ^ n31859 ^ 1'b0 ;
  assign n31862 = ~n23577 & n31861 ;
  assign n31863 = ( n4626 & ~n5774 ) | ( n4626 & n6413 ) | ( ~n5774 & n6413 ) ;
  assign n31864 = n31863 ^ n9896 ^ 1'b0 ;
  assign n31865 = n1195 & ~n31864 ;
  assign n31866 = n10739 | n18903 ;
  assign n31867 = ~n11952 & n31866 ;
  assign n31868 = n31867 ^ n12951 ^ 1'b0 ;
  assign n31869 = n31868 ^ n6028 ^ 1'b0 ;
  assign n31870 = n15153 & ~n25136 ;
  assign n31871 = n14198 & n20804 ;
  assign n31872 = n31871 ^ n20717 ^ 1'b0 ;
  assign n31873 = n1044 & ~n1666 ;
  assign n31874 = ~n6582 & n20971 ;
  assign n31875 = ~n15933 & n31874 ;
  assign n31876 = n1537 | n21458 ;
  assign n31877 = n17466 ^ n7630 ^ 1'b0 ;
  assign n31878 = n31761 ^ n23515 ^ 1'b0 ;
  assign n31879 = n28085 & ~n31878 ;
  assign n31880 = ~n29066 & n31879 ;
  assign n31881 = n12192 ^ n8612 ^ 1'b0 ;
  assign n31882 = ~n1914 & n31881 ;
  assign n31883 = n732 & ~n2731 ;
  assign n31884 = n22756 | n31883 ;
  assign n31885 = n1031 & n17607 ;
  assign n31886 = n31884 & n31885 ;
  assign n31887 = ~n1334 & n29022 ;
  assign n31888 = n9339 ^ n1027 ^ 1'b0 ;
  assign n31889 = n27575 & n31888 ;
  assign n31890 = n31889 ^ n17376 ^ 1'b0 ;
  assign n31891 = n16427 ^ n10877 ^ n401 ;
  assign n31892 = n2939 & n31891 ;
  assign n31893 = n17632 ^ n6215 ^ 1'b0 ;
  assign n31894 = n4134 & ~n27776 ;
  assign n31895 = n31576 & n31894 ;
  assign n31896 = n26022 ^ n2762 ^ 1'b0 ;
  assign n31897 = n2765 & ~n8553 ;
  assign n31898 = n6694 & n31897 ;
  assign n31899 = ( ~n3181 & n6339 ) | ( ~n3181 & n8453 ) | ( n6339 & n8453 ) ;
  assign n31900 = n13725 & n25037 ;
  assign n31901 = n5097 & ~n18842 ;
  assign n31902 = ~n22578 & n31901 ;
  assign n31903 = n5553 | n12691 ;
  assign n31904 = n2022 & ~n31903 ;
  assign n31905 = n9394 ^ n5215 ^ 1'b0 ;
  assign n31906 = n10885 ^ n9477 ^ 1'b0 ;
  assign n31907 = n9534 & n31906 ;
  assign n31908 = n10611 & n31907 ;
  assign n31909 = n31905 & n31908 ;
  assign n31910 = n22385 | n28948 ;
  assign n31911 = n17059 & ~n31910 ;
  assign n31912 = n12934 ^ n1075 ^ 1'b0 ;
  assign n31913 = n25101 & n31912 ;
  assign n31914 = x183 & ~n7718 ;
  assign n31915 = n1404 | n19555 ;
  assign n31916 = n9464 | n31915 ;
  assign n31917 = n1429 & ~n3736 ;
  assign n31918 = n20879 ^ x56 ^ 1'b0 ;
  assign n31919 = n31917 & ~n31918 ;
  assign n31920 = n6933 ^ n3527 ^ 1'b0 ;
  assign n31921 = n15640 ^ n3618 ^ 1'b0 ;
  assign n31922 = n4502 & ~n24528 ;
  assign n31923 = n31922 ^ n5308 ^ 1'b0 ;
  assign n31924 = ~n31921 & n31923 ;
  assign n31925 = n575 & ~n22672 ;
  assign n31926 = n1787 | n3779 ;
  assign n31927 = n23835 ^ n6556 ^ 1'b0 ;
  assign n31928 = n8616 & n11705 ;
  assign n31929 = ( n4179 & n4515 ) | ( n4179 & n31928 ) | ( n4515 & n31928 ) ;
  assign n31930 = ~n1216 & n4411 ;
  assign n31931 = n31930 ^ n12041 ^ 1'b0 ;
  assign n31932 = n31929 & n31931 ;
  assign n31933 = n2855 | n6735 ;
  assign n31934 = n12860 | n31933 ;
  assign n31935 = n2740 & n31934 ;
  assign n31936 = ~n15699 & n31935 ;
  assign n31937 = n24105 | n31936 ;
  assign n31938 = ( n2075 & n14409 ) | ( n2075 & ~n15667 ) | ( n14409 & ~n15667 ) ;
  assign n31939 = n1841 & n31938 ;
  assign n31940 = n15989 & n31939 ;
  assign n31941 = n657 & ~n31940 ;
  assign n31942 = ~n17684 & n26071 ;
  assign n31943 = n15233 ^ n540 ^ 1'b0 ;
  assign n31944 = n6951 & ~n21781 ;
  assign n31945 = n26542 & n31944 ;
  assign n31946 = n26537 ^ n3707 ^ 1'b0 ;
  assign n31947 = n29560 ^ n14470 ^ 1'b0 ;
  assign n31948 = n9393 & ~n13302 ;
  assign n31949 = n3678 & n31948 ;
  assign n31950 = ~n9394 & n30682 ;
  assign n31951 = n16072 ^ n1260 ^ 1'b0 ;
  assign n31952 = n2110 | n31951 ;
  assign n31954 = n22417 ^ n7491 ^ 1'b0 ;
  assign n31955 = n28795 & ~n31954 ;
  assign n31953 = n25437 ^ n21728 ^ 1'b0 ;
  assign n31956 = n31955 ^ n31953 ^ n29511 ;
  assign n31957 = n23519 ^ n3434 ^ 1'b0 ;
  assign n31958 = n23189 & ~n31957 ;
  assign n31959 = n5203 & n25857 ;
  assign n31960 = n31959 ^ n28123 ^ 1'b0 ;
  assign n31961 = n16728 ^ n4318 ^ 1'b0 ;
  assign n31962 = n8088 & n31961 ;
  assign n31963 = ~n18588 & n24223 ;
  assign n31964 = n3869 & ~n31963 ;
  assign n31965 = ~n3392 & n28343 ;
  assign n31966 = n31965 ^ n8094 ^ 1'b0 ;
  assign n31967 = n8907 & ~n31966 ;
  assign n31968 = n9559 & ~n31967 ;
  assign n31969 = n24024 ^ n22702 ^ n15720 ;
  assign n31970 = n20295 ^ n3758 ^ 1'b0 ;
  assign n31971 = n1361 & ~n31970 ;
  assign n31972 = n14069 ^ n3614 ^ 1'b0 ;
  assign n31973 = n1087 & n2188 ;
  assign n31974 = n26236 ^ n17304 ^ 1'b0 ;
  assign n31975 = n6285 ^ n4081 ^ 1'b0 ;
  assign n31976 = n5615 & n31975 ;
  assign n31978 = n1945 & n17072 ;
  assign n31979 = n31978 ^ n16103 ^ 1'b0 ;
  assign n31980 = n31216 ^ x219 ^ 1'b0 ;
  assign n31981 = n31979 | n31980 ;
  assign n31982 = n31981 ^ n5746 ^ 1'b0 ;
  assign n31977 = ~n16335 & n16777 ;
  assign n31983 = n31982 ^ n31977 ^ 1'b0 ;
  assign n31984 = n11565 ^ n4416 ^ 1'b0 ;
  assign n31985 = n12789 ^ x149 ^ 1'b0 ;
  assign n31986 = ~n11333 & n31985 ;
  assign n31987 = n16416 | n20211 ;
  assign n31988 = n1237 | n31987 ;
  assign n31989 = n31986 & ~n31988 ;
  assign n31990 = n2875 & n4978 ;
  assign n31991 = ( ~n11378 & n13557 ) | ( ~n11378 & n31990 ) | ( n13557 & n31990 ) ;
  assign n31992 = n31991 ^ n18895 ^ n12048 ;
  assign n31993 = n4149 | n14001 ;
  assign n31994 = n6693 & ~n31993 ;
  assign n31995 = ~n11082 & n13365 ;
  assign n31999 = ~x246 & n1725 ;
  assign n31996 = n278 | n8748 ;
  assign n31997 = n1263 | n31996 ;
  assign n31998 = ( n4054 & ~n28030 ) | ( n4054 & n31997 ) | ( ~n28030 & n31997 ) ;
  assign n32000 = n31999 ^ n31998 ^ 1'b0 ;
  assign n32001 = n6999 ^ n5852 ^ 1'b0 ;
  assign n32002 = ~n6238 & n32001 ;
  assign n32003 = n32002 ^ n8244 ^ 1'b0 ;
  assign n32004 = n21426 ^ n18046 ^ 1'b0 ;
  assign n32005 = n8202 & n9543 ;
  assign n32006 = ~n11719 & n32005 ;
  assign n32007 = n14238 ^ n5644 ^ 1'b0 ;
  assign n32008 = n11014 & n15698 ;
  assign n32009 = n20997 ^ n3054 ^ 1'b0 ;
  assign n32010 = ~n1896 & n32009 ;
  assign n32011 = n2071 | n6534 ;
  assign n32012 = n5417 | n32011 ;
  assign n32013 = n4532 | n32012 ;
  assign n32014 = n9902 ^ n5266 ^ 1'b0 ;
  assign n32015 = n3666 & ~n20328 ;
  assign n32016 = n7057 ^ n2507 ^ 1'b0 ;
  assign n32017 = n15524 ^ n10458 ^ 1'b0 ;
  assign n32018 = n9629 & n27578 ;
  assign n32019 = n9596 ^ n2044 ^ 1'b0 ;
  assign n32020 = n32019 ^ n9397 ^ 1'b0 ;
  assign n32021 = n5627 | n32020 ;
  assign n32022 = n25275 ^ n11371 ^ 1'b0 ;
  assign n32023 = n21959 ^ n4541 ^ n3140 ;
  assign n32024 = ( n5008 & n5617 ) | ( n5008 & n32023 ) | ( n5617 & n32023 ) ;
  assign n32025 = n16246 | n32024 ;
  assign n32026 = n5173 | n32025 ;
  assign n32027 = n18573 & ~n26225 ;
  assign n32028 = n3116 & n24877 ;
  assign n32029 = x86 & ~n666 ;
  assign n32030 = n13761 & n32029 ;
  assign n32031 = n18247 & n32030 ;
  assign n32032 = n12963 | n17891 ;
  assign n32033 = n6231 & n7679 ;
  assign n32034 = n4930 & n23454 ;
  assign n32035 = ~n8627 & n32034 ;
  assign n32036 = n32033 & ~n32035 ;
  assign n32037 = n32036 ^ n13109 ^ 1'b0 ;
  assign n32038 = n32032 | n32037 ;
  assign n32039 = n19199 | n21474 ;
  assign n32040 = n1815 | n32039 ;
  assign n32041 = n6821 & ~n17054 ;
  assign n32042 = n31631 ^ n8169 ^ 1'b0 ;
  assign n32043 = ~n13460 & n14993 ;
  assign n32044 = n2911 | n4499 ;
  assign n32045 = n3606 | n32044 ;
  assign n32046 = ~n2578 & n22524 ;
  assign n32047 = ~n32045 & n32046 ;
  assign n32048 = n31506 ^ n28766 ^ 1'b0 ;
  assign n32049 = n2723 & n32048 ;
  assign n32050 = n6146 & ~n25578 ;
  assign n32051 = ~n10316 & n32050 ;
  assign n32052 = n7624 ^ n562 ^ 1'b0 ;
  assign n32053 = n1743 | n32052 ;
  assign n32055 = n3755 & n9339 ;
  assign n32054 = n7689 ^ n1062 ^ 1'b0 ;
  assign n32056 = n32055 ^ n32054 ^ n3005 ;
  assign n32057 = ( n9548 & n32053 ) | ( n9548 & n32056 ) | ( n32053 & n32056 ) ;
  assign n32058 = n3774 & n4478 ;
  assign n32059 = n905 | n2861 ;
  assign n32060 = n17378 & ~n18457 ;
  assign n32061 = n5970 & n32060 ;
  assign n32062 = n32061 ^ n2470 ^ 1'b0 ;
  assign n32064 = ~n12317 & n23948 ;
  assign n32065 = n10822 & n32064 ;
  assign n32063 = n7265 | n10714 ;
  assign n32066 = n32065 ^ n32063 ^ n3521 ;
  assign n32067 = n3735 & n13521 ;
  assign n32068 = n18289 | n30952 ;
  assign n32069 = ~n707 & n5948 ;
  assign n32070 = n3252 | n7398 ;
  assign n32071 = n27668 | n32070 ;
  assign n32072 = n18159 & n32071 ;
  assign n32073 = n23393 & n25927 ;
  assign n32074 = n5373 ^ n1499 ^ 1'b0 ;
  assign n32075 = ~n8591 & n32074 ;
  assign n32076 = n32075 ^ n1678 ^ 1'b0 ;
  assign n32077 = n12440 ^ n294 ^ 1'b0 ;
  assign n32078 = n5564 & ~n32077 ;
  assign n32079 = n7798 ^ n2801 ^ 1'b0 ;
  assign n32080 = ~n18111 & n32079 ;
  assign n32081 = n23743 ^ n11191 ^ 1'b0 ;
  assign n32082 = ~n15203 & n32081 ;
  assign n32083 = n1397 & n15737 ;
  assign n32084 = n13673 ^ n8191 ^ 1'b0 ;
  assign n32085 = ~n5683 & n30104 ;
  assign n32086 = n32085 ^ n25780 ^ 1'b0 ;
  assign n32087 = n6396 & n32086 ;
  assign n32088 = n28740 ^ n1675 ^ 1'b0 ;
  assign n32089 = n20502 | n32088 ;
  assign n32090 = ~n666 & n11916 ;
  assign n32091 = n15089 ^ n12177 ^ 1'b0 ;
  assign n32092 = n22936 ^ n9327 ^ 1'b0 ;
  assign n32093 = n6797 ^ n269 ^ 1'b0 ;
  assign n32094 = n30498 ^ n19187 ^ 1'b0 ;
  assign n32095 = n12590 | n28946 ;
  assign n32096 = n18652 & n21735 ;
  assign n32097 = n1164 | n16454 ;
  assign n32098 = n16506 & ~n32097 ;
  assign n32099 = n32096 & n32098 ;
  assign n32100 = n6383 & ~n31144 ;
  assign n32101 = n32100 ^ n9454 ^ 1'b0 ;
  assign n32102 = ~n18465 & n24666 ;
  assign n32103 = n32101 & n32102 ;
  assign n32104 = ( ~n1483 & n13617 ) | ( ~n1483 & n18796 ) | ( n13617 & n18796 ) ;
  assign n32105 = n4428 & ~n32104 ;
  assign n32106 = n387 & n1942 ;
  assign n32107 = n32106 ^ n26067 ^ 1'b0 ;
  assign n32108 = n15233 & ~n30754 ;
  assign n32109 = n32108 ^ n13243 ^ 1'b0 ;
  assign n32110 = n16745 & ~n30678 ;
  assign n32111 = n32110 ^ n14823 ^ 1'b0 ;
  assign n32112 = x239 & n16868 ;
  assign n32113 = n32112 ^ n27106 ^ 1'b0 ;
  assign n32114 = ~n29069 & n32113 ;
  assign n32115 = n19373 | n21972 ;
  assign n32116 = n14545 & ~n32115 ;
  assign n32117 = n11694 ^ n4534 ^ 1'b0 ;
  assign n32118 = ( x187 & ~n7423 ) | ( x187 & n23061 ) | ( ~n7423 & n23061 ) ;
  assign n32119 = ~n7398 & n25252 ;
  assign n32120 = n27740 ^ n2380 ^ 1'b0 ;
  assign n32121 = n15227 & n26625 ;
  assign n32122 = ~n1788 & n14637 ;
  assign n32123 = ~n27681 & n32122 ;
  assign n32126 = n19273 | n30217 ;
  assign n32127 = n14071 & ~n32126 ;
  assign n32124 = n1399 | n21266 ;
  assign n32125 = n7890 | n32124 ;
  assign n32128 = n32127 ^ n32125 ^ n19746 ;
  assign n32129 = n15133 | n32128 ;
  assign n32130 = n32129 ^ n6427 ^ 1'b0 ;
  assign n32131 = n2326 & ~n20370 ;
  assign n32132 = ~n1679 & n32131 ;
  assign n32133 = n13904 | n15547 ;
  assign n32134 = ~n6413 & n18400 ;
  assign n32135 = n29594 ^ n9786 ^ 1'b0 ;
  assign n32136 = n32134 & ~n32135 ;
  assign n32137 = n7535 ^ n5378 ^ 1'b0 ;
  assign n32138 = ~n1175 & n32137 ;
  assign n32139 = n3745 ^ x26 ^ 1'b0 ;
  assign n32140 = ~n1165 & n32139 ;
  assign n32141 = x210 | n32140 ;
  assign n32142 = ~n14045 & n32141 ;
  assign n32143 = n32142 ^ n4787 ^ 1'b0 ;
  assign n32144 = ~n1723 & n18654 ;
  assign n32145 = n8411 & n29345 ;
  assign n32146 = n32145 ^ n17545 ^ 1'b0 ;
  assign n32147 = n2063 & n32146 ;
  assign n32148 = ~n32144 & n32147 ;
  assign n32149 = ~n11348 & n26586 ;
  assign n32150 = n17714 ^ n16466 ^ n5673 ;
  assign n32151 = n12478 ^ n10559 ^ 1'b0 ;
  assign n32152 = n11204 | n32151 ;
  assign n32153 = ~n9720 & n25853 ;
  assign n32154 = n32153 ^ n25454 ^ 1'b0 ;
  assign n32155 = ~n2042 & n8659 ;
  assign n32156 = ~n8314 & n32155 ;
  assign n32157 = n30166 | n32156 ;
  assign n32158 = n13854 & ~n32157 ;
  assign n32159 = n21328 ^ n4664 ^ 1'b0 ;
  assign n32160 = n21848 & n32159 ;
  assign n32161 = n23968 & n32160 ;
  assign n32162 = n12956 & n32161 ;
  assign n32163 = ~n17714 & n32162 ;
  assign n32166 = n1573 & ~n7395 ;
  assign n32167 = n13111 & n32166 ;
  assign n32164 = n10401 ^ n3578 ^ 1'b0 ;
  assign n32165 = n27374 & ~n32164 ;
  assign n32168 = n32167 ^ n32165 ^ 1'b0 ;
  assign n32169 = n32168 ^ n2169 ^ 1'b0 ;
  assign n32170 = n19335 ^ n14707 ^ 1'b0 ;
  assign n32171 = n9717 | n32170 ;
  assign n32172 = n8594 & n21246 ;
  assign n32173 = n32172 ^ n7223 ^ 1'b0 ;
  assign n32174 = n14504 & ~n17489 ;
  assign n32175 = ~n5501 & n24917 ;
  assign n32176 = ~n470 & n26886 ;
  assign n32177 = ~n8379 & n19865 ;
  assign n32178 = n14493 & ~n22707 ;
  assign n32179 = n1239 & n2591 ;
  assign n32180 = n5085 & ~n10477 ;
  assign n32181 = n5861 | n32180 ;
  assign n32182 = n18819 | n32181 ;
  assign n32183 = ~n9179 & n15746 ;
  assign n32184 = ( ~n666 & n14131 ) | ( ~n666 & n17497 ) | ( n14131 & n17497 ) ;
  assign n32185 = n10547 | n24031 ;
  assign n32186 = n29086 | n32185 ;
  assign n32187 = ~n3487 & n32186 ;
  assign n32188 = ( n22343 & n30592 ) | ( n22343 & n32187 ) | ( n30592 & n32187 ) ;
  assign n32190 = x111 & n608 ;
  assign n32189 = n7535 & n9560 ;
  assign n32191 = n32190 ^ n32189 ^ 1'b0 ;
  assign n32192 = n7593 & ~n32191 ;
  assign n32194 = n7554 & ~n23973 ;
  assign n32193 = n6583 & ~n17349 ;
  assign n32195 = n32194 ^ n32193 ^ 1'b0 ;
  assign n32196 = ~n3509 & n25274 ;
  assign n32198 = n15128 & ~n23325 ;
  assign n32199 = ~n753 & n32198 ;
  assign n32200 = ~n2425 & n32199 ;
  assign n32197 = ~n24025 & n28066 ;
  assign n32201 = n32200 ^ n32197 ^ 1'b0 ;
  assign n32202 = ~n4190 & n25579 ;
  assign n32203 = n32202 ^ n4169 ^ 1'b0 ;
  assign n32204 = n10270 & n23696 ;
  assign n32205 = n32204 ^ n8022 ^ 1'b0 ;
  assign n32206 = n20760 ^ n18796 ^ 1'b0 ;
  assign n32208 = ~n9229 & n15806 ;
  assign n32209 = n2371 & ~n32208 ;
  assign n32207 = n13118 & ~n18481 ;
  assign n32210 = n32209 ^ n32207 ^ 1'b0 ;
  assign n32211 = n24697 ^ n1926 ^ 1'b0 ;
  assign n32212 = ~n669 & n32211 ;
  assign n32213 = n32212 ^ n21941 ^ 1'b0 ;
  assign n32214 = n7709 & n18395 ;
  assign n32215 = n32214 ^ n16567 ^ 1'b0 ;
  assign n32216 = n2432 | n22906 ;
  assign n32217 = n32216 ^ n6785 ^ 1'b0 ;
  assign n32218 = n30003 ^ n5300 ^ 1'b0 ;
  assign n32219 = ~x235 & n13324 ;
  assign n32220 = n17841 ^ n1622 ^ 1'b0 ;
  assign n32221 = n26037 ^ n1488 ^ 1'b0 ;
  assign n32222 = n25432 ^ n8043 ^ 1'b0 ;
  assign n32223 = n32222 ^ n11915 ^ 1'b0 ;
  assign n32224 = n14288 | n32223 ;
  assign n32225 = n32221 | n32224 ;
  assign n32226 = n12008 ^ n8761 ^ n7079 ;
  assign n32229 = n15812 ^ n542 ^ 1'b0 ;
  assign n32230 = n11689 & n32229 ;
  assign n32231 = n18846 ^ n4400 ^ 1'b0 ;
  assign n32232 = n32230 & ~n32231 ;
  assign n32227 = n275 & ~n24808 ;
  assign n32228 = ~n27672 & n32227 ;
  assign n32233 = n32232 ^ n32228 ^ 1'b0 ;
  assign n32234 = n26169 | n32233 ;
  assign n32235 = n22641 ^ n13808 ^ 1'b0 ;
  assign n32236 = n4939 & n32235 ;
  assign n32237 = n3688 & n6440 ;
  assign n32238 = n32237 ^ n12721 ^ 1'b0 ;
  assign n32243 = ~n8957 & n11481 ;
  assign n32244 = ~n1795 & n32243 ;
  assign n32245 = n385 | n32244 ;
  assign n32246 = n32245 ^ n9807 ^ 1'b0 ;
  assign n32247 = n7251 | n32246 ;
  assign n32248 = n9734 | n32247 ;
  assign n32249 = n32248 ^ n31818 ^ 1'b0 ;
  assign n32239 = n23398 ^ n11001 ^ 1'b0 ;
  assign n32240 = n1232 | n25805 ;
  assign n32241 = n32239 | n32240 ;
  assign n32242 = n17046 & n32241 ;
  assign n32250 = n32249 ^ n32242 ^ 1'b0 ;
  assign n32251 = n17046 | n32250 ;
  assign n32252 = n22150 ^ n12559 ^ 1'b0 ;
  assign n32253 = ~n30926 & n32252 ;
  assign n32254 = n1164 & n11109 ;
  assign n32255 = n32254 ^ n12373 ^ 1'b0 ;
  assign n32256 = n2340 | n18402 ;
  assign n32257 = n32256 ^ n800 ^ 1'b0 ;
  assign n32258 = ~n7560 & n32257 ;
  assign n32259 = ~n27072 & n32258 ;
  assign n32260 = x87 & n7668 ;
  assign n32261 = ~n23749 & n32260 ;
  assign n32262 = n7928 ^ n4926 ^ 1'b0 ;
  assign n32263 = ~n32191 & n32262 ;
  assign n32264 = n15852 & n32263 ;
  assign n32265 = ~n11423 & n32264 ;
  assign n32266 = n26896 ^ n23244 ^ 1'b0 ;
  assign n32267 = n27367 & ~n32266 ;
  assign n32268 = n13813 ^ n8663 ^ 1'b0 ;
  assign n32269 = n3120 & ~n6900 ;
  assign n32270 = n32269 ^ n1630 ^ 1'b0 ;
  assign n32271 = n1405 & ~n10686 ;
  assign n32272 = n7649 | n32271 ;
  assign n32273 = n926 & ~n4891 ;
  assign n32274 = n2586 & ~n6283 ;
  assign n32275 = ~n32273 & n32274 ;
  assign n32276 = n32092 ^ n12652 ^ 1'b0 ;
  assign n32277 = n27187 & ~n30338 ;
  assign n32278 = n9482 ^ n9253 ^ 1'b0 ;
  assign n32279 = ~n30107 & n32278 ;
  assign n32280 = ~n6108 & n9589 ;
  assign n32281 = n31748 ^ n20797 ^ 1'b0 ;
  assign n32282 = n1111 & n6398 ;
  assign n32283 = n8333 & n32282 ;
  assign n32284 = n6089 | n22164 ;
  assign n32285 = ~n3695 & n3959 ;
  assign n32286 = n14941 & n32285 ;
  assign n32287 = n32286 ^ n13586 ^ 1'b0 ;
  assign n32288 = n15096 & n18448 ;
  assign n32289 = n5203 ^ n2897 ^ 1'b0 ;
  assign n32290 = n32288 & ~n32289 ;
  assign n32291 = n18215 & ~n30112 ;
  assign n32292 = n13619 ^ n3697 ^ 1'b0 ;
  assign n32293 = n3332 | n32292 ;
  assign n32294 = ~n4576 & n32012 ;
  assign n32295 = n4576 & n32294 ;
  assign n32296 = n32295 ^ n12094 ^ 1'b0 ;
  assign n32297 = ~n32293 & n32296 ;
  assign n32298 = ~n6116 & n23813 ;
  assign n32299 = n5577 & n32298 ;
  assign n32300 = n1397 & ~n32299 ;
  assign n32301 = n8977 & n32300 ;
  assign n32303 = n1658 & ~n9491 ;
  assign n32304 = n32303 ^ n11536 ^ 1'b0 ;
  assign n32302 = n967 & ~n1833 ;
  assign n32305 = n32304 ^ n32302 ^ 1'b0 ;
  assign n32306 = n2065 | n3342 ;
  assign n32307 = n32306 ^ n18441 ^ x76 ;
  assign n32308 = ~n2765 & n21386 ;
  assign n32309 = n32308 ^ n21014 ^ 1'b0 ;
  assign n32310 = n29801 & n32309 ;
  assign n32311 = ~n25335 & n32310 ;
  assign n32312 = n17172 ^ n4960 ^ 1'b0 ;
  assign n32313 = n13796 & ~n32312 ;
  assign n32314 = n13458 & n17979 ;
  assign n32315 = n5646 | n32314 ;
  assign n32316 = n6134 | n23159 ;
  assign n32317 = n17249 | n32316 ;
  assign n32318 = n17358 & n22279 ;
  assign n32319 = n20587 | n32318 ;
  assign n32320 = n26022 | n32319 ;
  assign n32321 = n3869 | n8550 ;
  assign n32322 = n12213 ^ n1249 ^ 1'b0 ;
  assign n32323 = n32321 & ~n32322 ;
  assign n32324 = n1407 & ~n22482 ;
  assign n32325 = n32324 ^ n7477 ^ 1'b0 ;
  assign n32326 = n9744 & ~n14907 ;
  assign n32327 = ~n1318 & n32326 ;
  assign n32328 = ~n6031 & n18088 ;
  assign n32329 = n23682 | n32328 ;
  assign n32330 = n32329 ^ n13373 ^ 1'b0 ;
  assign n32331 = ~n32327 & n32330 ;
  assign n32332 = n32331 ^ n2620 ^ 1'b0 ;
  assign n32333 = n32332 ^ n16079 ^ 1'b0 ;
  assign n32334 = n6932 & ~n32333 ;
  assign n32335 = ( n15824 & n32325 ) | ( n15824 & ~n32334 ) | ( n32325 & ~n32334 ) ;
  assign n32336 = ~n21579 & n25713 ;
  assign n32337 = n10963 ^ x67 ^ 1'b0 ;
  assign n32338 = ~n23337 & n32337 ;
  assign n32339 = ~n11705 & n32338 ;
  assign n32340 = n15694 & ~n16642 ;
  assign n32341 = n17038 ^ n14856 ^ 1'b0 ;
  assign n32345 = n9428 & n9885 ;
  assign n32346 = ~n20695 & n32345 ;
  assign n32342 = n13919 ^ n1366 ^ 1'b0 ;
  assign n32343 = x174 | n32342 ;
  assign n32344 = n13505 | n32343 ;
  assign n32347 = n32346 ^ n32344 ^ 1'b0 ;
  assign n32348 = n21041 ^ n6031 ^ 1'b0 ;
  assign n32349 = n32347 | n32348 ;
  assign n32350 = n2309 & ~n5248 ;
  assign n32351 = n32350 ^ n21297 ^ 1'b0 ;
  assign n32352 = n31990 & ~n32351 ;
  assign n32353 = n7355 | n32352 ;
  assign n32355 = n3376 & ~n24637 ;
  assign n32354 = ~n15556 & n26779 ;
  assign n32356 = n32355 ^ n32354 ^ 1'b0 ;
  assign n32357 = n743 | n2293 ;
  assign n32358 = n32357 ^ n30586 ^ 1'b0 ;
  assign n32359 = n5373 & n5973 ;
  assign n32360 = n32359 ^ n6051 ^ 1'b0 ;
  assign n32361 = n17614 ^ n3669 ^ 1'b0 ;
  assign n32362 = ~n651 & n32361 ;
  assign n32363 = ~n17068 & n24677 ;
  assign n32364 = ~n32362 & n32363 ;
  assign n32365 = n13617 & n18153 ;
  assign n32366 = n32365 ^ n27288 ^ 1'b0 ;
  assign n32367 = n11169 | n12726 ;
  assign n32368 = n8835 ^ n3634 ^ 1'b0 ;
  assign n32369 = n26136 & n32368 ;
  assign n32370 = n15003 ^ n7864 ^ n694 ;
  assign n32371 = n9470 & n10010 ;
  assign n32372 = ~n21676 & n32371 ;
  assign n32373 = ~n6154 & n25538 ;
  assign n32374 = ~n9382 & n32373 ;
  assign n32375 = n6513 & ~n12795 ;
  assign n32376 = n32375 ^ n3377 ^ 1'b0 ;
  assign n32377 = n1260 | n6934 ;
  assign n32378 = n32377 ^ n7032 ^ 1'b0 ;
  assign n32379 = n19595 | n23210 ;
  assign n32380 = n19364 & ~n32379 ;
  assign n32381 = n10751 | n14696 ;
  assign n32382 = n32381 ^ n1395 ^ 1'b0 ;
  assign n32385 = n2716 & ~n8754 ;
  assign n32383 = n8995 & ~n22237 ;
  assign n32384 = n32383 ^ n8683 ^ 1'b0 ;
  assign n32386 = n32385 ^ n32384 ^ 1'b0 ;
  assign n32387 = ( n7698 & n11851 ) | ( n7698 & ~n31881 ) | ( n11851 & ~n31881 ) ;
  assign n32388 = n14560 & ~n25241 ;
  assign n32389 = n21623 ^ n6182 ^ n2428 ;
  assign n32390 = n32389 ^ n19352 ^ 1'b0 ;
  assign n32391 = n415 & n6752 ;
  assign n32392 = n20085 ^ n12833 ^ 1'b0 ;
  assign n32393 = ~n1548 & n21487 ;
  assign n32394 = n12963 ^ n7113 ^ n4676 ;
  assign n32395 = n29460 & ~n32394 ;
  assign n32396 = n2776 | n3670 ;
  assign n32397 = n6715 & ~n29581 ;
  assign n32398 = n20903 & n32397 ;
  assign n32399 = ~n3416 & n17164 ;
  assign n32400 = n6317 & n32399 ;
  assign n32401 = n19911 | n32400 ;
  assign n32402 = n17370 | n32401 ;
  assign n32404 = n1859 & ~n5629 ;
  assign n32403 = n5292 & n9299 ;
  assign n32405 = n32404 ^ n32403 ^ 1'b0 ;
  assign n32406 = n32402 & ~n32405 ;
  assign n32407 = n32406 ^ n27712 ^ 1'b0 ;
  assign n32408 = n20992 | n30798 ;
  assign n32409 = n32408 ^ n3614 ^ 1'b0 ;
  assign n32410 = ~n994 & n13593 ;
  assign n32411 = ~n5185 & n32410 ;
  assign n32412 = n14951 | n32411 ;
  assign n32413 = n3093 | n32412 ;
  assign n32414 = n32413 ^ n23196 ^ 1'b0 ;
  assign n32415 = n7766 | n32414 ;
  assign n32416 = n921 & ~n32415 ;
  assign n32417 = n4991 & ~n22127 ;
  assign n32418 = n32417 ^ n17007 ^ 1'b0 ;
  assign n32419 = ~n290 & n14995 ;
  assign n32420 = n1514 & ~n6267 ;
  assign n32421 = n32420 ^ n904 ^ 1'b0 ;
  assign n32422 = n19021 ^ n1996 ^ 1'b0 ;
  assign n32423 = n3824 & n11363 ;
  assign n32424 = ~n18677 & n32423 ;
  assign n32425 = n2394 & ~n14901 ;
  assign n32426 = n32425 ^ n23196 ^ 1'b0 ;
  assign n32427 = ~n7876 & n13922 ;
  assign n32428 = n4091 & ~n32427 ;
  assign n32429 = ~n2266 & n26418 ;
  assign n32430 = ~n9744 & n32429 ;
  assign n32431 = n880 | n8977 ;
  assign n32432 = ~n1154 & n4177 ;
  assign n32433 = n7872 | n32432 ;
  assign n32434 = n32433 ^ n8568 ^ 1'b0 ;
  assign n32435 = n12394 & n32434 ;
  assign n32436 = n32435 ^ n24211 ^ n13943 ;
  assign n32437 = n3558 & ~n15781 ;
  assign n32438 = n723 & n32437 ;
  assign n32439 = n9133 ^ n4300 ^ 1'b0 ;
  assign n32440 = n3855 & ~n8977 ;
  assign n32441 = n20873 ^ n15617 ^ 1'b0 ;
  assign n32442 = n9620 & n32441 ;
  assign n32443 = n32442 ^ n30633 ^ 1'b0 ;
  assign n32446 = n25222 ^ n4512 ^ 1'b0 ;
  assign n32447 = x60 & n32446 ;
  assign n32445 = ~n3331 & n16797 ;
  assign n32448 = n32447 ^ n32445 ^ 1'b0 ;
  assign n32449 = n1661 & n32448 ;
  assign n32450 = n13675 & n32449 ;
  assign n32444 = ~n14822 & n29218 ;
  assign n32451 = n32450 ^ n32444 ^ 1'b0 ;
  assign n32452 = n7263 & n32451 ;
  assign n32453 = n17039 ^ n11899 ^ n8967 ;
  assign n32454 = n1656 & ~n32453 ;
  assign n32455 = n16446 ^ n888 ^ 1'b0 ;
  assign n32456 = n32454 & n32455 ;
  assign n32457 = n13370 ^ n10724 ^ 1'b0 ;
  assign n32458 = n14352 & n24656 ;
  assign n32459 = n3795 | n6437 ;
  assign n32460 = n32459 ^ n518 ^ 1'b0 ;
  assign n32461 = n32460 ^ n1974 ^ 1'b0 ;
  assign n32462 = n19432 & ~n32461 ;
  assign n32463 = n31720 & ~n32462 ;
  assign n32464 = ~n6154 & n12745 ;
  assign n32465 = n10790 & ~n32464 ;
  assign n32466 = n17085 & n32465 ;
  assign n32467 = n6745 ^ n5171 ^ 1'b0 ;
  assign n32468 = ( n11264 & n12259 ) | ( n11264 & ~n15306 ) | ( n12259 & ~n15306 ) ;
  assign n32469 = n32467 & n32468 ;
  assign n32470 = n9431 & n32146 ;
  assign n32471 = n32470 ^ n28087 ^ 1'b0 ;
  assign n32472 = n30950 ^ n28197 ^ 1'b0 ;
  assign n32473 = ~n3599 & n32472 ;
  assign n32474 = n10714 ^ n538 ^ 1'b0 ;
  assign n32475 = ~n2143 & n32474 ;
  assign n32476 = n32475 ^ n5503 ^ 1'b0 ;
  assign n32477 = n19474 & n32476 ;
  assign n32478 = n11498 ^ x31 ^ 1'b0 ;
  assign n32479 = n32478 ^ n3714 ^ 1'b0 ;
  assign n32480 = n4273 ^ n1732 ^ 1'b0 ;
  assign n32481 = ~n32479 & n32480 ;
  assign n32482 = n16503 & n21608 ;
  assign n32483 = n19833 ^ n6584 ^ 1'b0 ;
  assign n32484 = n25390 & ~n32483 ;
  assign n32485 = n8556 ^ n1622 ^ 1'b0 ;
  assign n32486 = n32485 ^ n8223 ^ x129 ;
  assign n32487 = n32486 ^ n285 ^ 1'b0 ;
  assign n32488 = n2100 & ~n17732 ;
  assign n32489 = n10327 ^ n5802 ^ 1'b0 ;
  assign n32490 = n17286 & ~n32489 ;
  assign n32491 = n271 & n32490 ;
  assign n32492 = n7416 & n32491 ;
  assign n32493 = n19796 ^ n8191 ^ 1'b0 ;
  assign n32494 = ~n25685 & n29221 ;
  assign n32495 = n19593 & n32494 ;
  assign n32496 = n9539 | n17575 ;
  assign n32497 = n21200 & ~n32496 ;
  assign n32498 = n894 | n23140 ;
  assign n32499 = n32497 & ~n32498 ;
  assign n32500 = n12594 ^ n2787 ^ 1'b0 ;
  assign n32501 = n32500 ^ n10777 ^ 1'b0 ;
  assign n32502 = n11565 & n23886 ;
  assign n32503 = n1361 & ~n17856 ;
  assign n32504 = n30918 | n32503 ;
  assign n32505 = n9895 & n12306 ;
  assign n32506 = n32505 ^ n15593 ^ 1'b0 ;
  assign n32507 = n10754 | n32506 ;
  assign n32508 = n1285 | n3662 ;
  assign n32509 = n3662 & ~n32508 ;
  assign n32510 = x60 & n32509 ;
  assign n32511 = n32510 ^ n1723 ^ 1'b0 ;
  assign n32512 = n1111 & ~n15187 ;
  assign n32513 = n32511 & n32512 ;
  assign n32514 = n13592 ^ n8880 ^ n2826 ;
  assign n32515 = n27132 ^ n18879 ^ 1'b0 ;
  assign n32516 = n32514 & n32515 ;
  assign n32517 = n4055 ^ n2373 ^ 1'b0 ;
  assign n32518 = ~x22 & n32517 ;
  assign n32519 = n8600 & ~n9589 ;
  assign n32520 = n10935 & n32519 ;
  assign n32521 = n3230 & n12536 ;
  assign n32522 = ~x1 & n838 ;
  assign n32523 = n821 & n32522 ;
  assign n32524 = n16181 ^ n15782 ^ 1'b0 ;
  assign n32525 = n32523 | n32524 ;
  assign n32526 = n1228 & n13812 ;
  assign n32527 = ~n10126 & n32526 ;
  assign n32528 = n32527 ^ n14795 ^ n1260 ;
  assign n32529 = n10638 ^ n7070 ^ 1'b0 ;
  assign n32530 = n6087 & ~n14344 ;
  assign n32531 = n1656 | n6350 ;
  assign n32532 = ( n11820 & ~n32530 ) | ( n11820 & n32531 ) | ( ~n32530 & n32531 ) ;
  assign n32533 = n32532 ^ n16389 ^ 1'b0 ;
  assign n32534 = n2241 & ~n32533 ;
  assign n32535 = n923 & n11220 ;
  assign n32536 = ~n4455 & n9881 ;
  assign n32537 = n32536 ^ n5929 ^ 1'b0 ;
  assign n32538 = n13822 & n31053 ;
  assign n32539 = ~n3581 & n32538 ;
  assign n32540 = ~n21753 & n32539 ;
  assign n32541 = ( n715 & n8460 ) | ( n715 & ~n29930 ) | ( n8460 & ~n29930 ) ;
  assign n32542 = ~n17167 & n20149 ;
  assign n32543 = ~n5840 & n32542 ;
  assign n32544 = n1512 & ~n22733 ;
  assign n32545 = ~n32543 & n32544 ;
  assign n32546 = ( n8148 & n18917 ) | ( n8148 & ~n26064 ) | ( n18917 & ~n26064 ) ;
  assign n32547 = ~n5835 & n10801 ;
  assign n32548 = ( n286 & n9430 ) | ( n286 & n32547 ) | ( n9430 & n32547 ) ;
  assign n32549 = n32548 ^ n21497 ^ 1'b0 ;
  assign n32550 = n32546 & ~n32549 ;
  assign n32551 = n2250 & ~n11887 ;
  assign n32552 = ~n32550 & n32551 ;
  assign n32553 = n15048 ^ n2671 ^ 1'b0 ;
  assign n32554 = n4323 ^ x174 ^ 1'b0 ;
  assign n32555 = n11259 & n22363 ;
  assign n32556 = n28332 ^ n26728 ^ n7569 ;
  assign n32557 = n5458 | n20738 ;
  assign n32558 = n13157 & n21975 ;
  assign n32559 = x61 | n16690 ;
  assign n32560 = n1646 & ~n3842 ;
  assign n32561 = n18973 | n26403 ;
  assign n32562 = ~n7411 & n10591 ;
  assign n32563 = n32562 ^ n9947 ^ 1'b0 ;
  assign n32564 = n20401 ^ n7253 ^ 1'b0 ;
  assign n32565 = ~n32563 & n32564 ;
  assign n32566 = n22109 & n32447 ;
  assign n32567 = n19727 & n32566 ;
  assign n32568 = ~n5116 & n14866 ;
  assign n32569 = n25388 | n32568 ;
  assign n32570 = ~n3165 & n5987 ;
  assign n32571 = ~n5083 & n32570 ;
  assign n32572 = n6394 | n32571 ;
  assign n32573 = n15090 ^ n11574 ^ 1'b0 ;
  assign n32574 = n25576 & ~n32573 ;
  assign n32575 = n6584 & ~n32574 ;
  assign n32576 = n29789 ^ x207 ^ 1'b0 ;
  assign n32577 = n2185 | n6938 ;
  assign n32578 = n27665 ^ n19621 ^ 1'b0 ;
  assign n32579 = n18972 ^ n13904 ^ n10432 ;
  assign n32580 = x201 | n13818 ;
  assign n32581 = ~n11443 & n15297 ;
  assign n32582 = n16443 & ~n32581 ;
  assign n32583 = n13714 ^ n8876 ^ 1'b0 ;
  assign n32584 = ~n20232 & n32583 ;
  assign n32585 = n32584 ^ n16055 ^ n4920 ;
  assign n32586 = n31773 ^ n8093 ^ 1'b0 ;
  assign n32587 = n2048 & ~n5883 ;
  assign n32589 = n13330 ^ n9122 ^ 1'b0 ;
  assign n32588 = ~n3319 & n20796 ;
  assign n32590 = n32589 ^ n32588 ^ 1'b0 ;
  assign n32591 = n26630 ^ n11500 ^ 1'b0 ;
  assign n32594 = n8239 & ~n8369 ;
  assign n32592 = ~n17475 & n22388 ;
  assign n32593 = ~n9333 & n32592 ;
  assign n32595 = n32594 ^ n32593 ^ 1'b0 ;
  assign n32596 = n9076 & ~n16211 ;
  assign n32597 = n3308 & n32596 ;
  assign n32598 = n32597 ^ n5864 ^ 1'b0 ;
  assign n32599 = n31238 ^ n14089 ^ 1'b0 ;
  assign n32603 = n30183 ^ n9807 ^ x95 ;
  assign n32604 = n10875 ^ n5675 ^ 1'b0 ;
  assign n32605 = ~n32603 & n32604 ;
  assign n32606 = ( ~n18063 & n30220 ) | ( ~n18063 & n32605 ) | ( n30220 & n32605 ) ;
  assign n32600 = n8261 | n8606 ;
  assign n32601 = n3739 | n32600 ;
  assign n32602 = n7668 & ~n32601 ;
  assign n32607 = n32606 ^ n32602 ^ 1'b0 ;
  assign n32608 = n26316 ^ n9449 ^ 1'b0 ;
  assign n32609 = n28930 ^ n9564 ^ 1'b0 ;
  assign n32610 = n26538 ^ n16561 ^ 1'b0 ;
  assign n32611 = ~n21706 & n32610 ;
  assign n32612 = n2861 | n12452 ;
  assign n32613 = n20151 & ~n32612 ;
  assign n32614 = n6517 & n17627 ;
  assign n32615 = n4874 & n32614 ;
  assign n32616 = ~n2264 & n5203 ;
  assign n32617 = n14471 & n32616 ;
  assign n32619 = n6750 & n26100 ;
  assign n32620 = n32619 ^ n16792 ^ 1'b0 ;
  assign n32621 = n29626 ^ n18875 ^ 1'b0 ;
  assign n32622 = ~n32620 & n32621 ;
  assign n32618 = n21753 & ~n24999 ;
  assign n32623 = n32622 ^ n32618 ^ 1'b0 ;
  assign n32624 = n3186 | n20918 ;
  assign n32625 = n25759 ^ n19921 ^ 1'b0 ;
  assign n32626 = n12172 | n32625 ;
  assign n32627 = n2336 | n15743 ;
  assign n32628 = n14438 ^ n6563 ^ 1'b0 ;
  assign n32629 = x163 & ~n19967 ;
  assign n32630 = ~n32628 & n32629 ;
  assign n32631 = n5424 & n11194 ;
  assign n32632 = n3576 & n32631 ;
  assign n32633 = n32632 ^ n9113 ^ 1'b0 ;
  assign n32634 = ~n956 & n11453 ;
  assign n32635 = n11899 & n32634 ;
  assign n32636 = n4888 | n32635 ;
  assign n32637 = n32636 ^ n521 ^ 1'b0 ;
  assign n32638 = n32633 & n32637 ;
  assign n32639 = n32638 ^ n19639 ^ 1'b0 ;
  assign n32640 = n29125 ^ n10154 ^ 1'b0 ;
  assign n32641 = n10120 & ~n32640 ;
  assign n32642 = n32641 ^ n11856 ^ 1'b0 ;
  assign n32643 = ~n5476 & n26921 ;
  assign n32644 = n31557 ^ n9389 ^ 1'b0 ;
  assign n32645 = n32643 | n32644 ;
  assign n32646 = n415 & n13956 ;
  assign n32647 = n32646 ^ n13912 ^ 1'b0 ;
  assign n32648 = n15565 & ~n26518 ;
  assign n32649 = n11506 & n32648 ;
  assign n32650 = n25785 | n27904 ;
  assign n32651 = ~n20784 & n22974 ;
  assign n32652 = n6469 ^ n6285 ^ 1'b0 ;
  assign n32653 = n17819 & n31055 ;
  assign n32654 = n30923 ^ n1683 ^ 1'b0 ;
  assign n32655 = ~n4859 & n32304 ;
  assign n32656 = n28849 & ~n32655 ;
  assign n32657 = n32656 ^ n13089 ^ 1'b0 ;
  assign n32658 = n2537 & ~n6196 ;
  assign n32659 = n5692 & n32658 ;
  assign n32660 = x3 & n32659 ;
  assign n32661 = n19203 ^ n9454 ^ 1'b0 ;
  assign n32662 = n20139 ^ n1345 ^ 1'b0 ;
  assign n32663 = n32488 ^ n21884 ^ 1'b0 ;
  assign n32664 = ~n22814 & n32663 ;
  assign n32665 = n9762 ^ n7046 ^ n5585 ;
  assign n32666 = n32665 ^ n30181 ^ 1'b0 ;
  assign n32667 = n30373 & n32666 ;
  assign n32668 = ~n2510 & n12291 ;
  assign n32669 = n32668 ^ n27904 ^ n2476 ;
  assign n32670 = n32669 ^ n16767 ^ 1'b0 ;
  assign n32671 = ~n690 & n11302 ;
  assign n32672 = ~n9382 & n32671 ;
  assign n32673 = n12404 | n32672 ;
  assign n32674 = n32673 ^ n9160 ^ 1'b0 ;
  assign n32675 = ~x24 & n17410 ;
  assign n32676 = n17014 ^ n1991 ^ 1'b0 ;
  assign n32677 = n3618 & ~n27049 ;
  assign n32678 = n32676 & ~n32677 ;
  assign n32679 = n12035 & ~n32207 ;
  assign n32680 = n12975 & ~n20954 ;
  assign n32681 = n27212 & n32680 ;
  assign n32682 = ~n2318 & n32681 ;
  assign n32683 = n1321 & n4356 ;
  assign n32684 = ~n5902 & n32683 ;
  assign n32685 = n27218 | n29547 ;
  assign n32686 = n11623 ^ n2861 ^ 1'b0 ;
  assign n32687 = n5835 ^ n5045 ^ 1'b0 ;
  assign n32688 = n3046 & ~n32687 ;
  assign n32689 = n10488 ^ n6271 ^ 1'b0 ;
  assign n32690 = n32688 & n32689 ;
  assign n32691 = ~n11695 & n32690 ;
  assign n32692 = n13606 & ~n15235 ;
  assign n32693 = ~n1442 & n32692 ;
  assign n32694 = ~n3207 & n13277 ;
  assign n32695 = n12833 & n26249 ;
  assign n32702 = n1031 | n1326 ;
  assign n32703 = n1326 & ~n32702 ;
  assign n32696 = n1427 | n3223 ;
  assign n32697 = n3223 & ~n32696 ;
  assign n32698 = n6493 & ~n32697 ;
  assign n32699 = ~n6493 & n32698 ;
  assign n32700 = n3286 | n32699 ;
  assign n32701 = n1039 | n32700 ;
  assign n32704 = n32703 ^ n32701 ^ 1'b0 ;
  assign n32705 = n4791 & ~n9624 ;
  assign n32706 = ~n4426 & n32705 ;
  assign n32707 = n17767 ^ n7709 ^ 1'b0 ;
  assign n32708 = ~n23729 & n32707 ;
  assign n32709 = ~n32706 & n32708 ;
  assign n32710 = n32704 & n32709 ;
  assign n32711 = n387 & ~n32453 ;
  assign n32712 = n17136 & n32711 ;
  assign n32713 = n16110 | n32712 ;
  assign n32714 = n25526 ^ n9773 ^ n3599 ;
  assign n32715 = n6049 | n32714 ;
  assign n32716 = ~n1809 & n11961 ;
  assign n32717 = n9186 ^ n2035 ^ 1'b0 ;
  assign n32718 = n32717 ^ n6516 ^ n2235 ;
  assign n32719 = n32718 ^ n2733 ^ 1'b0 ;
  assign n32720 = n20576 & n25034 ;
  assign n32721 = ~n9059 & n20793 ;
  assign n32722 = n809 & n13811 ;
  assign n32723 = ~n265 & n32722 ;
  assign n32724 = ~n23499 & n32723 ;
  assign n32726 = n16931 & n27985 ;
  assign n32727 = n32726 ^ n9697 ^ 1'b0 ;
  assign n32725 = n12018 | n25244 ;
  assign n32728 = n32727 ^ n32725 ^ 1'b0 ;
  assign n32729 = n12389 ^ n3187 ^ 1'b0 ;
  assign n32730 = n13661 & n32729 ;
  assign n32731 = n32730 ^ n23489 ^ n11695 ;
  assign n32732 = n7440 & n19265 ;
  assign n32733 = n23322 ^ n5942 ^ 1'b0 ;
  assign n32734 = n8192 & n10623 ;
  assign n32735 = n10758 & n21371 ;
  assign n32736 = n32735 ^ n3766 ^ 1'b0 ;
  assign n32737 = n32736 ^ n4444 ^ 1'b0 ;
  assign n32738 = ~n2371 & n17192 ;
  assign n32739 = ~n32737 & n32738 ;
  assign n32740 = n28947 ^ n23034 ^ 1'b0 ;
  assign n32741 = n31622 | n32740 ;
  assign n32742 = ~n3870 & n9149 ;
  assign n32743 = ~n18392 & n32742 ;
  assign n32744 = n15436 | n32743 ;
  assign n32745 = n10521 ^ n6587 ^ x240 ;
  assign n32746 = n19972 & n32745 ;
  assign n32747 = n548 & ~n10422 ;
  assign n32748 = ~n2040 & n32747 ;
  assign n32749 = n31757 ^ n1079 ^ 1'b0 ;
  assign n32750 = n23630 & n32749 ;
  assign n32751 = ~n720 & n5112 ;
  assign n32752 = ~n16284 & n32751 ;
  assign n32753 = n7269 | n16288 ;
  assign n32754 = n32753 ^ n1988 ^ 1'b0 ;
  assign n32755 = n32754 ^ n23387 ^ 1'b0 ;
  assign n32756 = ( ~n9861 & n16063 ) | ( ~n9861 & n32755 ) | ( n16063 & n32755 ) ;
  assign n32757 = n12535 & ~n21198 ;
  assign n32758 = ~n4094 & n32757 ;
  assign n32759 = n510 | n29582 ;
  assign n32760 = ( n3865 & ~n4021 ) | ( n3865 & n21319 ) | ( ~n4021 & n21319 ) ;
  assign n32761 = n19774 | n32760 ;
  assign n32762 = n9168 ^ n1133 ^ 1'b0 ;
  assign n32763 = n21377 ^ n8258 ^ 1'b0 ;
  assign n32764 = ~n1361 & n32763 ;
  assign n32765 = ~n28622 & n29816 ;
  assign n32766 = n32765 ^ n10192 ^ 1'b0 ;
  assign n32767 = n32766 ^ n23416 ^ 1'b0 ;
  assign n32768 = n20612 | n29978 ;
  assign n32769 = n19090 & ~n32768 ;
  assign n32770 = n15382 ^ n536 ^ 1'b0 ;
  assign n32771 = n31340 & ~n32770 ;
  assign n32772 = n32771 ^ n8290 ^ 1'b0 ;
  assign n32773 = n820 & n10509 ;
  assign n32774 = n5726 ^ n3314 ^ x178 ;
  assign n32775 = n17247 | n32774 ;
  assign n32776 = n23893 | n32775 ;
  assign n32777 = ~n3561 & n8729 ;
  assign n32778 = ~n32776 & n32777 ;
  assign n32779 = n32773 & ~n32778 ;
  assign n32780 = ~n32772 & n32779 ;
  assign n32781 = ~n4063 & n30742 ;
  assign n32782 = ~n8827 & n16747 ;
  assign n32783 = ~n444 & n32782 ;
  assign n32784 = n9783 & n15886 ;
  assign n32785 = n32784 ^ n744 ^ 1'b0 ;
  assign n32786 = n32783 | n32785 ;
  assign n32787 = n20617 ^ n6355 ^ 1'b0 ;
  assign n32788 = n1390 & ~n9105 ;
  assign n32789 = ~n343 & n32788 ;
  assign n32790 = n17192 & ~n30639 ;
  assign n32791 = n32789 & n32790 ;
  assign n32792 = n7755 ^ n2315 ^ 1'b0 ;
  assign n32793 = n32792 ^ n27710 ^ 1'b0 ;
  assign n32794 = ~n25252 & n32793 ;
  assign n32795 = n3359 & n10873 ;
  assign n32796 = ~n13291 & n32795 ;
  assign n32797 = n7953 & ~n16593 ;
  assign n32798 = ~n12237 & n24113 ;
  assign n32799 = ~n1693 & n22180 ;
  assign n32800 = n32799 ^ n30044 ^ 1'b0 ;
  assign n32801 = n25703 ^ n24635 ^ 1'b0 ;
  assign n32802 = ~n3678 & n32801 ;
  assign n32805 = n3669 & ~n4149 ;
  assign n32804 = n14331 & n27714 ;
  assign n32806 = n32805 ^ n32804 ^ 1'b0 ;
  assign n32803 = n13115 & n18665 ;
  assign n32807 = n32806 ^ n32803 ^ 1'b0 ;
  assign n32808 = n14157 ^ n11063 ^ 1'b0 ;
  assign n32809 = n3047 ^ n1337 ^ 1'b0 ;
  assign n32810 = n32808 & ~n32809 ;
  assign n32811 = n6311 ^ x86 ^ 1'b0 ;
  assign n32812 = n22104 & ~n32811 ;
  assign n32813 = n21445 ^ x158 ^ 1'b0 ;
  assign n32814 = n32812 & n32813 ;
  assign n32815 = n32814 ^ n1792 ^ 1'b0 ;
  assign n32816 = ~n18219 & n32815 ;
  assign n32817 = n6279 & n32816 ;
  assign n32818 = n9904 & ~n26383 ;
  assign n32819 = n956 | n15263 ;
  assign n32820 = n32819 ^ n12690 ^ 1'b0 ;
  assign n32821 = n29103 ^ n10281 ^ 1'b0 ;
  assign n32822 = n5073 & ~n32821 ;
  assign n32823 = n31955 ^ n30054 ^ 1'b0 ;
  assign n32824 = n3870 | n24351 ;
  assign n32825 = n32824 ^ n7531 ^ 1'b0 ;
  assign n32826 = n21825 & n32825 ;
  assign n32827 = ( n841 & n4925 ) | ( n841 & n11920 ) | ( n4925 & n11920 ) ;
  assign n32828 = n6343 & n32827 ;
  assign n32829 = n30865 ^ n3303 ^ 1'b0 ;
  assign n32830 = n25196 ^ n3216 ^ 1'b0 ;
  assign n32831 = n7809 ^ n5473 ^ 1'b0 ;
  assign n32832 = n9176 | n32831 ;
  assign n32833 = ~n7527 & n10813 ;
  assign n32834 = n32832 & n32833 ;
  assign n32835 = ~n17150 & n23831 ;
  assign n32836 = ~n4879 & n20784 ;
  assign n32837 = n2887 & n32836 ;
  assign n32838 = n20503 ^ n15780 ^ 1'b0 ;
  assign n32839 = ~n2718 & n31053 ;
  assign n32840 = ~n26621 & n32839 ;
  assign n32841 = ~n4261 & n9592 ;
  assign n32842 = n7440 & ~n32841 ;
  assign n32843 = n27658 & n28822 ;
  assign n32844 = n16967 ^ n11714 ^ 1'b0 ;
  assign n32845 = n4943 & ~n32754 ;
  assign n32846 = n32845 ^ n16377 ^ 1'b0 ;
  assign n32847 = n5943 | n8832 ;
  assign n32848 = n22811 & n32847 ;
  assign n32849 = ~n29662 & n32848 ;
  assign n32850 = n934 & n14610 ;
  assign n32851 = n32055 ^ n17199 ^ 1'b0 ;
  assign n32852 = n13585 | n32851 ;
  assign n32853 = n8341 | n12427 ;
  assign n32854 = n32853 ^ n9137 ^ 1'b0 ;
  assign n32855 = n32854 ^ n3362 ^ 1'b0 ;
  assign n32856 = ~n5004 & n16694 ;
  assign n32857 = ~n24009 & n32856 ;
  assign n32858 = ~n21786 & n32857 ;
  assign n32859 = n26825 ^ n8665 ^ 1'b0 ;
  assign n32860 = n13049 & n32859 ;
  assign n32861 = n651 & ~n2752 ;
  assign n32862 = ~n3779 & n30170 ;
  assign n32863 = ~n15025 & n32862 ;
  assign n32864 = n15993 & ~n32863 ;
  assign n32865 = n12835 & n32864 ;
  assign n32866 = ~n13725 & n29570 ;
  assign n32867 = n5977 | n32866 ;
  assign n32868 = n4433 | n32867 ;
  assign n32869 = ~n3731 & n12789 ;
  assign n32870 = ~n18389 & n20469 ;
  assign n32871 = ~n24774 & n32870 ;
  assign n32872 = ~x23 & n4385 ;
  assign n32873 = ~n2457 & n32872 ;
  assign n32874 = n20488 & n32873 ;
  assign n32875 = n7888 | n9380 ;
  assign n32876 = n29114 & ~n32875 ;
  assign n32877 = n32876 ^ n30388 ^ 1'b0 ;
  assign n32878 = ~n677 & n11268 ;
  assign n32879 = n32878 ^ n19220 ^ 1'b0 ;
  assign n32880 = n20787 & n29623 ;
  assign n32881 = n3280 & ~n32880 ;
  assign n32882 = n4201 ^ n824 ^ 1'b0 ;
  assign n32883 = n32882 ^ n20398 ^ 1'b0 ;
  assign n32884 = ~n6147 & n24820 ;
  assign n32885 = n6250 & n6809 ;
  assign n32890 = n5896 | n15665 ;
  assign n32891 = n5896 & ~n32890 ;
  assign n32886 = n4875 & ~n4899 ;
  assign n32887 = n4899 & n32886 ;
  assign n32888 = ( n12671 & ~n18723 ) | ( n12671 & n32887 ) | ( ~n18723 & n32887 ) ;
  assign n32889 = n11210 | n32888 ;
  assign n32892 = n32891 ^ n32889 ^ 1'b0 ;
  assign n32893 = n11669 & ~n28011 ;
  assign n32894 = n32893 ^ n996 ^ 1'b0 ;
  assign n32895 = n32894 ^ n13671 ^ 1'b0 ;
  assign n32896 = ( n3558 & n21404 ) | ( n3558 & n32222 ) | ( n21404 & n32222 ) ;
  assign n32897 = ~n26927 & n32637 ;
  assign n32898 = n32897 ^ n10731 ^ 1'b0 ;
  assign n32899 = n10646 | n11119 ;
  assign n32900 = n26083 & n32899 ;
  assign n32901 = n12738 | n18302 ;
  assign n32902 = n32901 ^ n9886 ^ n9335 ;
  assign n32903 = x152 & n32902 ;
  assign n32904 = n32903 ^ n1372 ^ 1'b0 ;
  assign n32905 = ~x236 & n1978 ;
  assign n32906 = n9331 & n18627 ;
  assign n32907 = n32906 ^ n10284 ^ n854 ;
  assign n32908 = n12535 & ~n20087 ;
  assign n32909 = n20277 ^ n2667 ^ 1'b0 ;
  assign n32910 = n21564 & ~n32909 ;
  assign n32911 = n19792 & n25701 ;
  assign n32912 = n28381 & n32911 ;
  assign n32913 = n305 | n15418 ;
  assign n32914 = n31152 ^ n26625 ^ 1'b0 ;
  assign n32915 = n22631 & ~n32914 ;
  assign n32916 = ~n20325 & n27975 ;
  assign n32917 = x84 | n2476 ;
  assign n32918 = n2476 & ~n32917 ;
  assign n32923 = ~n2435 & n3444 ;
  assign n32924 = n2435 & n32923 ;
  assign n32925 = n17656 | n32924 ;
  assign n32926 = n32924 & ~n32925 ;
  assign n32920 = ~n3678 & n3945 ;
  assign n32921 = n32920 ^ n1400 ^ 1'b0 ;
  assign n32919 = n10095 ^ n9458 ^ 1'b0 ;
  assign n32922 = n32921 ^ n32919 ^ n10929 ;
  assign n32927 = n32926 ^ n32922 ^ 1'b0 ;
  assign n32928 = ~n32918 & n32927 ;
  assign n32929 = ~n3645 & n5774 ;
  assign n32930 = n4643 & ~n6391 ;
  assign n32931 = ~n454 & n32930 ;
  assign n32932 = ~n13868 & n19791 ;
  assign n32933 = ~n2217 & n22430 ;
  assign n32934 = ( ~n339 & n534 ) | ( ~n339 & n32933 ) | ( n534 & n32933 ) ;
  assign n32935 = n32934 ^ n31242 ^ 1'b0 ;
  assign n32937 = n7609 ^ n3503 ^ 1'b0 ;
  assign n32938 = ~n14071 & n32937 ;
  assign n32939 = x25 & ~n23489 ;
  assign n32940 = ~n32938 & n32939 ;
  assign n32936 = n6659 & ~n7700 ;
  assign n32941 = n32940 ^ n32936 ^ 1'b0 ;
  assign n32942 = n4860 & ~n21146 ;
  assign n32943 = n32942 ^ n20412 ^ 1'b0 ;
  assign n32944 = n32943 ^ n1492 ^ 1'b0 ;
  assign n32945 = n24434 ^ n18736 ^ 1'b0 ;
  assign n32946 = ~n26146 & n32945 ;
  assign n32947 = n296 | n2124 ;
  assign n32948 = n4298 | n6504 ;
  assign n32949 = n9720 & ~n32948 ;
  assign n32950 = n13040 & ~n32949 ;
  assign n32951 = n4209 ^ n1368 ^ 1'b0 ;
  assign n32954 = ~n3625 & n15106 ;
  assign n32952 = n4237 | n5869 ;
  assign n32953 = n32952 ^ n23026 ^ 1'b0 ;
  assign n32955 = n32954 ^ n32953 ^ 1'b0 ;
  assign n32956 = n5824 & n32955 ;
  assign n32957 = n12170 & n17251 ;
  assign n32958 = n1847 | n24612 ;
  assign n32961 = n1410 & n11241 ;
  assign n32959 = n14020 ^ n1814 ^ 1'b0 ;
  assign n32960 = n381 | n32959 ;
  assign n32962 = n32961 ^ n32960 ^ 1'b0 ;
  assign n32963 = n13750 ^ n5192 ^ 1'b0 ;
  assign n32964 = n32962 | n32963 ;
  assign n32965 = n29473 ^ n3503 ^ 1'b0 ;
  assign n32966 = n21063 & ~n31330 ;
  assign n32967 = n28490 & n32966 ;
  assign n32968 = n528 | n32967 ;
  assign n32969 = ~n21929 & n32968 ;
  assign n32970 = n7386 ^ n7016 ^ 1'b0 ;
  assign n32971 = n1920 ^ x47 ^ 1'b0 ;
  assign n32972 = n607 & n32971 ;
  assign n32973 = ~n32970 & n32972 ;
  assign n32974 = ~n21411 & n29204 ;
  assign n32975 = n11645 & ~n26335 ;
  assign n32976 = n9212 | n21581 ;
  assign n32977 = n9663 ^ x130 ^ 1'b0 ;
  assign n32978 = n23162 & ~n32977 ;
  assign n32979 = n32978 ^ n14376 ^ 1'b0 ;
  assign n32986 = n28551 ^ n10467 ^ 1'b0 ;
  assign n32983 = n12527 ^ n6394 ^ 1'b0 ;
  assign n32984 = n637 & n4825 ;
  assign n32985 = n32983 & n32984 ;
  assign n32987 = n32986 ^ n32985 ^ 1'b0 ;
  assign n32980 = ~n12745 & n17391 ;
  assign n32981 = n9389 & n32980 ;
  assign n32982 = n15427 | n32981 ;
  assign n32988 = n32987 ^ n32982 ^ 1'b0 ;
  assign n32989 = n12666 ^ n8663 ^ 1'b0 ;
  assign n32990 = n12402 | n32989 ;
  assign n32991 = n32990 ^ n2210 ^ 1'b0 ;
  assign n32992 = ~n7185 & n15998 ;
  assign n32993 = n32992 ^ n8637 ^ 1'b0 ;
  assign n32994 = n10492 & n32993 ;
  assign n32995 = n32994 ^ n19717 ^ 1'b0 ;
  assign n32996 = n5412 | n17176 ;
  assign n32997 = n32996 ^ n11589 ^ 1'b0 ;
  assign n32998 = n4988 & ~n7049 ;
  assign n32999 = n6097 & ~n32998 ;
  assign n33000 = ~n32997 & n32999 ;
  assign n33001 = n10915 | n16198 ;
  assign n33002 = n9620 & ~n20707 ;
  assign n33003 = ~n24628 & n33002 ;
  assign n33004 = ~n6646 & n12861 ;
  assign n33005 = ~n21998 & n33004 ;
  assign n33006 = n21387 | n33005 ;
  assign n33007 = n11241 & ~n22567 ;
  assign n33008 = n4755 & ~n12030 ;
  assign n33009 = n33008 ^ n4456 ^ 1'b0 ;
  assign n33010 = ~n2711 & n6590 ;
  assign n33011 = n17542 & n33010 ;
  assign n33012 = n1701 | n3000 ;
  assign n33013 = n25015 ^ n22783 ^ 1'b0 ;
  assign n33014 = n33012 & n33013 ;
  assign n33018 = n2100 ^ n659 ^ 1'b0 ;
  assign n33015 = n2146 | n13647 ;
  assign n33016 = n33015 ^ n19130 ^ n13945 ;
  assign n33017 = n10498 & n33016 ;
  assign n33019 = n33018 ^ n33017 ^ 1'b0 ;
  assign n33020 = n3331 ^ n2180 ^ 1'b0 ;
  assign n33021 = n1630 ^ n1320 ^ 1'b0 ;
  assign n33022 = ~n715 & n33021 ;
  assign n33023 = n33022 ^ n7131 ^ 1'b0 ;
  assign n33024 = n4251 & ~n33023 ;
  assign n33025 = n3549 & n25413 ;
  assign n33026 = n1302 & n33025 ;
  assign n33027 = ~n33024 & n33026 ;
  assign n33028 = ~n18243 & n31289 ;
  assign n33029 = n15178 | n24363 ;
  assign n33030 = n33029 ^ n3895 ^ 1'b0 ;
  assign n33031 = ~n2072 & n5701 ;
  assign n33032 = n33031 ^ n3625 ^ 1'b0 ;
  assign n33033 = n18095 ^ n13225 ^ 1'b0 ;
  assign n33034 = n4412 ^ n532 ^ 1'b0 ;
  assign n33035 = n5350 & n33034 ;
  assign n33036 = ( n6061 & n9178 ) | ( n6061 & ~n19800 ) | ( n9178 & ~n19800 ) ;
  assign n33037 = n9135 | n33036 ;
  assign n33038 = ~n10629 & n19309 ;
  assign n33039 = ~n7206 & n26260 ;
  assign n33040 = n1897 ^ n1725 ^ 1'b0 ;
  assign n33041 = n9178 & n33040 ;
  assign n33042 = n33041 ^ n13543 ^ n9344 ;
  assign n33043 = n1507 | n4575 ;
  assign n33044 = n13918 | n33043 ;
  assign n33045 = n33044 ^ n29401 ^ 1'b0 ;
  assign n33046 = n33045 ^ n26004 ^ n18437 ;
  assign n33047 = ~n3694 & n23534 ;
  assign n33048 = ~n26366 & n33047 ;
  assign n33049 = n10042 ^ n5897 ^ 1'b0 ;
  assign n33050 = n33048 | n33049 ;
  assign n33051 = n4304 ^ n3854 ^ 1'b0 ;
  assign n33052 = n10979 & ~n33051 ;
  assign n33053 = n2296 & n33052 ;
  assign n33054 = n1769 | n33028 ;
  assign n33055 = n15825 & ~n33054 ;
  assign n33056 = n1096 & n1572 ;
  assign n33057 = n3272 | n12627 ;
  assign n33058 = x20 | n33057 ;
  assign n33059 = n33056 & ~n33058 ;
  assign n33060 = n29547 ^ n9946 ^ 1'b0 ;
  assign n33061 = n4138 & n6054 ;
  assign n33062 = n15394 & ~n33061 ;
  assign n33063 = n644 & n1402 ;
  assign n33064 = n4074 & ~n20418 ;
  assign n33065 = n33064 ^ n13513 ^ 1'b0 ;
  assign n33066 = n25772 ^ n3473 ^ 1'b0 ;
  assign n33067 = n5207 & ~n5369 ;
  assign n33068 = n8008 ^ n643 ^ 1'b0 ;
  assign n33069 = n7232 | n14580 ;
  assign n33070 = n4203 & ~n23327 ;
  assign n33071 = n9724 | n33070 ;
  assign n33072 = n33071 ^ n545 ^ 1'b0 ;
  assign n33073 = n9108 & n21096 ;
  assign n33074 = n3748 & n32351 ;
  assign n33075 = ( n8277 & ~n28297 ) | ( n8277 & n29856 ) | ( ~n28297 & n29856 ) ;
  assign n33076 = n10185 ^ x25 ^ 1'b0 ;
  assign n33077 = n5768 | n18462 ;
  assign n33078 = n33077 ^ n12360 ^ 1'b0 ;
  assign n33079 = n7924 & ~n9231 ;
  assign n33080 = n5275 & ~n19704 ;
  assign n33081 = n33080 ^ n8801 ^ 1'b0 ;
  assign n33082 = n13756 ^ n9317 ^ 1'b0 ;
  assign n33083 = n8956 | n16246 ;
  assign n33084 = n10500 & ~n33083 ;
  assign n33085 = n33084 ^ n13746 ^ 1'b0 ;
  assign n33086 = n18660 | n22667 ;
  assign n33087 = n5564 & ~n28380 ;
  assign n33088 = n5593 ^ x213 ^ 1'b0 ;
  assign n33089 = n14786 ^ n10432 ^ 1'b0 ;
  assign n33090 = n31785 & ~n33089 ;
  assign n33091 = ~n13503 & n19213 ;
  assign n33092 = ~n10214 & n33091 ;
  assign n33093 = n626 & ~n8068 ;
  assign n33094 = n33093 ^ n1845 ^ 1'b0 ;
  assign n33095 = n23898 & n33094 ;
  assign n33096 = n6372 & ~n7398 ;
  assign n33097 = n33096 ^ n2035 ^ 1'b0 ;
  assign n33098 = n33097 ^ n5163 ^ 1'b0 ;
  assign n33099 = n3756 | n33098 ;
  assign n33100 = n5012 | n32681 ;
  assign n33101 = n21682 ^ n9269 ^ 1'b0 ;
  assign n33102 = n14591 ^ n9561 ^ n5160 ;
  assign n33103 = n33101 & ~n33102 ;
  assign n33104 = ~n788 & n16472 ;
  assign n33105 = n3163 & ~n17290 ;
  assign n33106 = n13926 & n33105 ;
  assign n33107 = n4625 | n11011 ;
  assign n33108 = n5176 & n14643 ;
  assign n33109 = n33108 ^ n11533 ^ 1'b0 ;
  assign n33110 = n20220 & ~n33109 ;
  assign n33111 = ~n33107 & n33110 ;
  assign n33112 = n26136 & ~n33111 ;
  assign n33113 = n1693 & n33112 ;
  assign n33114 = x95 | n24607 ;
  assign n33115 = x7 | n33114 ;
  assign n33116 = n33115 ^ n9808 ^ 1'b0 ;
  assign n33117 = n33116 ^ n9916 ^ 1'b0 ;
  assign n33118 = n5824 | n28376 ;
  assign n33119 = n11713 & ~n33118 ;
  assign n33120 = n33119 ^ n1451 ^ 1'b0 ;
  assign n33121 = n2465 & ~n33120 ;
  assign n33123 = n8691 & ~n26927 ;
  assign n33122 = n9939 & ~n13978 ;
  assign n33124 = n33123 ^ n33122 ^ 1'b0 ;
  assign n33125 = n29806 & ~n33124 ;
  assign n33126 = n7749 & n16829 ;
  assign n33127 = n9156 ^ n4258 ^ 1'b0 ;
  assign n33128 = n33126 & ~n33127 ;
  assign n33129 = ~n9279 & n31261 ;
  assign n33130 = n4678 | n10935 ;
  assign n33131 = n2225 & ~n33130 ;
  assign n33132 = n6649 & n9590 ;
  assign n33133 = n33131 & n33132 ;
  assign n33134 = ~n3045 & n29745 ;
  assign n33135 = n2910 & ~n20898 ;
  assign n33136 = n9060 & ~n31060 ;
  assign n33137 = n23538 & n33136 ;
  assign n33138 = n13734 | n16843 ;
  assign n33139 = n4467 & ~n7624 ;
  assign n33140 = ~n33138 & n33139 ;
  assign n33141 = ~n2892 & n33140 ;
  assign n33142 = n12744 ^ n11013 ^ n6484 ;
  assign n33143 = n1102 | n1295 ;
  assign n33144 = n29742 ^ n9741 ^ 1'b0 ;
  assign n33145 = n33144 ^ n18750 ^ 1'b0 ;
  assign n33146 = n24396 ^ n18767 ^ n10143 ;
  assign n33147 = n2652 & n33146 ;
  assign n33148 = n8811 & ~n18128 ;
  assign n33149 = n33148 ^ n20144 ^ 1'b0 ;
  assign n33150 = n2122 | n27718 ;
  assign n33151 = n33150 ^ n21293 ^ 1'b0 ;
  assign n33152 = n33151 ^ n5500 ^ 1'b0 ;
  assign n33153 = n17552 ^ n12387 ^ 1'b0 ;
  assign n33154 = n27533 ^ n24301 ^ 1'b0 ;
  assign n33155 = ~n9985 & n33154 ;
  assign n33156 = n33155 ^ n552 ^ 1'b0 ;
  assign n33157 = ~n13560 & n14610 ;
  assign n33158 = ~n33156 & n33157 ;
  assign n33159 = n19118 ^ n2766 ^ n924 ;
  assign n33163 = n21544 ^ n14629 ^ 1'b0 ;
  assign n33164 = n27729 & ~n33163 ;
  assign n33160 = n9339 & n12675 ;
  assign n33161 = n14807 & n33160 ;
  assign n33162 = n4417 & ~n33161 ;
  assign n33165 = n33164 ^ n33162 ^ 1'b0 ;
  assign n33166 = x170 & n3629 ;
  assign n33167 = n2977 ^ n1210 ^ 1'b0 ;
  assign n33168 = n33167 ^ n6742 ^ 1'b0 ;
  assign n33169 = n33166 & n33168 ;
  assign n33170 = n27427 ^ n25922 ^ 1'b0 ;
  assign n33171 = n31928 & ~n33170 ;
  assign n33172 = n1613 ^ n452 ^ 1'b0 ;
  assign n33173 = n9185 & n33172 ;
  assign n33174 = n3045 & n10760 ;
  assign n33175 = n27530 & n33174 ;
  assign n33176 = n8631 ^ n1435 ^ 1'b0 ;
  assign n33177 = ~n33175 & n33176 ;
  assign n33178 = n8720 ^ n1588 ^ 1'b0 ;
  assign n33179 = n15555 & ~n33178 ;
  assign n33180 = n13734 ^ n3878 ^ 1'b0 ;
  assign n33181 = n33179 & ~n33180 ;
  assign n33182 = n25837 | n33175 ;
  assign n33183 = n23430 & ~n33182 ;
  assign n33184 = n14654 & n25926 ;
  assign n33185 = n16174 & n33184 ;
  assign n33186 = n15904 | n33185 ;
  assign n33189 = n10333 ^ n2793 ^ 1'b0 ;
  assign n33190 = n2569 & ~n33189 ;
  assign n33187 = n9933 & ~n18015 ;
  assign n33188 = n8082 & n33187 ;
  assign n33191 = n33190 ^ n33188 ^ 1'b0 ;
  assign n33192 = n7434 & n7937 ;
  assign n33193 = ~n14595 & n20873 ;
  assign n33194 = ~n33192 & n33193 ;
  assign n33195 = n17812 & ~n33194 ;
  assign n33196 = n29827 ^ n8453 ^ 1'b0 ;
  assign n33197 = n5225 & ~n33196 ;
  assign n33198 = n9832 & ~n33197 ;
  assign n33199 = n7410 | n32542 ;
  assign n33200 = n785 & ~n33199 ;
  assign n33201 = n33200 ^ n313 ^ 1'b0 ;
  assign n33202 = n5506 | n33201 ;
  assign n33203 = n3566 | n25239 ;
  assign n33204 = n465 | n33203 ;
  assign n33205 = ~n4055 & n31170 ;
  assign n33206 = n33205 ^ n13647 ^ 1'b0 ;
  assign n33207 = n618 & n33206 ;
  assign n33208 = n11128 | n23779 ;
  assign n33209 = n3574 & ~n33208 ;
  assign n33210 = n1806 | n3307 ;
  assign n33211 = n12825 & n30068 ;
  assign n33213 = n6078 | n17258 ;
  assign n33214 = n33213 ^ n26766 ^ 1'b0 ;
  assign n33212 = ~n9811 & n12314 ;
  assign n33215 = n33214 ^ n33212 ^ 1'b0 ;
  assign n33216 = n20073 & ~n24662 ;
  assign n33217 = ~n20905 & n33216 ;
  assign n33218 = n387 & n17952 ;
  assign n33219 = n33218 ^ n1738 ^ 1'b0 ;
  assign n33220 = n19236 ^ n12023 ^ 1'b0 ;
  assign n33221 = n10808 ^ n2668 ^ 1'b0 ;
  assign n33222 = n957 & n18092 ;
  assign n33223 = n33222 ^ n3888 ^ 1'b0 ;
  assign n33226 = n17073 ^ n4684 ^ 1'b0 ;
  assign n33224 = n8636 | n14354 ;
  assign n33225 = x123 | n33224 ;
  assign n33227 = n33226 ^ n33225 ^ 1'b0 ;
  assign n33228 = n9657 | n21019 ;
  assign n33229 = n17358 ^ n11157 ^ 1'b0 ;
  assign n33230 = n33228 | n33229 ;
  assign n33231 = n18751 ^ n4322 ^ 1'b0 ;
  assign n33232 = ~n33230 & n33231 ;
  assign n33233 = n3451 & ~n12273 ;
  assign n33234 = n22820 ^ n4777 ^ 1'b0 ;
  assign n33235 = n18454 | n33234 ;
  assign n33236 = n6456 ^ x140 ^ 1'b0 ;
  assign n33237 = n713 | n10747 ;
  assign n33238 = n16789 | n33237 ;
  assign n33239 = n11663 | n18134 ;
  assign n33240 = n5676 | n33239 ;
  assign n33241 = n33238 | n33240 ;
  assign n33242 = n10398 ^ n1815 ^ 1'b0 ;
  assign n33243 = n17350 | n33242 ;
  assign n33244 = n3163 & ~n28280 ;
  assign n33245 = x87 & n22292 ;
  assign n33246 = ~n516 & n2225 ;
  assign n33247 = n3314 | n6792 ;
  assign n33248 = n14992 | n33247 ;
  assign n33249 = n5808 | n33248 ;
  assign n33250 = n26640 & ~n33249 ;
  assign n33251 = n8275 ^ n6464 ^ 1'b0 ;
  assign n33252 = ~n3899 & n14560 ;
  assign n33253 = n16132 ^ n7388 ^ 1'b0 ;
  assign n33254 = n497 | n4358 ;
  assign n33255 = n33254 ^ n12197 ^ 1'b0 ;
  assign n33256 = n33255 ^ n29551 ^ 1'b0 ;
  assign n33257 = n16432 ^ n8843 ^ 1'b0 ;
  assign n33258 = ~n7323 & n31514 ;
  assign n33259 = n28223 & n33258 ;
  assign n33260 = n1455 | n33259 ;
  assign n33261 = n33260 ^ n16007 ^ 1'b0 ;
  assign n33262 = ~n28129 & n33261 ;
  assign n33263 = n4140 & ~n8730 ;
  assign n33264 = n33263 ^ n9961 ^ 1'b0 ;
  assign n33265 = ~n1302 & n33264 ;
  assign n33266 = ( n1381 & n2744 ) | ( n1381 & n3281 ) | ( n2744 & n3281 ) ;
  assign n33267 = n2970 & n33266 ;
  assign n33268 = ~n8902 & n13875 ;
  assign n33269 = ~n33267 & n33268 ;
  assign n33270 = n25214 ^ n15123 ^ 1'b0 ;
  assign n33271 = n26488 & ~n29792 ;
  assign n33272 = n15719 | n33194 ;
  assign n33273 = n298 & ~n11802 ;
  assign n33274 = ~n3349 & n33273 ;
  assign n33275 = n33264 ^ n19710 ^ 1'b0 ;
  assign n33276 = n6587 ^ n3802 ^ 1'b0 ;
  assign n33277 = ~n33275 & n33276 ;
  assign n33278 = n12981 & n33277 ;
  assign n33279 = ( n607 & n2818 ) | ( n607 & ~n33278 ) | ( n2818 & ~n33278 ) ;
  assign n33280 = n18380 & ~n29498 ;
  assign n33281 = n31647 ^ n18857 ^ n13776 ;
  assign n33282 = n16962 & ~n33281 ;
  assign n33283 = n33282 ^ n21255 ^ 1'b0 ;
  assign n33284 = n4029 & ~n19420 ;
  assign n33285 = n33284 ^ n2904 ^ 1'b0 ;
  assign n33286 = n5879 & ~n20808 ;
  assign n33287 = ~n12140 & n21076 ;
  assign n33288 = ~n33286 & n33287 ;
  assign n33289 = ( n10330 & n18164 ) | ( n10330 & n33288 ) | ( n18164 & n33288 ) ;
  assign n33290 = n22663 ^ n2145 ^ 1'b0 ;
  assign n33291 = ~n1843 & n23353 ;
  assign n33292 = n23256 & n33291 ;
  assign n33293 = n9371 ^ n1675 ^ 1'b0 ;
  assign n33294 = n16505 ^ n5328 ^ 1'b0 ;
  assign n33295 = n1729 | n3442 ;
  assign n33297 = x11 & ~n5980 ;
  assign n33298 = ~n21397 & n33297 ;
  assign n33296 = n21340 ^ n11040 ^ 1'b0 ;
  assign n33299 = n33298 ^ n33296 ^ n32622 ;
  assign n33300 = n29860 ^ n3881 ^ 1'b0 ;
  assign n33301 = n1131 & n33300 ;
  assign n33302 = n33301 ^ n13256 ^ 1'b0 ;
  assign n33303 = n22323 ^ n14771 ^ 1'b0 ;
  assign n33304 = n17214 & ~n33303 ;
  assign n33305 = n21811 & ~n28286 ;
  assign n33306 = n33305 ^ n31253 ^ 1'b0 ;
  assign n33307 = ~n1314 & n12926 ;
  assign n33308 = n33307 ^ n2916 ^ 1'b0 ;
  assign n33309 = n28721 ^ n12436 ^ 1'b0 ;
  assign n33310 = n33308 & ~n33309 ;
  assign n33311 = n26622 ^ n17225 ^ 1'b0 ;
  assign n33312 = ~n9475 & n33311 ;
  assign n33313 = n33312 ^ n9251 ^ 1'b0 ;
  assign n33314 = n12443 & ~n23886 ;
  assign n33315 = n1081 | n33314 ;
  assign n33316 = n27967 ^ n7296 ^ 1'b0 ;
  assign n33317 = ~n9589 & n33316 ;
  assign n33318 = n25470 ^ n8651 ^ 1'b0 ;
  assign n33319 = n4021 | n33318 ;
  assign n33320 = n9278 | n21566 ;
  assign n33321 = n10090 & ~n33320 ;
  assign n33322 = ( n6684 & n10130 ) | ( n6684 & ~n10398 ) | ( n10130 & ~n10398 ) ;
  assign n33323 = n7181 | n30713 ;
  assign n33326 = n9956 ^ n5875 ^ 1'b0 ;
  assign n33324 = n1205 | n21398 ;
  assign n33325 = n20359 & ~n33324 ;
  assign n33327 = n33326 ^ n33325 ^ 1'b0 ;
  assign n33328 = ~n5173 & n9589 ;
  assign n33329 = n11226 & n31236 ;
  assign n33330 = n33329 ^ n6756 ^ 1'b0 ;
  assign n33331 = n6020 & n9022 ;
  assign n33332 = n3009 ^ n1444 ^ 1'b0 ;
  assign n33333 = n25443 ^ n12745 ^ 1'b0 ;
  assign n33334 = n9057 ^ n1028 ^ 1'b0 ;
  assign n33335 = n33333 & ~n33334 ;
  assign n33336 = x3 & n33335 ;
  assign n33337 = n18162 ^ n17540 ^ n12172 ;
  assign n33338 = n33337 ^ n2146 ^ 1'b0 ;
  assign n33339 = n8597 & n24414 ;
  assign n33340 = n3823 | n13420 ;
  assign n33341 = ( n2293 & ~n11052 ) | ( n2293 & n12767 ) | ( ~n11052 & n12767 ) ;
  assign n33342 = n26775 & n31796 ;
  assign n33343 = ~n26775 & n33342 ;
  assign n33344 = n4758 ^ n3026 ^ 1'b0 ;
  assign n33345 = n12516 & ~n33344 ;
  assign n33346 = ~n18059 & n33345 ;
  assign n33347 = n10422 ^ n3367 ^ 1'b0 ;
  assign n33348 = ~n7984 & n13996 ;
  assign n33349 = n6724 & n33348 ;
  assign n33350 = n25054 & ~n33349 ;
  assign n33351 = n2571 & n33350 ;
  assign n33352 = n3090 ^ n1648 ^ 1'b0 ;
  assign n33353 = ( n15705 & n25505 ) | ( n15705 & n33352 ) | ( n25505 & n33352 ) ;
  assign n33354 = n33353 ^ n23873 ^ 1'b0 ;
  assign n33355 = n7869 | n13621 ;
  assign n33356 = n11987 & ~n26368 ;
  assign n33357 = n33355 & n33356 ;
  assign n33358 = ~n6176 & n12783 ;
  assign n33359 = n31671 | n33358 ;
  assign n33360 = n1651 & ~n8692 ;
  assign n33361 = n30004 ^ n18311 ^ 1'b0 ;
  assign n33362 = n33360 & n33361 ;
  assign n33363 = x86 | n15065 ;
  assign n33364 = n12948 | n28959 ;
  assign n33365 = n13511 | n32074 ;
  assign n33366 = ~n11249 & n33365 ;
  assign n33367 = ~n8419 & n20211 ;
  assign n33368 = ~n1369 & n1633 ;
  assign n33369 = n2760 & n11338 ;
  assign n33370 = n33369 ^ n5136 ^ 1'b0 ;
  assign n33371 = n33368 & ~n33370 ;
  assign n33372 = n18213 ^ n6308 ^ 1'b0 ;
  assign n33373 = n4382 ^ n3132 ^ 1'b0 ;
  assign n33374 = n6578 & n33373 ;
  assign n33375 = n2991 & ~n33374 ;
  assign n33376 = n12813 | n15463 ;
  assign n33377 = n21839 | n33376 ;
  assign n33378 = n33192 ^ n13515 ^ 1'b0 ;
  assign n33379 = ~n1379 & n6610 ;
  assign n33380 = n3328 | n3343 ;
  assign n33381 = n33379 & ~n33380 ;
  assign n33382 = n23657 ^ n7689 ^ 1'b0 ;
  assign n33383 = n6905 ^ n2082 ^ 1'b0 ;
  assign n33384 = n1139 & n33383 ;
  assign n33385 = ~n14425 & n33384 ;
  assign n33386 = n3071 | n14261 ;
  assign n33387 = n33385 & ~n33386 ;
  assign n33388 = n32482 ^ n5366 ^ 1'b0 ;
  assign n33389 = ~n1104 & n33388 ;
  assign n33390 = n15673 | n19635 ;
  assign n33391 = ~x28 & n7436 ;
  assign n33392 = n10130 ^ n7519 ^ 1'b0 ;
  assign n33393 = n8456 | n13696 ;
  assign n33394 = n33393 ^ n8223 ^ 1'b0 ;
  assign n33395 = n9220 ^ n7338 ^ 1'b0 ;
  assign n33396 = n27283 | n33395 ;
  assign n33397 = ~n5808 & n12610 ;
  assign n33398 = ~n11763 & n33397 ;
  assign n33399 = n805 | n16868 ;
  assign n33400 = n14442 ^ n4388 ^ 1'b0 ;
  assign n33401 = n1447 | n33400 ;
  assign n33402 = n1620 & n11474 ;
  assign n33403 = n11491 | n33402 ;
  assign n33404 = n33403 ^ n8182 ^ 1'b0 ;
  assign n33405 = n33404 ^ n8118 ^ 1'b0 ;
  assign n33406 = n33401 | n33405 ;
  assign n33407 = ~n13786 & n25470 ;
  assign n33408 = n33407 ^ n29746 ^ 1'b0 ;
  assign n33409 = n15737 & n24693 ;
  assign n33410 = n15561 ^ n666 ^ 1'b0 ;
  assign n33411 = n22872 ^ n22025 ^ 1'b0 ;
  assign n33412 = n452 & ~n33411 ;
  assign n33413 = ~n28680 & n28922 ;
  assign n33414 = n4764 & ~n7263 ;
  assign n33415 = n9794 & ~n18609 ;
  assign n33416 = n33415 ^ n7833 ^ 1'b0 ;
  assign n33417 = ( n307 & n1501 ) | ( n307 & ~n7997 ) | ( n1501 & ~n7997 ) ;
  assign n33423 = n1578 & ~n13118 ;
  assign n33418 = ~n4846 & n8684 ;
  assign n33419 = n11857 & n33418 ;
  assign n33420 = n33419 ^ n21938 ^ 1'b0 ;
  assign n33421 = n9881 | n33420 ;
  assign n33422 = n27440 & n33421 ;
  assign n33424 = n33423 ^ n33422 ^ 1'b0 ;
  assign n33425 = n11066 & ~n15346 ;
  assign n33426 = n2150 & ~n28991 ;
  assign n33427 = n15723 & n33426 ;
  assign n33428 = n4059 | n33427 ;
  assign n33429 = n33428 ^ n27510 ^ 1'b0 ;
  assign n33430 = n18318 | n33429 ;
  assign n33431 = n13389 | n18658 ;
  assign n33432 = n21995 | n33431 ;
  assign n33433 = n2078 ^ n661 ^ 1'b0 ;
  assign n33434 = n2909 | n5015 ;
  assign n33435 = n33434 ^ n14133 ^ 1'b0 ;
  assign n33436 = ~n12379 & n33435 ;
  assign n33437 = n33433 | n33436 ;
  assign n33438 = n2394 & n3381 ;
  assign n33439 = ( ~n2531 & n3633 ) | ( ~n2531 & n21956 ) | ( n3633 & n21956 ) ;
  assign n33440 = n13087 & n33439 ;
  assign n33441 = n15264 | n21012 ;
  assign n33442 = n33441 ^ n19340 ^ 1'b0 ;
  assign n33443 = ( ~x28 & n602 ) | ( ~x28 & n12595 ) | ( n602 & n12595 ) ;
  assign n33444 = n7244 | n33443 ;
  assign n33445 = n33444 ^ n1773 ^ 1'b0 ;
  assign n33446 = x65 & n2835 ;
  assign n33447 = n26100 | n27220 ;
  assign n33448 = n33447 ^ n31570 ^ n23622 ;
  assign n33449 = n3473 & n33448 ;
  assign n33450 = n16659 ^ n3946 ^ 1'b0 ;
  assign n33451 = n5727 | n33450 ;
  assign n33452 = n33451 ^ n6840 ^ 1'b0 ;
  assign n33453 = n7212 & ~n28204 ;
  assign n33454 = n11143 & n33453 ;
  assign n33455 = n3768 & n9220 ;
  assign n33456 = n20469 | n33455 ;
  assign n33457 = n29701 & n33456 ;
  assign n33458 = n4129 & ~n6222 ;
  assign n33459 = ~n2546 & n27840 ;
  assign n33460 = n19837 ^ n7252 ^ 1'b0 ;
  assign n33461 = n32712 ^ n4968 ^ 1'b0 ;
  assign n33462 = n5485 & ~n7411 ;
  assign n33463 = n33462 ^ n5107 ^ 1'b0 ;
  assign n33464 = n2263 & ~n33463 ;
  assign n33465 = n10241 | n19359 ;
  assign n33466 = n633 & ~n1344 ;
  assign n33467 = ~n7785 & n33466 ;
  assign n33468 = n32995 ^ n21611 ^ 1'b0 ;
  assign n33470 = n3903 ^ n3469 ^ 1'b0 ;
  assign n33471 = n14055 | n33470 ;
  assign n33472 = n26230 & ~n33471 ;
  assign n33469 = n18719 ^ n387 ^ 1'b0 ;
  assign n33473 = n33472 ^ n33469 ^ 1'b0 ;
  assign n33474 = n18933 ^ n9522 ^ 1'b0 ;
  assign n33475 = n25754 ^ n20012 ^ 1'b0 ;
  assign n33476 = n1736 & ~n33475 ;
  assign n33479 = n286 | n4957 ;
  assign n33480 = n3199 | n33479 ;
  assign n33477 = n13845 & ~n14065 ;
  assign n33478 = ~n10979 & n33477 ;
  assign n33481 = n33480 ^ n33478 ^ 1'b0 ;
  assign n33482 = n3948 | n9362 ;
  assign n33483 = n33482 ^ n23777 ^ 1'b0 ;
  assign n33484 = n4920 & ~n33483 ;
  assign n33485 = n32184 ^ n17694 ^ 1'b0 ;
  assign n33486 = n31850 ^ n11388 ^ 1'b0 ;
  assign n33487 = n21712 | n33486 ;
  assign n33488 = ~n3588 & n9444 ;
  assign n33489 = n10220 | n19508 ;
  assign n33490 = n33489 ^ n365 ^ 1'b0 ;
  assign n33491 = n17309 ^ n691 ^ 1'b0 ;
  assign n33492 = n4927 | n33491 ;
  assign n33493 = n9349 ^ n1256 ^ 1'b0 ;
  assign n33494 = n33492 | n33493 ;
  assign n33495 = n4586 & ~n16718 ;
  assign n33496 = n33495 ^ n4512 ^ 1'b0 ;
  assign n33497 = n2990 & ~n19707 ;
  assign n33498 = n33497 ^ n20364 ^ 1'b0 ;
  assign n33499 = n10787 ^ n2597 ^ 1'b0 ;
  assign n33500 = ~n5382 & n18134 ;
  assign n33501 = n6152 & n33500 ;
  assign n33502 = n19084 ^ n16206 ^ 1'b0 ;
  assign n33503 = n5715 & n21794 ;
  assign n33504 = ~n9994 & n33503 ;
  assign n33505 = n33504 ^ n896 ^ 1'b0 ;
  assign n33506 = n33502 & ~n33505 ;
  assign n33507 = ~n5398 & n6165 ;
  assign n33508 = n6357 & ~n16822 ;
  assign n33509 = n5094 & n7316 ;
  assign n33510 = n15306 & n25140 ;
  assign n33511 = n4368 | n4488 ;
  assign n33512 = n33511 ^ n6416 ^ 1'b0 ;
  assign n33513 = n5904 | n33512 ;
  assign n33514 = ( n5021 & n13519 ) | ( n5021 & n33513 ) | ( n13519 & n33513 ) ;
  assign n33515 = n33514 ^ n30137 ^ 1'b0 ;
  assign n33516 = n15233 & n17192 ;
  assign n33517 = n33516 ^ n1608 ^ 1'b0 ;
  assign n33518 = n28086 ^ n13711 ^ 1'b0 ;
  assign n33519 = n1765 & ~n33518 ;
  assign n33520 = ~n13052 & n15900 ;
  assign n33521 = n7694 & n33520 ;
  assign n33524 = n2237 & n8706 ;
  assign n33525 = ~n4680 & n33524 ;
  assign n33526 = n6033 | n33525 ;
  assign n33527 = n33526 ^ n21878 ^ 1'b0 ;
  assign n33522 = n28336 ^ n6884 ^ 1'b0 ;
  assign n33523 = ~n3709 & n33522 ;
  assign n33528 = n33527 ^ n33523 ^ 1'b0 ;
  assign n33529 = n31364 ^ n13952 ^ n10222 ;
  assign n33530 = n33529 ^ n8842 ^ 1'b0 ;
  assign n33531 = n33528 & ~n33530 ;
  assign n33532 = n756 & ~n16928 ;
  assign n33533 = n4549 & n10891 ;
  assign n33534 = ~n33532 & n33533 ;
  assign n33535 = n1560 & n3030 ;
  assign n33536 = n6343 & n33535 ;
  assign n33537 = n30824 ^ n16233 ^ 1'b0 ;
  assign n33538 = n27947 & ~n33537 ;
  assign n33539 = n4204 ^ x86 ^ 1'b0 ;
  assign n33540 = ~n8796 & n33539 ;
  assign n33541 = ~n3536 & n33540 ;
  assign n33542 = ~n8825 & n12631 ;
  assign n33543 = ~n3676 & n6670 ;
  assign n33544 = n23376 & n23893 ;
  assign n33545 = ~n1786 & n33544 ;
  assign n33546 = ( n9068 & n33543 ) | ( n9068 & ~n33545 ) | ( n33543 & ~n33545 ) ;
  assign n33547 = n28930 ^ n19597 ^ 1'b0 ;
  assign n33548 = n22402 ^ n10773 ^ 1'b0 ;
  assign n33549 = ~n11802 & n33548 ;
  assign n33550 = n33549 ^ n5496 ^ 1'b0 ;
  assign n33551 = n1435 | n29705 ;
  assign n33552 = n32250 & ~n33551 ;
  assign n33553 = n5457 & n10094 ;
  assign n33554 = n23722 & ~n32640 ;
  assign n33555 = n28994 ^ n6878 ^ n6487 ;
  assign n33556 = n10016 | n31159 ;
  assign n33557 = n7800 ^ n5125 ^ 1'b0 ;
  assign n33558 = n15757 ^ n15050 ^ 1'b0 ;
  assign n33559 = n24322 ^ x220 ^ 1'b0 ;
  assign n33561 = n13040 | n20563 ;
  assign n33560 = n15959 ^ n5504 ^ n3260 ;
  assign n33562 = n33561 ^ n33560 ^ 1'b0 ;
  assign n33563 = n21919 ^ n1589 ^ 1'b0 ;
  assign n33564 = n12046 & n14639 ;
  assign n33565 = ~n482 & n33564 ;
  assign n33566 = n5372 & n20156 ;
  assign n33567 = ~n11509 & n33566 ;
  assign n33568 = n33567 ^ n3181 ^ 1'b0 ;
  assign n33569 = n33565 & n33568 ;
  assign n33570 = n22189 | n30340 ;
  assign n33571 = n7171 & ~n33570 ;
  assign n33572 = ~n10744 & n18159 ;
  assign n33573 = n16777 ^ n10507 ^ 1'b0 ;
  assign n33574 = n7406 | n33573 ;
  assign n33575 = n8341 | n14520 ;
  assign n33576 = n1847 | n25062 ;
  assign n33577 = n22824 | n33576 ;
  assign n33578 = n20340 | n33577 ;
  assign n33579 = ~n1914 & n25960 ;
  assign n33580 = n12140 & n12889 ;
  assign n33581 = ~n8529 & n33580 ;
  assign n33582 = n5442 | n6446 ;
  assign n33583 = n33582 ^ n32276 ^ 1'b0 ;
  assign n33584 = n33581 & ~n33583 ;
  assign n33585 = n1268 & n9978 ;
  assign n33586 = n33585 ^ n805 ^ 1'b0 ;
  assign n33587 = n2435 & ~n3625 ;
  assign n33588 = n1779 & n33587 ;
  assign n33589 = ~n33586 & n33588 ;
  assign n33590 = n29794 & n33589 ;
  assign n33591 = n2097 & ~n7603 ;
  assign n33592 = n29626 & n33591 ;
  assign n33593 = ~n2547 & n27463 ;
  assign n33594 = n13616 ^ n7300 ^ 1'b0 ;
  assign n33595 = n10537 & ~n33594 ;
  assign n33596 = n5503 & n12148 ;
  assign n33597 = n8944 & n33596 ;
  assign n33598 = n7824 | n27638 ;
  assign n33599 = n4553 & n4849 ;
  assign n33600 = ( n6273 & n33598 ) | ( n6273 & ~n33599 ) | ( n33598 & ~n33599 ) ;
  assign n33601 = n4819 & ~n14352 ;
  assign n33602 = n2382 & n33601 ;
  assign n33603 = n33602 ^ n15123 ^ 1'b0 ;
  assign n33604 = n33600 | n33603 ;
  assign n33605 = n13418 ^ n5798 ^ 1'b0 ;
  assign n33606 = n33605 ^ n11628 ^ 1'b0 ;
  assign n33607 = n257 & n9113 ;
  assign n33608 = n33607 ^ n13956 ^ 1'b0 ;
  assign n33609 = n1762 & ~n27168 ;
  assign n33610 = n20938 ^ n12095 ^ 1'b0 ;
  assign n33611 = n9206 & n14974 ;
  assign n33612 = n33611 ^ n10228 ^ 1'b0 ;
  assign n33613 = ~n11427 & n25963 ;
  assign n33614 = ~n33612 & n33613 ;
  assign n33615 = n7642 & ~n17741 ;
  assign n33616 = n33615 ^ n3348 ^ 1'b0 ;
  assign n33617 = n11729 & ~n32023 ;
  assign n33618 = ~n30102 & n33617 ;
  assign n33619 = n5563 | n33618 ;
  assign n33620 = n33619 ^ n26672 ^ 1'b0 ;
  assign n33621 = n6863 ^ n4179 ^ 1'b0 ;
  assign n33622 = n2063 & n33621 ;
  assign n33623 = n33622 ^ n19254 ^ 1'b0 ;
  assign n33624 = n29204 ^ n25456 ^ 1'b0 ;
  assign n33625 = x43 & ~n33624 ;
  assign n33626 = n6106 & n24831 ;
  assign n33627 = n15497 ^ n6511 ^ n1299 ;
  assign n33628 = n15568 & n16752 ;
  assign n33629 = n18611 ^ n7187 ^ 1'b0 ;
  assign n33630 = n17294 & n17826 ;
  assign n33631 = n10363 ^ n9066 ^ 1'b0 ;
  assign n33633 = n4545 ^ n1521 ^ 1'b0 ;
  assign n33634 = n3595 | n9077 ;
  assign n33635 = n33633 | n33634 ;
  assign n33632 = ~n14680 & n26389 ;
  assign n33636 = n33635 ^ n33632 ^ 1'b0 ;
  assign n33637 = n11376 | n24892 ;
  assign n33638 = n30802 | n33637 ;
  assign n33639 = n24232 & ~n33638 ;
  assign n33640 = ~n3601 & n7655 ;
  assign n33641 = n16628 ^ n7694 ^ 1'b0 ;
  assign n33642 = n26038 | n33641 ;
  assign n33643 = n9413 ^ n3280 ^ 1'b0 ;
  assign n33644 = ~n5120 & n25708 ;
  assign n33645 = n19650 & n27144 ;
  assign n33646 = n15630 & ~n33645 ;
  assign n33647 = ~n3364 & n33646 ;
  assign n33648 = n33647 ^ n15975 ^ 1'b0 ;
  assign n33649 = ~n7860 & n33648 ;
  assign n33650 = ~n23540 & n29969 ;
  assign n33651 = n33650 ^ n12734 ^ 1'b0 ;
  assign n33652 = n3891 & n9810 ;
  assign n33654 = ~n6082 & n11710 ;
  assign n33655 = n13755 & n33654 ;
  assign n33653 = x100 & n31969 ;
  assign n33656 = n33655 ^ n33653 ^ 1'b0 ;
  assign n33657 = n15651 & ~n20697 ;
  assign n33658 = n3109 | n3549 ;
  assign n33659 = n3109 & ~n33658 ;
  assign n33660 = ~n1360 & n32019 ;
  assign n33661 = n1360 & n33660 ;
  assign n33662 = n33659 | n33661 ;
  assign n33663 = n33659 & ~n33662 ;
  assign n33664 = n25835 | n33663 ;
  assign n33665 = n9551 | n33664 ;
  assign n33666 = ~n22965 & n25140 ;
  assign n33667 = n33398 & n33666 ;
  assign n33668 = n7397 & n25489 ;
  assign n33669 = ~n25489 & n33668 ;
  assign n33670 = ~n9234 & n27003 ;
  assign n33671 = n23754 & n33670 ;
  assign n33672 = n15912 ^ n3258 ^ 1'b0 ;
  assign n33673 = n14381 | n33672 ;
  assign n33675 = n7723 | n24785 ;
  assign n33674 = n2715 | n11427 ;
  assign n33676 = n33675 ^ n33674 ^ 1'b0 ;
  assign n33677 = n23624 ^ n5422 ^ 1'b0 ;
  assign n33678 = n33676 | n33677 ;
  assign n33679 = n33678 ^ n33070 ^ 1'b0 ;
  assign n33680 = n8840 & ~n16659 ;
  assign n33681 = n33680 ^ n8473 ^ 1'b0 ;
  assign n33682 = n6134 | n10826 ;
  assign n33683 = n33681 & ~n33682 ;
  assign n33684 = n33538 ^ n31299 ^ 1'b0 ;
  assign n33685 = n18824 | n33684 ;
  assign n33686 = n9806 & ~n33349 ;
  assign n33687 = n4880 & n31559 ;
  assign n33688 = n33687 ^ n9177 ^ 1'b0 ;
  assign n33689 = n33688 ^ n18455 ^ 1'b0 ;
  assign n33690 = n28577 ^ n580 ^ 1'b0 ;
  assign n33691 = ~n833 & n10316 ;
  assign n33692 = n833 & n33691 ;
  assign n33693 = n2112 & n2655 ;
  assign n33694 = n33692 & n33693 ;
  assign n33695 = n33694 ^ n4645 ^ n3753 ;
  assign n33696 = n33695 ^ n5955 ^ 1'b0 ;
  assign n33697 = n33696 ^ n14451 ^ 1'b0 ;
  assign n33698 = n4730 & ~n17062 ;
  assign n33699 = n11871 & n33698 ;
  assign n33700 = n17475 ^ n8967 ^ 1'b0 ;
  assign n33701 = n25880 ^ n9575 ^ 1'b0 ;
  assign n33702 = n33119 ^ n15665 ^ 1'b0 ;
  assign n33703 = n7118 | n13435 ;
  assign n33704 = n24487 | n27842 ;
  assign n33705 = n10829 ^ n1626 ^ 1'b0 ;
  assign n33706 = n5061 & n33705 ;
  assign n33707 = ~n6381 & n33706 ;
  assign n33708 = ~n1368 & n33707 ;
  assign n33709 = n7599 & ~n11181 ;
  assign n33710 = n14583 & n28082 ;
  assign n33711 = ~n3983 & n9013 ;
  assign n33712 = n14895 ^ n6311 ^ 1'b0 ;
  assign n33713 = n8008 ^ n320 ^ 1'b0 ;
  assign n33714 = n13592 ^ n1521 ^ 1'b0 ;
  assign n33715 = n16600 & ~n33714 ;
  assign n33716 = n9661 & ~n23754 ;
  assign n33717 = n12441 | n33716 ;
  assign n33718 = n10054 & ~n22425 ;
  assign n33719 = n33718 ^ n24561 ^ 1'b0 ;
  assign n33720 = n7644 ^ n4538 ^ 1'b0 ;
  assign n33721 = n33719 & n33720 ;
  assign n33722 = n3854 | n29043 ;
  assign n33723 = n33722 ^ n5761 ^ 1'b0 ;
  assign n33724 = n26846 | n33723 ;
  assign n33725 = n26970 ^ n7333 ^ 1'b0 ;
  assign n33726 = ~n6147 & n33725 ;
  assign n33727 = n20021 ^ n4412 ^ 1'b0 ;
  assign n33728 = ~n8011 & n8892 ;
  assign n33729 = ~n28212 & n33728 ;
  assign n33730 = n13225 ^ n5372 ^ n1608 ;
  assign n33731 = n24832 ^ n2150 ^ 1'b0 ;
  assign n33732 = ( ~n445 & n11705 ) | ( ~n445 & n12932 ) | ( n11705 & n12932 ) ;
  assign n33733 = n18116 & ~n33732 ;
  assign n33734 = n33733 ^ n5475 ^ 1'b0 ;
  assign n33735 = n1928 & n5948 ;
  assign n33736 = n32479 & n33735 ;
  assign n33737 = x132 & ~n11226 ;
  assign n33738 = n4993 & ~n24529 ;
  assign n33739 = ( n2566 & n29127 ) | ( n2566 & n33738 ) | ( n29127 & n33738 ) ;
  assign n33740 = ~n3688 & n5714 ;
  assign n33741 = n33740 ^ n15025 ^ 1'b0 ;
  assign n33742 = n7297 & n10168 ;
  assign n33745 = x90 & ~n10434 ;
  assign n33746 = n33745 ^ n894 ^ 1'b0 ;
  assign n33743 = n7471 & n10135 ;
  assign n33744 = ~n32922 & n33743 ;
  assign n33747 = n33746 ^ n33744 ^ 1'b0 ;
  assign n33748 = n681 & n12860 ;
  assign n33749 = n7519 & ~n33567 ;
  assign n33750 = ~n13983 & n16061 ;
  assign n33751 = n33750 ^ n9012 ^ 1'b0 ;
  assign n33752 = n33749 | n33751 ;
  assign n33753 = n19022 ^ n6548 ^ 1'b0 ;
  assign n33754 = n11891 ^ n610 ^ 1'b0 ;
  assign n33755 = n33754 ^ n25643 ^ 1'b0 ;
  assign n33756 = ~n2305 & n8387 ;
  assign n33757 = n3294 & n8821 ;
  assign n33758 = n33757 ^ n1660 ^ 1'b0 ;
  assign n33759 = n33756 | n33758 ;
  assign n33760 = n14930 ^ n5017 ^ 1'b0 ;
  assign n33761 = n11902 & ~n33760 ;
  assign n33762 = n15853 & n33761 ;
  assign n33763 = n13972 & n33762 ;
  assign n33764 = n10635 & n15919 ;
  assign n33765 = n33764 ^ n14969 ^ 1'b0 ;
  assign n33766 = ( n3746 & n5133 ) | ( n3746 & n33765 ) | ( n5133 & n33765 ) ;
  assign n33767 = n18268 ^ n11506 ^ 1'b0 ;
  assign n33768 = ~n7907 & n33767 ;
  assign n33769 = ~n4694 & n23900 ;
  assign n33770 = n11751 ^ n10844 ^ 1'b0 ;
  assign n33771 = ~n19098 & n33770 ;
  assign n33772 = n12207 | n20259 ;
  assign n33773 = n25169 ^ n22702 ^ 1'b0 ;
  assign n33774 = n12177 ^ n6012 ^ 1'b0 ;
  assign n33775 = n271 & n14391 ;
  assign n33776 = n2047 | n33775 ;
  assign n33777 = ( n8902 & n33774 ) | ( n8902 & n33776 ) | ( n33774 & n33776 ) ;
  assign n33778 = n28563 | n31084 ;
  assign n33779 = n4473 & n13970 ;
  assign n33780 = n28437 & n33779 ;
  assign n33781 = n10692 ^ n6496 ^ 1'b0 ;
  assign n33782 = ~n15124 & n33781 ;
  assign n33783 = n5993 & ~n22331 ;
  assign n33784 = n33783 ^ n13651 ^ 1'b0 ;
  assign n33785 = n2723 & n3911 ;
  assign n33786 = ~n30297 & n33785 ;
  assign n33788 = n8508 ^ n390 ^ 1'b0 ;
  assign n33787 = n17172 | n24470 ;
  assign n33789 = n33788 ^ n33787 ^ 1'b0 ;
  assign n33790 = n2359 & ~n12419 ;
  assign n33791 = n21090 & n33790 ;
  assign n33792 = n30537 ^ n17109 ^ 1'b0 ;
  assign n33793 = n27497 ^ n6553 ^ 1'b0 ;
  assign n33794 = n31054 ^ n27438 ^ n587 ;
  assign n33795 = n24545 & n31863 ;
  assign n33796 = n5386 | n6025 ;
  assign n33797 = n33796 ^ n17552 ^ 1'b0 ;
  assign n33798 = n1704 | n2454 ;
  assign n33799 = n33798 ^ n10854 ^ 1'b0 ;
  assign n33800 = n3060 | n33799 ;
  assign n33801 = n397 & ~n33800 ;
  assign n33802 = n33801 ^ n16037 ^ 1'b0 ;
  assign n33803 = n6455 ^ n1521 ^ 1'b0 ;
  assign n33804 = n8487 & n28455 ;
  assign n33805 = ~n33803 & n33804 ;
  assign n33806 = ~n21712 & n33805 ;
  assign n33807 = ~n15860 & n16601 ;
  assign n33808 = n33807 ^ n14568 ^ 1'b0 ;
  assign n33809 = n2618 & n3014 ;
  assign n33810 = ~n9139 & n20519 ;
  assign n33811 = n33810 ^ n4328 ^ 1'b0 ;
  assign n33812 = n22820 ^ n8541 ^ 1'b0 ;
  assign n33813 = n33811 | n33812 ;
  assign n33814 = n1031 | n33813 ;
  assign n33815 = n8589 & ~n33814 ;
  assign n33816 = n33815 ^ n3045 ^ 1'b0 ;
  assign n33817 = ~n33031 & n33816 ;
  assign n33819 = ~n895 & n11245 ;
  assign n33820 = n33819 ^ n22498 ^ 1'b0 ;
  assign n33818 = ~n875 & n13882 ;
  assign n33821 = n33820 ^ n33818 ^ 1'b0 ;
  assign n33822 = ~n3074 & n24257 ;
  assign n33823 = n26595 ^ n10166 ^ 1'b0 ;
  assign n33824 = ( n9580 & ~n27306 ) | ( n9580 & n33823 ) | ( ~n27306 & n33823 ) ;
  assign n33826 = n6442 & ~n7690 ;
  assign n33827 = n5832 & n33826 ;
  assign n33825 = ~n10329 & n28949 ;
  assign n33828 = n33827 ^ n33825 ^ 1'b0 ;
  assign n33829 = n9256 ^ n2463 ^ 1'b0 ;
  assign n33830 = n14071 | n20316 ;
  assign n33831 = n5845 & ~n14919 ;
  assign n33832 = n15739 ^ n8543 ^ 1'b0 ;
  assign n33833 = n27808 ^ n25835 ^ 1'b0 ;
  assign n33834 = n33832 & n33833 ;
  assign n33835 = n22524 & ~n22746 ;
  assign n33836 = ~n8511 & n33835 ;
  assign n33837 = n33836 ^ n1847 ^ 1'b0 ;
  assign n33838 = n1976 ^ n1299 ^ 1'b0 ;
  assign n33839 = ~n11720 & n33838 ;
  assign n33840 = ~n21045 & n33839 ;
  assign n33841 = n10030 & n16061 ;
  assign n33842 = n17362 & ~n27194 ;
  assign n33843 = n33842 ^ n24363 ^ 1'b0 ;
  assign n33844 = n9479 & n16096 ;
  assign n33845 = n22286 & n33844 ;
  assign n33846 = n3902 | n4576 ;
  assign n33847 = n2875 & n12608 ;
  assign n33848 = ~n1346 & n33847 ;
  assign n33849 = n2099 & n7912 ;
  assign n33850 = n1815 | n24694 ;
  assign n33851 = n33850 ^ n18453 ^ 1'b0 ;
  assign n33852 = n19017 ^ n4398 ^ 1'b0 ;
  assign n33853 = n15545 & ~n33852 ;
  assign n33854 = ~n13080 & n15927 ;
  assign n33855 = n33854 ^ n6511 ^ 1'b0 ;
  assign n33856 = n5160 & ~n18038 ;
  assign n33857 = n33856 ^ n22599 ^ n2276 ;
  assign n33858 = n26270 ^ n1629 ^ 1'b0 ;
  assign n33859 = n13460 | n16652 ;
  assign n33860 = n18530 ^ n11276 ^ 1'b0 ;
  assign n33861 = n4009 | n33860 ;
  assign n33862 = n6948 | n33861 ;
  assign n33863 = n2397 & n5047 ;
  assign n33864 = n29338 ^ n2013 ^ 1'b0 ;
  assign n33865 = n1906 & n33864 ;
  assign n33866 = ~x37 & n19697 ;
  assign n33867 = n31953 ^ n18687 ^ 1'b0 ;
  assign n33868 = ~n26440 & n33867 ;
  assign n33869 = ( n3127 & n3842 ) | ( n3127 & ~n33868 ) | ( n3842 & ~n33868 ) ;
  assign n33870 = n9553 | n27179 ;
  assign n33871 = n33870 ^ n15223 ^ 1'b0 ;
  assign n33872 = ~n13228 & n33871 ;
  assign n33873 = n19429 ^ n9060 ^ 1'b0 ;
  assign n33874 = n23752 ^ n3908 ^ 1'b0 ;
  assign n33875 = n9264 | n31444 ;
  assign n33876 = n33874 & ~n33875 ;
  assign n33877 = n9144 ^ n6391 ^ 1'b0 ;
  assign n33878 = ~n22999 & n33877 ;
  assign n33879 = n33878 ^ n5235 ^ 1'b0 ;
  assign n33880 = n15739 & n33879 ;
  assign n33881 = n10329 | n21018 ;
  assign n33882 = n6745 | n33881 ;
  assign n33883 = n33880 & ~n33882 ;
  assign n33884 = n33883 ^ n12931 ^ 1'b0 ;
  assign n33885 = n33884 ^ n10457 ^ 1'b0 ;
  assign n33886 = n18068 ^ n5704 ^ 1'b0 ;
  assign n33887 = n7325 & n33886 ;
  assign n33888 = n33887 ^ n1383 ^ 1'b0 ;
  assign n33889 = ( n4460 & ~n20158 ) | ( n4460 & n23797 ) | ( ~n20158 & n23797 ) ;
  assign n33890 = ~n14007 & n33889 ;
  assign n33891 = ( ~n1139 & n5371 ) | ( ~n1139 & n5763 ) | ( n5371 & n5763 ) ;
  assign n33892 = n9212 ^ n2107 ^ 1'b0 ;
  assign n33893 = n2868 | n33892 ;
  assign n33894 = n9369 & ~n33893 ;
  assign n33895 = n33891 & n33894 ;
  assign n33896 = n16996 ^ n3978 ^ 1'b0 ;
  assign n33897 = n3768 & ~n16090 ;
  assign n33898 = n16193 | n33897 ;
  assign n33899 = n3955 & ~n28717 ;
  assign n33900 = n31345 & n33899 ;
  assign n33901 = ~n1411 & n14687 ;
  assign n33902 = n2677 & n33901 ;
  assign n33903 = n17594 | n33902 ;
  assign n33904 = n14360 ^ n3265 ^ 1'b0 ;
  assign n33905 = n33903 & n33904 ;
  assign n33906 = n33905 ^ n18648 ^ 1'b0 ;
  assign n33907 = n2718 | n15057 ;
  assign n33908 = n19490 ^ n833 ^ 1'b0 ;
  assign n33909 = n2120 | n33908 ;
  assign n33910 = n5712 & n33909 ;
  assign n33911 = n4063 & n33910 ;
  assign n33912 = n21319 ^ n485 ^ 1'b0 ;
  assign n33913 = n635 & ~n33912 ;
  assign n33914 = ~n5201 & n11696 ;
  assign n33915 = n33914 ^ n16349 ^ 1'b0 ;
  assign n33916 = n7431 & ~n33915 ;
  assign n33917 = n9483 & ~n10105 ;
  assign n33921 = n11551 ^ x204 ^ 1'b0 ;
  assign n33922 = n24753 & ~n33921 ;
  assign n33918 = x63 & ~n2568 ;
  assign n33919 = ~x63 & n33918 ;
  assign n33920 = n1672 | n33919 ;
  assign n33923 = n33922 ^ n33920 ^ 1'b0 ;
  assign n33924 = ~n8964 & n33923 ;
  assign n33925 = ~n9817 & n33924 ;
  assign n33926 = n936 ^ n378 ^ 1'b0 ;
  assign n33927 = ~n18641 & n33926 ;
  assign n33928 = n17015 ^ n14812 ^ 1'b0 ;
  assign n33929 = n17301 | n33928 ;
  assign n33930 = ~n5169 & n27665 ;
  assign n33931 = n14482 | n33930 ;
  assign n33932 = n10637 & ~n33931 ;
  assign n33933 = n33932 ^ n341 ^ 1'b0 ;
  assign n33936 = n27687 ^ n18753 ^ 1'b0 ;
  assign n33934 = n5983 | n9990 ;
  assign n33935 = ~n27738 & n33934 ;
  assign n33937 = n33936 ^ n33935 ^ 1'b0 ;
  assign n33944 = ~n4188 & n22370 ;
  assign n33945 = ~n257 & n33944 ;
  assign n33941 = n7961 ^ n5015 ^ 1'b0 ;
  assign n33938 = n812 & ~n4243 ;
  assign n33939 = n8449 & ~n33938 ;
  assign n33940 = n33939 ^ n19437 ^ 1'b0 ;
  assign n33942 = n33941 ^ n33940 ^ n30315 ;
  assign n33943 = n15974 | n33942 ;
  assign n33946 = n33945 ^ n33943 ^ 1'b0 ;
  assign n33947 = n10168 ^ n8578 ^ 1'b0 ;
  assign n33948 = n5423 & ~n33947 ;
  assign n33949 = n33948 ^ n22389 ^ 1'b0 ;
  assign n33950 = n17909 | n33949 ;
  assign n33951 = n10473 ^ n5186 ^ 1'b0 ;
  assign n33952 = ~n30918 & n33951 ;
  assign n33953 = n33600 ^ n14198 ^ n6555 ;
  assign n33954 = n6585 ^ n4224 ^ 1'b0 ;
  assign n33955 = n7259 ^ n1473 ^ 1'b0 ;
  assign n33956 = n20085 | n33955 ;
  assign n33957 = x134 & n8045 ;
  assign n33958 = n5447 & n33957 ;
  assign n33959 = n4417 & n33958 ;
  assign n33960 = n27237 ^ n23449 ^ 1'b0 ;
  assign n33961 = n28415 & n33960 ;
  assign n33962 = n19439 ^ n5229 ^ 1'b0 ;
  assign n33963 = x213 & n33962 ;
  assign n33964 = n3140 & ~n21435 ;
  assign n33965 = n32343 & n33964 ;
  assign n33966 = n7805 ^ n786 ^ 1'b0 ;
  assign n33967 = n14093 & ~n33966 ;
  assign n33968 = n21246 & ~n29585 ;
  assign n33969 = ~n33967 & n33968 ;
  assign n33970 = n33969 ^ n5931 ^ 1'b0 ;
  assign n33971 = n17317 | n33970 ;
  assign n33972 = n27411 ^ n2747 ^ 1'b0 ;
  assign n33973 = n16817 & n33972 ;
  assign n33974 = n10545 | n31780 ;
  assign n33975 = n2589 & ~n24016 ;
  assign n33976 = ( n438 & ~n33974 ) | ( n438 & n33975 ) | ( ~n33974 & n33975 ) ;
  assign n33977 = x150 & n562 ;
  assign n33978 = ~n22396 & n22689 ;
  assign n33979 = ~n33977 & n33978 ;
  assign n33980 = n3794 & ~n7509 ;
  assign n33981 = n19024 ^ n14349 ^ 1'b0 ;
  assign n33982 = n4843 & ~n33981 ;
  assign n33983 = n19041 | n23506 ;
  assign n33984 = n13844 ^ n3945 ^ 1'b0 ;
  assign n33985 = ~n8340 & n33984 ;
  assign n33986 = n33985 ^ n33022 ^ n18658 ;
  assign n33987 = n1283 & ~n33986 ;
  assign n33988 = n1177 & n8145 ;
  assign n33989 = n33988 ^ n16110 ^ 1'b0 ;
  assign n33990 = n4414 & n19388 ;
  assign n33991 = n33990 ^ n7214 ^ n4001 ;
  assign n33992 = n30828 ^ n19052 ^ 1'b0 ;
  assign n33993 = n8821 & ~n33992 ;
  assign n33994 = n11457 & n28866 ;
  assign n33995 = n33994 ^ x48 ^ 1'b0 ;
  assign n33996 = n21630 ^ n8427 ^ n2975 ;
  assign n33997 = n5880 | n33996 ;
  assign n33998 = n259 & n18069 ;
  assign n33999 = n33998 ^ n3334 ^ 1'b0 ;
  assign n34000 = n33999 ^ n31048 ^ n18913 ;
  assign n34001 = n5064 ^ n3703 ^ 1'b0 ;
  assign n34002 = n9375 | n34001 ;
  assign n34003 = n13808 & n34002 ;
  assign n34004 = n978 & ~n8127 ;
  assign n34005 = n20612 ^ n7282 ^ 1'b0 ;
  assign n34006 = n19320 | n34005 ;
  assign n34007 = n32445 ^ n16211 ^ n4388 ;
  assign n34008 = n360 ^ x76 ^ 1'b0 ;
  assign n34009 = n21522 ^ n5896 ^ 1'b0 ;
  assign n34010 = n14000 & ~n34009 ;
  assign n34011 = n34010 ^ n18676 ^ 1'b0 ;
  assign n34012 = n6715 & n16052 ;
  assign n34013 = ~n31637 & n34012 ;
  assign n34014 = n5207 | n15876 ;
  assign n34015 = n19187 & n34014 ;
  assign n34016 = n20419 ^ n20261 ^ 1'b0 ;
  assign n34017 = n34016 ^ n24351 ^ 1'b0 ;
  assign n34018 = n5985 | n9769 ;
  assign n34019 = n3768 & ~n5210 ;
  assign n34020 = n16160 & n34019 ;
  assign n34021 = ( n13335 & n25710 ) | ( n13335 & ~n26125 ) | ( n25710 & ~n26125 ) ;
  assign n34022 = n15723 ^ n14252 ^ 1'b0 ;
  assign n34023 = n1728 & ~n4671 ;
  assign n34024 = n1038 & ~n34023 ;
  assign n34025 = ~n34022 & n34024 ;
  assign n34026 = n17168 ^ n12309 ^ 1'b0 ;
  assign n34027 = ~n1299 & n4490 ;
  assign n34028 = n7252 & n34027 ;
  assign n34029 = n16750 | n20650 ;
  assign n34030 = ~n11210 & n20019 ;
  assign n34031 = n3643 ^ n1773 ^ 1'b0 ;
  assign n34032 = n10162 & n34031 ;
  assign n34033 = n20606 ^ n5088 ^ 1'b0 ;
  assign n34034 = n20975 ^ n18096 ^ 1'b0 ;
  assign n34035 = x212 & ~n7931 ;
  assign n34036 = n6661 | n19363 ;
  assign n34037 = n9728 | n33298 ;
  assign n34038 = ~n532 & n34037 ;
  assign n34039 = ~n1361 & n24388 ;
  assign n34040 = n9527 ^ x46 ^ 1'b0 ;
  assign n34041 = ~n397 & n34040 ;
  assign n34042 = n774 & n34041 ;
  assign n34043 = n6233 ^ n4016 ^ 1'b0 ;
  assign n34044 = n34042 & ~n34043 ;
  assign n34045 = n415 | n10328 ;
  assign n34046 = n33119 & ~n34045 ;
  assign n34047 = n16841 ^ n13757 ^ 1'b0 ;
  assign n34048 = n10691 ^ n6764 ^ 1'b0 ;
  assign n34049 = n34047 | n34048 ;
  assign n34050 = ~n577 & n20630 ;
  assign n34051 = n34050 ^ n4108 ^ 1'b0 ;
  assign n34052 = n34051 ^ n21751 ^ 1'b0 ;
  assign n34053 = n5728 & n34052 ;
  assign n34054 = ~n2029 & n3407 ;
  assign n34055 = ~n10214 & n34054 ;
  assign n34056 = n34055 ^ n7136 ^ 1'b0 ;
  assign n34057 = n21111 ^ n17750 ^ 1'b0 ;
  assign n34058 = n20274 & ~n34057 ;
  assign n34059 = ~n3176 & n15339 ;
  assign n34060 = ~n14022 & n34059 ;
  assign n34061 = n34060 ^ n22481 ^ 1'b0 ;
  assign n34062 = n28732 ^ n6558 ^ 1'b0 ;
  assign n34063 = n9864 ^ n1646 ^ 1'b0 ;
  assign n34064 = ~n3855 & n34063 ;
  assign n34065 = n34064 ^ n1236 ^ 1'b0 ;
  assign n34066 = n34062 & ~n34065 ;
  assign n34067 = n34066 ^ n20078 ^ 1'b0 ;
  assign n34068 = n12147 & ~n34067 ;
  assign n34069 = n527 | n2623 ;
  assign n34070 = ( n21019 & n25167 ) | ( n21019 & n34069 ) | ( n25167 & n34069 ) ;
  assign n34071 = n22105 & ~n29747 ;
  assign n34072 = n34071 ^ n13697 ^ 1'b0 ;
  assign n34073 = ( n1714 & n6412 ) | ( n1714 & ~n33335 ) | ( n6412 & ~n33335 ) ;
  assign n34074 = n6940 | n7729 ;
  assign n34075 = n13850 ^ n3649 ^ 1'b0 ;
  assign n34076 = n17046 & ~n34075 ;
  assign n34077 = n34074 & n34076 ;
  assign n34078 = n30890 & n34077 ;
  assign n34079 = n5396 | n14525 ;
  assign n34080 = n4524 | n34079 ;
  assign n34081 = n25728 & n34080 ;
  assign n34082 = n2122 & n34081 ;
  assign n34083 = n5446 & n9534 ;
  assign n34084 = ~n11443 & n34083 ;
  assign n34085 = n34084 ^ n458 ^ x134 ;
  assign n34086 = ( n6020 & n22133 ) | ( n6020 & n34085 ) | ( n22133 & n34085 ) ;
  assign n34087 = n14981 ^ n10025 ^ 1'b0 ;
  assign n34088 = n6938 & ~n31645 ;
  assign n34092 = n13813 ^ n10619 ^ 1'b0 ;
  assign n34093 = n19278 | n34092 ;
  assign n34089 = n944 & ~n7169 ;
  assign n34090 = n34089 ^ n8708 ^ 1'b0 ;
  assign n34091 = n343 & n34090 ;
  assign n34094 = n34093 ^ n34091 ^ 1'b0 ;
  assign n34095 = n14498 & n25604 ;
  assign n34096 = n34095 ^ n13953 ^ 1'b0 ;
  assign n34097 = x124 | n2725 ;
  assign n34098 = n3266 | n7074 ;
  assign n34099 = n34098 ^ n19588 ^ 1'b0 ;
  assign n34100 = n32819 & ~n34099 ;
  assign n34101 = x101 | n16818 ;
  assign n34102 = n8919 ^ n6838 ^ 1'b0 ;
  assign n34103 = n10058 ^ n2761 ^ 1'b0 ;
  assign n34104 = n30843 ^ n15918 ^ 1'b0 ;
  assign n34105 = n1610 & n3086 ;
  assign n34106 = n18236 ^ n3965 ^ 1'b0 ;
  assign n34107 = n13362 & ~n23329 ;
  assign n34108 = n7882 & n34107 ;
  assign n34109 = n15212 & n18796 ;
  assign n34110 = ~n8257 & n23574 ;
  assign n34111 = n23898 & n34110 ;
  assign n34112 = n5774 & n19652 ;
  assign n34113 = n32855 & n34112 ;
  assign n34114 = n3018 & ~n24459 ;
  assign n34115 = n13052 & n34114 ;
  assign n34116 = n3221 & n7259 ;
  assign n34117 = ~n4523 & n34116 ;
  assign n34118 = n7126 & n9558 ;
  assign n34119 = n34117 & n34118 ;
  assign n34120 = n13076 ^ n7925 ^ 1'b0 ;
  assign n34121 = n9911 & n34120 ;
  assign n34122 = x177 & ~n8317 ;
  assign n34123 = ( n6802 & n34121 ) | ( n6802 & ~n34122 ) | ( n34121 & ~n34122 ) ;
  assign n34124 = ( n11274 & n32845 ) | ( n11274 & ~n34123 ) | ( n32845 & ~n34123 ) ;
  assign n34125 = n12194 & ~n34124 ;
  assign n34126 = n14210 | n14525 ;
  assign n34127 = n23308 ^ n10263 ^ 1'b0 ;
  assign n34128 = n34126 & ~n34127 ;
  assign n34129 = n3057 ^ n828 ^ 1'b0 ;
  assign n34130 = n10458 | n34129 ;
  assign n34131 = n34130 ^ n27570 ^ n5965 ;
  assign n34132 = n937 & ~n22776 ;
  assign n34133 = n26122 | n28601 ;
  assign n34134 = n2060 & ~n12194 ;
  assign n34135 = ~n1444 & n34134 ;
  assign n34136 = x80 & n6747 ;
  assign n34137 = n30073 & n34136 ;
  assign n34138 = n22296 ^ n7169 ^ 1'b0 ;
  assign n34139 = ( n844 & n9366 ) | ( n844 & ~n34138 ) | ( n9366 & ~n34138 ) ;
  assign n34140 = n20144 & n34139 ;
  assign n34141 = n34140 ^ n31948 ^ 1'b0 ;
  assign n34142 = n9607 | n29658 ;
  assign n34143 = n2012 ^ n605 ^ 1'b0 ;
  assign n34144 = n16264 & n24016 ;
  assign n34145 = n4013 & n34144 ;
  assign n34146 = ~n10980 & n15935 ;
  assign n34147 = n22725 ^ n12417 ^ n738 ;
  assign n34148 = n8127 & ~n12601 ;
  assign n34149 = n34148 ^ n14197 ^ 1'b0 ;
  assign n34150 = n5965 & n9652 ;
  assign n34151 = n1605 | n4815 ;
  assign n34152 = n4791 & ~n15232 ;
  assign n34153 = n8849 & ~n34152 ;
  assign n34154 = n28280 ^ n21644 ^ 1'b0 ;
  assign n34155 = n3055 | n34154 ;
  assign n34156 = n7491 & ~n10626 ;
  assign n34157 = n4065 & n34156 ;
  assign n34158 = n34157 ^ n2849 ^ 1'b0 ;
  assign n34159 = n24028 ^ n11374 ^ 1'b0 ;
  assign n34160 = n4935 & n7669 ;
  assign n34161 = n1154 & ~n9356 ;
  assign n34162 = n12916 & n34161 ;
  assign n34163 = n12390 | n34162 ;
  assign n34164 = n34160 | n34163 ;
  assign n34165 = ~n11869 & n13595 ;
  assign n34166 = ~n15641 & n34165 ;
  assign n34168 = n17542 | n25713 ;
  assign n34167 = n1658 | n25442 ;
  assign n34169 = n34168 ^ n34167 ^ 1'b0 ;
  assign n34170 = n3877 & n18157 ;
  assign n34171 = ~n32970 & n34170 ;
  assign n34172 = n34171 ^ n305 ^ 1'b0 ;
  assign n34173 = ~x123 & n34172 ;
  assign n34174 = ( n34166 & ~n34169 ) | ( n34166 & n34173 ) | ( ~n34169 & n34173 ) ;
  assign n34175 = n21975 ^ n7966 ^ 1'b0 ;
  assign n34176 = x254 | n34175 ;
  assign n34177 = n7340 & ~n28985 ;
  assign n34178 = n1809 & n14842 ;
  assign n34179 = n34178 ^ n28855 ^ 1'b0 ;
  assign n34180 = n13821 & ~n18680 ;
  assign n34181 = n34180 ^ n9276 ^ 1'b0 ;
  assign n34182 = n1134 & ~n26064 ;
  assign n34183 = ~n26886 & n34182 ;
  assign n34184 = n30783 ^ n25169 ^ 1'b0 ;
  assign n34185 = n5996 & ~n7251 ;
  assign n34187 = n24088 & ~n31729 ;
  assign n34186 = n13377 & n13627 ;
  assign n34188 = n34187 ^ n34186 ^ 1'b0 ;
  assign n34189 = n3229 | n9339 ;
  assign n34190 = n1302 & n25888 ;
  assign n34191 = n17307 | n30843 ;
  assign n34192 = n4347 & ~n34191 ;
  assign n34193 = n34192 ^ n22899 ^ n2464 ;
  assign n34194 = n14982 ^ n6934 ^ 1'b0 ;
  assign n34195 = n28733 ^ n12577 ^ 1'b0 ;
  assign n34196 = n34194 | n34195 ;
  assign n34197 = n29811 | n34196 ;
  assign n34198 = n7824 | n7841 ;
  assign n34200 = n2700 | n22095 ;
  assign n34201 = n7628 | n34200 ;
  assign n34199 = n4211 ^ n3509 ^ 1'b0 ;
  assign n34202 = n34201 ^ n34199 ^ 1'b0 ;
  assign n34203 = n1472 | n28294 ;
  assign n34204 = ~n1751 & n34203 ;
  assign n34205 = n34204 ^ n2903 ^ 1'b0 ;
  assign n34206 = n3140 & n13395 ;
  assign n34207 = n13745 & ~n32405 ;
  assign n34208 = n951 & ~n16332 ;
  assign n34209 = ~n3758 & n34208 ;
  assign n34210 = n34209 ^ n15529 ^ 1'b0 ;
  assign n34212 = ~n2166 & n16357 ;
  assign n34211 = ~n13603 & n26864 ;
  assign n34213 = n34212 ^ n34211 ^ 1'b0 ;
  assign n34214 = n21059 ^ n16750 ^ 1'b0 ;
  assign n34215 = n22659 ^ n13413 ^ 1'b0 ;
  assign n34216 = n4767 & ~n6572 ;
  assign n34217 = n34216 ^ n30953 ^ 1'b0 ;
  assign n34218 = n1654 | n5100 ;
  assign n34219 = n9388 & n34218 ;
  assign n34220 = n34219 ^ n7484 ^ 1'b0 ;
  assign n34221 = n6760 & ~n14073 ;
  assign n34222 = n31099 ^ n9793 ^ n651 ;
  assign n34223 = n13293 | n18278 ;
  assign n34224 = n16090 ^ n11800 ^ 1'b0 ;
  assign n34225 = ~n747 & n34224 ;
  assign n34226 = n34225 ^ n2970 ^ 1'b0 ;
  assign n34227 = n4375 & n34226 ;
  assign n34228 = ~n3395 & n11339 ;
  assign n34229 = n3395 & n34228 ;
  assign n34230 = n1451 | n34229 ;
  assign n34231 = n1451 & ~n34230 ;
  assign n34232 = n8719 & ~n11486 ;
  assign n34233 = n34231 & n34232 ;
  assign n34234 = n23165 | n34233 ;
  assign n34235 = n7571 & ~n34234 ;
  assign n34236 = n552 & n16734 ;
  assign n34237 = n480 & ~n1219 ;
  assign n34238 = x194 & n2718 ;
  assign n34239 = ~n2718 & n34238 ;
  assign n34240 = ~n15682 & n34239 ;
  assign n34241 = n34240 ^ n20477 ^ 1'b0 ;
  assign n34242 = n34237 & ~n34241 ;
  assign n34243 = x43 & ~n3288 ;
  assign n34244 = ~n4733 & n34243 ;
  assign n34245 = ( n4118 & n4600 ) | ( n4118 & ~n6411 ) | ( n4600 & ~n6411 ) ;
  assign n34246 = n16364 & ~n34245 ;
  assign n34247 = n23493 & n34246 ;
  assign n34248 = ~n4982 & n28196 ;
  assign n34249 = n34248 ^ n22591 ^ 1'b0 ;
  assign n34250 = n12943 & n16357 ;
  assign n34252 = n16163 ^ n9176 ^ 1'b0 ;
  assign n34251 = n1353 & n17096 ;
  assign n34253 = n34252 ^ n34251 ^ 1'b0 ;
  assign n34254 = n25896 ^ n4538 ^ 1'b0 ;
  assign n34255 = ~n32359 & n34254 ;
  assign n34256 = ~n24286 & n34255 ;
  assign n34257 = n3187 & n34256 ;
  assign n34258 = n34257 ^ n17960 ^ 1'b0 ;
  assign n34259 = n11370 & ~n17344 ;
  assign n34260 = n16337 ^ n2392 ^ 1'b0 ;
  assign n34261 = n20469 | n34260 ;
  assign n34262 = n2243 | n26817 ;
  assign n34263 = n34262 ^ n16154 ^ 1'b0 ;
  assign n34264 = x141 & n28812 ;
  assign n34265 = n34264 ^ n10668 ^ 1'b0 ;
  assign n34266 = n34265 ^ n26884 ^ 1'b0 ;
  assign n34267 = n17660 & ~n34266 ;
  assign n34268 = ~n7720 & n11280 ;
  assign n34269 = n21744 & ~n34268 ;
  assign n34270 = n2901 & ~n34269 ;
  assign n34271 = n34270 ^ n3440 ^ 1'b0 ;
  assign n34272 = n2185 & n24320 ;
  assign n34273 = n34272 ^ n1925 ^ 1'b0 ;
  assign n34276 = n3773 | n14451 ;
  assign n34277 = n34276 ^ n5865 ^ 1'b0 ;
  assign n34274 = ~n13916 & n20454 ;
  assign n34275 = n8261 & ~n34274 ;
  assign n34278 = n34277 ^ n34275 ^ 1'b0 ;
  assign n34279 = n34278 ^ n24134 ^ 1'b0 ;
  assign n34280 = n21103 ^ n5828 ^ 1'b0 ;
  assign n34281 = n1829 & n34280 ;
  assign n34282 = n4695 | n17536 ;
  assign n34283 = n33038 ^ n1724 ^ 1'b0 ;
  assign n34284 = n34282 & n34283 ;
  assign n34285 = ~n9558 & n21338 ;
  assign n34286 = ~n19299 & n34285 ;
  assign n34287 = n16627 & n34286 ;
  assign n34288 = n6295 & ~n34287 ;
  assign n34289 = n1361 & n1368 ;
  assign n34290 = n34289 ^ n1740 ^ 1'b0 ;
  assign n34291 = n34290 ^ n12707 ^ n1859 ;
  assign n34292 = n34291 ^ n20708 ^ n4294 ;
  assign n34295 = n5692 ^ n703 ^ 1'b0 ;
  assign n34293 = ~n3628 & n10016 ;
  assign n34294 = n14561 & n34293 ;
  assign n34296 = n34295 ^ n34294 ^ 1'b0 ;
  assign n34297 = n34296 ^ n11119 ^ 1'b0 ;
  assign n34298 = n27640 & n34297 ;
  assign n34299 = ( n681 & ~n3753 ) | ( n681 & n11385 ) | ( ~n3753 & n11385 ) ;
  assign n34300 = n12982 ^ n7257 ^ 1'b0 ;
  assign n34301 = n25570 ^ n2860 ^ 1'b0 ;
  assign n34302 = ~n24638 & n34301 ;
  assign n34303 = n11486 | n21714 ;
  assign n34304 = n3624 & ~n34303 ;
  assign n34305 = n12230 & ~n30410 ;
  assign n34306 = ~n2307 & n34305 ;
  assign n34307 = n34304 | n34306 ;
  assign n34308 = n34307 ^ n28432 ^ 1'b0 ;
  assign n34309 = n34308 ^ n2350 ^ 1'b0 ;
  assign n34310 = n34309 ^ n8322 ^ 1'b0 ;
  assign n34311 = n22677 & ~n34310 ;
  assign n34312 = n14524 ^ n10570 ^ 1'b0 ;
  assign n34313 = ~n2060 & n2320 ;
  assign n34314 = n29333 ^ n11341 ^ 1'b0 ;
  assign n34315 = n6562 & n15028 ;
  assign n34316 = ~x76 & n23347 ;
  assign n34317 = n34316 ^ n15711 ^ n7475 ;
  assign n34318 = n34315 & n34317 ;
  assign n34319 = n14522 ^ n12750 ^ 1'b0 ;
  assign n34320 = n1264 & n3116 ;
  assign n34321 = ~n2664 & n34320 ;
  assign n34322 = n14783 | n34321 ;
  assign n34325 = n22999 ^ n17710 ^ n10568 ;
  assign n34324 = n14780 | n22041 ;
  assign n34326 = n34325 ^ n34324 ^ 1'b0 ;
  assign n34327 = x225 & ~n34326 ;
  assign n34328 = n34327 ^ n5250 ^ 1'b0 ;
  assign n34323 = n15535 & ~n17254 ;
  assign n34329 = n34328 ^ n34323 ^ 1'b0 ;
  assign n34330 = n8609 ^ n1926 ^ 1'b0 ;
  assign n34331 = n12142 | n34330 ;
  assign n34332 = n8627 ^ n5470 ^ n602 ;
  assign n34333 = n4641 & ~n17716 ;
  assign n34334 = ~n17370 & n34333 ;
  assign n34335 = ~n22290 & n31922 ;
  assign n34336 = n18831 ^ n3193 ^ n1629 ;
  assign n34337 = x0 & ~n19780 ;
  assign n34338 = n27208 ^ n16478 ^ 1'b0 ;
  assign n34339 = n2892 | n5445 ;
  assign n34340 = n34339 ^ n18068 ^ n5913 ;
  assign n34341 = n460 | n956 ;
  assign n34342 = n33308 ^ n26590 ^ 1'b0 ;
  assign n34343 = n34341 | n34342 ;
  assign n34344 = n5354 & ~n34343 ;
  assign n34345 = n34344 ^ n6267 ^ 1'b0 ;
  assign n34346 = n859 & n15907 ;
  assign n34347 = ~n23230 & n34346 ;
  assign n34348 = ~n9589 & n19911 ;
  assign n34349 = n34348 ^ n27204 ^ 1'b0 ;
  assign n34350 = n20229 ^ n7633 ^ 1'b0 ;
  assign n34351 = n1784 & ~n34350 ;
  assign n34352 = ~n9207 & n34351 ;
  assign n34353 = n14424 ^ n5678 ^ n2324 ;
  assign n34354 = n30501 ^ n11226 ^ 1'b0 ;
  assign n34355 = n3295 & ~n34354 ;
  assign n34356 = n25418 ^ n16495 ^ 1'b0 ;
  assign n34357 = n3988 & n6471 ;
  assign n34358 = n5413 & ~n34357 ;
  assign n34359 = n3181 & n8687 ;
  assign n34360 = n34359 ^ n33238 ^ 1'b0 ;
  assign n34361 = n15039 | n19858 ;
  assign n34362 = n4413 | n7982 ;
  assign n34363 = n3714 | n34362 ;
  assign n34364 = n34363 ^ n8294 ^ 1'b0 ;
  assign n34365 = ~n16815 & n34364 ;
  assign n34366 = x213 & n3552 ;
  assign n34367 = ~n34365 & n34366 ;
  assign n34368 = n34367 ^ n3714 ^ 1'b0 ;
  assign n34369 = n15295 ^ n3836 ^ 1'b0 ;
  assign n34370 = x78 & n34369 ;
  assign n34371 = n34370 ^ n12827 ^ 1'b0 ;
  assign n34372 = n12660 ^ n9986 ^ 1'b0 ;
  assign n34373 = n34372 ^ n21012 ^ n4961 ;
  assign n34374 = n34373 ^ n26833 ^ 1'b0 ;
  assign n34375 = n8014 | n34374 ;
  assign n34376 = n1825 & n2672 ;
  assign n34377 = n34376 ^ n24396 ^ 1'b0 ;
  assign n34378 = n19977 ^ n10939 ^ 1'b0 ;
  assign n34379 = n5242 & n34378 ;
  assign n34380 = n34379 ^ n7578 ^ 1'b0 ;
  assign n34381 = n15178 & ~n23966 ;
  assign n34382 = ~n7281 & n34381 ;
  assign n34383 = n14531 & ~n34382 ;
  assign n34384 = n25432 ^ n9092 ^ 1'b0 ;
  assign n34385 = n32708 ^ n1859 ^ 1'b0 ;
  assign n34386 = n3009 & ~n34385 ;
  assign n34387 = ~n10952 & n18630 ;
  assign n34388 = n34387 ^ n22722 ^ 1'b0 ;
  assign n34389 = n16204 & ~n21121 ;
  assign n34390 = n1295 & n34389 ;
  assign n34391 = n11221 ^ n8002 ^ 1'b0 ;
  assign n34392 = ( ~n23894 & n25856 ) | ( ~n23894 & n34391 ) | ( n25856 & n34391 ) ;
  assign n34393 = n9165 | n18122 ;
  assign n34394 = n13321 | n34393 ;
  assign n34395 = n12064 & ~n34394 ;
  assign n34397 = n21542 ^ n8622 ^ 1'b0 ;
  assign n34398 = ~n16892 & n29753 ;
  assign n34399 = n34397 & n34398 ;
  assign n34396 = ~n4658 & n10213 ;
  assign n34400 = n34399 ^ n34396 ^ 1'b0 ;
  assign n34401 = n4972 & ~n13077 ;
  assign n34402 = n34401 ^ n760 ^ 1'b0 ;
  assign n34403 = n741 | n34402 ;
  assign n34404 = n34403 ^ n15751 ^ 1'b0 ;
  assign n34405 = n12966 ^ n11763 ^ 1'b0 ;
  assign n34406 = n8803 | n34405 ;
  assign n34407 = n15607 & n24853 ;
  assign n34408 = ~n8049 & n34407 ;
  assign n34409 = n16207 | n25671 ;
  assign n34410 = n29409 | n34409 ;
  assign n34411 = ~n8180 & n32019 ;
  assign n34413 = n5904 ^ n3169 ^ 1'b0 ;
  assign n34412 = x222 & ~n12744 ;
  assign n34414 = n34413 ^ n34412 ^ 1'b0 ;
  assign n34415 = n34414 ^ n4348 ^ 1'b0 ;
  assign n34416 = n16649 ^ n7575 ^ 1'b0 ;
  assign n34417 = n11075 & ~n34416 ;
  assign n34418 = ~n2247 & n34417 ;
  assign n34419 = n2793 | n34418 ;
  assign n34420 = n34415 | n34419 ;
  assign n34421 = ~n14025 & n34420 ;
  assign n34422 = ~n34411 & n34421 ;
  assign n34423 = n15411 & n22820 ;
  assign n34424 = n14459 ^ n2366 ^ 1'b0 ;
  assign n34425 = n34423 & n34424 ;
  assign n34426 = n4802 & ~n10728 ;
  assign n34427 = n34426 ^ n17788 ^ 1'b0 ;
  assign n34428 = n29524 | n34427 ;
  assign n34429 = n10936 & n20812 ;
  assign n34430 = n9835 ^ n1805 ^ 1'b0 ;
  assign n34431 = n2569 ^ x127 ^ 1'b0 ;
  assign n34432 = n34430 & n34431 ;
  assign n34433 = n2518 & n34432 ;
  assign n34434 = n34429 & n34433 ;
  assign n34435 = n5351 ^ n3794 ^ 1'b0 ;
  assign n34436 = n9809 & ~n34435 ;
  assign n34437 = n15208 ^ n2883 ^ 1'b0 ;
  assign n34438 = n6527 & n20519 ;
  assign n34439 = ~n445 & n34438 ;
  assign n34440 = n26056 ^ n10195 ^ 1'b0 ;
  assign n34441 = n21995 & ~n34440 ;
  assign n34442 = ~n19465 & n25735 ;
  assign n34443 = n8200 & n34442 ;
  assign n34444 = n34443 ^ n14871 ^ 1'b0 ;
  assign n34445 = n19468 ^ n3695 ^ 1'b0 ;
  assign n34446 = n34445 ^ n14294 ^ 1'b0 ;
  assign n34447 = ~n11433 & n34446 ;
  assign n34448 = ~n34444 & n34447 ;
  assign n34449 = n485 & n6843 ;
  assign n34450 = n15320 ^ n14316 ^ 1'b0 ;
  assign n34451 = n27803 & ~n34450 ;
  assign n34452 = n22431 ^ n19082 ^ 1'b0 ;
  assign n34453 = n4177 & n6419 ;
  assign n34454 = n26064 ^ n6312 ^ 1'b0 ;
  assign n34455 = x90 & n34454 ;
  assign n34456 = n15184 & n20292 ;
  assign n34457 = ~n3546 & n11920 ;
  assign n34458 = n26257 ^ n5506 ^ 1'b0 ;
  assign n34459 = n4922 | n34458 ;
  assign n34460 = ~n2185 & n19819 ;
  assign n34461 = n19685 & ~n26197 ;
  assign n34462 = n15584 & n34461 ;
  assign n34463 = n27443 & n34462 ;
  assign n34464 = ~n4358 & n16789 ;
  assign n34465 = n34464 ^ n13373 ^ 1'b0 ;
  assign n34466 = ~n5728 & n34465 ;
  assign n34467 = n34466 ^ n9193 ^ 1'b0 ;
  assign n34468 = n1009 | n1919 ;
  assign n34469 = n27862 & ~n34468 ;
  assign n34470 = x87 & n34469 ;
  assign n34471 = n686 & ~n34470 ;
  assign n34472 = ~n22296 & n34471 ;
  assign n34473 = n1920 | n34472 ;
  assign n34474 = n5999 & ~n28176 ;
  assign n34475 = n16429 & n34474 ;
  assign n34476 = n3957 ^ n1900 ^ 1'b0 ;
  assign n34477 = n6527 | n16591 ;
  assign n34478 = ~n2374 & n34477 ;
  assign n34479 = n10357 & n34478 ;
  assign n34480 = n8449 | n34479 ;
  assign n34481 = ~n354 & n12756 ;
  assign n34482 = n8345 & n27164 ;
  assign n34483 = n10612 & ~n12349 ;
  assign n34484 = n34483 ^ n6372 ^ 1'b0 ;
  assign n34485 = n7183 & ~n24569 ;
  assign n34486 = n34485 ^ n15701 ^ 1'b0 ;
  assign n34487 = n14401 & n29539 ;
  assign n34488 = n34487 ^ n27242 ^ 1'b0 ;
  assign n34489 = n17324 ^ n16343 ^ 1'b0 ;
  assign n34490 = ~n5798 & n12364 ;
  assign n34491 = ~n29640 & n34490 ;
  assign n34492 = n13046 | n32143 ;
  assign n34493 = n28585 & ~n34492 ;
  assign n34494 = n11176 | n34282 ;
  assign n34495 = n10792 | n31467 ;
  assign n34496 = n34495 ^ n21012 ^ 1'b0 ;
  assign n34498 = n15707 ^ n12923 ^ 1'b0 ;
  assign n34497 = n8218 & n9579 ;
  assign n34499 = n34498 ^ n34497 ^ 1'b0 ;
  assign n34500 = n27532 & ~n34499 ;
  assign n34501 = n3441 & n34500 ;
  assign n34502 = ~n6146 & n6443 ;
  assign n34503 = n34502 ^ n4398 ^ 1'b0 ;
  assign n34504 = ~n4808 & n34503 ;
  assign n34505 = n1190 | n1473 ;
  assign n34506 = n34505 ^ n2778 ^ 1'b0 ;
  assign n34507 = n13420 ^ n3807 ^ 1'b0 ;
  assign n34508 = n20993 & ~n34507 ;
  assign n34509 = n28388 ^ n2180 ^ 1'b0 ;
  assign n34510 = n34508 & n34509 ;
  assign n34511 = n2602 ^ x98 ^ 1'b0 ;
  assign n34512 = ~n8175 & n34511 ;
  assign n34513 = n1444 & n27627 ;
  assign n34514 = ~n19189 & n34513 ;
  assign n34515 = n4819 & n10517 ;
  assign n34516 = n34515 ^ x249 ^ 1'b0 ;
  assign n34517 = n34516 ^ n16787 ^ n6573 ;
  assign n34518 = ~n3100 & n10364 ;
  assign n34519 = n23905 & n34518 ;
  assign n34520 = n3191 ^ n880 ^ 1'b0 ;
  assign n34521 = n13696 & ~n17182 ;
  assign n34522 = n34521 ^ n16456 ^ n9400 ;
  assign n34523 = n12763 & ~n31857 ;
  assign n34524 = n34523 ^ n478 ^ 1'b0 ;
  assign n34525 = n34522 & ~n34524 ;
  assign n34526 = n9562 | n14185 ;
  assign n34527 = n6231 | n11269 ;
  assign n34528 = n5465 | n34527 ;
  assign n34529 = n298 & ~n34528 ;
  assign n34530 = ( n6927 & n16144 ) | ( n6927 & n34529 ) | ( n16144 & n34529 ) ;
  assign n34531 = n8520 | n14805 ;
  assign n34532 = n3979 | n34531 ;
  assign n34533 = n6288 & n34532 ;
  assign n34534 = n34533 ^ n7484 ^ 1'b0 ;
  assign n34535 = ~n602 & n6644 ;
  assign n34536 = ~n8223 & n17497 ;
  assign n34537 = n27850 & n34536 ;
  assign n34538 = n34537 ^ n25885 ^ 1'b0 ;
  assign n34539 = n11101 & ~n34538 ;
  assign n34540 = ~n4091 & n24354 ;
  assign n34541 = n10145 | n18126 ;
  assign n34542 = n3865 | n28339 ;
  assign n34543 = n20412 | n34542 ;
  assign n34544 = n34543 ^ n5847 ^ 1'b0 ;
  assign n34545 = n11330 ^ n1736 ^ 1'b0 ;
  assign n34546 = n34545 ^ n23252 ^ 1'b0 ;
  assign n34547 = ~n9029 & n34546 ;
  assign n34548 = n8841 & n26534 ;
  assign n34549 = n3754 & ~n20692 ;
  assign n34550 = n29014 ^ n21115 ^ 1'b0 ;
  assign n34551 = ~n4892 & n34550 ;
  assign n34552 = ~n11854 & n24879 ;
  assign n34553 = n16982 ^ n10166 ^ 1'b0 ;
  assign n34554 = n14448 & n34553 ;
  assign n34555 = n11130 ^ n9311 ^ 1'b0 ;
  assign n34556 = n24433 ^ n7005 ^ 1'b0 ;
  assign n34557 = n6505 & ~n31271 ;
  assign n34558 = n15361 & n34557 ;
  assign n34559 = ~n10269 & n34558 ;
  assign n34560 = n3469 & n22164 ;
  assign n34561 = n33234 ^ n13027 ^ 1'b0 ;
  assign n34562 = ~n22032 & n34561 ;
  assign n34563 = ~n19777 & n34562 ;
  assign n34564 = n10650 ^ n4411 ^ 1'b0 ;
  assign n34565 = n3746 & n13627 ;
  assign n34566 = ~n12238 & n34565 ;
  assign n34567 = n1402 & ~n10005 ;
  assign n34568 = ~n24477 & n34567 ;
  assign n34569 = n34568 ^ n17111 ^ 1'b0 ;
  assign n34570 = n8397 & n34569 ;
  assign n34571 = n784 | n34570 ;
  assign n34572 = n14302 ^ n7713 ^ 1'b0 ;
  assign n34573 = n34572 ^ n28310 ^ n5236 ;
  assign n34574 = n12997 ^ n8470 ^ 1'b0 ;
  assign n34575 = ~n4712 & n28545 ;
  assign n34577 = n5679 ^ n5452 ^ 1'b0 ;
  assign n34578 = n1976 | n34577 ;
  assign n34576 = n4445 & ~n10006 ;
  assign n34579 = n34578 ^ n34576 ^ 1'b0 ;
  assign n34580 = n25001 | n34579 ;
  assign n34581 = n3805 | n26415 ;
  assign n34582 = n15354 | n34581 ;
  assign n34583 = n4736 ^ n4695 ^ 1'b0 ;
  assign n34584 = n30502 ^ n11240 ^ n3154 ;
  assign n34585 = n3534 & ~n12772 ;
  assign n34586 = ~n13492 & n34585 ;
  assign n34587 = n8830 | n23544 ;
  assign n34588 = n16814 & n34587 ;
  assign n34589 = n16206 & n22901 ;
  assign n34590 = ~n3159 & n25630 ;
  assign n34591 = n7677 & n34590 ;
  assign n34592 = n19253 ^ n7509 ^ 1'b0 ;
  assign n34593 = n10750 & n34592 ;
  assign n34594 = n13962 & ~n19797 ;
  assign n34595 = n600 & n34594 ;
  assign n34596 = ~x232 & n26240 ;
  assign n34597 = n30007 | n34596 ;
  assign n34598 = n34597 ^ n21608 ^ n4476 ;
  assign n34599 = n6703 & ~n11119 ;
  assign n34600 = n31368 ^ n17869 ^ 1'b0 ;
  assign n34601 = n15993 & ~n34600 ;
  assign n34602 = n34601 ^ n31119 ^ 1'b0 ;
  assign n34603 = n8756 & ~n15000 ;
  assign n34604 = n9908 & n34603 ;
  assign n34605 = n7993 | n8665 ;
  assign n34606 = n11061 | n13182 ;
  assign n34607 = n34606 ^ n8950 ^ 1'b0 ;
  assign n34608 = n34607 ^ n4617 ^ 1'b0 ;
  assign n34609 = ~n34605 & n34608 ;
  assign n34610 = n1762 ^ n556 ^ 1'b0 ;
  assign n34611 = n9408 ^ n3756 ^ n1120 ;
  assign n34612 = n7431 | n22417 ;
  assign n34613 = n13109 ^ n10567 ^ 1'b0 ;
  assign n34614 = n34613 ^ n22616 ^ n21404 ;
  assign n34615 = n26746 ^ n12691 ^ 1'b0 ;
  assign n34616 = n34615 ^ n16627 ^ 1'b0 ;
  assign n34617 = n32556 & ~n34616 ;
  assign n34618 = n4475 ^ n1325 ^ 1'b0 ;
  assign n34619 = n23965 & ~n34618 ;
  assign n34620 = n34619 ^ n20514 ^ 1'b0 ;
  assign n34621 = ~n26818 & n34620 ;
  assign n34622 = n16326 | n20996 ;
  assign n34623 = n11758 & ~n13271 ;
  assign n34624 = n16705 ^ n1660 ^ 1'b0 ;
  assign n34627 = n1039 & n22621 ;
  assign n34625 = n24668 & n28770 ;
  assign n34626 = ~n20588 & n34625 ;
  assign n34628 = n34627 ^ n34626 ^ 1'b0 ;
  assign n34629 = ~n298 & n14131 ;
  assign n34630 = n8974 ^ n3718 ^ 1'b0 ;
  assign n34631 = n25977 ^ n11654 ^ n10844 ;
  assign n34634 = n16742 ^ n5801 ^ 1'b0 ;
  assign n34632 = n32931 ^ n28727 ^ 1'b0 ;
  assign n34633 = n11492 | n34632 ;
  assign n34635 = n34634 ^ n34633 ^ 1'b0 ;
  assign n34636 = n7498 & n27410 ;
  assign n34637 = n8087 & n34636 ;
  assign n34638 = n25185 & n34637 ;
  assign n34639 = n15907 & ~n16647 ;
  assign n34640 = n3614 & n34639 ;
  assign n34641 = ~n11191 & n14637 ;
  assign n34642 = ( n5297 & n18819 ) | ( n5297 & n29057 ) | ( n18819 & n29057 ) ;
  assign n34643 = n32921 ^ n29948 ^ 1'b0 ;
  assign n34644 = n23412 ^ n1158 ^ 1'b0 ;
  assign n34645 = n15589 ^ n6281 ^ 1'b0 ;
  assign n34646 = n22235 & n23425 ;
  assign n34647 = n34646 ^ n15489 ^ 1'b0 ;
  assign n34648 = n12132 & n13949 ;
  assign n34649 = n15908 & ~n20729 ;
  assign n34650 = n8773 ^ n482 ^ 1'b0 ;
  assign n34651 = n4810 & n34650 ;
  assign n34652 = n21595 & n34651 ;
  assign n34653 = ( ~n11675 & n12564 ) | ( ~n11675 & n34652 ) | ( n12564 & n34652 ) ;
  assign n34654 = ~n4063 & n16843 ;
  assign n34655 = n7716 & n34654 ;
  assign n34656 = n34655 ^ n4095 ^ 1'b0 ;
  assign n34657 = n12803 & n34656 ;
  assign n34658 = n19771 ^ n2078 ^ 1'b0 ;
  assign n34659 = x42 | n34658 ;
  assign n34660 = n5882 | n34659 ;
  assign n34661 = ~n24169 & n34660 ;
  assign n34662 = n9995 | n34568 ;
  assign n34663 = n34662 ^ n15487 ^ 1'b0 ;
  assign n34664 = n5833 & n34663 ;
  assign n34665 = n34661 & n34664 ;
  assign n34666 = n8919 ^ n2451 ^ 1'b0 ;
  assign n34667 = n6433 ^ n4328 ^ 1'b0 ;
  assign n34668 = n3304 & n11903 ;
  assign n34669 = n34668 ^ n18783 ^ 1'b0 ;
  assign n34670 = n23462 ^ n4718 ^ 1'b0 ;
  assign n34671 = ~n26776 & n34670 ;
  assign n34673 = n5597 & ~n10236 ;
  assign n34674 = ~n4719 & n34673 ;
  assign n34672 = n5504 | n5759 ;
  assign n34675 = n34674 ^ n34672 ^ 1'b0 ;
  assign n34676 = n7973 & n8324 ;
  assign n34677 = ~n1787 & n34676 ;
  assign n34678 = n12853 | n21404 ;
  assign n34679 = n34678 ^ n1727 ^ 1'b0 ;
  assign n34680 = n20528 ^ n9540 ^ 1'b0 ;
  assign n34681 = n34679 | n34680 ;
  assign n34682 = n34677 | n34681 ;
  assign n34683 = n31586 & n34682 ;
  assign n34685 = ~n2315 & n12855 ;
  assign n34686 = n34685 ^ n10111 ^ 1'b0 ;
  assign n34687 = ~n5135 & n34686 ;
  assign n34684 = ~x195 & n7920 ;
  assign n34688 = n34687 ^ n34684 ^ 1'b0 ;
  assign n34689 = n6494 & ~n21882 ;
  assign n34690 = n25036 ^ n5788 ^ 1'b0 ;
  assign n34691 = n33756 ^ n11744 ^ 1'b0 ;
  assign n34692 = ~n30913 & n34691 ;
  assign n34693 = n2568 & ~n34413 ;
  assign n34694 = n4549 & ~n34693 ;
  assign n34695 = n34694 ^ n34659 ^ 1'b0 ;
  assign n34696 = x237 & n30921 ;
  assign n34697 = n27103 ^ n19990 ^ n15179 ;
  assign n34698 = ~n6195 & n9836 ;
  assign n34699 = n34698 ^ n4853 ^ 1'b0 ;
  assign n34700 = n14000 & n34699 ;
  assign n34701 = n34700 ^ n21796 ^ 1'b0 ;
  assign n34702 = ~n22274 & n32899 ;
  assign n34703 = n28419 ^ n9778 ^ 1'b0 ;
  assign n34704 = n8215 ^ x144 ^ 1'b0 ;
  assign n34705 = n34703 & n34704 ;
  assign n34706 = n34705 ^ n21416 ^ n3451 ;
  assign n34707 = x221 & ~n3750 ;
  assign n34708 = n4076 & ~n12511 ;
  assign n34709 = n13473 & n34708 ;
  assign n34710 = ~n6337 & n28932 ;
  assign n34711 = n3184 & n26666 ;
  assign n34712 = ~n2391 & n10328 ;
  assign n34713 = n14300 & ~n24150 ;
  assign n34714 = n34712 & n34713 ;
  assign n34715 = ~n1851 & n9587 ;
  assign n34716 = n4731 & n34715 ;
  assign n34717 = n34716 ^ n27869 ^ 1'b0 ;
  assign n34718 = n10613 & n30871 ;
  assign n34719 = n7021 ^ n5484 ^ 1'b0 ;
  assign n34720 = n1851 | n34719 ;
  assign n34721 = n2689 & ~n34720 ;
  assign n34722 = n12790 ^ n5639 ^ 1'b0 ;
  assign n34723 = n34722 ^ n18754 ^ 1'b0 ;
  assign n34724 = n11207 | n13414 ;
  assign n34725 = n10346 | n34724 ;
  assign n34726 = n15035 ^ n11829 ^ 1'b0 ;
  assign n34727 = n17672 | n34726 ;
  assign n34728 = n5426 & ~n34727 ;
  assign n34729 = ~n6311 & n12448 ;
  assign n34732 = n15314 | n16346 ;
  assign n34733 = n3358 | n34732 ;
  assign n34730 = n2185 | n20961 ;
  assign n34731 = n20601 & ~n34730 ;
  assign n34734 = n34733 ^ n34731 ^ n956 ;
  assign n34735 = n6706 & ~n23932 ;
  assign n34736 = n1075 & n3608 ;
  assign n34737 = n19098 & n34736 ;
  assign n34738 = n8821 ^ n3820 ^ 1'b0 ;
  assign n34739 = ~n5207 & n34738 ;
  assign n34740 = n9661 & n34739 ;
  assign n34741 = n3906 & n34740 ;
  assign n34742 = n13561 & ~n34741 ;
  assign n34743 = n34742 ^ n28011 ^ 1'b0 ;
  assign n34744 = n3062 & n15241 ;
  assign n34745 = n8354 ^ n6729 ^ 1'b0 ;
  assign n34746 = n2153 & ~n20211 ;
  assign n34747 = n34746 ^ n18746 ^ 1'b0 ;
  assign n34748 = n14043 ^ n3310 ^ 1'b0 ;
  assign n34749 = ~n31146 & n34748 ;
  assign n34750 = n3568 | n34749 ;
  assign n34751 = n3563 & n34750 ;
  assign n34752 = n19570 ^ n6712 ^ 1'b0 ;
  assign n34753 = n1255 & ~n22977 ;
  assign n34754 = n34753 ^ n9097 ^ 1'b0 ;
  assign n34755 = n7032 | n19915 ;
  assign n34756 = n34755 ^ n28282 ^ 1'b0 ;
  assign n34757 = ~n3963 & n34756 ;
  assign n34758 = n34757 ^ n19996 ^ 1'b0 ;
  assign n34759 = n32462 ^ n8291 ^ 1'b0 ;
  assign n34760 = n26841 & n34759 ;
  assign n34761 = n34758 & n34760 ;
  assign n34762 = n9431 ^ n417 ^ 1'b0 ;
  assign n34763 = ~n6149 & n34762 ;
  assign n34764 = n34194 ^ n16671 ^ 1'b0 ;
  assign n34765 = n34763 & ~n34764 ;
  assign n34766 = n1562 | n24924 ;
  assign n34767 = n23279 & ~n34766 ;
  assign n34768 = n21041 & ~n27781 ;
  assign n34769 = n7406 & ~n31801 ;
  assign n34770 = n11865 ^ n4747 ^ 1'b0 ;
  assign n34771 = n26985 & n34770 ;
  assign n34772 = n4904 & ~n30848 ;
  assign n34773 = n29498 & n34772 ;
  assign n34774 = n22830 ^ n8804 ^ 1'b0 ;
  assign n34775 = n5506 | n34774 ;
  assign n34776 = ~x154 & n34775 ;
  assign n34777 = n14501 ^ n3667 ^ 1'b0 ;
  assign n34778 = n22305 | n34777 ;
  assign n34779 = ( x200 & n25094 ) | ( x200 & ~n32970 ) | ( n25094 & ~n32970 ) ;
  assign n34780 = n21867 & ~n32900 ;
  assign n34781 = n34780 ^ n11582 ^ 1'b0 ;
  assign n34782 = x94 & ~n9497 ;
  assign n34783 = n34782 ^ n10278 ^ 1'b0 ;
  assign n34784 = n10157 ^ n1291 ^ 1'b0 ;
  assign n34785 = n6288 & n34784 ;
  assign n34786 = ~n1071 & n30677 ;
  assign n34787 = ~n2227 & n34786 ;
  assign n34788 = n17226 ^ n421 ^ 1'b0 ;
  assign n34789 = n17270 ^ n14299 ^ 1'b0 ;
  assign n34790 = ( ~n614 & n667 ) | ( ~n614 & n6976 ) | ( n667 & n6976 ) ;
  assign n34791 = n29265 & n34790 ;
  assign n34792 = ~n34789 & n34791 ;
  assign n34793 = n17680 ^ n355 ^ 1'b0 ;
  assign n34794 = n3670 & ~n34793 ;
  assign n34795 = ~n10526 & n34794 ;
  assign n34796 = ~x210 & n34795 ;
  assign n34797 = n18864 | n25467 ;
  assign n34798 = n8718 ^ n1818 ^ 1'b0 ;
  assign n34799 = ( n663 & ~n8118 ) | ( n663 & n30071 ) | ( ~n8118 & n30071 ) ;
  assign n34800 = x47 & n9988 ;
  assign n34801 = ~n32327 & n34800 ;
  assign n34802 = n5991 | n6487 ;
  assign n34803 = n13775 & n14466 ;
  assign n34805 = ~x52 & n9240 ;
  assign n34804 = n3641 | n29106 ;
  assign n34806 = n34805 ^ n34804 ^ 1'b0 ;
  assign n34807 = n832 & ~n14830 ;
  assign n34808 = n2445 & n34807 ;
  assign n34809 = n4201 | n34808 ;
  assign n34810 = n34809 ^ n6032 ^ 1'b0 ;
  assign n34811 = n32404 ^ n5754 ^ 1'b0 ;
  assign n34812 = n502 | n3540 ;
  assign n34813 = n6737 ^ x198 ^ 1'b0 ;
  assign n34814 = ~n28835 & n34813 ;
  assign n34815 = n25365 ^ n1216 ^ 1'b0 ;
  assign n34816 = x3 & n10302 ;
  assign n34817 = n3216 | n13324 ;
  assign n34818 = n34816 | n34817 ;
  assign n34819 = n30911 ^ n7696 ^ 1'b0 ;
  assign n34820 = n15061 & ~n34819 ;
  assign n34821 = n34820 ^ n5023 ^ 1'b0 ;
  assign n34822 = n32251 & n34821 ;
  assign n34823 = n4333 ^ n3988 ^ 1'b0 ;
  assign n34824 = n15298 & n34823 ;
  assign n34825 = n6693 & n33830 ;
  assign n34826 = n34825 ^ n17966 ^ 1'b0 ;
  assign n34827 = ~n18877 & n34579 ;
  assign n34828 = n34827 ^ n9638 ^ 1'b0 ;
  assign n34829 = ~n3412 & n8193 ;
  assign n34830 = n34829 ^ n8016 ^ 1'b0 ;
  assign n34831 = n23754 ^ n20468 ^ 1'b0 ;
  assign n34832 = ~n34830 & n34831 ;
  assign n34833 = n2465 ^ n1847 ^ 1'b0 ;
  assign n34834 = n34832 & ~n34833 ;
  assign n34835 = n13395 & n13412 ;
  assign n34836 = n33314 & n34835 ;
  assign n34837 = n34836 ^ n18625 ^ 1'b0 ;
  assign n34838 = n34837 ^ n31796 ^ 1'b0 ;
  assign n34839 = n15724 & ~n33161 ;
  assign n34840 = n14815 & n34839 ;
  assign n34841 = n5984 | n16062 ;
  assign n34842 = n13926 | n34841 ;
  assign n34843 = n11276 | n32301 ;
  assign n34844 = n34843 ^ n28312 ^ 1'b0 ;
  assign n34846 = n3333 & n4719 ;
  assign n34847 = n34846 ^ n3966 ^ 1'b0 ;
  assign n34845 = ~n1064 & n17383 ;
  assign n34848 = n34847 ^ n34845 ^ 1'b0 ;
  assign n34850 = x226 | n27156 ;
  assign n34849 = n354 & n8383 ;
  assign n34851 = n34850 ^ n34849 ^ 1'b0 ;
  assign n34852 = n587 & ~n2744 ;
  assign n34853 = n24138 ^ x153 ^ 1'b0 ;
  assign n34854 = n16456 ^ n4655 ^ 1'b0 ;
  assign n34855 = n34854 ^ n6592 ^ 1'b0 ;
  assign n34856 = n18047 | n34855 ;
  assign n34857 = x89 & n12790 ;
  assign n34858 = n34857 ^ n7703 ^ 1'b0 ;
  assign n34859 = n5368 | n33018 ;
  assign n34860 = n13972 & n34859 ;
  assign n34861 = ~n6118 & n17046 ;
  assign n34862 = n34861 ^ n17009 ^ 1'b0 ;
  assign n34863 = n24095 ^ n8381 ^ 1'b0 ;
  assign n34864 = n22073 & ~n34863 ;
  assign n34865 = n34864 ^ n21346 ^ 1'b0 ;
  assign n34866 = n4530 & n9874 ;
  assign n34867 = n7668 & ~n14117 ;
  assign n34868 = n9616 ^ n6431 ^ 1'b0 ;
  assign n34869 = ~n2929 & n34868 ;
  assign n34870 = ~n589 & n5177 ;
  assign n34871 = ~n34869 & n34870 ;
  assign n34872 = n34867 & n34871 ;
  assign n34876 = n553 | n2853 ;
  assign n34877 = n34876 ^ n3153 ^ 1'b0 ;
  assign n34873 = ~n788 & n2107 ;
  assign n34874 = n18877 & n34873 ;
  assign n34875 = n26080 | n34874 ;
  assign n34878 = n34877 ^ n34875 ^ 1'b0 ;
  assign n34879 = ~n395 & n10206 ;
  assign n34880 = n31883 & ~n34879 ;
  assign n34881 = n34880 ^ n33824 ^ 1'b0 ;
  assign n34882 = n12570 | n23489 ;
  assign n34883 = n1360 & ~n22573 ;
  assign n34884 = n2744 & ~n14445 ;
  assign n34885 = ~n34883 & n34884 ;
  assign n34886 = n3531 & ~n31423 ;
  assign n34887 = n16001 ^ n14809 ^ 1'b0 ;
  assign n34888 = n16312 ^ n10239 ^ 1'b0 ;
  assign n34889 = n8772 ^ n6799 ^ 1'b0 ;
  assign n34890 = n20565 & n34889 ;
  assign n34891 = ~n15362 & n19719 ;
  assign n34892 = n34891 ^ n13348 ^ 1'b0 ;
  assign n34893 = ( ~n5382 & n15106 ) | ( ~n5382 & n34892 ) | ( n15106 & n34892 ) ;
  assign n34894 = n3984 & n26658 ;
  assign n34895 = n1524 & ~n28113 ;
  assign n34896 = n1901 & ~n12405 ;
  assign n34897 = n8115 ^ n2249 ^ 1'b0 ;
  assign n34898 = n34896 | n34897 ;
  assign n34899 = n12888 & n34898 ;
  assign n34900 = n1578 & ~n33269 ;
  assign n34901 = n34900 ^ n22055 ^ 1'b0 ;
  assign n34902 = n1345 & n12441 ;
  assign n34903 = ~n9688 & n34902 ;
  assign n34904 = n30947 | n34903 ;
  assign n34905 = n1079 | n23677 ;
  assign n34906 = n34904 & ~n34905 ;
  assign n34907 = n6191 | n8242 ;
  assign n34908 = n34393 & ~n34907 ;
  assign n34909 = n31392 ^ n5283 ^ 1'b0 ;
  assign n34910 = n11712 ^ n6866 ^ 1'b0 ;
  assign n34911 = n5791 | n18784 ;
  assign n34912 = n10918 & ~n34911 ;
  assign n34913 = ~n6375 & n18311 ;
  assign n34914 = n8112 & n34913 ;
  assign n34915 = n16229 & ~n34914 ;
  assign n34916 = n34912 & n34915 ;
  assign n34917 = n623 & n1847 ;
  assign n34918 = ~n1847 & n34917 ;
  assign n34919 = ( ~n8637 & n34620 ) | ( ~n8637 & n34918 ) | ( n34620 & n34918 ) ;
  assign n34920 = n13358 & n34919 ;
  assign n34921 = n5481 & n34920 ;
  assign n34922 = n19235 ^ n13742 ^ 1'b0 ;
  assign n34923 = n24936 | n34922 ;
  assign n34924 = n34923 ^ n7968 ^ 1'b0 ;
  assign n34925 = n22970 | n24653 ;
  assign n34926 = n23510 & ~n34925 ;
  assign n34927 = n34237 & n34304 ;
  assign n34928 = n8767 & n10650 ;
  assign n34929 = ~n1499 & n34928 ;
  assign n34930 = n1239 | n20841 ;
  assign n34931 = n3725 & ~n34930 ;
  assign n34932 = n34931 ^ n20272 ^ 1'b0 ;
  assign n34933 = n3356 & n10403 ;
  assign n34934 = n34933 ^ n9319 ^ 1'b0 ;
  assign n34935 = n5859 & n34934 ;
  assign n34936 = n8384 | n34935 ;
  assign n34937 = n34936 ^ n27460 ^ 1'b0 ;
  assign n34938 = n30581 ^ n5323 ^ 1'b0 ;
  assign n34939 = n5529 & n26944 ;
  assign n34940 = n34939 ^ n8693 ^ 1'b0 ;
  assign n34942 = n6554 & ~n16982 ;
  assign n34941 = ~n1361 & n13172 ;
  assign n34943 = n34942 ^ n34941 ^ 1'b0 ;
  assign n34944 = ~n4955 & n17182 ;
  assign n34945 = n34944 ^ n2417 ^ 1'b0 ;
  assign n34946 = n11517 & n34945 ;
  assign n34947 = n34946 ^ n1207 ^ 1'b0 ;
  assign n34948 = ~x204 & n1546 ;
  assign n34949 = n27069 ^ n11294 ^ 1'b0 ;
  assign n34950 = x3 & n34949 ;
  assign n34951 = ~n34745 & n34950 ;
  assign n34952 = ~n14272 & n34951 ;
  assign n34954 = n2846 & n5198 ;
  assign n34953 = n1733 | n31856 ;
  assign n34955 = n34954 ^ n34953 ^ 1'b0 ;
  assign n34956 = n16709 ^ n1286 ^ 1'b0 ;
  assign n34957 = n16712 & ~n34956 ;
  assign n34958 = n9946 & ~n34957 ;
  assign n34959 = n10740 ^ n6305 ^ 1'b0 ;
  assign n34961 = n22055 ^ n18072 ^ 1'b0 ;
  assign n34962 = n23266 | n34961 ;
  assign n34963 = ~n13778 & n34962 ;
  assign n34960 = n444 & ~n31191 ;
  assign n34964 = n34963 ^ n34960 ^ 1'b0 ;
  assign n34965 = n24464 | n32603 ;
  assign n34966 = n2034 & ~n34965 ;
  assign n34967 = n3740 | n18273 ;
  assign n34968 = n8935 ^ n8873 ^ n1926 ;
  assign n34969 = n4116 & n4188 ;
  assign n34970 = ( n3095 & ~n31521 ) | ( n3095 & n34969 ) | ( ~n31521 & n34969 ) ;
  assign n34972 = n4075 & n8293 ;
  assign n34971 = ~n4075 & n12080 ;
  assign n34973 = n34972 ^ n34971 ^ 1'b0 ;
  assign n34974 = n1383 | n3169 ;
  assign n34975 = n11749 | n34974 ;
  assign n34976 = n5085 & ~n34975 ;
  assign n34977 = n6484 | n18254 ;
  assign n34978 = n32074 ^ n19285 ^ 1'b0 ;
  assign n34979 = n14929 | n34978 ;
  assign n34980 = ~n12250 & n18508 ;
  assign n34981 = n8258 & ~n28286 ;
  assign n34982 = n8919 & n34981 ;
  assign n34983 = n21182 ^ n11339 ^ 1'b0 ;
  assign n34984 = n1277 & n23076 ;
  assign n34985 = n5828 ^ n1974 ^ 1'b0 ;
  assign n34986 = ~n32830 & n34985 ;
  assign n34988 = n3287 & n13821 ;
  assign n34989 = n842 & n34988 ;
  assign n34990 = n9387 & ~n27711 ;
  assign n34991 = n34989 & n34990 ;
  assign n34987 = n8148 & ~n9076 ;
  assign n34992 = n34991 ^ n34987 ^ 1'b0 ;
  assign n34994 = n956 & n9108 ;
  assign n34993 = n1141 | n5207 ;
  assign n34995 = n34994 ^ n34993 ^ 1'b0 ;
  assign n34996 = n6222 & n22174 ;
  assign n34997 = n15179 | n34996 ;
  assign n34998 = ~n34995 & n34997 ;
  assign n34999 = n20474 | n28407 ;
  assign n35000 = n34999 ^ n6791 ^ 1'b0 ;
  assign n35001 = ~n25758 & n35000 ;
  assign n35002 = n11150 ^ n2165 ^ 1'b0 ;
  assign n35003 = n30482 & ~n35002 ;
  assign n35004 = n9083 | n18241 ;
  assign n35005 = n3414 & ~n35004 ;
  assign n35006 = ~n5072 & n7749 ;
  assign n35007 = n21398 ^ n9907 ^ 1'b0 ;
  assign n35008 = n6362 | n35007 ;
  assign n35009 = ~n3114 & n34722 ;
  assign n35010 = ( n2673 & n24653 ) | ( n2673 & n35009 ) | ( n24653 & n35009 ) ;
  assign n35011 = n2443 | n34197 ;
  assign n35012 = n35011 ^ n13593 ^ 1'b0 ;
  assign n35013 = ~n7128 & n13627 ;
  assign n35014 = n35013 ^ n28210 ^ n5978 ;
  assign n35015 = n9835 | n35014 ;
  assign n35016 = n29037 ^ n2315 ^ 1'b0 ;
  assign n35017 = ~n3125 & n9560 ;
  assign n35018 = n20624 & n35017 ;
  assign n35019 = n35018 ^ n6558 ^ 1'b0 ;
  assign n35020 = ~n16591 & n35019 ;
  assign n35021 = n2301 | n3024 ;
  assign n35022 = n35021 ^ n9341 ^ 1'b0 ;
  assign n35023 = ( ~x25 & n6523 ) | ( ~x25 & n14845 ) | ( n6523 & n14845 ) ;
  assign n35024 = ~n1638 & n3573 ;
  assign n35025 = n35024 ^ x76 ^ 1'b0 ;
  assign n35026 = n1146 | n7133 ;
  assign n35027 = n35026 ^ n19275 ^ 1'b0 ;
  assign n35028 = ~n11266 & n35027 ;
  assign n35029 = n1239 & n5435 ;
  assign n35030 = ~n4699 & n35029 ;
  assign n35031 = ~n12845 & n35030 ;
  assign n35032 = n18296 & n35031 ;
  assign n35033 = n3794 & ~n15510 ;
  assign n35034 = n708 & n22323 ;
  assign n35035 = n35034 ^ n18128 ^ 1'b0 ;
  assign n35036 = n23130 & ~n35035 ;
  assign n35037 = n35036 ^ n15481 ^ 1'b0 ;
  assign n35038 = ~n3915 & n11596 ;
  assign n35039 = n28831 ^ n8990 ^ 1'b0 ;
  assign n35040 = n4118 & ~n35039 ;
  assign n35041 = n2371 & n35040 ;
  assign n35042 = n21240 ^ n19613 ^ 1'b0 ;
  assign n35043 = n14244 & ~n35042 ;
  assign n35044 = n6942 & n23697 ;
  assign n35045 = n27220 ^ x170 ^ 1'b0 ;
  assign n35046 = n12022 | n35045 ;
  assign n35047 = n2310 & n24574 ;
  assign n35048 = n35047 ^ n33543 ^ 1'b0 ;
  assign n35049 = n5704 & ~n32640 ;
  assign n35050 = n18788 | n28800 ;
  assign n35051 = n14236 ^ x182 ^ 1'b0 ;
  assign n35052 = ~n12811 & n35051 ;
  assign n35054 = ~n3685 & n5872 ;
  assign n35055 = ~n5097 & n35054 ;
  assign n35053 = ~n8091 & n10708 ;
  assign n35056 = n35055 ^ n35053 ^ 1'b0 ;
  assign n35057 = ~n4824 & n7842 ;
  assign n35058 = n35057 ^ n25896 ^ 1'b0 ;
  assign n35059 = n10774 | n35058 ;
  assign n35060 = n12526 & n21338 ;
  assign n35061 = n35060 ^ n21387 ^ 1'b0 ;
  assign n35062 = ~n1487 & n23852 ;
  assign n35063 = n35062 ^ n22292 ^ 1'b0 ;
  assign n35064 = n16689 ^ n15033 ^ n10030 ;
  assign n35065 = n35063 & n35064 ;
  assign n35066 = ( n4783 & n4806 ) | ( n4783 & ~n10310 ) | ( n4806 & ~n10310 ) ;
  assign n35067 = n22035 & ~n35066 ;
  assign n35068 = n35067 ^ n5027 ^ 1'b0 ;
  assign n35069 = n35068 ^ n23315 ^ n1236 ;
  assign n35071 = n6191 ^ n1557 ^ 1'b0 ;
  assign n35072 = ~n1291 & n35071 ;
  assign n35070 = ~n11632 & n11669 ;
  assign n35073 = n35072 ^ n35070 ^ 1'b0 ;
  assign n35074 = ~n2143 & n17182 ;
  assign n35075 = n35074 ^ n8137 ^ 1'b0 ;
  assign n35076 = n35073 | n35075 ;
  assign n35077 = ~n2711 & n13155 ;
  assign n35078 = n35077 ^ n8948 ^ 1'b0 ;
  assign n35079 = n12604 & ~n12903 ;
  assign n35080 = n2267 ^ n1028 ^ 1'b0 ;
  assign n35081 = n35079 & n35080 ;
  assign n35082 = n35081 ^ n31461 ^ 1'b0 ;
  assign n35083 = n1444 & n16221 ;
  assign n35084 = n5742 ^ n2655 ^ 1'b0 ;
  assign n35085 = n1725 | n35084 ;
  assign n35086 = n13538 | n17367 ;
  assign n35087 = n13084 & ~n24730 ;
  assign n35088 = n35086 & n35087 ;
  assign n35089 = n1266 ^ n623 ^ 1'b0 ;
  assign n35090 = ~n19684 & n35089 ;
  assign n35091 = n5170 & n35090 ;
  assign n35092 = n4402 & ~n29437 ;
  assign n35093 = ~n18038 & n21034 ;
  assign n35094 = n35093 ^ n15191 ^ 1'b0 ;
  assign n35095 = n4061 & ~n25940 ;
  assign n35096 = n35095 ^ n25350 ^ 1'b0 ;
  assign n35097 = n28206 ^ n3820 ^ 1'b0 ;
  assign n35098 = n19191 ^ n1815 ^ 1'b0 ;
  assign n35099 = n17480 & ~n35098 ;
  assign n35100 = n3184 & n18553 ;
  assign n35101 = n571 & ~n2223 ;
  assign n35102 = ~n7137 & n33580 ;
  assign n35103 = n6220 | n35102 ;
  assign n35104 = n35103 ^ n23297 ^ 1'b0 ;
  assign n35105 = n30941 ^ n4784 ^ 1'b0 ;
  assign n35107 = n1044 & ~n4358 ;
  assign n35108 = n35107 ^ n14061 ^ 1'b0 ;
  assign n35106 = n6940 | n21796 ;
  assign n35109 = n35108 ^ n35106 ^ 1'b0 ;
  assign n35110 = n35109 ^ n7993 ^ 1'b0 ;
  assign n35111 = n7578 | n8674 ;
  assign n35112 = n35111 ^ n16043 ^ 1'b0 ;
  assign n35113 = n6012 & n16364 ;
  assign n35114 = n21022 ^ n9592 ^ 1'b0 ;
  assign n35115 = n35113 & ~n35114 ;
  assign n35116 = n35115 ^ n11673 ^ 1'b0 ;
  assign n35117 = n7457 & n35116 ;
  assign n35118 = x28 | n6702 ;
  assign n35119 = n1743 ^ n1111 ^ 1'b0 ;
  assign n35120 = n22710 & n35119 ;
  assign n35121 = ~n35118 & n35120 ;
  assign n35122 = n14197 ^ n8004 ^ 1'b0 ;
  assign n35123 = n3166 & n35122 ;
  assign n35124 = n35123 ^ n32981 ^ 1'b0 ;
  assign n35125 = n553 & n2593 ;
  assign n35126 = n35125 ^ n2715 ^ 1'b0 ;
  assign n35127 = ~n35124 & n35126 ;
  assign n35128 = n2110 | n21708 ;
  assign n35129 = n14910 | n17290 ;
  assign n35134 = n12906 | n20926 ;
  assign n35135 = n7133 | n35134 ;
  assign n35130 = n8033 ^ n5348 ^ 1'b0 ;
  assign n35131 = n1814 & n35130 ;
  assign n35132 = n35131 ^ n19435 ^ 1'b0 ;
  assign n35133 = n8628 & n35132 ;
  assign n35136 = n35135 ^ n35133 ^ 1'b0 ;
  assign n35137 = n24658 & ~n35136 ;
  assign n35138 = n12260 ^ n11851 ^ 1'b0 ;
  assign n35139 = n22141 | n35138 ;
  assign n35140 = ~n614 & n8750 ;
  assign n35141 = n860 & n28962 ;
  assign n35142 = n35140 & n35141 ;
  assign n35143 = n15600 & ~n35142 ;
  assign n35144 = n35143 ^ n11072 ^ 1'b0 ;
  assign n35145 = ~n3540 & n29569 ;
  assign n35146 = n23852 & n30801 ;
  assign n35147 = ~n9860 & n24261 ;
  assign n35148 = x226 & n35147 ;
  assign n35149 = n22207 ^ n5366 ^ 1'b0 ;
  assign n35150 = ~n16813 & n29066 ;
  assign n35151 = n35150 ^ n19279 ^ 1'b0 ;
  assign n35152 = n1117 & ~n35151 ;
  assign n35153 = n8417 ^ n7594 ^ 1'b0 ;
  assign n35154 = n5835 & ~n35153 ;
  assign n35155 = n11004 & n16075 ;
  assign n35156 = n9122 ^ n5999 ^ 1'b0 ;
  assign n35157 = n21999 ^ n15197 ^ 1'b0 ;
  assign n35158 = n35156 | n35157 ;
  assign n35160 = n12990 ^ n8752 ^ 1'b0 ;
  assign n35161 = n9651 & n35160 ;
  assign n35159 = n27364 & ~n27529 ;
  assign n35162 = n35161 ^ n35159 ^ 1'b0 ;
  assign n35163 = n26836 & ~n35162 ;
  assign n35164 = n23859 ^ n13717 ^ 1'b0 ;
  assign n35165 = n6590 & n35164 ;
  assign n35166 = n14163 & ~n35165 ;
  assign n35167 = n32708 ^ n7680 ^ 1'b0 ;
  assign n35168 = n3750 & n10345 ;
  assign n35169 = ~n4223 & n12232 ;
  assign n35170 = n35169 ^ n2248 ^ 1'b0 ;
  assign n35174 = ~n13453 & n26304 ;
  assign n35171 = n14076 | n21822 ;
  assign n35172 = n26921 | n35171 ;
  assign n35173 = ~n7674 & n35172 ;
  assign n35175 = n35174 ^ n35173 ^ 1'b0 ;
  assign n35176 = ( n6432 & ~n7310 ) | ( n6432 & n18084 ) | ( ~n7310 & n18084 ) ;
  assign n35177 = n21771 ^ n19998 ^ 1'b0 ;
  assign n35178 = n3003 & n7361 ;
  assign n35179 = n28172 ^ n6398 ^ 1'b0 ;
  assign n35180 = n35178 | n35179 ;
  assign n35181 = n26400 ^ n1073 ^ 1'b0 ;
  assign n35182 = ~n17169 & n35181 ;
  assign n35183 = n35182 ^ n23856 ^ 1'b0 ;
  assign n35184 = n15295 | n25247 ;
  assign n35185 = n11589 | n35184 ;
  assign n35186 = n3424 | n11612 ;
  assign n35187 = n7434 & ~n13042 ;
  assign n35188 = n651 & ~n6050 ;
  assign n35189 = n7028 & n35188 ;
  assign n35190 = n34660 | n35189 ;
  assign n35191 = ~n11661 & n13943 ;
  assign n35192 = ~n20788 & n35191 ;
  assign n35193 = ~n26250 & n35192 ;
  assign n35194 = n27717 ^ n3974 ^ 1'b0 ;
  assign n35195 = n7595 & n25995 ;
  assign n35196 = ~n19041 & n35195 ;
  assign n35197 = n12974 & ~n35196 ;
  assign n35198 = n7648 & n35197 ;
  assign n35199 = n1646 | n5826 ;
  assign n35200 = n7650 & ~n35199 ;
  assign n35201 = n6850 ^ n1775 ^ 1'b0 ;
  assign n35202 = n22944 & n35201 ;
  assign n35203 = n35202 ^ n15242 ^ 1'b0 ;
  assign n35204 = ~n1651 & n3743 ;
  assign n35205 = ~n30742 & n34312 ;
  assign n35206 = n8217 & n11371 ;
  assign n35207 = ~n35205 & n35206 ;
  assign n35208 = ~n3229 & n30769 ;
  assign n35209 = x27 & n35208 ;
  assign n35210 = n11426 & n14803 ;
  assign n35211 = n14554 & n35210 ;
  assign n35212 = n8218 | n26054 ;
  assign n35213 = n35211 & ~n35212 ;
  assign n35214 = n29236 ^ n13496 ^ 1'b0 ;
  assign n35215 = ~n35213 & n35214 ;
  assign n35216 = n6344 & ~n13742 ;
  assign n35217 = n19438 & n35216 ;
  assign n35218 = n4047 ^ n590 ^ 1'b0 ;
  assign n35219 = ~n35217 & n35218 ;
  assign n35220 = ~n19968 & n35219 ;
  assign n35221 = n9660 | n20496 ;
  assign n35222 = n11322 | n24821 ;
  assign n35223 = n553 & ~n35222 ;
  assign n35224 = n3837 & n18464 ;
  assign n35225 = n35224 ^ n22035 ^ 1'b0 ;
  assign n35226 = n12048 | n21168 ;
  assign n35227 = n2185 | n35226 ;
  assign n35228 = n33116 ^ n3062 ^ 1'b0 ;
  assign n35229 = n22379 ^ n13996 ^ n5138 ;
  assign n35230 = n7361 ^ n5904 ^ 1'b0 ;
  assign n35231 = n12093 | n35230 ;
  assign n35232 = n16337 ^ n10433 ^ 1'b0 ;
  assign n35233 = n4636 | n18783 ;
  assign n35234 = n16347 ^ n4703 ^ 1'b0 ;
  assign n35235 = n1964 | n35234 ;
  assign n35236 = n8628 ^ n5767 ^ 1'b0 ;
  assign n35237 = n2517 & ~n6048 ;
  assign n35238 = ~n35236 & n35237 ;
  assign n35239 = n1736 & ~n6245 ;
  assign n35240 = n35239 ^ n20387 ^ 1'b0 ;
  assign n35241 = n11400 ^ n6189 ^ 1'b0 ;
  assign n35242 = n644 & ~n35241 ;
  assign n35243 = n2358 & ~n35242 ;
  assign n35244 = n6532 & ~n35243 ;
  assign n35245 = n35244 ^ n4953 ^ 1'b0 ;
  assign n35246 = n6792 ^ n1697 ^ 1'b0 ;
  assign n35247 = n10571 ^ x33 ^ 1'b0 ;
  assign n35248 = n8693 & ~n10593 ;
  assign n35249 = n26309 & n31522 ;
  assign n35250 = n35249 ^ n30843 ^ 1'b0 ;
  assign n35251 = n12023 | n29079 ;
  assign n35252 = n6372 & ~n12713 ;
  assign n35253 = ~n16074 & n35252 ;
  assign n35254 = n10094 | n14431 ;
  assign n35255 = n4376 | n35254 ;
  assign n35256 = n12772 ^ n4711 ^ 1'b0 ;
  assign n35257 = ~n2098 & n35256 ;
  assign n35258 = n4826 & ~n15019 ;
  assign n35259 = n35258 ^ n3267 ^ 1'b0 ;
  assign n35260 = n2681 & n35259 ;
  assign n35261 = n35257 & ~n35260 ;
  assign n35262 = n17429 ^ n6461 ^ 1'b0 ;
  assign n35263 = n1656 | n7473 ;
  assign n35264 = n1656 & ~n35263 ;
  assign n35265 = n35264 ^ n10140 ^ 1'b0 ;
  assign n35266 = ~n35262 & n35265 ;
  assign n35267 = n35266 ^ n19212 ^ 1'b0 ;
  assign n35268 = n16749 ^ n10152 ^ 1'b0 ;
  assign n35269 = x245 | n35268 ;
  assign n35270 = n20411 & ~n35269 ;
  assign n35271 = n3791 & ~n4523 ;
  assign n35272 = n35271 ^ n22925 ^ n15167 ;
  assign n35273 = n18232 & n35272 ;
  assign n35274 = ~n3213 & n9011 ;
  assign n35275 = n9225 & ~n35274 ;
  assign n35276 = n4227 & ~n19547 ;
  assign n35277 = ~n7508 & n35276 ;
  assign n35278 = n7882 | n35277 ;
  assign n35279 = n33605 | n35278 ;
  assign n35280 = ~n17073 & n23076 ;
  assign n35281 = n35280 ^ n623 ^ 1'b0 ;
  assign n35282 = n14498 ^ n4128 ^ 1'b0 ;
  assign n35283 = n6149 | n6962 ;
  assign n35284 = n10629 | n35283 ;
  assign n35285 = n35284 ^ n20721 ^ 1'b0 ;
  assign n35286 = n22467 ^ n5869 ^ 1'b0 ;
  assign n35287 = ~n7124 & n35286 ;
  assign n35288 = n35287 ^ x220 ^ 1'b0 ;
  assign n35289 = ~n20926 & n35288 ;
  assign n35290 = n35289 ^ n5860 ^ 1'b0 ;
  assign n35291 = n3441 & ~n15517 ;
  assign n35292 = n4901 & ~n19521 ;
  assign n35293 = n22161 & n35292 ;
  assign n35294 = n4870 | n35293 ;
  assign n35295 = n15743 & n15947 ;
  assign n35296 = n35295 ^ n15627 ^ 1'b0 ;
  assign n35297 = n35296 ^ n8150 ^ 1'b0 ;
  assign n35298 = n13800 & ~n15094 ;
  assign n35299 = n23026 & n35298 ;
  assign n35300 = n35299 ^ n7908 ^ 1'b0 ;
  assign n35301 = n32789 ^ n22820 ^ 1'b0 ;
  assign n35302 = n5027 & ~n35301 ;
  assign n35303 = n8082 | n9106 ;
  assign n35304 = n35302 & ~n35303 ;
  assign n35305 = ~n14933 & n20996 ;
  assign n35306 = n6489 & n23582 ;
  assign n35308 = n4068 & ~n18329 ;
  assign n35309 = n35308 ^ n3102 ^ 1'b0 ;
  assign n35307 = n10575 & ~n13001 ;
  assign n35310 = n35309 ^ n35307 ^ 1'b0 ;
  assign n35311 = ~n17495 & n35310 ;
  assign n35312 = n35311 ^ n15593 ^ 1'b0 ;
  assign n35313 = n35312 ^ n3308 ^ 1'b0 ;
  assign n35314 = n9557 & ~n19438 ;
  assign n35315 = n3009 & ~n31184 ;
  assign n35316 = ~n28234 & n35315 ;
  assign n35317 = n2333 | n28434 ;
  assign n35318 = n25861 & ~n35317 ;
  assign n35319 = n31312 ^ n20988 ^ 1'b0 ;
  assign n35320 = n35319 ^ n21025 ^ 1'b0 ;
  assign n35321 = x160 & ~n4122 ;
  assign n35322 = n5272 & ~n11267 ;
  assign n35323 = ( n18944 & ~n35321 ) | ( n18944 & n35322 ) | ( ~n35321 & n35322 ) ;
  assign n35324 = n16439 ^ n6458 ^ 1'b0 ;
  assign n35325 = n17056 ^ n10997 ^ n4241 ;
  assign n35326 = n8089 & n35325 ;
  assign n35327 = n1641 & ~n1758 ;
  assign n35328 = ~n12748 & n35327 ;
  assign n35329 = n35328 ^ n30602 ^ 1'b0 ;
  assign n35330 = n35326 & ~n35329 ;
  assign n35331 = n3800 & n35330 ;
  assign n35332 = n35331 ^ n6817 ^ 1'b0 ;
  assign n35333 = n23006 | n35332 ;
  assign n35334 = n35333 ^ n12417 ^ 1'b0 ;
  assign n35335 = n7162 ^ n3661 ^ 1'b0 ;
  assign n35336 = n22705 ^ n10724 ^ 1'b0 ;
  assign n35337 = ~n17490 & n35336 ;
  assign n35338 = n16616 & ~n26164 ;
  assign n35340 = ~n1588 & n2466 ;
  assign n35339 = ~n12088 & n21361 ;
  assign n35341 = n35340 ^ n35339 ^ 1'b0 ;
  assign n35342 = n22135 ^ n5029 ^ n801 ;
  assign n35343 = n2370 | n35342 ;
  assign n35344 = n4813 | n11789 ;
  assign n35345 = ~n2529 & n14359 ;
  assign n35346 = n34712 ^ n29800 ^ 1'b0 ;
  assign n35347 = n5557 & n11057 ;
  assign n35348 = ~n9744 & n35347 ;
  assign n35349 = n8532 | n21516 ;
  assign n35350 = n1117 & ~n35349 ;
  assign n35351 = ~n10859 & n12655 ;
  assign n35352 = ~n23996 & n35351 ;
  assign n35353 = ~n16435 & n31436 ;
  assign n35354 = n10340 & ~n17766 ;
  assign n35355 = n15430 ^ n10294 ^ 1'b0 ;
  assign n35356 = n10630 & ~n35355 ;
  assign n35357 = ~n21955 & n27894 ;
  assign n35359 = n11046 & ~n26351 ;
  assign n35360 = ~n6745 & n35359 ;
  assign n35358 = n5085 | n33602 ;
  assign n35361 = n35360 ^ n35358 ^ 1'b0 ;
  assign n35362 = ( n5720 & n20661 ) | ( n5720 & ~n23096 ) | ( n20661 & ~n23096 ) ;
  assign n35363 = ( n2869 & n3768 ) | ( n2869 & n35362 ) | ( n3768 & n35362 ) ;
  assign n35364 = n22655 | n35363 ;
  assign n35365 = n11004 & ~n14784 ;
  assign n35366 = n32949 ^ n3158 ^ 1'b0 ;
  assign n35367 = n2219 | n35366 ;
  assign n35368 = n20336 ^ n10031 ^ 1'b0 ;
  assign n35369 = n24853 & ~n35368 ;
  assign n35370 = n31815 & n35369 ;
  assign n35371 = n11196 | n27583 ;
  assign n35372 = n29745 ^ n29106 ^ 1'b0 ;
  assign n35373 = n35371 & ~n35372 ;
  assign n35374 = n23057 | n23677 ;
  assign n35375 = n3962 & n11621 ;
  assign n35376 = ~n35374 & n35375 ;
  assign n35377 = ~n2047 & n4793 ;
  assign n35378 = ~x234 & n35377 ;
  assign n35379 = n17864 & ~n35378 ;
  assign n35380 = n35379 ^ n2618 ^ 1'b0 ;
  assign n35381 = n6617 | n8722 ;
  assign n35382 = n1939 | n7420 ;
  assign n35383 = n6546 & ~n35382 ;
  assign n35385 = x64 & n21385 ;
  assign n35384 = ~n6362 & n10114 ;
  assign n35386 = n35385 ^ n35384 ^ 1'b0 ;
  assign n35387 = n28196 ^ n1326 ^ 1'b0 ;
  assign n35388 = n32453 ^ n2676 ^ 1'b0 ;
  assign n35389 = n1710 & n35388 ;
  assign n35390 = n298 & n35389 ;
  assign n35391 = n8667 ^ n3938 ^ 1'b0 ;
  assign n35392 = n1076 | n35391 ;
  assign n35393 = n21867 | n35392 ;
  assign n35394 = n1014 & n4562 ;
  assign n35395 = ~n35393 & n35394 ;
  assign n35396 = n35395 ^ n23199 ^ 1'b0 ;
  assign n35397 = x9 & ~n30018 ;
  assign n35398 = ~n22997 & n35397 ;
  assign n35399 = n24200 ^ n3378 ^ 1'b0 ;
  assign n35400 = n18588 & n33094 ;
  assign n35401 = n23788 ^ n2725 ^ 1'b0 ;
  assign n35402 = n13543 & ~n26370 ;
  assign n35403 = n7181 & n35402 ;
  assign n35404 = n7136 | n7878 ;
  assign n35405 = n11778 ^ n1339 ^ 1'b0 ;
  assign n35406 = ~n12901 & n35405 ;
  assign n35407 = n6502 | n8099 ;
  assign n35408 = ~n22907 & n30432 ;
  assign n35409 = n2975 & ~n19476 ;
  assign n35410 = n35409 ^ n18828 ^ 1'b0 ;
  assign n35411 = n23281 ^ n13602 ^ 1'b0 ;
  assign n35412 = n16948 & ~n26468 ;
  assign n35413 = ~n7196 & n35412 ;
  assign n35414 = n12581 & ~n15242 ;
  assign n35415 = n35414 ^ n6985 ^ 1'b0 ;
  assign n35416 = n29412 ^ n1419 ^ 1'b0 ;
  assign n35417 = n35415 | n35416 ;
  assign n35418 = n3496 & ~n35417 ;
  assign n35419 = n7924 ^ n6060 ^ 1'b0 ;
  assign n35420 = n25100 ^ n22729 ^ 1'b0 ;
  assign n35421 = ~n35419 & n35420 ;
  assign n35422 = n31053 ^ n22914 ^ n18705 ;
  assign n35423 = n29052 ^ n2409 ^ 1'b0 ;
  assign n35424 = n2061 ^ n1227 ^ 1'b0 ;
  assign n35425 = ~n5560 & n35424 ;
  assign n35426 = ~n14233 & n31820 ;
  assign n35427 = n35426 ^ n30258 ^ 1'b0 ;
  assign n35428 = n24442 & n33089 ;
  assign n35429 = n1754 & n35428 ;
  assign n35430 = ~n2495 & n27443 ;
  assign n35431 = n35430 ^ n24351 ^ 1'b0 ;
  assign n35432 = ~n35429 & n35431 ;
  assign n35433 = n519 & ~n11521 ;
  assign n35434 = n19575 ^ n12451 ^ 1'b0 ;
  assign n35435 = n9907 & n26372 ;
  assign n35436 = ~n35434 & n35435 ;
  assign n35437 = n709 | n2248 ;
  assign n35438 = n35437 ^ n19249 ^ 1'b0 ;
  assign n35439 = ~n2609 & n22659 ;
  assign n35440 = n15964 ^ n1038 ^ 1'b0 ;
  assign n35441 = n8107 & n35440 ;
  assign n35442 = n35441 ^ n9541 ^ 1'b0 ;
  assign n35443 = ~n4215 & n18494 ;
  assign n35444 = n2335 & ~n17548 ;
  assign n35445 = n6553 | n35444 ;
  assign n35446 = n921 | n28241 ;
  assign n35447 = n23763 ^ n9976 ^ 1'b0 ;
  assign n35448 = ~n25556 & n35447 ;
  assign n35449 = n5203 | n6365 ;
  assign n35450 = n7715 & ~n35449 ;
  assign n35451 = n11973 ^ n552 ^ 1'b0 ;
  assign n35452 = n7713 & n35451 ;
  assign n35453 = ~n35450 & n35452 ;
  assign n35454 = n35453 ^ n11346 ^ 1'b0 ;
  assign n35455 = n17706 ^ n6368 ^ 1'b0 ;
  assign n35456 = n35454 & n35455 ;
  assign n35457 = n10436 & ~n13232 ;
  assign n35458 = n20151 ^ n9652 ^ 1'b0 ;
  assign n35459 = n26225 | n27977 ;
  assign n35460 = n20783 | n35459 ;
  assign n35461 = ~n8113 & n10865 ;
  assign n35462 = x28 & n8843 ;
  assign n35463 = n35462 ^ n7112 ^ 1'b0 ;
  assign n35464 = n1939 | n35463 ;
  assign n35465 = n35461 & ~n35464 ;
  assign n35466 = n3033 & ~n23279 ;
  assign n35467 = n290 | n19122 ;
  assign n35468 = ~n1248 & n23721 ;
  assign n35469 = ~n12965 & n35468 ;
  assign n35470 = ~n15081 & n16200 ;
  assign n35471 = n35470 ^ n10302 ^ 1'b0 ;
  assign n35472 = n33036 ^ n27704 ^ 1'b0 ;
  assign n35473 = ~n35471 & n35472 ;
  assign n35474 = ~n2436 & n2714 ;
  assign n35475 = n17552 ^ n3473 ^ 1'b0 ;
  assign n35476 = n11171 & ~n35475 ;
  assign n35477 = x237 & n29086 ;
  assign n35478 = n1656 | n8584 ;
  assign n35479 = n35478 ^ n17461 ^ 1'b0 ;
  assign n35480 = n15210 & n34748 ;
  assign n35481 = n25050 | n25227 ;
  assign n35482 = x6 & ~n6523 ;
  assign n35483 = ~n968 & n20358 ;
  assign n35484 = ~n35482 & n35483 ;
  assign n35485 = n23449 & n24993 ;
  assign n35486 = n28079 ^ n13712 ^ 1'b0 ;
  assign n35487 = n7967 & ~n35486 ;
  assign n35488 = ~n6449 & n17372 ;
  assign n35489 = n21233 | n22760 ;
  assign n35490 = n15032 & ~n35489 ;
  assign n35491 = n4500 & ~n12809 ;
  assign n35492 = n32745 ^ n31773 ^ n28640 ;
  assign n35493 = n4326 & n7640 ;
  assign n35494 = n33074 ^ n2785 ^ 1'b0 ;
  assign n35495 = n8773 & n18077 ;
  assign n35496 = ~n2310 & n35495 ;
  assign n35497 = n35496 ^ n28640 ^ 1'b0 ;
  assign n35498 = n13093 & n14332 ;
  assign n35499 = n4039 & n35498 ;
  assign n35500 = n4707 ^ x100 ^ 1'b0 ;
  assign n35501 = n10394 | n35500 ;
  assign n35502 = n35501 ^ n1247 ^ 1'b0 ;
  assign n35503 = n27733 & ~n35502 ;
  assign n35504 = n2589 & ~n3879 ;
  assign n35505 = ( n663 & n4490 ) | ( n663 & ~n35504 ) | ( n4490 & ~n35504 ) ;
  assign n35506 = n8646 ^ n1195 ^ 1'b0 ;
  assign n35507 = n10298 & n29317 ;
  assign n35508 = n20790 ^ n5018 ^ 1'b0 ;
  assign n35509 = n24661 & n35508 ;
  assign n35510 = n8387 ^ n7054 ^ 1'b0 ;
  assign n35511 = n26588 | n35510 ;
  assign n35512 = ~n15051 & n21497 ;
  assign n35513 = n2181 | n4655 ;
  assign n35514 = n561 | n35513 ;
  assign n35515 = ~n3793 & n21474 ;
  assign n35516 = n1389 & ~n10383 ;
  assign n35517 = n6862 & n31423 ;
  assign n35518 = n5728 | n21943 ;
  assign n35519 = n11385 | n14038 ;
  assign n35520 = n9776 | n35519 ;
  assign n35524 = ~n5691 & n16269 ;
  assign n35525 = n35524 ^ n1637 ^ 1'b0 ;
  assign n35523 = n10523 ^ n825 ^ 1'b0 ;
  assign n35526 = n35525 ^ n35523 ^ 1'b0 ;
  assign n35521 = ~n4671 & n6094 ;
  assign n35522 = n35521 ^ n29556 ^ 1'b0 ;
  assign n35527 = n35526 ^ n35522 ^ 1'b0 ;
  assign n35528 = n25290 ^ n16122 ^ 1'b0 ;
  assign n35529 = n10340 & ~n35528 ;
  assign n35531 = n31101 ^ n26962 ^ 1'b0 ;
  assign n35530 = n1773 & ~n34397 ;
  assign n35532 = n35531 ^ n35530 ^ 1'b0 ;
  assign n35533 = n8518 | n35532 ;
  assign n35534 = ~n7253 & n12928 ;
  assign n35535 = n20751 ^ n18671 ^ 1'b0 ;
  assign n35536 = n14509 & n35535 ;
  assign n35537 = n6045 & ~n13503 ;
  assign n35538 = n35537 ^ n2433 ^ 1'b0 ;
  assign n35539 = ~n12030 & n35538 ;
  assign n35540 = n9857 & n35539 ;
  assign n35541 = n14236 ^ x132 ^ 1'b0 ;
  assign n35542 = n3377 & ~n35541 ;
  assign n35543 = n21097 & n35542 ;
  assign n35544 = n35543 ^ n7646 ^ 1'b0 ;
  assign n35545 = n20563 & ~n30851 ;
  assign n35546 = n17480 & n26489 ;
  assign n35547 = n19725 & n35546 ;
  assign n35548 = n9919 & ~n18668 ;
  assign n35552 = x2 | n11687 ;
  assign n35549 = n926 & n23929 ;
  assign n35550 = ~n2684 & n35549 ;
  assign n35551 = n35514 | n35550 ;
  assign n35553 = n35552 ^ n35551 ^ 1'b0 ;
  assign n35554 = n26343 ^ n25238 ^ 1'b0 ;
  assign n35555 = n29926 & ~n32981 ;
  assign n35556 = n11856 ^ n6399 ^ 1'b0 ;
  assign n35557 = n16489 | n35556 ;
  assign n35558 = n2818 | n12041 ;
  assign n35559 = n35558 ^ n13285 ^ 1'b0 ;
  assign n35560 = ~n2737 & n35559 ;
  assign n35561 = n16568 & ~n28161 ;
  assign n35562 = ~n35560 & n35561 ;
  assign n35563 = n23417 ^ n6498 ^ 1'b0 ;
  assign n35564 = ~n9944 & n35563 ;
  assign n35565 = n26239 & n27153 ;
  assign n35566 = n19681 ^ n1588 ^ 1'b0 ;
  assign n35567 = n21105 | n30246 ;
  assign n35568 = ~n8730 & n19089 ;
  assign n35569 = ~n1657 & n3054 ;
  assign n35570 = ~n942 & n35569 ;
  assign n35571 = n11204 | n21729 ;
  assign n35572 = n35571 ^ n815 ^ 1'b0 ;
  assign n35573 = n35572 ^ n2841 ^ 1'b0 ;
  assign n35574 = n1703 & n35573 ;
  assign n35575 = n4159 | n34247 ;
  assign n35576 = n4334 & ~n35575 ;
  assign n35577 = n9745 & n34880 ;
  assign n35578 = n25100 ^ n1488 ^ 1'b0 ;
  assign n35579 = x57 & ~n3521 ;
  assign n35580 = n19780 & n35579 ;
  assign n35581 = n20716 ^ n16855 ^ 1'b0 ;
  assign n35582 = n17609 ^ n6851 ^ 1'b0 ;
  assign n35583 = n13978 ^ n337 ^ 1'b0 ;
  assign n35584 = ~n9654 & n35583 ;
  assign n35585 = n5698 | n32327 ;
  assign n35586 = n11945 & ~n35585 ;
  assign n35587 = n35586 ^ n10149 ^ 1'b0 ;
  assign n35588 = n35587 ^ n24702 ^ 1'b0 ;
  assign n35589 = n15614 & ~n26243 ;
  assign n35590 = n19908 ^ n2378 ^ 1'b0 ;
  assign n35591 = n11323 & ~n22168 ;
  assign n35592 = n35591 ^ n4538 ^ 1'b0 ;
  assign n35593 = n15478 ^ n10626 ^ n3322 ;
  assign n35594 = n26067 | n35593 ;
  assign n35595 = n32681 & ~n35594 ;
  assign n35596 = n26554 & ~n35595 ;
  assign n35597 = n35596 ^ n4701 ^ 1'b0 ;
  assign n35598 = n3026 & ~n3169 ;
  assign n35599 = n35598 ^ n11335 ^ 1'b0 ;
  assign n35600 = n6997 & ~n35599 ;
  assign n35601 = n3603 & n35600 ;
  assign n35602 = n5790 | n22641 ;
  assign n35603 = n12525 ^ n5958 ^ 1'b0 ;
  assign n35604 = n35602 & n35603 ;
  assign n35605 = n11570 ^ n2078 ^ 1'b0 ;
  assign n35606 = ~n3611 & n14449 ;
  assign n35607 = n25337 & ~n35606 ;
  assign n35608 = n27657 ^ n12514 ^ 1'b0 ;
  assign n35609 = ~n11442 & n14525 ;
  assign n35610 = n31243 & ~n35609 ;
  assign n35611 = n35608 & ~n35610 ;
  assign n35612 = ~n8054 & n32556 ;
  assign n35613 = n23952 ^ n11950 ^ 1'b0 ;
  assign n35614 = n21361 & n35613 ;
  assign n35616 = n16588 ^ n6039 ^ 1'b0 ;
  assign n35617 = ~n17935 & n35616 ;
  assign n35615 = n7454 & n27457 ;
  assign n35618 = n35617 ^ n35615 ^ 1'b0 ;
  assign n35619 = n35618 ^ n13311 ^ 1'b0 ;
  assign n35620 = n35614 & n35619 ;
  assign n35621 = n14299 & n33312 ;
  assign n35626 = n17800 | n28835 ;
  assign n35627 = n14994 & ~n35626 ;
  assign n35624 = n2861 | n9707 ;
  assign n35622 = n22977 ^ n9360 ^ 1'b0 ;
  assign n35623 = n4265 & n35622 ;
  assign n35625 = n35624 ^ n35623 ^ 1'b0 ;
  assign n35628 = n35627 ^ n35625 ^ n6343 ;
  assign n35629 = ( n1605 & n2870 ) | ( n1605 & ~n24426 ) | ( n2870 & ~n24426 ) ;
  assign n35630 = ~n2519 & n35629 ;
  assign n35631 = ~n14102 & n35630 ;
  assign n35632 = n3015 & n22160 ;
  assign n35633 = n14261 & n35632 ;
  assign n35634 = n21342 ^ n5560 ^ 1'b0 ;
  assign n35635 = n20283 & n35634 ;
  assign n35636 = ~n1623 & n18092 ;
  assign n35637 = n35636 ^ n28886 ^ 1'b0 ;
  assign n35638 = n307 | n27747 ;
  assign n35639 = n1977 ^ n1488 ^ 1'b0 ;
  assign n35640 = ~n15104 & n21669 ;
  assign n35641 = n35640 ^ n35082 ^ 1'b0 ;
  assign n35642 = n35639 | n35641 ;
  assign n35643 = n2561 & ~n5146 ;
  assign n35644 = n35643 ^ n6372 ^ 1'b0 ;
  assign n35645 = n4622 | n10877 ;
  assign n35646 = n6054 & ~n35645 ;
  assign n35647 = n35646 ^ n25805 ^ 1'b0 ;
  assign n35648 = n17477 | n35647 ;
  assign n35649 = n3158 & n10423 ;
  assign n35650 = n2333 & n35649 ;
  assign n35651 = n6211 ^ n1661 ^ 1'b0 ;
  assign n35652 = n15363 | n35651 ;
  assign n35653 = ~n2709 & n22669 ;
  assign n35654 = n25124 ^ n10709 ^ 1'b0 ;
  assign n35655 = n23653 ^ n1912 ^ n934 ;
  assign n35656 = n6443 ^ n1181 ^ 1'b0 ;
  assign n35657 = ~n8837 & n35656 ;
  assign n35658 = n21825 ^ n2296 ^ 1'b0 ;
  assign n35659 = n28689 ^ n8816 ^ 1'b0 ;
  assign n35660 = ~n35658 & n35659 ;
  assign n35661 = n35660 ^ n956 ^ 1'b0 ;
  assign n35662 = n11655 & ~n15552 ;
  assign n35664 = n17864 ^ n17114 ^ 1'b0 ;
  assign n35665 = n4549 & ~n35664 ;
  assign n35663 = ~n7588 & n27917 ;
  assign n35666 = n35665 ^ n35663 ^ 1'b0 ;
  assign n35670 = n1622 & ~n6811 ;
  assign n35667 = n5500 & n9353 ;
  assign n35668 = n35667 ^ n415 ^ 1'b0 ;
  assign n35669 = n2872 | n35668 ;
  assign n35671 = n35670 ^ n35669 ^ 1'b0 ;
  assign n35674 = ~n381 & n7738 ;
  assign n35672 = n8116 ^ n3437 ^ 1'b0 ;
  assign n35673 = n4152 & n35672 ;
  assign n35675 = n35674 ^ n35673 ^ n1815 ;
  assign n35676 = ~n2053 & n10387 ;
  assign n35677 = n16161 | n35676 ;
  assign n35678 = n666 & ~n10381 ;
  assign n35679 = ~n1553 & n10937 ;
  assign n35680 = n35679 ^ n14400 ^ 1'b0 ;
  assign n35681 = n25960 & ~n35680 ;
  assign n35682 = n35681 ^ n11915 ^ 1'b0 ;
  assign n35683 = n8403 | n14506 ;
  assign n35684 = n35683 ^ n23042 ^ 1'b0 ;
  assign n35685 = n35684 ^ n17130 ^ n4796 ;
  assign n35686 = n25189 ^ n7465 ^ n2849 ;
  assign n35687 = n11751 | n26447 ;
  assign n35688 = ~n15024 & n35687 ;
  assign n35689 = n3091 & n9907 ;
  assign n35690 = ~n26331 & n35689 ;
  assign n35691 = ~n8242 & n9276 ;
  assign n35692 = ~n5470 & n35691 ;
  assign n35693 = n35692 ^ n18913 ^ 1'b0 ;
  assign n35694 = n16337 ^ n3830 ^ 1'b0 ;
  assign n35695 = n10456 ^ n9606 ^ 1'b0 ;
  assign n35696 = ~n26187 & n27904 ;
  assign n35697 = n25216 ^ n20272 ^ 1'b0 ;
  assign n35700 = n3454 | n28560 ;
  assign n35701 = n4367 | n35700 ;
  assign n35698 = n3053 & ~n7495 ;
  assign n35699 = ~n16939 & n35698 ;
  assign n35702 = n35701 ^ n35699 ^ 1'b0 ;
  assign n35703 = ( n5070 & n26301 ) | ( n5070 & ~n28297 ) | ( n26301 & ~n28297 ) ;
  assign n35704 = n20208 ^ n556 ^ 1'b0 ;
  assign n35705 = n26152 ^ n4566 ^ 1'b0 ;
  assign n35706 = n4953 & n35705 ;
  assign n35707 = n27596 & n30760 ;
  assign n35708 = n21321 ^ n7045 ^ 1'b0 ;
  assign n35709 = ~n3950 & n35708 ;
  assign n35710 = ~n32487 & n35709 ;
  assign n35711 = n35710 ^ n18916 ^ 1'b0 ;
  assign n35712 = n35429 ^ n21329 ^ n15374 ;
  assign n35713 = n27704 ^ n14084 ^ 1'b0 ;
  assign n35714 = ~n5634 & n31627 ;
  assign n35715 = n2466 & n3428 ;
  assign n35716 = ~n14350 & n35715 ;
  assign n35717 = n16733 ^ n5646 ^ 1'b0 ;
  assign n35718 = n35716 & ~n35717 ;
  assign n35719 = n19475 ^ n6433 ^ 1'b0 ;
  assign n35720 = n6311 & ~n35719 ;
  assign n35721 = n4204 & ~n17783 ;
  assign n35722 = ~n18148 & n35721 ;
  assign n35723 = n2515 & ~n3100 ;
  assign n35724 = n35723 ^ x170 ^ 1'b0 ;
  assign n35725 = n392 | n35724 ;
  assign n35726 = n19549 ^ n5097 ^ 1'b0 ;
  assign n35727 = ~n1512 & n35726 ;
  assign n35728 = n3175 | n4108 ;
  assign n35729 = n35728 ^ n16142 ^ 1'b0 ;
  assign n35730 = n28357 | n33743 ;
  assign n35731 = n35730 ^ n19508 ^ 1'b0 ;
  assign n35735 = n1671 & ~n2237 ;
  assign n35732 = n4608 & ~n7278 ;
  assign n35733 = ~n4238 & n35732 ;
  assign n35734 = n35733 ^ n2938 ^ 1'b0 ;
  assign n35736 = n35735 ^ n35734 ^ n28240 ;
  assign n35737 = n19300 | n23985 ;
  assign n35738 = n2616 | n35737 ;
  assign n35739 = n17579 ^ n17132 ^ 1'b0 ;
  assign n35740 = n23402 & n35739 ;
  assign n35741 = n35740 ^ n25417 ^ 1'b0 ;
  assign n35742 = n35738 & ~n35741 ;
  assign n35743 = ~n19273 & n23463 ;
  assign n35744 = n35743 ^ n3774 ^ 1'b0 ;
  assign n35745 = n19216 | n28412 ;
  assign n35746 = n35744 | n35745 ;
  assign n35747 = n4094 & n8844 ;
  assign n35748 = ~n444 & n35747 ;
  assign n35749 = n16134 ^ n14518 ^ 1'b0 ;
  assign n35750 = n11455 & n35749 ;
  assign n35751 = ( n14353 & n29324 ) | ( n14353 & ~n35750 ) | ( n29324 & ~n35750 ) ;
  assign n35752 = n19052 ^ n15306 ^ 1'b0 ;
  assign n35753 = n19299 ^ n10225 ^ 1'b0 ;
  assign n35754 = ~n6440 & n12855 ;
  assign n35755 = n12389 ^ n10135 ^ 1'b0 ;
  assign n35756 = ~n35754 & n35755 ;
  assign n35757 = n10222 & n35756 ;
  assign n35758 = n35753 & n35757 ;
  assign n35760 = ~n11904 & n16676 ;
  assign n35759 = n10288 & ~n15583 ;
  assign n35761 = n35760 ^ n35759 ^ 1'b0 ;
  assign n35762 = n15991 & ~n23165 ;
  assign n35763 = n35762 ^ n593 ^ 1'b0 ;
  assign n35764 = n35763 ^ n10376 ^ 1'b0 ;
  assign n35765 = n10155 | n35764 ;
  assign n35766 = n22245 ^ n17443 ^ 1'b0 ;
  assign n35767 = n2578 & n35766 ;
  assign n35768 = n35767 ^ n8733 ^ n6932 ;
  assign n35769 = n35768 ^ n13034 ^ 1'b0 ;
  assign n35770 = n24908 & ~n35769 ;
  assign n35771 = n11108 & n35770 ;
  assign n35772 = n35771 ^ n30100 ^ 1'b0 ;
  assign n35773 = n20729 ^ n1568 ^ 1'b0 ;
  assign n35774 = n1027 & ~n35773 ;
  assign n35775 = n11919 ^ n3625 ^ 1'b0 ;
  assign n35776 = n25094 ^ n1579 ^ 1'b0 ;
  assign n35777 = n5774 & ~n35776 ;
  assign n35778 = n16391 & ~n34893 ;
  assign n35779 = ~n35777 & n35778 ;
  assign n35781 = n16893 ^ n1228 ^ 1'b0 ;
  assign n35780 = n23480 ^ n4464 ^ 1'b0 ;
  assign n35782 = n35781 ^ n35780 ^ n33089 ;
  assign n35783 = n5748 | n11568 ;
  assign n35784 = n562 & ~n35783 ;
  assign n35785 = ~n15416 & n18196 ;
  assign n35786 = ~n3475 & n25395 ;
  assign n35787 = n4728 | n22286 ;
  assign n35788 = n14590 & ~n35260 ;
  assign n35789 = n1275 & n8417 ;
  assign n35790 = n28369 & n35789 ;
  assign n35791 = n2807 & n7931 ;
  assign n35792 = ~n10886 & n21786 ;
  assign n35793 = n35792 ^ n744 ^ 1'b0 ;
  assign n35794 = n10330 | n28478 ;
  assign n35795 = x25 & ~n35794 ;
  assign n35796 = ~n2711 & n35795 ;
  assign n35797 = ~n17896 & n35796 ;
  assign n35798 = n10328 & n35797 ;
  assign n35799 = n4217 ^ n2239 ^ 1'b0 ;
  assign n35800 = x112 | n3336 ;
  assign n35802 = n1701 & ~n10829 ;
  assign n35801 = n20275 | n30498 ;
  assign n35803 = n35802 ^ n35801 ^ 1'b0 ;
  assign n35804 = n35803 ^ n23593 ^ 1'b0 ;
  assign n35805 = n3721 & n4811 ;
  assign n35806 = ~n672 & n2040 ;
  assign n35807 = n35806 ^ n5664 ^ 1'b0 ;
  assign n35808 = ( ~n540 & n21545 ) | ( ~n540 & n25730 ) | ( n21545 & n25730 ) ;
  assign n35809 = ~n7028 & n10827 ;
  assign n35810 = n9897 & n35809 ;
  assign n35811 = n16832 ^ n747 ^ 1'b0 ;
  assign n35812 = n24262 ^ n2138 ^ 1'b0 ;
  assign n35813 = n3844 & ~n35812 ;
  assign n35814 = ~n4919 & n12941 ;
  assign n35815 = n35814 ^ n1256 ^ 1'b0 ;
  assign n35816 = n12248 | n35815 ;
  assign n35817 = n35816 ^ n10469 ^ 1'b0 ;
  assign n35818 = n7268 & ~n18835 ;
  assign n35819 = n20608 | n35818 ;
  assign n35820 = n35817 | n35819 ;
  assign n35822 = n2790 ^ n1568 ^ 1'b0 ;
  assign n35823 = n2218 & ~n35822 ;
  assign n35821 = n20884 & n22663 ;
  assign n35824 = n35823 ^ n35821 ^ 1'b0 ;
  assign n35825 = n5512 & n18796 ;
  assign n35826 = n35825 ^ n1691 ^ 1'b0 ;
  assign n35827 = ~x22 & n25162 ;
  assign n35828 = n28249 ^ n807 ^ 1'b0 ;
  assign n35829 = n963 | n33845 ;
  assign n35830 = n7777 ^ n7195 ^ 1'b0 ;
  assign n35831 = n411 | n35830 ;
  assign n35832 = n35831 ^ n15486 ^ 1'b0 ;
  assign n35833 = ~n10437 & n25800 ;
  assign n35834 = n15328 ^ n12213 ^ 1'b0 ;
  assign n35835 = n9590 & n9989 ;
  assign n35836 = n11488 & ~n24429 ;
  assign n35837 = n35836 ^ n20085 ^ 1'b0 ;
  assign n35838 = n7427 | n14078 ;
  assign n35839 = n12559 & ~n35838 ;
  assign n35840 = n27281 ^ n1018 ^ 1'b0 ;
  assign n35841 = n26838 | n35840 ;
  assign n35842 = ~n6389 & n21969 ;
  assign n35843 = ( ~n987 & n3181 ) | ( ~n987 & n35842 ) | ( n3181 & n35842 ) ;
  assign n35844 = n22604 ^ n10273 ^ 1'b0 ;
  assign n35845 = ~n15429 & n35844 ;
  assign n35846 = n19130 & n21182 ;
  assign n35847 = n3532 & ~n30610 ;
  assign n35848 = n35847 ^ n3487 ^ 1'b0 ;
  assign n35849 = n12498 | n35848 ;
  assign n35850 = n35846 & ~n35849 ;
  assign n35851 = n1071 & ~n35850 ;
  assign n35852 = ~n35845 & n35851 ;
  assign n35853 = n18254 & n21820 ;
  assign n35854 = n13532 | n24676 ;
  assign n35855 = n28299 | n35854 ;
  assign n35856 = ~n325 & n4026 ;
  assign n35857 = n2707 & n35856 ;
  assign n35858 = n35857 ^ n34250 ^ 1'b0 ;
  assign n35859 = ~n5574 & n29753 ;
  assign n35860 = n12058 & n35859 ;
  assign n35861 = n35860 ^ n32986 ^ 1'b0 ;
  assign n35862 = n19907 & ~n30563 ;
  assign n35863 = n35862 ^ n29872 ^ n1515 ;
  assign n35864 = n19754 ^ n16174 ^ 1'b0 ;
  assign n35865 = n1970 & n35864 ;
  assign n35866 = n320 & n6822 ;
  assign n35867 = n820 & n35866 ;
  assign n35868 = n15825 | n26565 ;
  assign n35869 = n1441 & n16657 ;
  assign n35870 = ~n24073 & n35869 ;
  assign n35871 = n7555 & n35870 ;
  assign n35872 = n35871 ^ n24502 ^ 1'b0 ;
  assign n35873 = n14472 | n35872 ;
  assign n35874 = n10826 | n20488 ;
  assign n35875 = ~n12924 & n30537 ;
  assign n35876 = ~n9562 & n35875 ;
  assign n35877 = n13895 | n17240 ;
  assign n35878 = n32194 ^ n16376 ^ 1'b0 ;
  assign n35879 = n5880 & n27380 ;
  assign n35880 = n6735 | n35879 ;
  assign n35881 = ~n1882 & n11567 ;
  assign n35882 = n12151 ^ n5462 ^ 1'b0 ;
  assign n35883 = ~n2591 & n35882 ;
  assign n35885 = n12131 ^ n718 ^ 1'b0 ;
  assign n35884 = n9923 ^ n2378 ^ x253 ;
  assign n35886 = n35885 ^ n35884 ^ n20717 ;
  assign n35887 = n27532 ^ n3530 ^ 1'b0 ;
  assign n35888 = n30894 ^ n8951 ^ n3171 ;
  assign n35889 = n33559 ^ n21930 ^ 1'b0 ;
  assign n35890 = ( n6595 & n7196 ) | ( n6595 & n26520 ) | ( n7196 & n26520 ) ;
  assign n35891 = n2486 & ~n20619 ;
  assign n35892 = n6812 & n13262 ;
  assign n35893 = n35892 ^ n9304 ^ 1'b0 ;
  assign n35894 = n15381 ^ x146 ^ 1'b0 ;
  assign n35895 = n27411 & n35894 ;
  assign n35896 = ~n2114 & n35895 ;
  assign n35897 = ~n33512 & n35896 ;
  assign n35898 = n35897 ^ n4370 ^ 1'b0 ;
  assign n35899 = n17260 ^ n7000 ^ 1'b0 ;
  assign n35900 = n28692 & ~n35899 ;
  assign n35901 = ~n9990 & n35900 ;
  assign n35902 = n490 & ~n7757 ;
  assign n35903 = ~n31341 & n33872 ;
  assign n35904 = n35903 ^ n10488 ^ 1'b0 ;
  assign n35905 = n4380 & ~n17046 ;
  assign n35906 = n15054 | n17182 ;
  assign n35907 = n4429 & n13982 ;
  assign n35908 = n17593 ^ n11732 ^ n7400 ;
  assign n35909 = n3635 | n35908 ;
  assign n35910 = n16157 ^ n9246 ^ 1'b0 ;
  assign n35911 = n18231 ^ n7710 ^ 1'b0 ;
  assign n35912 = ~n25622 & n35911 ;
  assign n35913 = ~n19110 & n35912 ;
  assign n35914 = ~n32787 & n35913 ;
  assign n35915 = n35914 ^ n27212 ^ 1'b0 ;
  assign n35916 = x200 | n4708 ;
  assign n35917 = n26208 & ~n35916 ;
  assign n35918 = ~n3378 & n18937 ;
  assign n35919 = ~n35917 & n35918 ;
  assign n35920 = n12161 & n14344 ;
  assign n35921 = n5443 ^ n4169 ^ 1'b0 ;
  assign n35922 = n9562 & n12402 ;
  assign n35923 = n35922 ^ n4095 ^ 1'b0 ;
  assign n35924 = n35923 ^ n19966 ^ 1'b0 ;
  assign n35925 = n35921 & ~n35924 ;
  assign n35926 = ~n14907 & n27967 ;
  assign n35927 = n35926 ^ n9188 ^ 1'b0 ;
  assign n35928 = n10126 ^ n2087 ^ 1'b0 ;
  assign n35929 = n8088 & ~n35928 ;
  assign n35930 = n11341 ^ n4711 ^ 1'b0 ;
  assign n35931 = ~n13075 & n35930 ;
  assign n35932 = ( n23874 & n35929 ) | ( n23874 & n35931 ) | ( n35929 & n35931 ) ;
  assign n35933 = n3740 ^ n1361 ^ 1'b0 ;
  assign n35934 = n35933 ^ n30648 ^ 1'b0 ;
  assign n35935 = n22572 ^ n21812 ^ 1'b0 ;
  assign n35936 = n15089 & n35935 ;
  assign n35937 = ~n18041 & n35936 ;
  assign n35938 = n14474 ^ n2591 ^ 1'b0 ;
  assign n35939 = n16782 ^ n14852 ^ 1'b0 ;
  assign n35940 = n3203 & ~n6162 ;
  assign n35941 = ~n17726 & n34145 ;
  assign n35942 = n32582 & ~n35941 ;
  assign n35943 = ~n5484 & n12354 ;
  assign n35944 = ~n24850 & n35943 ;
  assign n35945 = n2242 & ~n29028 ;
  assign n35946 = ~n18192 & n35945 ;
  assign n35947 = n35946 ^ n14301 ^ 1'b0 ;
  assign n35948 = n35944 & n35947 ;
  assign n35951 = n5298 ^ n1855 ^ 1'b0 ;
  assign n35952 = n6034 & ~n35951 ;
  assign n35950 = n10697 & ~n18527 ;
  assign n35953 = n35952 ^ n35950 ^ 1'b0 ;
  assign n35949 = n5932 & n17536 ;
  assign n35954 = n35953 ^ n35949 ^ 1'b0 ;
  assign n35955 = n24363 & ~n28115 ;
  assign n35956 = n15715 ^ n10146 ^ 1'b0 ;
  assign n35957 = n11093 & n35956 ;
  assign n35958 = ~n30290 & n34017 ;
  assign n35959 = n14669 & ~n17255 ;
  assign n35960 = n22439 & ~n32097 ;
  assign n35961 = n35960 ^ n13206 ^ 1'b0 ;
  assign n35962 = n21577 & n32388 ;
  assign n35963 = ~n4325 & n17590 ;
  assign n35964 = n35963 ^ n27433 ^ 1'b0 ;
  assign n35965 = n1321 | n2462 ;
  assign n35966 = n16238 ^ n13850 ^ 1'b0 ;
  assign n35967 = n17746 ^ n7384 ^ 1'b0 ;
  assign n35968 = n35966 & n35967 ;
  assign n35969 = n19138 & n32953 ;
  assign n35970 = n14703 & ~n26625 ;
  assign n35971 = n13288 | n17531 ;
  assign n35972 = n35971 ^ n10567 ^ 1'b0 ;
  assign n35973 = n480 | n5758 ;
  assign n35974 = n20619 | n35973 ;
  assign n35975 = n7021 & ~n35974 ;
  assign n35976 = n35975 ^ n2076 ^ 1'b0 ;
  assign n35977 = n26216 & n35976 ;
  assign n35978 = ~n20430 & n21636 ;
  assign n35979 = n6368 | n35978 ;
  assign n35980 = n35979 ^ n10944 ^ 1'b0 ;
  assign n35981 = n1937 ^ n1857 ^ 1'b0 ;
  assign n35982 = n858 | n35981 ;
  assign n35984 = n9547 & ~n31637 ;
  assign n35983 = ~n13818 & n15421 ;
  assign n35985 = n35984 ^ n35983 ^ 1'b0 ;
  assign n35986 = n2870 & ~n5048 ;
  assign n35987 = n18609 | n26199 ;
  assign n35988 = n35987 ^ n24119 ^ 1'b0 ;
  assign n35989 = n4048 & n12162 ;
  assign n35990 = ~n5615 & n9269 ;
  assign n35991 = n4159 | n6557 ;
  assign n35992 = n4932 ^ n354 ^ 1'b0 ;
  assign n35993 = n35991 & n35992 ;
  assign n35994 = n10575 ^ n6355 ^ 1'b0 ;
  assign n35995 = n11100 & n19130 ;
  assign n35996 = ( n10931 & n19442 ) | ( n10931 & n30003 ) | ( n19442 & n30003 ) ;
  assign n35997 = n5728 ^ n4537 ^ 1'b0 ;
  assign n35998 = ~n21939 & n35997 ;
  assign n35999 = n13217 | n18512 ;
  assign n36000 = n17807 ^ n1784 ^ 1'b0 ;
  assign n36001 = n2715 & n36000 ;
  assign n36002 = n33374 ^ n3140 ^ 1'b0 ;
  assign n36003 = n1441 & ~n17584 ;
  assign n36004 = n13630 ^ n10239 ^ 1'b0 ;
  assign n36005 = n2293 | n31074 ;
  assign n36006 = n36005 ^ n22667 ^ 1'b0 ;
  assign n36007 = n1212 | n14923 ;
  assign n36008 = n36007 ^ n5750 ^ 1'b0 ;
  assign n36009 = n4826 & ~n24816 ;
  assign n36010 = n35037 ^ n26074 ^ 1'b0 ;
  assign n36011 = n2853 & n36010 ;
  assign n36012 = ~n7683 & n14525 ;
  assign n36013 = x36 & ~n10192 ;
  assign n36014 = n36013 ^ n35791 ^ n2083 ;
  assign n36015 = n8049 & ~n18947 ;
  assign n36016 = n36015 ^ n31967 ^ 1'b0 ;
  assign n36017 = ~n5440 & n8223 ;
  assign n36018 = n1056 | n11738 ;
  assign n36019 = n36017 | n36018 ;
  assign n36020 = n10488 | n36019 ;
  assign n36021 = n11615 | n18407 ;
  assign n36022 = n36021 ^ n3531 ^ 1'b0 ;
  assign n36023 = n7646 | n36022 ;
  assign n36026 = n19774 ^ n19696 ^ n12988 ;
  assign n36024 = n5852 & ~n9463 ;
  assign n36025 = ~n14216 & n36024 ;
  assign n36027 = n36026 ^ n36025 ^ 1'b0 ;
  assign n36028 = n6869 | n19033 ;
  assign n36029 = n12512 | n20672 ;
  assign n36030 = n4005 | n36029 ;
  assign n36031 = n35102 ^ n384 ^ 1'b0 ;
  assign n36032 = n17134 & n24244 ;
  assign n36033 = n32778 & n36032 ;
  assign n36034 = n5566 | n14472 ;
  assign n36035 = n36034 ^ n6978 ^ 1'b0 ;
  assign n36036 = n36035 ^ n33308 ^ 1'b0 ;
  assign n36037 = n4891 & n34208 ;
  assign n36038 = n5998 | n18070 ;
  assign n36039 = n19966 ^ n6945 ^ 1'b0 ;
  assign n36040 = n2221 & ~n12238 ;
  assign n36041 = n8126 & n20314 ;
  assign n36042 = n8216 & n36041 ;
  assign n36043 = n27529 ^ n3364 ^ 1'b0 ;
  assign n36044 = n1260 & ~n1383 ;
  assign n36045 = n11082 | n36044 ;
  assign n36046 = n1914 & n2276 ;
  assign n36047 = n36046 ^ n4576 ^ 1'b0 ;
  assign n36048 = n26312 ^ n4197 ^ 1'b0 ;
  assign n36049 = x27 & n28427 ;
  assign n36050 = ~n36048 & n36049 ;
  assign n36051 = x66 & n3097 ;
  assign n36052 = ~n3741 & n10238 ;
  assign n36053 = n36052 ^ n35072 ^ 1'b0 ;
  assign n36054 = n15389 & ~n28339 ;
  assign n36055 = ~n4132 & n27211 ;
  assign n36056 = n36055 ^ n17926 ^ 1'b0 ;
  assign n36057 = n13116 & n36056 ;
  assign n36058 = n36057 ^ n21527 ^ 1'b0 ;
  assign n36059 = n9057 & ~n20337 ;
  assign n36060 = n4972 & n36059 ;
  assign n36061 = n11885 | n16733 ;
  assign n36062 = n35961 ^ n8489 ^ 1'b0 ;
  assign n36063 = n7437 & n36062 ;
  assign n36064 = n10218 & ~n29858 ;
  assign n36065 = n36064 ^ n8047 ^ 1'b0 ;
  assign n36066 = n6355 ^ n3549 ^ 1'b0 ;
  assign n36067 = n36066 ^ n20185 ^ 1'b0 ;
  assign n36068 = ~n7415 & n15971 ;
  assign n36069 = n36068 ^ n16561 ^ 1'b0 ;
  assign n36070 = ~n30475 & n31259 ;
  assign n36071 = n16083 ^ n9548 ^ 1'b0 ;
  assign n36072 = ~n11968 & n23647 ;
  assign n36073 = n36071 & n36072 ;
  assign n36074 = n3933 & ~n16246 ;
  assign n36075 = n36074 ^ n2431 ^ x78 ;
  assign n36076 = n13169 & n26592 ;
  assign n36077 = n36076 ^ n34188 ^ 1'b0 ;
  assign n36078 = n21230 & ~n36077 ;
  assign n36079 = n11520 ^ n1356 ^ 1'b0 ;
  assign n36080 = n34121 & n36079 ;
  assign n36081 = n20692 & n30491 ;
  assign n36082 = ~n36080 & n36081 ;
  assign n36083 = n20553 ^ n1710 ^ 1'b0 ;
  assign n36084 = ~n3243 & n8442 ;
  assign n36085 = ~n36083 & n36084 ;
  assign n36086 = n4993 | n8647 ;
  assign n36087 = n8454 & n36086 ;
  assign n36088 = ~n1952 & n36087 ;
  assign n36089 = n28750 ^ n3060 ^ 1'b0 ;
  assign n36090 = n3356 & ~n36089 ;
  assign n36091 = n36090 ^ n10188 ^ 1'b0 ;
  assign n36092 = n17199 ^ n12163 ^ 1'b0 ;
  assign n36093 = n20938 ^ n5867 ^ 1'b0 ;
  assign n36094 = n26642 & n36093 ;
  assign n36095 = ~n5336 & n7400 ;
  assign n36096 = n16466 & n36095 ;
  assign n36097 = n23874 ^ n19316 ^ 1'b0 ;
  assign n36098 = n10488 ^ n1523 ^ 1'b0 ;
  assign n36099 = n6792 & ~n36098 ;
  assign n36100 = n4005 ^ x31 ^ 1'b0 ;
  assign n36101 = ~n13416 & n36100 ;
  assign n36102 = n12207 & n36101 ;
  assign n36103 = ~n8792 & n36102 ;
  assign n36104 = n10384 & ~n16552 ;
  assign n36105 = n13027 & n17342 ;
  assign n36106 = n36105 ^ n30581 ^ 1'b0 ;
  assign n36107 = n2587 & n3483 ;
  assign n36108 = n2492 | n9807 ;
  assign n36109 = n21172 & ~n36108 ;
  assign n36110 = n36109 ^ n16319 ^ n12346 ;
  assign n36112 = ~n7049 & n7392 ;
  assign n36113 = n36112 ^ n8456 ^ 1'b0 ;
  assign n36114 = n4037 & n36113 ;
  assign n36115 = n1485 & n36114 ;
  assign n36116 = n9035 & n36115 ;
  assign n36111 = ~n3825 & n9250 ;
  assign n36117 = n36116 ^ n36111 ^ 1'b0 ;
  assign n36118 = n7793 ^ n2968 ^ 1'b0 ;
  assign n36119 = ~n14246 & n36118 ;
  assign n36120 = n5911 ^ n2548 ^ 1'b0 ;
  assign n36121 = ~n2857 & n36120 ;
  assign n36122 = ~n4035 & n10762 ;
  assign n36123 = n10100 ^ n3883 ^ 1'b0 ;
  assign n36124 = n8679 & ~n16952 ;
  assign n36125 = ~x27 & n36124 ;
  assign n36126 = n19725 ^ n7888 ^ 1'b0 ;
  assign n36127 = n20302 & n29432 ;
  assign n36128 = n36127 ^ n2541 ^ 1'b0 ;
  assign n36129 = ~n18611 & n36128 ;
  assign n36130 = n8049 & n36129 ;
  assign n36131 = n14072 ^ n3542 ^ 1'b0 ;
  assign n36132 = ~n9175 & n36131 ;
  assign n36133 = n677 & n36132 ;
  assign n36134 = ~n20450 & n25619 ;
  assign n36135 = ~n10501 & n36134 ;
  assign n36136 = n33413 & ~n36135 ;
  assign n36137 = n36136 ^ n32632 ^ 1'b0 ;
  assign n36138 = n1635 & ~n2061 ;
  assign n36139 = ~n3421 & n14041 ;
  assign n36140 = n12014 ^ n6330 ^ 1'b0 ;
  assign n36141 = n5175 & n36140 ;
  assign n36142 = n36141 ^ n1644 ^ 1'b0 ;
  assign n36143 = n36142 ^ n5189 ^ 1'b0 ;
  assign n36144 = n13383 & ~n28197 ;
  assign n36145 = ~n17525 & n36144 ;
  assign n36146 = n36145 ^ n17097 ^ 1'b0 ;
  assign n36147 = n33986 & ~n36146 ;
  assign n36148 = n22012 ^ n12145 ^ n2526 ;
  assign n36149 = n35695 ^ n35419 ^ 1'b0 ;
  assign n36150 = n5850 & n20876 ;
  assign n36151 = ~n4032 & n6526 ;
  assign n36152 = n36151 ^ n1098 ^ 1'b0 ;
  assign n36153 = ~n1859 & n12392 ;
  assign n36154 = n36152 & n36153 ;
  assign n36155 = n18274 | n36154 ;
  assign n36156 = n36155 ^ n16460 ^ 1'b0 ;
  assign n36157 = ~n30912 & n36156 ;
  assign n36158 = n36157 ^ x170 ^ 1'b0 ;
  assign n36159 = n36158 ^ n15391 ^ 1'b0 ;
  assign n36160 = n19555 & ~n36159 ;
  assign n36161 = ~n27517 & n32065 ;
  assign n36162 = n14841 ^ n3142 ^ 1'b0 ;
  assign n36163 = n9590 ^ n5569 ^ 1'b0 ;
  assign n36164 = ~n7195 & n36163 ;
  assign n36165 = ( n7395 & ~n11974 ) | ( n7395 & n36164 ) | ( ~n11974 & n36164 ) ;
  assign n36166 = n1754 & n36165 ;
  assign n36167 = n1271 & ~n24892 ;
  assign n36168 = n7161 ^ n849 ^ 1'b0 ;
  assign n36169 = n36168 ^ n17693 ^ 1'b0 ;
  assign n36170 = ~n1920 & n10440 ;
  assign n36171 = n36105 ^ n21103 ^ 1'b0 ;
  assign n36172 = n16598 | n36171 ;
  assign n36173 = n36172 ^ n33688 ^ 1'b0 ;
  assign n36174 = ~n6194 & n6542 ;
  assign n36175 = n36174 ^ n27017 ^ 1'b0 ;
  assign n36176 = ~n5403 & n6749 ;
  assign n36177 = x60 | n36019 ;
  assign n36182 = n796 | n32464 ;
  assign n36183 = n29157 & ~n36182 ;
  assign n36178 = n2689 | n4940 ;
  assign n36179 = n36178 ^ n3532 ^ 1'b0 ;
  assign n36180 = n36179 ^ n545 ^ 1'b0 ;
  assign n36181 = ~n21261 & n36180 ;
  assign n36184 = n36183 ^ n36181 ^ n4696 ;
  assign n36185 = n21221 & n36184 ;
  assign n36186 = n36185 ^ n19128 ^ 1'b0 ;
  assign n36187 = n20387 ^ n1154 ^ 1'b0 ;
  assign n36188 = n17294 ^ n2858 ^ 1'b0 ;
  assign n36189 = n438 & ~n36188 ;
  assign n36190 = ( ~n5376 & n13517 ) | ( ~n5376 & n31374 ) | ( n13517 & n31374 ) ;
  assign n36191 = n27564 | n33413 ;
  assign n36192 = n1658 & n6427 ;
  assign n36193 = n2019 & n36192 ;
  assign n36194 = n5703 | n23029 ;
  assign n36195 = n36194 ^ n10666 ^ 1'b0 ;
  assign n36196 = n36193 | n36195 ;
  assign n36197 = n10833 & n34443 ;
  assign n36198 = x113 | n16517 ;
  assign n36199 = n36198 ^ n10387 ^ 1'b0 ;
  assign n36200 = x232 | n17750 ;
  assign n36201 = n36200 ^ n3492 ^ 1'b0 ;
  assign n36202 = n5707 & n36201 ;
  assign n36203 = n20677 | n36202 ;
  assign n36204 = x180 & ~n36203 ;
  assign n36205 = n36204 ^ n18122 ^ 1'b0 ;
  assign n36206 = n22429 ^ n15866 ^ n11914 ;
  assign n36209 = n6637 & n13738 ;
  assign n36207 = n26160 ^ n6283 ^ 1'b0 ;
  assign n36208 = n33278 & n36207 ;
  assign n36210 = n36209 ^ n36208 ^ 1'b0 ;
  assign n36211 = n31883 ^ n22338 ^ 1'b0 ;
  assign n36212 = n13918 | n36211 ;
  assign n36213 = ~n1890 & n16015 ;
  assign n36214 = n10833 & ~n31119 ;
  assign n36215 = n36213 & n36214 ;
  assign n36216 = n13846 | n35138 ;
  assign n36217 = ~n917 & n5817 ;
  assign n36218 = n16132 ^ n10344 ^ 1'b0 ;
  assign n36219 = x128 & n32209 ;
  assign n36220 = n715 | n5286 ;
  assign n36221 = n36220 ^ n504 ^ 1'b0 ;
  assign n36222 = n34615 ^ n8963 ^ 1'b0 ;
  assign n36223 = n1591 | n12529 ;
  assign n36224 = n21504 | n36223 ;
  assign n36225 = ~n1898 & n4565 ;
  assign n36226 = ~n5648 & n28240 ;
  assign n36227 = ~n20708 & n25189 ;
  assign n36228 = n4701 ^ n4087 ^ 1'b0 ;
  assign n36229 = n631 & n8660 ;
  assign n36230 = n36229 ^ n1535 ^ 1'b0 ;
  assign n36231 = n11358 | n25614 ;
  assign n36232 = ~n532 & n3294 ;
  assign n36233 = n36232 ^ n14956 ^ 1'b0 ;
  assign n36234 = n12154 | n17722 ;
  assign n36235 = n36234 ^ x232 ^ 1'b0 ;
  assign n36236 = ~n36233 & n36235 ;
  assign n36237 = ~n2072 & n29852 ;
  assign n36238 = n36237 ^ n32655 ^ 1'b0 ;
  assign n36239 = n1974 | n29024 ;
  assign n36240 = n26090 ^ n9477 ^ 1'b0 ;
  assign n36241 = n8309 | n36240 ;
  assign n36242 = n31436 ^ n6375 ^ 1'b0 ;
  assign n36243 = n1635 | n24856 ;
  assign n36244 = n36243 ^ n5670 ^ 1'b0 ;
  assign n36245 = ~n8038 & n33513 ;
  assign n36246 = ~n3824 & n36245 ;
  assign n36247 = n1387 ^ n859 ^ 1'b0 ;
  assign n36248 = n6788 & ~n36247 ;
  assign n36249 = n36248 ^ n29478 ^ 1'b0 ;
  assign n36250 = n21427 | n36249 ;
  assign n36251 = n985 | n36250 ;
  assign n36252 = ( n3726 & n7621 ) | ( n3726 & n16646 ) | ( n7621 & n16646 ) ;
  assign n36253 = n17298 | n36252 ;
  assign n36254 = ~n1883 & n8824 ;
  assign n36255 = n36254 ^ n23132 ^ 1'b0 ;
  assign n36256 = ~n720 & n2764 ;
  assign n36257 = n36256 ^ n21443 ^ 1'b0 ;
  assign n36258 = n15323 & ~n36257 ;
  assign n36259 = ~n13913 & n36258 ;
  assign n36260 = n24099 ^ n6974 ^ 1'b0 ;
  assign n36261 = ~n1195 & n9314 ;
  assign n36262 = n18131 | n26465 ;
  assign n36263 = n36261 & ~n36262 ;
  assign n36264 = n15782 ^ n3153 ^ 1'b0 ;
  assign n36265 = n36264 ^ n29887 ^ 1'b0 ;
  assign n36266 = ~n3260 & n10306 ;
  assign n36267 = n23307 & n36266 ;
  assign n36268 = n7864 & n7910 ;
  assign n36269 = n36268 ^ n13167 ^ 1'b0 ;
  assign n36270 = n36269 ^ n30458 ^ n911 ;
  assign n36271 = n29504 ^ n5938 ^ 1'b0 ;
  assign n36272 = n6412 & n36271 ;
  assign n36273 = ~n18883 & n21416 ;
  assign n36274 = n13381 ^ n11074 ^ 1'b0 ;
  assign n36275 = ~n26828 & n36274 ;
  assign n36276 = n27744 ^ n5189 ^ 1'b0 ;
  assign n36277 = n20804 & n33507 ;
  assign n36278 = n3914 & n5471 ;
  assign n36279 = n4875 & ~n5027 ;
  assign n36280 = n29380 ^ n16463 ^ 1'b0 ;
  assign n36281 = ~n36279 & n36280 ;
  assign n36282 = ~n22986 & n26389 ;
  assign n36283 = n36282 ^ n25637 ^ 1'b0 ;
  assign n36284 = n10840 & n36283 ;
  assign n36285 = n1717 ^ n1573 ^ 1'b0 ;
  assign n36286 = ~n10014 & n15650 ;
  assign n36287 = n7761 ^ n5844 ^ n5190 ;
  assign n36288 = n4257 | n36287 ;
  assign n36289 = n6402 & ~n10182 ;
  assign n36290 = ~n9423 & n36289 ;
  assign n36291 = n1714 & ~n36290 ;
  assign n36292 = n36291 ^ n2091 ^ 1'b0 ;
  assign n36293 = ~n5923 & n11159 ;
  assign n36294 = n17218 ^ n10400 ^ 1'b0 ;
  assign n36295 = n3933 & ~n19913 ;
  assign n36296 = ~n5651 & n36295 ;
  assign n36297 = n16750 ^ n11149 ^ 1'b0 ;
  assign n36298 = n492 | n7721 ;
  assign n36299 = n11720 & n36298 ;
  assign n36300 = n12855 & ~n13252 ;
  assign n36301 = ~n1977 & n36300 ;
  assign n36302 = n18457 ^ n13845 ^ 1'b0 ;
  assign n36303 = n36301 | n36302 ;
  assign n36304 = n34414 ^ n14084 ^ 1'b0 ;
  assign n36305 = n15392 & n24645 ;
  assign n36306 = ~n19439 & n36305 ;
  assign n36307 = n4747 | n36306 ;
  assign n36308 = x121 ^ x65 ^ 1'b0 ;
  assign n36309 = n8474 ^ n4260 ^ 1'b0 ;
  assign n36310 = n8644 | n36309 ;
  assign n36311 = n1271 & n36310 ;
  assign n36312 = n36311 ^ n11085 ^ 1'b0 ;
  assign n36313 = ~n3166 & n14487 ;
  assign n36314 = n36313 ^ n19409 ^ 1'b0 ;
  assign n36315 = n1531 | n31157 ;
  assign n36316 = n36315 ^ n7907 ^ 1'b0 ;
  assign n36317 = n2275 & n18468 ;
  assign n36318 = n18191 & n36317 ;
  assign n36319 = n20895 ^ n15998 ^ 1'b0 ;
  assign n36320 = n34991 ^ n29040 ^ 1'b0 ;
  assign n36321 = n13455 ^ n7076 ^ n6222 ;
  assign n36322 = ~n3022 & n36321 ;
  assign n36323 = ~n35953 & n36322 ;
  assign n36324 = n2035 & n36120 ;
  assign n36325 = n36323 & n36324 ;
  assign n36326 = n2063 & ~n29507 ;
  assign n36327 = ~n3878 & n36326 ;
  assign n36328 = ~n9990 & n21645 ;
  assign n36329 = n36327 | n36328 ;
  assign n36330 = n1324 & n8742 ;
  assign n36331 = ~n8811 & n36330 ;
  assign n36332 = ~x245 & n15239 ;
  assign n36333 = n444 & ~n1239 ;
  assign n36334 = n36333 ^ n25702 ^ 1'b0 ;
  assign n36335 = n36334 ^ n13295 ^ n7074 ;
  assign n36336 = n19762 & n36335 ;
  assign n36337 = n4688 & n28367 ;
  assign n36338 = x95 & n14234 ;
  assign n36339 = n36338 ^ n12781 ^ 1'b0 ;
  assign n36340 = ~n18246 & n22068 ;
  assign n36341 = n36340 ^ n4534 ^ 1'b0 ;
  assign n36342 = n36339 & ~n36341 ;
  assign n36343 = n19439 ^ n2034 ^ 1'b0 ;
  assign n36344 = n397 & n36343 ;
  assign n36345 = n13473 | n16409 ;
  assign n36346 = n36344 | n36345 ;
  assign n36347 = n30866 & n36346 ;
  assign n36348 = n20089 ^ n14158 ^ 1'b0 ;
  assign n36349 = ~n10584 & n36348 ;
  assign n36350 = n14509 & n23042 ;
  assign n36351 = ~n36349 & n36350 ;
  assign n36352 = n9428 | n26858 ;
  assign n36353 = n5288 | n29831 ;
  assign n36354 = n36353 ^ n14424 ^ 1'b0 ;
  assign n36355 = n768 | n5867 ;
  assign n36356 = n14586 | n36355 ;
  assign n36357 = n13101 | n36356 ;
  assign n36358 = n12616 ^ n11004 ^ 1'b0 ;
  assign n36359 = n16357 & n19452 ;
  assign n36360 = ~n4246 & n36359 ;
  assign n36361 = n36360 ^ n18750 ^ 1'b0 ;
  assign n36362 = n5610 & ~n36361 ;
  assign n36363 = ~n18385 & n19319 ;
  assign n36364 = n27236 & ~n36363 ;
  assign n36365 = n26450 ^ n20414 ^ 1'b0 ;
  assign n36366 = n20015 | n36365 ;
  assign n36367 = n36366 ^ n12781 ^ 1'b0 ;
  assign n36368 = x67 & ~n36367 ;
  assign n36369 = n10389 ^ n1232 ^ 1'b0 ;
  assign n36370 = n36369 ^ n9430 ^ 1'b0 ;
  assign n36371 = n14580 | n36370 ;
  assign n36372 = ~n9324 & n21845 ;
  assign n36373 = ~n3348 & n36372 ;
  assign n36374 = ( n9786 & ~n9832 ) | ( n9786 & n10221 ) | ( ~n9832 & n10221 ) ;
  assign n36375 = n36374 ^ x64 ^ 1'b0 ;
  assign n36377 = n3974 ^ n2307 ^ 1'b0 ;
  assign n36376 = ~n8320 & n34798 ;
  assign n36378 = n36377 ^ n36376 ^ 1'b0 ;
  assign n36379 = n6935 & ~n22616 ;
  assign n36380 = ~n15644 & n15693 ;
  assign n36381 = n36380 ^ n6740 ^ 1'b0 ;
  assign n36382 = n13907 | n14689 ;
  assign n36383 = n11144 ^ n4733 ^ 1'b0 ;
  assign n36384 = n36382 | n36383 ;
  assign n36385 = n27448 | n36384 ;
  assign n36386 = ( n7214 & n8315 ) | ( n7214 & n22791 ) | ( n8315 & n22791 ) ;
  assign n36387 = n21040 | n36386 ;
  assign n36388 = x252 & ~n3437 ;
  assign n36389 = n36388 ^ n25882 ^ n3300 ;
  assign n36390 = ~n7003 & n15326 ;
  assign n36391 = n36390 ^ n13912 ^ 1'b0 ;
  assign n36392 = ~n2076 & n6343 ;
  assign n36393 = n6149 & n18882 ;
  assign n36394 = n8555 & n11373 ;
  assign n36395 = n36394 ^ n498 ^ 1'b0 ;
  assign n36396 = n1091 & ~n12757 ;
  assign n36397 = n1075 & ~n5909 ;
  assign n36398 = n19693 & n36397 ;
  assign n36399 = n36398 ^ n11519 ^ 1'b0 ;
  assign n36400 = n4882 ^ n3611 ^ 1'b0 ;
  assign n36401 = ~n6104 & n36400 ;
  assign n36402 = n36401 ^ n7308 ^ n6499 ;
  assign n36403 = ~n1667 & n3083 ;
  assign n36404 = ~n12590 & n36403 ;
  assign n36405 = n7703 & ~n36404 ;
  assign n36406 = n2711 & n36405 ;
  assign n36407 = n12148 ^ n6362 ^ 1'b0 ;
  assign n36408 = ~n13771 & n36407 ;
  assign n36409 = n19604 ^ n6883 ^ 1'b0 ;
  assign n36410 = n3368 & n34705 ;
  assign n36411 = n36410 ^ n9941 ^ 1'b0 ;
  assign n36412 = ( n18357 & n34498 ) | ( n18357 & ~n36411 ) | ( n34498 & ~n36411 ) ;
  assign n36413 = n21638 | n36334 ;
  assign n36416 = n14675 & n30706 ;
  assign n36417 = n36416 ^ n3437 ^ 1'b0 ;
  assign n36414 = n27581 ^ n6554 ^ 1'b0 ;
  assign n36415 = n5963 | n36414 ;
  assign n36418 = n36417 ^ n36415 ^ 1'b0 ;
  assign n36419 = n5983 ^ n4976 ^ n2920 ;
  assign n36420 = n36419 ^ n17412 ^ 1'b0 ;
  assign n36421 = n23539 ^ n14813 ^ n11685 ;
  assign n36422 = n36421 ^ n36033 ^ 1'b0 ;
  assign n36423 = x238 & n22412 ;
  assign n36424 = ~n11004 & n20572 ;
  assign n36425 = n36424 ^ n18286 ^ 1'b0 ;
  assign n36426 = n36425 ^ n17297 ^ 1'b0 ;
  assign n36427 = n1521 & ~n7331 ;
  assign n36428 = n36427 ^ n20528 ^ 1'b0 ;
  assign n36429 = n13763 & ~n36428 ;
  assign n36430 = x159 & ~n16184 ;
  assign n36431 = n1423 | n22961 ;
  assign n36432 = n10241 & n21967 ;
  assign n36433 = n26495 & ~n33031 ;
  assign n36434 = ( n4296 & n14680 ) | ( n4296 & n36433 ) | ( n14680 & n36433 ) ;
  assign n36435 = n25721 ^ n21226 ^ 1'b0 ;
  assign n36436 = n34016 | n36435 ;
  assign n36437 = n13437 | n36436 ;
  assign n36438 = n20358 ^ n7452 ^ n4283 ;
  assign n36439 = n4620 & n32903 ;
  assign n36440 = n25645 ^ n13968 ^ 1'b0 ;
  assign n36441 = ~n782 & n5952 ;
  assign n36442 = n10888 | n36441 ;
  assign n36443 = n20956 ^ n3529 ^ 1'b0 ;
  assign n36444 = n24781 & n36443 ;
  assign n36445 = ( n14397 & ~n15601 ) | ( n14397 & n18910 ) | ( ~n15601 & n18910 ) ;
  assign n36446 = ~n9778 & n34027 ;
  assign n36447 = n36446 ^ n5317 ^ 1'b0 ;
  assign n36448 = ~n10302 & n33264 ;
  assign n36449 = n14101 & ~n22431 ;
  assign n36450 = ( n8747 & n14023 ) | ( n8747 & ~n14707 ) | ( n14023 & ~n14707 ) ;
  assign n36451 = n36450 ^ n8507 ^ 1'b0 ;
  assign n36452 = n31392 | n36451 ;
  assign n36453 = n1623 & ~n32986 ;
  assign n36454 = ( n4796 & n10759 ) | ( n4796 & ~n14726 ) | ( n10759 & ~n14726 ) ;
  assign n36455 = ~n17782 & n36454 ;
  assign n36456 = n18619 ^ n6933 ^ 1'b0 ;
  assign n36457 = n1009 ^ x124 ^ 1'b0 ;
  assign n36458 = n7461 | n17014 ;
  assign n36459 = n36458 ^ n4955 ^ 1'b0 ;
  assign n36460 = n35595 ^ n2469 ^ 1'b0 ;
  assign n36461 = n6025 & ~n36460 ;
  assign n36462 = n17930 & ~n21241 ;
  assign n36463 = n19374 & n36462 ;
  assign n36464 = ~n3057 & n31830 ;
  assign n36465 = ~n4233 & n36464 ;
  assign n36466 = n9463 | n20788 ;
  assign n36467 = n36466 ^ n8668 ^ 1'b0 ;
  assign n36468 = n11616 & ~n13945 ;
  assign n36469 = ~n28439 & n36468 ;
  assign n36470 = ~n11115 & n36469 ;
  assign n36471 = n23837 ^ n10456 ^ 1'b0 ;
  assign n36472 = n23627 & ~n36471 ;
  assign n36473 = n3432 | n5197 ;
  assign n36474 = n36473 ^ n1643 ^ 1'b0 ;
  assign n36475 = n8331 & n36474 ;
  assign n36476 = n36475 ^ n8412 ^ 1'b0 ;
  assign n36477 = n1474 & ~n31414 ;
  assign n36478 = ~n3573 & n36477 ;
  assign n36480 = ~n11285 & n15690 ;
  assign n36479 = x63 & ~n10437 ;
  assign n36481 = n36480 ^ n36479 ^ 1'b0 ;
  assign n36482 = n33828 ^ x202 ^ 1'b0 ;
  assign n36484 = n19754 | n25314 ;
  assign n36485 = n36484 ^ n14871 ^ 1'b0 ;
  assign n36483 = n22393 ^ n17528 ^ 1'b0 ;
  assign n36486 = n36485 ^ n36483 ^ 1'b0 ;
  assign n36487 = n33732 | n36486 ;
  assign n36488 = n33470 ^ n5135 ^ 1'b0 ;
  assign n36489 = n994 & n13184 ;
  assign n36490 = n36489 ^ n5564 ^ 1'b0 ;
  assign n36491 = n16818 | n19643 ;
  assign n36492 = n4726 & n5619 ;
  assign n36493 = n30269 & n36492 ;
  assign n36494 = ~n4995 & n36493 ;
  assign n36495 = n32478 ^ n22715 ^ n16824 ;
  assign n36496 = n12427 & n36495 ;
  assign n36497 = ~n6590 & n36496 ;
  assign n36498 = n15122 & ~n15743 ;
  assign n36499 = n36498 ^ n23888 ^ 1'b0 ;
  assign n36500 = n17463 & ~n36499 ;
  assign n36501 = n7794 & ~n15304 ;
  assign n36502 = n3237 | n36501 ;
  assign n36503 = n36502 ^ n6205 ^ 1'b0 ;
  assign n36504 = n12205 ^ n9105 ^ 1'b0 ;
  assign n36505 = n1880 & n36504 ;
  assign n36506 = n36505 ^ n9432 ^ 1'b0 ;
  assign n36507 = n10705 ^ n1709 ^ 1'b0 ;
  assign n36508 = n36506 | n36507 ;
  assign n36509 = n36508 ^ n29640 ^ 1'b0 ;
  assign n36510 = n36503 | n36509 ;
  assign n36511 = ~n6001 & n23856 ;
  assign n36514 = x55 & n630 ;
  assign n36515 = ~n630 & n36514 ;
  assign n36516 = n1575 | n36515 ;
  assign n36517 = n36515 & ~n36516 ;
  assign n36518 = n32998 & ~n36517 ;
  assign n36526 = x74 & n575 ;
  assign n36527 = n12109 & n36526 ;
  assign n36519 = ~n608 & n14723 ;
  assign n36520 = n2266 | n3931 ;
  assign n36521 = n3931 & ~n36520 ;
  assign n36522 = n1713 & ~n36521 ;
  assign n36523 = n36521 & n36522 ;
  assign n36524 = ~n8765 & n36523 ;
  assign n36525 = ~n36519 & n36524 ;
  assign n36528 = n36527 ^ n36525 ^ 1'b0 ;
  assign n36529 = ~n6994 & n36528 ;
  assign n36530 = n36518 & n36529 ;
  assign n36531 = n36530 ^ x132 ^ 1'b0 ;
  assign n36512 = ~n7771 & n8438 ;
  assign n36513 = n19468 & ~n36512 ;
  assign n36532 = n36531 ^ n36513 ^ 1'b0 ;
  assign n36533 = n1988 & n25343 ;
  assign n36534 = n33239 ^ n30631 ^ 1'b0 ;
  assign n36535 = n9580 | n19515 ;
  assign n36536 = n35236 | n36535 ;
  assign n36537 = n36536 ^ n9133 ^ 1'b0 ;
  assign n36538 = n10162 ^ n4980 ^ 1'b0 ;
  assign n36539 = n8916 | n36264 ;
  assign n36540 = ~n846 & n4596 ;
  assign n36541 = n36540 ^ n6766 ^ 1'b0 ;
  assign n36542 = n36541 ^ n4366 ^ 1'b0 ;
  assign n36543 = ~n5869 & n28585 ;
  assign n36545 = n15737 & ~n18760 ;
  assign n36544 = n16968 | n28652 ;
  assign n36546 = n36545 ^ n36544 ^ 1'b0 ;
  assign n36550 = n16968 & ~n31343 ;
  assign n36547 = n8087 | n8890 ;
  assign n36548 = n36512 | n36547 ;
  assign n36549 = n7350 & ~n36548 ;
  assign n36551 = n36550 ^ n36549 ^ 1'b0 ;
  assign n36552 = n10383 & n14590 ;
  assign n36553 = n36552 ^ n1240 ^ 1'b0 ;
  assign n36554 = n923 | n25188 ;
  assign n36555 = n36554 ^ n18471 ^ 1'b0 ;
  assign n36556 = n5656 | n10553 ;
  assign n36557 = n36555 & ~n36556 ;
  assign n36558 = n2225 ^ n1863 ^ 1'b0 ;
  assign n36559 = n12287 & n36558 ;
  assign n36560 = ( n13265 & n31217 ) | ( n13265 & n36559 ) | ( n31217 & n36559 ) ;
  assign n36561 = n28829 | n36560 ;
  assign n36562 = n36557 & ~n36561 ;
  assign n36563 = n1499 | n19856 ;
  assign n36564 = n23892 & ~n36563 ;
  assign n36565 = n28861 & ~n36564 ;
  assign n36566 = n15101 ^ n8543 ^ 1'b0 ;
  assign n36567 = x162 & n36566 ;
  assign n36568 = n24286 ^ x174 ^ 1'b0 ;
  assign n36569 = n15243 & n36057 ;
  assign n36570 = n36569 ^ n2335 ^ 1'b0 ;
  assign n36571 = n17331 & n36321 ;
  assign n36572 = n4824 & n36571 ;
  assign n36573 = n26774 ^ n9364 ^ 1'b0 ;
  assign n36574 = n16072 ^ n1239 ^ 1'b0 ;
  assign n36575 = n3933 & n36574 ;
  assign n36576 = n11659 | n36575 ;
  assign n36577 = n14820 | n19229 ;
  assign n36578 = n9386 & ~n36577 ;
  assign n36579 = n10762 & ~n29343 ;
  assign n36580 = n36579 ^ n7278 ^ 1'b0 ;
  assign n36581 = n36580 ^ n815 ^ 1'b0 ;
  assign n36582 = n10492 & ~n36581 ;
  assign n36583 = n36582 ^ n10689 ^ 1'b0 ;
  assign n36584 = n4327 | n31881 ;
  assign n36585 = n25960 | n36584 ;
  assign n36586 = n29285 & ~n30002 ;
  assign n36587 = n36586 ^ n35800 ^ 1'b0 ;
  assign n36590 = n9977 ^ n2696 ^ 1'b0 ;
  assign n36588 = n21064 ^ n978 ^ 1'b0 ;
  assign n36589 = n951 & n36588 ;
  assign n36591 = n36590 ^ n36589 ^ n16862 ;
  assign n36592 = n1473 | n1974 ;
  assign n36593 = n1974 & ~n36592 ;
  assign n36594 = n1485 | n36593 ;
  assign n36595 = n36594 ^ n28073 ^ 1'b0 ;
  assign n36596 = n3405 & ~n36595 ;
  assign n36597 = ~n10803 & n36596 ;
  assign n36598 = n23773 & n29762 ;
  assign n36599 = n36598 ^ n3979 ^ 1'b0 ;
  assign n36600 = n13629 | n24434 ;
  assign n36601 = n12792 ^ n816 ^ 1'b0 ;
  assign n36602 = n10883 | n15800 ;
  assign n36603 = n25545 & ~n36602 ;
  assign n36604 = n14605 ^ n11873 ^ 1'b0 ;
  assign n36605 = n1111 & ~n36604 ;
  assign n36606 = n14404 & n33513 ;
  assign n36607 = n36047 & n36606 ;
  assign n36608 = ~n36605 & n36607 ;
  assign n36610 = ~n3939 & n8127 ;
  assign n36609 = n1507 & ~n23833 ;
  assign n36611 = n36610 ^ n36609 ^ 1'b0 ;
  assign n36612 = n36611 ^ n27100 ^ n4862 ;
  assign n36613 = n29678 ^ n2778 ^ 1'b0 ;
  assign n36615 = ~n4940 & n10314 ;
  assign n36614 = x106 & ~n1304 ;
  assign n36616 = n36615 ^ n36614 ^ 1'b0 ;
  assign n36617 = ~n3574 & n20408 ;
  assign n36618 = n36617 ^ n34651 ^ 1'b0 ;
  assign n36619 = n36259 & ~n36618 ;
  assign n36620 = ~n15913 & n36619 ;
  assign n36621 = n31402 ^ n26110 ^ 1'b0 ;
  assign n36622 = n14953 & ~n36621 ;
  assign n36623 = n19479 & n25708 ;
  assign n36624 = n1337 & n32136 ;
  assign n36625 = n36624 ^ n20871 ^ 1'b0 ;
  assign n36626 = n36090 ^ n1507 ^ 1'b0 ;
  assign n36627 = ~n19227 & n36626 ;
  assign n36630 = n12645 & ~n15351 ;
  assign n36629 = ~n7892 & n10376 ;
  assign n36631 = n36630 ^ n36629 ^ 1'b0 ;
  assign n36628 = n17470 & ~n34898 ;
  assign n36632 = n36631 ^ n36628 ^ 1'b0 ;
  assign n36633 = ~n27894 & n36495 ;
  assign n36634 = n36633 ^ n9057 ^ 1'b0 ;
  assign n36635 = n36634 ^ n28491 ^ 1'b0 ;
  assign n36636 = n27209 & n36635 ;
  assign n36637 = n30598 ^ n20351 ^ n15014 ;
  assign n36638 = ~n36636 & n36637 ;
  assign n36639 = n3516 & n14959 ;
  assign n36640 = n3097 | n6028 ;
  assign n36641 = n36640 ^ n12901 ^ 1'b0 ;
  assign n36642 = n3143 & ~n36641 ;
  assign n36643 = n623 & n36642 ;
  assign n36644 = n1658 | n36156 ;
  assign n36645 = n7662 ^ n4021 ^ 1'b0 ;
  assign n36646 = n6635 | n36645 ;
  assign n36648 = n559 & ~n31340 ;
  assign n36649 = n36648 ^ n6772 ^ 1'b0 ;
  assign n36647 = n27835 & ~n36437 ;
  assign n36650 = n36649 ^ n36647 ^ 1'b0 ;
  assign n36651 = ~n4327 & n20228 ;
  assign n36652 = n36651 ^ n7081 ^ 1'b0 ;
  assign n36653 = n5140 & n36652 ;
  assign n36654 = n6522 & n36653 ;
  assign n36655 = n11461 & ~n15430 ;
  assign n36656 = n36655 ^ n13104 ^ 1'b0 ;
  assign n36657 = n7959 ^ n1872 ^ n1237 ;
  assign n36658 = n36657 ^ n4059 ^ 1'b0 ;
  assign n36659 = n9143 & ~n10458 ;
  assign n36660 = n36659 ^ n16927 ^ 1'b0 ;
  assign n36661 = n7153 | n9178 ;
  assign n36662 = n31698 ^ n2955 ^ 1'b0 ;
  assign n36663 = n7749 & n22287 ;
  assign n36664 = n3565 | n4738 ;
  assign n36665 = n36664 ^ n3566 ^ 1'b0 ;
  assign n36666 = n36665 ^ n10294 ^ 1'b0 ;
  assign n36667 = n11111 | n17488 ;
  assign n36668 = ~n20241 & n36667 ;
  assign n36669 = n18519 ^ x251 ^ 1'b0 ;
  assign n36670 = n14974 ^ n1693 ^ 1'b0 ;
  assign n36671 = n36669 | n36670 ;
  assign n36672 = n21927 & ~n36671 ;
  assign n36673 = ~n5974 & n36672 ;
  assign n36674 = ~n7383 & n16856 ;
  assign n36675 = ~n4095 & n5368 ;
  assign n36676 = n1214 & n6342 ;
  assign n36677 = ~n18157 & n36676 ;
  assign n36678 = n36677 ^ n31941 ^ 1'b0 ;
  assign n36679 = ~n7411 & n36678 ;
  assign n36680 = n4791 & ~n17549 ;
  assign n36681 = n4804 & n36680 ;
  assign n36682 = n23761 & ~n36681 ;
  assign n36683 = n34181 ^ n24796 ^ 1'b0 ;
  assign n36684 = n36682 & n36683 ;
  assign n36685 = n16907 ^ n6834 ^ n5398 ;
  assign n36686 = n5122 | n6845 ;
  assign n36687 = n19211 & n36686 ;
  assign n36688 = n587 | n12557 ;
  assign n36689 = n36688 ^ n27747 ^ 1'b0 ;
  assign n36690 = n6969 | n17752 ;
  assign n36691 = n36690 ^ n5375 ^ 1'b0 ;
  assign n36692 = n36071 ^ n7189 ^ 1'b0 ;
  assign n36693 = n36691 | n36692 ;
  assign n36695 = n12504 & n14834 ;
  assign n36694 = n5619 & ~n35638 ;
  assign n36696 = n36695 ^ n36694 ^ 1'b0 ;
  assign n36697 = n35399 ^ n20538 ^ 1'b0 ;
  assign n36698 = n32146 ^ n6019 ^ 1'b0 ;
  assign n36699 = n12520 & ~n18453 ;
  assign n36700 = ~n36698 & n36699 ;
  assign n36701 = n27169 & ~n36700 ;
  assign n36702 = ~n7781 & n22641 ;
  assign n36703 = n27587 & n36702 ;
  assign n36704 = n34660 ^ n7376 ^ n2225 ;
  assign n36705 = n2371 | n6210 ;
  assign n36706 = n4881 & n35172 ;
  assign n36707 = n36705 & n36706 ;
  assign n36708 = n298 & n8033 ;
  assign n36709 = n9458 ^ n8169 ^ 1'b0 ;
  assign n36710 = n1740 & n1926 ;
  assign n36711 = n36710 ^ n5896 ^ 1'b0 ;
  assign n36712 = n395 | n840 ;
  assign n36713 = n36712 ^ n3318 ^ n860 ;
  assign n36714 = n36711 | n36713 ;
  assign n36715 = n26263 & n36714 ;
  assign n36716 = n3652 & n14417 ;
  assign n36717 = n12763 | n36716 ;
  assign n36718 = n8612 & ~n36717 ;
  assign n36719 = n5670 & ~n8028 ;
  assign n36720 = n36718 & n36719 ;
  assign n36721 = n13455 & ~n25269 ;
  assign n36722 = n22494 ^ n19059 ^ 1'b0 ;
  assign n36723 = n18783 & n36722 ;
  assign n36724 = n1588 | n36723 ;
  assign n36725 = n36721 | n36724 ;
  assign n36726 = n4506 ^ n2541 ^ 1'b0 ;
  assign n36727 = n36726 ^ n34408 ^ 1'b0 ;
  assign n36728 = n10382 | n36727 ;
  assign n36729 = n19250 & ~n28095 ;
  assign n36730 = n18492 ^ n7533 ^ 1'b0 ;
  assign n36731 = n36729 | n36730 ;
  assign n36732 = n18820 ^ n16305 ^ 1'b0 ;
  assign n36734 = n5496 & n5909 ;
  assign n36733 = ~n3593 & n6486 ;
  assign n36735 = n36734 ^ n36733 ^ 1'b0 ;
  assign n36736 = n11770 | n18854 ;
  assign n36737 = n36736 ^ n8298 ^ 1'b0 ;
  assign n36738 = n36737 ^ n20444 ^ 1'b0 ;
  assign n36739 = ~n7813 & n10210 ;
  assign n36740 = n3980 & n36739 ;
  assign n36742 = n8665 & ~n10647 ;
  assign n36743 = ~n10657 & n36742 ;
  assign n36741 = n28032 & ~n33428 ;
  assign n36744 = n36743 ^ n36741 ^ 1'b0 ;
  assign n36748 = n2411 & n11454 ;
  assign n36749 = n36748 ^ n12041 ^ 1'b0 ;
  assign n36750 = ( n8443 & n29928 ) | ( n8443 & n36749 ) | ( n29928 & n36749 ) ;
  assign n36751 = ( x106 & n13697 ) | ( x106 & ~n36750 ) | ( n13697 & ~n36750 ) ;
  assign n36745 = ~n4575 & n26145 ;
  assign n36746 = n3935 & n36745 ;
  assign n36747 = n16555 | n36746 ;
  assign n36752 = n36751 ^ n36747 ^ 1'b0 ;
  assign n36753 = n6836 | n10904 ;
  assign n36754 = n36753 ^ n26985 ^ 1'b0 ;
  assign n36755 = ~n9870 & n36750 ;
  assign n36756 = n2482 & n13854 ;
  assign n36757 = n36756 ^ x140 ^ 1'b0 ;
  assign n36758 = ~n3973 & n36757 ;
  assign n36759 = n23862 ^ n12184 ^ 1'b0 ;
  assign n36760 = ~n27163 & n36759 ;
  assign n36761 = n1697 & n36760 ;
  assign n36762 = n12329 & n23691 ;
  assign n36763 = n36762 ^ n5000 ^ 1'b0 ;
  assign n36764 = n10220 ^ x26 ^ 1'b0 ;
  assign n36765 = ~n30607 & n36764 ;
  assign n36766 = n12825 ^ n5574 ^ 1'b0 ;
  assign n36767 = n36765 & n36766 ;
  assign n36768 = n2013 & ~n7204 ;
  assign n36769 = ~n4961 & n36768 ;
  assign n36770 = n3914 & ~n12051 ;
  assign n36771 = n36770 ^ n11580 ^ 1'b0 ;
  assign n36772 = ~n3910 & n36771 ;
  assign n36773 = n703 | n7364 ;
  assign n36774 = n15139 | n19821 ;
  assign n36775 = ~n10888 & n16627 ;
  assign n36776 = n3953 & ~n3963 ;
  assign n36777 = n5756 ^ n2310 ^ 1'b0 ;
  assign n36778 = n36776 & n36777 ;
  assign n36779 = ~n16523 & n36778 ;
  assign n36780 = n1964 | n15258 ;
  assign n36781 = n1964 & ~n36780 ;
  assign n36782 = n13072 | n33792 ;
  assign n36783 = n10092 ^ n5691 ^ 1'b0 ;
  assign n36784 = n373 & ~n1199 ;
  assign n36785 = n8080 | n8094 ;
  assign n36786 = n1239 & ~n36785 ;
  assign n36787 = ~n36784 & n36786 ;
  assign n36788 = n11965 & n36787 ;
  assign n36789 = n4432 ^ n1812 ^ 1'b0 ;
  assign n36790 = n1841 & ~n36789 ;
  assign n36791 = n36790 ^ n22885 ^ n10638 ;
  assign n36792 = n4814 & ~n23371 ;
  assign n36793 = n5456 & ~n8181 ;
  assign n36794 = n14803 & ~n32706 ;
  assign n36795 = ~n36793 & n36794 ;
  assign n36796 = ~n10357 & n11402 ;
  assign n36797 = n6360 | n16870 ;
  assign n36798 = n32160 ^ n3984 ^ 1'b0 ;
  assign n36799 = n19275 | n32943 ;
  assign n36800 = n13696 ^ n4400 ^ 1'b0 ;
  assign n36801 = n1399 & ~n3666 ;
  assign n36802 = n32487 ^ n16152 ^ 1'b0 ;
  assign n36803 = n36801 | n36802 ;
  assign n36804 = ~n18926 & n24404 ;
  assign n36805 = n36804 ^ n3950 ^ 1'b0 ;
  assign n36806 = n21297 & ~n36805 ;
  assign n36807 = n36806 ^ n20220 ^ 1'b0 ;
  assign n36808 = ~n6025 & n7567 ;
  assign n36809 = n36808 ^ n19674 ^ 1'b0 ;
  assign n36810 = ~n7109 & n7953 ;
  assign n36811 = n36810 ^ n23648 ^ 1'b0 ;
  assign n36812 = ~n2037 & n27890 ;
  assign n36813 = ~n1091 & n36812 ;
  assign n36814 = n2757 | n15965 ;
  assign n36815 = n21827 & ~n36814 ;
  assign n36816 = n11439 | n36815 ;
  assign n36817 = n12144 | n29572 ;
  assign n36818 = n2227 & ~n5690 ;
  assign n36819 = n4112 | n35818 ;
  assign n36820 = n36819 ^ n10022 ^ 1'b0 ;
  assign n36821 = n20257 ^ n15453 ^ 1'b0 ;
  assign n36822 = n21815 ^ n7736 ^ 1'b0 ;
  assign n36823 = n36821 & n36822 ;
  assign n36824 = n12093 ^ n11373 ^ 1'b0 ;
  assign n36825 = n7996 & ~n31061 ;
  assign n36826 = n36649 ^ n3963 ^ 1'b0 ;
  assign n36827 = n6516 & n6983 ;
  assign n36828 = ~n15185 & n36827 ;
  assign n36829 = n5507 | n12865 ;
  assign n36830 = n8293 & ~n36829 ;
  assign n36831 = n16007 | n36830 ;
  assign n36832 = ~n4688 & n10980 ;
  assign n36833 = n8704 & ~n12671 ;
  assign n36834 = n5840 & n36833 ;
  assign n36835 = n36834 ^ n6005 ^ 1'b0 ;
  assign n36836 = n10068 | n19273 ;
  assign n36837 = n4497 | n33861 ;
  assign n36838 = n36837 ^ n22588 ^ 1'b0 ;
  assign n36839 = n7414 & ~n15136 ;
  assign n36840 = ~n3281 & n36839 ;
  assign n36841 = n12813 & ~n29012 ;
  assign n36844 = ~n951 & n31261 ;
  assign n36845 = n15618 & n36844 ;
  assign n36842 = ~n1205 & n5588 ;
  assign n36843 = ~n21274 & n36842 ;
  assign n36846 = n36845 ^ n36843 ^ 1'b0 ;
  assign n36847 = ( n3645 & n6443 ) | ( n3645 & n23995 ) | ( n6443 & n23995 ) ;
  assign n36848 = n1079 | n21376 ;
  assign n36849 = n36848 ^ n5983 ^ 1'b0 ;
  assign n36850 = n21527 ^ n6872 ^ n2087 ;
  assign n36851 = n2078 & ~n36850 ;
  assign n36852 = n257 & ~n25774 ;
  assign n36853 = n31551 & ~n36852 ;
  assign n36854 = n27121 ^ n12324 ^ 1'b0 ;
  assign n36855 = n34447 ^ n25172 ^ 1'b0 ;
  assign n36856 = n2068 & n28186 ;
  assign n36857 = n16842 & ~n30340 ;
  assign n36858 = n3473 & n12247 ;
  assign n36859 = n2078 & n36858 ;
  assign n36860 = n36859 ^ n17605 ^ 1'b0 ;
  assign n36861 = ~n14157 & n23275 ;
  assign n36862 = n33485 | n36861 ;
  assign n36863 = n36860 | n36862 ;
  assign n36864 = ( n17897 & n36857 ) | ( n17897 & ~n36863 ) | ( n36857 & ~n36863 ) ;
  assign n36865 = n32771 ^ n3134 ^ 1'b0 ;
  assign n36866 = ~n7323 & n36865 ;
  assign n36867 = x112 & ~n9256 ;
  assign n36868 = n36867 ^ n12193 ^ 1'b0 ;
  assign n36869 = n1707 & ~n2669 ;
  assign n36870 = n3346 & ~n36869 ;
  assign n36871 = ( n2449 & n26527 ) | ( n2449 & n36870 ) | ( n26527 & n36870 ) ;
  assign n36872 = n19544 ^ n1808 ^ 1'b0 ;
  assign n36873 = n8092 | n11134 ;
  assign n36874 = n20253 | n36873 ;
  assign n36875 = ~n13629 & n36874 ;
  assign n36876 = ~n29162 & n36875 ;
  assign n36877 = n2119 & ~n20569 ;
  assign n36878 = n16019 ^ n8089 ^ 1'b0 ;
  assign n36879 = n36877 & ~n36878 ;
  assign n36880 = n31554 ^ n20808 ^ 1'b0 ;
  assign n36881 = n2055 & ~n36880 ;
  assign n36882 = n6281 ^ n5723 ^ 1'b0 ;
  assign n36883 = n36881 & ~n36882 ;
  assign n36884 = n22926 ^ n3583 ^ 1'b0 ;
  assign n36885 = n14298 | n36884 ;
  assign n36886 = ~n32219 & n36885 ;
  assign n36888 = n18477 ^ n3948 ^ x31 ;
  assign n36887 = n15204 ^ n4657 ^ n4416 ;
  assign n36889 = n36888 ^ n36887 ^ n19774 ;
  assign n36890 = n15260 & ~n15824 ;
  assign n36891 = ~n36495 & n36890 ;
  assign n36892 = n11514 | n32184 ;
  assign n36893 = n7113 | n15624 ;
  assign n36894 = n11890 & n36893 ;
  assign n36895 = ~n13698 & n36894 ;
  assign n36896 = n21093 ^ n9857 ^ 1'b0 ;
  assign n36897 = n562 | n36896 ;
  assign n36898 = n11136 & ~n25785 ;
  assign n36899 = ~n20094 & n36898 ;
  assign n36900 = ~n4214 & n23815 ;
  assign n36901 = ( n15315 & n15537 ) | ( n15315 & n27398 ) | ( n15537 & n27398 ) ;
  assign n36902 = n15673 ^ n4051 ^ 1'b0 ;
  assign n36903 = n2106 & ~n36902 ;
  assign n36904 = ~n21967 & n36903 ;
  assign n36905 = n9590 & n36904 ;
  assign n36906 = n36905 ^ n13934 ^ 1'b0 ;
  assign n36907 = n741 | n36906 ;
  assign n36908 = n36907 ^ n29047 ^ 1'b0 ;
  assign n36909 = n31450 ^ n20024 ^ n12352 ;
  assign n36910 = n34194 & n36909 ;
  assign n36911 = n5188 & n27695 ;
  assign n36912 = n2861 & n36911 ;
  assign n36913 = n8412 | n20145 ;
  assign n36914 = n7824 & n25738 ;
  assign n36915 = n17449 ^ n4647 ^ 1'b0 ;
  assign n36916 = n16939 | n36915 ;
  assign n36919 = n6031 ^ n3666 ^ 1'b0 ;
  assign n36917 = n12448 & n32901 ;
  assign n36918 = n36917 ^ n7368 ^ 1'b0 ;
  assign n36920 = n36919 ^ n36918 ^ 1'b0 ;
  assign n36921 = ~n18812 & n36920 ;
  assign n36924 = ~n2753 & n4787 ;
  assign n36925 = n7415 ^ n4293 ^ 1'b0 ;
  assign n36926 = n36924 | n36925 ;
  assign n36922 = n3966 ^ n2860 ^ 1'b0 ;
  assign n36923 = ~n21033 & n36922 ;
  assign n36927 = n36926 ^ n36923 ^ 1'b0 ;
  assign n36928 = n27212 ^ n17748 ^ 1'b0 ;
  assign n36929 = n6264 & n23696 ;
  assign n36930 = ~n36928 & n36929 ;
  assign n36931 = n807 & ~n5277 ;
  assign n36932 = n6091 & ~n16337 ;
  assign n36933 = n36932 ^ n19604 ^ 1'b0 ;
  assign n36934 = ~n2846 & n8703 ;
  assign n36935 = n36934 ^ n20183 ^ n13572 ;
  assign n36936 = n6570 & n8818 ;
  assign n36937 = x170 & n32813 ;
  assign n36938 = n36937 ^ n8770 ^ 1'b0 ;
  assign n36939 = n25643 ^ n8673 ^ 1'b0 ;
  assign n36940 = n17586 ^ n6647 ^ 1'b0 ;
  assign n36941 = n9033 & ~n36940 ;
  assign n36942 = n36941 ^ n14876 ^ 1'b0 ;
  assign n36943 = n1512 & ~n2983 ;
  assign n36944 = ~n36942 & n36943 ;
  assign n36945 = n24695 ^ n22895 ^ 1'b0 ;
  assign n36946 = ~n18840 & n36945 ;
  assign n36947 = n16188 & ~n36946 ;
  assign n36948 = ~n19265 & n36947 ;
  assign n36949 = n10403 ^ n2589 ^ 1'b0 ;
  assign n36950 = n3187 & ~n5988 ;
  assign n36951 = n20782 ^ n11205 ^ 1'b0 ;
  assign n36952 = n16390 | n19976 ;
  assign n36953 = n19533 & n36952 ;
  assign n36954 = n32546 ^ n1950 ^ 1'b0 ;
  assign n36955 = ~n14359 & n36954 ;
  assign n36956 = n4721 & ~n16954 ;
  assign n36957 = ~n15018 & n36956 ;
  assign n36958 = n14867 ^ n5026 ^ 1'b0 ;
  assign n36959 = ~n11058 & n36958 ;
  assign n36960 = ~n17255 & n36959 ;
  assign n36961 = n14587 & n36960 ;
  assign n36962 = n36961 ^ n19506 ^ 1'b0 ;
  assign n36963 = n4499 ^ n546 ^ 1'b0 ;
  assign n36964 = n2068 & n36963 ;
  assign n36965 = ~n7179 & n36964 ;
  assign n36966 = n8401 ^ n602 ^ 1'b0 ;
  assign n36967 = n1326 | n2892 ;
  assign n36968 = n5056 & ~n36967 ;
  assign n36969 = ~n18854 & n36968 ;
  assign n36970 = ( n17179 & n22180 ) | ( n17179 & n36969 ) | ( n22180 & n36969 ) ;
  assign n36971 = ~n14861 & n16716 ;
  assign n36972 = ~n1062 & n36971 ;
  assign n36973 = n3045 & ~n36972 ;
  assign n36974 = n35332 & n36973 ;
  assign n36975 = ~n1628 & n26392 ;
  assign n36976 = n18502 & n36975 ;
  assign n36977 = n6553 & ~n31854 ;
  assign n36978 = n36976 & n36977 ;
  assign n36980 = n8263 | n9966 ;
  assign n36979 = ~n23279 & n26679 ;
  assign n36981 = n36980 ^ n36979 ^ 1'b0 ;
  assign n36982 = n3963 ^ n302 ^ 1'b0 ;
  assign n36983 = n15589 | n36982 ;
  assign n36984 = n33069 | n36983 ;
  assign n36985 = ~n3574 & n6065 ;
  assign n36986 = n36985 ^ n10443 ^ 1'b0 ;
  assign n36987 = n36986 ^ n9256 ^ n1643 ;
  assign n36988 = ~n22616 & n35123 ;
  assign n36989 = n32225 & n36988 ;
  assign n36990 = ~n25003 & n36989 ;
  assign n36991 = n2296 | n18028 ;
  assign n36992 = n36991 ^ n10663 ^ 1'b0 ;
  assign n36996 = n35209 ^ n8333 ^ 1'b0 ;
  assign n36993 = n5305 | n22885 ;
  assign n36994 = n19774 | n36993 ;
  assign n36995 = n15854 & n36994 ;
  assign n36997 = n36996 ^ n36995 ^ 1'b0 ;
  assign n37000 = n14549 ^ n1038 ^ 1'b0 ;
  assign n36998 = n11894 & ~n26104 ;
  assign n36999 = n8464 & n36998 ;
  assign n37001 = n37000 ^ n36999 ^ 1'b0 ;
  assign n37002 = ~n7049 & n12714 ;
  assign n37003 = n9191 ^ n8225 ^ 1'b0 ;
  assign n37004 = n28640 & n32866 ;
  assign n37005 = x92 & n30104 ;
  assign n37006 = n1278 & n21042 ;
  assign n37007 = n37006 ^ n3817 ^ 1'b0 ;
  assign n37008 = n8532 & ~n37007 ;
  assign n37009 = ~n1566 & n34153 ;
  assign n37010 = n37008 & n37009 ;
  assign n37011 = n23084 ^ n19774 ^ 1'b0 ;
  assign n37012 = n3740 | n37011 ;
  assign n37013 = n10560 | n11143 ;
  assign n37014 = n1764 | n37013 ;
  assign n37015 = n27271 ^ n4289 ^ 1'b0 ;
  assign n37016 = n16375 & ~n37015 ;
  assign n37017 = n37016 ^ n16197 ^ 1'b0 ;
  assign n37018 = n11865 ^ n9118 ^ n2324 ;
  assign n37019 = n13867 | n37018 ;
  assign n37020 = n4372 | n16045 ;
  assign n37021 = n35966 ^ n8088 ^ 1'b0 ;
  assign n37022 = n30962 ^ n20713 ^ 1'b0 ;
  assign n37023 = n1825 & ~n6531 ;
  assign n37024 = n10579 ^ x196 ^ 1'b0 ;
  assign n37025 = x88 & n37024 ;
  assign n37026 = n6017 | n25094 ;
  assign n37027 = ( n2212 & n32505 ) | ( n2212 & ~n37026 ) | ( n32505 & ~n37026 ) ;
  assign n37028 = n1252 & n20657 ;
  assign n37029 = n7937 & n12904 ;
  assign n37030 = n35850 & n37029 ;
  assign n37031 = ~n2643 & n12888 ;
  assign n37032 = ~n13837 & n33989 ;
  assign n37033 = ~n37031 & n37032 ;
  assign n37034 = n20685 ^ n5903 ^ 1'b0 ;
  assign n37035 = n14430 & ~n15678 ;
  assign n37036 = n22995 & n29938 ;
  assign n37037 = n19275 ^ n18061 ^ 1'b0 ;
  assign n37038 = n33587 ^ n14247 ^ 1'b0 ;
  assign n37039 = n6882 & n10525 ;
  assign n37040 = n37038 & n37039 ;
  assign n37041 = n37037 & ~n37040 ;
  assign n37042 = n1048 & ~n37041 ;
  assign n37043 = ~n683 & n31766 ;
  assign n37044 = ~n7163 & n37043 ;
  assign n37045 = n6298 | n22331 ;
  assign n37046 = n29064 & ~n37045 ;
  assign n37047 = n7796 & ~n8481 ;
  assign n37048 = ~n4191 & n37047 ;
  assign n37049 = n17217 ^ n11284 ^ 1'b0 ;
  assign n37050 = ~n15359 & n37049 ;
  assign n37051 = ~n10757 & n30813 ;
  assign n37052 = n37051 ^ n36615 ^ 1'b0 ;
  assign n37053 = n13796 | n27462 ;
  assign n37054 = n37053 ^ n8574 ^ 1'b0 ;
  assign n37055 = n4315 & n31926 ;
  assign n37059 = n10418 ^ n4539 ^ 1'b0 ;
  assign n37060 = n16377 | n37059 ;
  assign n37061 = n37060 ^ n2011 ^ 1'b0 ;
  assign n37056 = n2906 & n6781 ;
  assign n37057 = n11465 & n37056 ;
  assign n37058 = n20153 | n37057 ;
  assign n37062 = n37061 ^ n37058 ^ 1'b0 ;
  assign n37063 = n3055 | n18193 ;
  assign n37064 = n15719 ^ n1606 ^ 1'b0 ;
  assign n37065 = n10164 & ~n13290 ;
  assign n37066 = n37065 ^ n4690 ^ 1'b0 ;
  assign n37067 = n10000 | n20617 ;
  assign n37068 = ( n11815 & n16514 ) | ( n11815 & n22342 ) | ( n16514 & n22342 ) ;
  assign n37069 = ~n36494 & n37068 ;
  assign n37070 = ~n10697 & n37069 ;
  assign n37071 = n24996 & ~n32467 ;
  assign n37072 = n2718 & ~n37071 ;
  assign n37073 = ( ~n5569 & n7644 ) | ( ~n5569 & n17116 ) | ( n7644 & n17116 ) ;
  assign n37074 = n14377 & n37073 ;
  assign n37075 = n11400 & n18061 ;
  assign n37076 = n5891 ^ n460 ^ 1'b0 ;
  assign n37077 = n23443 | n37076 ;
  assign n37078 = n11205 & ~n37077 ;
  assign n37079 = x226 & n37078 ;
  assign n37080 = n415 & n2848 ;
  assign n37081 = n31773 & ~n37080 ;
  assign n37082 = n30950 ^ n4592 ^ 1'b0 ;
  assign n37083 = n29311 & ~n30783 ;
  assign n37084 = n14646 & ~n15605 ;
  assign n37085 = n37084 ^ n4584 ^ 1'b0 ;
  assign n37086 = n1920 | n3884 ;
  assign n37087 = n37086 ^ n1588 ^ 1'b0 ;
  assign n37088 = ( n2510 & n37085 ) | ( n2510 & ~n37087 ) | ( n37085 & ~n37087 ) ;
  assign n37089 = n28635 ^ n9000 ^ 1'b0 ;
  assign n37090 = x7 & n28013 ;
  assign n37091 = n37089 & n37090 ;
  assign n37092 = n26400 ^ n5874 ^ 1'b0 ;
  assign n37093 = n21558 ^ x65 ^ 1'b0 ;
  assign n37094 = n16024 | n37093 ;
  assign n37095 = n1227 | n1356 ;
  assign n37096 = n37095 ^ n9974 ^ 1'b0 ;
  assign n37097 = n13111 | n13267 ;
  assign n37098 = n27435 & ~n37097 ;
  assign n37099 = n8902 | n22731 ;
  assign n37100 = n33138 | n37099 ;
  assign n37101 = n20353 ^ n12355 ^ 1'b0 ;
  assign n37102 = n5112 & ~n5328 ;
  assign n37103 = n37102 ^ n16489 ^ n10107 ;
  assign n37104 = n34341 ^ n15481 ^ 1'b0 ;
  assign n37105 = n37103 | n37104 ;
  assign n37106 = ~n15315 & n20870 ;
  assign n37107 = n28070 ^ n11518 ^ 1'b0 ;
  assign n37108 = n5959 & n14566 ;
  assign n37109 = ~n8228 & n30790 ;
  assign n37110 = ~n2386 & n8829 ;
  assign n37111 = n29972 ^ n17546 ^ 1'b0 ;
  assign n37112 = ~n19988 & n37111 ;
  assign n37113 = n19036 | n32367 ;
  assign n37114 = n6801 | n8710 ;
  assign n37115 = ~n17980 & n19896 ;
  assign n37116 = n20186 ^ n17694 ^ 1'b0 ;
  assign n37117 = n24472 & n37116 ;
  assign n37118 = n5748 & ~n20982 ;
  assign n37119 = ~n23573 & n37118 ;
  assign n37120 = n37119 ^ n11292 ^ 1'b0 ;
  assign n37121 = n9559 & ~n32566 ;
  assign n37122 = n37121 ^ n10571 ^ 1'b0 ;
  assign n37123 = n8809 ^ n399 ^ 1'b0 ;
  assign n37124 = n2356 & n37123 ;
  assign n37125 = ( n3390 & n17736 ) | ( n3390 & ~n37124 ) | ( n17736 & ~n37124 ) ;
  assign n37126 = n15243 & n37125 ;
  assign n37127 = n7792 | n17499 ;
  assign n37131 = n3128 & ~n6854 ;
  assign n37132 = ~n3128 & n37131 ;
  assign n37128 = n2975 & n3140 ;
  assign n37129 = ~n3140 & n37128 ;
  assign n37130 = n6523 | n37129 ;
  assign n37133 = n37132 ^ n37130 ^ 1'b0 ;
  assign n37134 = n37133 ^ n8298 ^ 1'b0 ;
  assign n37135 = x95 & ~n37134 ;
  assign n37136 = ~n6315 & n37135 ;
  assign n37137 = ~n15261 & n37136 ;
  assign n37138 = ~n5890 & n11419 ;
  assign n37139 = n32640 & n37138 ;
  assign n37140 = n4615 | n36483 ;
  assign n37141 = n16001 & n24713 ;
  assign n37142 = n19699 & n37141 ;
  assign n37143 = ~n1298 & n5494 ;
  assign n37144 = n6003 & n37143 ;
  assign n37145 = ~n1009 & n37144 ;
  assign n37146 = n36830 ^ n16829 ^ 1'b0 ;
  assign n37147 = n18557 ^ n10114 ^ 1'b0 ;
  assign n37148 = n36319 ^ n6017 ^ 1'b0 ;
  assign n37149 = ~n2394 & n3956 ;
  assign n37150 = n15515 ^ n6093 ^ 1'b0 ;
  assign n37151 = ~n22402 & n23364 ;
  assign n37152 = n5509 | n10855 ;
  assign n37153 = n37152 ^ n16186 ^ 1'b0 ;
  assign n37154 = n2772 & ~n37153 ;
  assign n37155 = ~n13420 & n22570 ;
  assign n37156 = n1152 | n18263 ;
  assign n37157 = n31869 ^ n24253 ^ 1'b0 ;
  assign n37158 = ~n29099 & n33232 ;
  assign n37159 = n37158 ^ n10094 ^ 1'b0 ;
  assign n37160 = n11914 ^ n10844 ^ 1'b0 ;
  assign n37161 = n23519 ^ n15250 ^ 1'b0 ;
  assign n37162 = n13184 & n37161 ;
  assign n37163 = x243 & n26418 ;
  assign n37164 = n37163 ^ n17841 ^ 1'b0 ;
  assign n37165 = ( ~n7210 & n12912 ) | ( ~n7210 & n14997 ) | ( n12912 & n14997 ) ;
  assign n37166 = n6308 ^ n3419 ^ 1'b0 ;
  assign n37167 = n5177 ^ n1339 ^ 1'b0 ;
  assign n37168 = n24899 | n29914 ;
  assign n37169 = n37167 & n37168 ;
  assign n37170 = n10217 & ~n37169 ;
  assign n37171 = ~n12594 & n34644 ;
  assign n37172 = n37171 ^ n36055 ^ 1'b0 ;
  assign n37173 = n24200 ^ n2053 ^ 1'b0 ;
  assign n37174 = n20926 ^ n2790 ^ 1'b0 ;
  assign n37175 = n37174 ^ n23936 ^ n18578 ;
  assign n37176 = n10815 ^ n4412 ^ 1'b0 ;
  assign n37177 = n10735 ^ n1335 ^ 1'b0 ;
  assign n37178 = n4691 & n37177 ;
  assign n37179 = n32708 ^ n7028 ^ 1'b0 ;
  assign n37180 = n9177 & n37179 ;
  assign n37181 = n6786 & ~n24925 ;
  assign n37182 = n36805 ^ n24612 ^ n17833 ;
  assign n37183 = ~n829 & n29979 ;
  assign n37184 = n37183 ^ n6991 ^ 1'b0 ;
  assign n37185 = n639 & ~n15221 ;
  assign n37186 = n31773 ^ n14823 ^ 1'b0 ;
  assign n37187 = n33188 ^ n1610 ^ 1'b0 ;
  assign n37188 = n10836 ^ n1485 ^ 1'b0 ;
  assign n37189 = n30309 ^ n1093 ^ 1'b0 ;
  assign n37190 = ~n5015 & n37189 ;
  assign n37191 = n14440 ^ n1914 ^ n452 ;
  assign n37192 = n415 & n37191 ;
  assign n37193 = n7898 ^ n1404 ^ 1'b0 ;
  assign n37194 = ~n7578 & n37193 ;
  assign n37195 = n3328 ^ n1170 ^ 1'b0 ;
  assign n37196 = x67 & n18145 ;
  assign n37197 = n37196 ^ n9994 ^ 1'b0 ;
  assign n37198 = n7934 & n9239 ;
  assign n37199 = ~n10525 & n37198 ;
  assign n37200 = n37199 ^ n31883 ^ 1'b0 ;
  assign n37201 = n11068 & n29759 ;
  assign n37202 = ~n23162 & n37201 ;
  assign n37203 = ~n618 & n9423 ;
  assign n37204 = n10969 & n37203 ;
  assign n37205 = n34002 | n37204 ;
  assign n37206 = n6399 & n18069 ;
  assign n37207 = n11802 & n37206 ;
  assign n37208 = x228 & n7340 ;
  assign n37209 = ~n16039 & n37208 ;
  assign n37210 = n37209 ^ n27450 ^ 1'b0 ;
  assign n37211 = n5686 | n10931 ;
  assign n37212 = ~n9454 & n14060 ;
  assign n37213 = ~n37211 & n37212 ;
  assign n37214 = n15690 ^ n8702 ^ 1'b0 ;
  assign n37215 = ~n5667 & n25267 ;
  assign n37216 = n37215 ^ n25456 ^ 1'b0 ;
  assign n37217 = n29040 ^ n4569 ^ 1'b0 ;
  assign n37218 = n7350 & ~n37217 ;
  assign n37219 = n1546 & n32896 ;
  assign n37220 = n26809 | n34700 ;
  assign n37221 = n37220 ^ n1405 ^ 1'b0 ;
  assign n37222 = n11689 ^ n1856 ^ 1'b0 ;
  assign n37223 = ( n18588 & n19609 ) | ( n18588 & n37222 ) | ( n19609 & n37222 ) ;
  assign n37224 = n15692 | n17521 ;
  assign n37225 = n25620 & ~n37224 ;
  assign n37226 = n8589 & n15578 ;
  assign n37227 = n1429 & n22573 ;
  assign n37228 = n10611 & ~n27612 ;
  assign n37229 = n27756 ^ n1027 ^ 1'b0 ;
  assign n37230 = n844 & n37229 ;
  assign n37231 = ~n21512 & n21901 ;
  assign n37232 = n13413 & n23546 ;
  assign n37233 = n37232 ^ n23035 ^ 1'b0 ;
  assign n37234 = n19699 ^ n8474 ^ 1'b0 ;
  assign n37235 = n23077 ^ n17223 ^ 1'b0 ;
  assign n37237 = n11702 ^ n6014 ^ 1'b0 ;
  assign n37238 = n14982 | n37237 ;
  assign n37236 = n4989 & n26271 ;
  assign n37239 = n37238 ^ n37236 ^ 1'b0 ;
  assign n37240 = n10898 & ~n17874 ;
  assign n37241 = n37240 ^ n4518 ^ 1'b0 ;
  assign n37242 = n21886 ^ n5852 ^ n4526 ;
  assign n37243 = n3459 ^ n261 ^ 1'b0 ;
  assign n37244 = n21232 ^ n5578 ^ 1'b0 ;
  assign n37245 = ~n1920 & n6759 ;
  assign n37246 = n37245 ^ n18433 ^ 1'b0 ;
  assign n37247 = n2022 & ~n28051 ;
  assign n37248 = n8409 & n37247 ;
  assign n37249 = ( n8570 & n20967 ) | ( n8570 & n26716 ) | ( n20967 & n26716 ) ;
  assign n37250 = ~n14592 & n22096 ;
  assign n37251 = n16608 & n37250 ;
  assign n37252 = n9817 & n37251 ;
  assign n37253 = n17798 & n18890 ;
  assign n37254 = n4764 ^ n4398 ^ 1'b0 ;
  assign n37255 = n37253 & n37254 ;
  assign n37256 = n5671 ^ n2106 ^ 1'b0 ;
  assign n37257 = n13939 & ~n16656 ;
  assign n37258 = n37257 ^ n12959 ^ 1'b0 ;
  assign n37259 = ~n4936 & n37258 ;
  assign n37260 = ~n6025 & n37259 ;
  assign n37261 = ~n18882 & n37260 ;
  assign n37262 = ( ~n25068 & n37256 ) | ( ~n25068 & n37261 ) | ( n37256 & n37261 ) ;
  assign n37263 = n15995 & ~n24286 ;
  assign n37264 = n1810 & n37263 ;
  assign n37265 = n30117 & n35995 ;
  assign n37266 = n36071 ^ n2382 ^ 1'b0 ;
  assign n37267 = n35543 & n37266 ;
  assign n37268 = n25139 ^ n16908 ^ 1'b0 ;
  assign n37269 = n36163 | n37268 ;
  assign n37270 = n1361 & ~n5904 ;
  assign n37271 = n9326 | n11219 ;
  assign n37272 = n37270 | n37271 ;
  assign n37273 = n5021 & ~n30501 ;
  assign n37274 = ~n37272 & n37273 ;
  assign n37276 = n8657 ^ n5256 ^ 1'b0 ;
  assign n37277 = n8677 | n37276 ;
  assign n37275 = ~n6245 & n11148 ;
  assign n37278 = n37277 ^ n37275 ^ 1'b0 ;
  assign n37279 = n2970 & n37278 ;
  assign n37280 = n2687 | n14830 ;
  assign n37281 = n37280 ^ n6164 ^ 1'b0 ;
  assign n37283 = n4529 ^ n3263 ^ 1'b0 ;
  assign n37282 = n10090 | n18281 ;
  assign n37284 = n37283 ^ n37282 ^ 1'b0 ;
  assign n37285 = n6076 & ~n20712 ;
  assign n37286 = n13514 ^ n5642 ^ 1'b0 ;
  assign n37287 = ~n5988 & n28056 ;
  assign n37288 = n37287 ^ n7878 ^ 1'b0 ;
  assign n37289 = ~n4166 & n28880 ;
  assign n37290 = n37289 ^ n5518 ^ 1'b0 ;
  assign n37291 = n14344 & ~n37290 ;
  assign n37292 = n21173 & ~n33942 ;
  assign n37293 = n37292 ^ n8047 ^ 1'b0 ;
  assign n37294 = n10645 ^ n472 ^ 1'b0 ;
  assign n37295 = n5356 & ~n21482 ;
  assign n37296 = n18232 | n37295 ;
  assign n37297 = n28280 ^ n8750 ^ n6331 ;
  assign n37298 = ~n17811 & n37297 ;
  assign n37299 = ~n9022 & n37298 ;
  assign n37300 = ~n21796 & n37299 ;
  assign n37301 = n21031 ^ n13763 ^ 1'b0 ;
  assign n37302 = n27643 & n37301 ;
  assign n37303 = n8438 | n16355 ;
  assign n37304 = n12805 & n13613 ;
  assign n37305 = n24978 & n31158 ;
  assign n37306 = n20892 & n37305 ;
  assign n37307 = n15920 ^ n10888 ^ 1'b0 ;
  assign n37308 = n360 & n9173 ;
  assign n37309 = n23026 ^ n16000 ^ 1'b0 ;
  assign n37310 = ~n22696 & n37309 ;
  assign n37311 = n32320 & n33224 ;
  assign n37312 = n19622 & ~n23325 ;
  assign n37313 = ~n27532 & n37312 ;
  assign n37318 = n15241 | n29099 ;
  assign n37319 = n16862 | n37318 ;
  assign n37314 = n5287 & n25351 ;
  assign n37315 = n24990 ^ n1746 ^ 1'b0 ;
  assign n37316 = ~n37314 & n37315 ;
  assign n37317 = n1952 & n37316 ;
  assign n37320 = n37319 ^ n37317 ^ 1'b0 ;
  assign n37321 = n4059 & ~n17905 ;
  assign n37322 = n37320 & n37321 ;
  assign n37323 = n22256 ^ n10146 ^ n2399 ;
  assign n37324 = n26177 & ~n37323 ;
  assign n37325 = n13721 & ~n37324 ;
  assign n37326 = n37325 ^ n1395 ^ 1'b0 ;
  assign n37327 = n4810 & ~n17050 ;
  assign n37328 = n21879 | n37327 ;
  assign n37329 = n24341 & n28936 ;
  assign n37330 = n12346 & ~n13551 ;
  assign n37331 = n3727 ^ n1280 ^ 1'b0 ;
  assign n37332 = n629 & n37331 ;
  assign n37333 = n977 | n37332 ;
  assign n37334 = n22753 | n37333 ;
  assign n37335 = n37334 ^ n28762 ^ 1'b0 ;
  assign n37336 = n1757 & n19488 ;
  assign n37337 = ~n37335 & n37336 ;
  assign n37338 = n37337 ^ n9019 ^ 1'b0 ;
  assign n37339 = ~n15748 & n37338 ;
  assign n37340 = ~n798 & n37339 ;
  assign n37341 = ~n15423 & n37340 ;
  assign n37342 = n6322 | n15601 ;
  assign n37343 = n23251 ^ n11977 ^ 1'b0 ;
  assign n37344 = ~n16750 & n37343 ;
  assign n37345 = n8468 & n10147 ;
  assign n37346 = ~n2701 & n37345 ;
  assign n37347 = n37346 ^ n33034 ^ n18314 ;
  assign n37348 = ~n8120 & n31275 ;
  assign n37349 = n3589 & ~n37348 ;
  assign n37350 = n18874 ^ n1773 ^ 1'b0 ;
  assign n37351 = ~n17393 & n37350 ;
  assign n37352 = n37351 ^ n24496 ^ 1'b0 ;
  assign n37353 = n1423 & n6165 ;
  assign n37354 = n4173 & n37353 ;
  assign n37355 = n11964 ^ n4321 ^ 1'b0 ;
  assign n37356 = ~n1646 & n37355 ;
  assign n37357 = n4301 | n8025 ;
  assign n37358 = n14078 & ~n37357 ;
  assign n37359 = n5091 & ~n11978 ;
  assign n37360 = n24234 ^ n14472 ^ n1179 ;
  assign n37361 = n35330 ^ n29210 ^ 1'b0 ;
  assign n37362 = n2757 | n34009 ;
  assign n37363 = n13542 | n20103 ;
  assign n37364 = n37363 ^ n29155 ^ 1'b0 ;
  assign n37365 = n16967 ^ n13982 ^ 1'b0 ;
  assign n37366 = n37364 | n37365 ;
  assign n37367 = n29708 ^ n27575 ^ n20948 ;
  assign n37368 = n10792 ^ n2143 ^ 1'b0 ;
  assign n37369 = n10292 & ~n37368 ;
  assign n37370 = n37369 ^ n31164 ^ 1'b0 ;
  assign n37371 = n12877 & ~n27994 ;
  assign n37372 = x44 & n1242 ;
  assign n37373 = n21767 & n37372 ;
  assign n37374 = n8406 | n8830 ;
  assign n37375 = n6878 & ~n37374 ;
  assign n37376 = ( n34655 & ~n37373 ) | ( n34655 & n37375 ) | ( ~n37373 & n37375 ) ;
  assign n37377 = n12346 & n14947 ;
  assign n37378 = ~n5390 & n37377 ;
  assign n37379 = n19209 ^ n3750 ^ 1'b0 ;
  assign n37380 = n22791 & ~n37379 ;
  assign n37381 = n37178 ^ n9831 ^ 1'b0 ;
  assign n37382 = n18213 & n37381 ;
  assign n37383 = ~n9374 & n22342 ;
  assign n37384 = n5442 & n37383 ;
  assign n37385 = n8935 & ~n28562 ;
  assign n37386 = n7636 ^ n4656 ^ 1'b0 ;
  assign n37387 = n18939 | n37386 ;
  assign n37388 = n1321 & ~n7533 ;
  assign n37389 = n12414 & ~n18152 ;
  assign n37390 = n25753 & n37389 ;
  assign n37391 = ( n37387 & n37388 ) | ( n37387 & n37390 ) | ( n37388 & n37390 ) ;
  assign n37392 = ~n14022 & n23281 ;
  assign n37393 = n1457 & n8286 ;
  assign n37394 = n2883 | n4957 ;
  assign n37395 = n37394 ^ n17712 ^ 1'b0 ;
  assign n37396 = n7337 & n19959 ;
  assign n37397 = ~n28528 & n35340 ;
  assign n37398 = n4104 & ~n29776 ;
  assign n37399 = n37398 ^ n458 ^ 1'b0 ;
  assign n37400 = n28919 ^ n25618 ^ 1'b0 ;
  assign n37401 = n37399 | n37400 ;
  assign n37402 = ( n11001 & n37397 ) | ( n11001 & n37401 ) | ( n37397 & n37401 ) ;
  assign n37403 = ~n7860 & n7894 ;
  assign n37404 = ~n12781 & n37403 ;
  assign n37405 = n22229 ^ n4238 ^ 1'b0 ;
  assign n37406 = n14436 & ~n37405 ;
  assign n37407 = ~n28445 & n37406 ;
  assign n37408 = n23932 & n37407 ;
  assign n37409 = n37408 ^ n15908 ^ 1'b0 ;
  assign n37410 = n9160 & n24852 ;
  assign n37411 = n24044 & n37410 ;
  assign n37412 = n3970 | n20583 ;
  assign n37413 = n37412 ^ n19083 ^ 1'b0 ;
  assign n37414 = ~n37411 & n37413 ;
  assign n37415 = n18672 ^ n17594 ^ n5583 ;
  assign n37416 = n32899 ^ n31742 ^ 1'b0 ;
  assign n37417 = ~n4300 & n19218 ;
  assign n37418 = n37417 ^ n34716 ^ 1'b0 ;
  assign n37419 = n7928 & n37418 ;
  assign n37420 = n19265 & n37419 ;
  assign n37421 = n1793 & ~n9955 ;
  assign n37422 = n19479 & n37421 ;
  assign n37423 = ~n14093 & n37422 ;
  assign n37424 = n37423 ^ n18310 ^ 1'b0 ;
  assign n37425 = ~n29813 & n37424 ;
  assign n37426 = n37425 ^ n23131 ^ 1'b0 ;
  assign n37427 = n37426 ^ n35898 ^ 1'b0 ;
  assign n37428 = n6370 & ~n10024 ;
  assign n37429 = n37427 | n37428 ;
  assign n37430 = n32593 ^ n27283 ^ 1'b0 ;
  assign n37431 = n9831 & n21411 ;
  assign n37432 = ~n37430 & n37431 ;
  assign n37433 = n1205 & ~n28478 ;
  assign n37434 = n2310 & n37433 ;
  assign n37435 = ~n33633 & n37434 ;
  assign n37436 = ( n1996 & n7971 ) | ( n1996 & n19229 ) | ( n7971 & n19229 ) ;
  assign n37437 = ( n3017 & ~n37435 ) | ( n3017 & n37436 ) | ( ~n37435 & n37436 ) ;
  assign n37438 = n10553 ^ n7798 ^ 1'b0 ;
  assign n37439 = n26003 ^ n8853 ^ n2274 ;
  assign n37440 = n4478 & ~n18476 ;
  assign n37441 = n37440 ^ n3874 ^ 1'b0 ;
  assign n37442 = n5833 & ~n9283 ;
  assign n37443 = n36105 ^ n18895 ^ n3134 ;
  assign n37444 = n10808 ^ n7051 ^ 1'b0 ;
  assign n37445 = n2350 | n37444 ;
  assign n37446 = n37445 ^ n7601 ^ 1'b0 ;
  assign n37447 = ~n29705 & n37446 ;
  assign n37448 = n5475 | n20017 ;
  assign n37449 = n3001 & ~n32218 ;
  assign n37450 = n11683 ^ n1727 ^ 1'b0 ;
  assign n37451 = n17219 ^ n4172 ^ 1'b0 ;
  assign n37452 = n37451 ^ n19848 ^ 1'b0 ;
  assign n37453 = n6662 & ~n36811 ;
  assign n37454 = ~n2342 & n37453 ;
  assign n37455 = ~n9553 & n29545 ;
  assign n37456 = n28997 & n37455 ;
  assign n37457 = n37456 ^ n15444 ^ 1'b0 ;
  assign n37458 = n5203 & n13631 ;
  assign n37459 = n37458 ^ n21867 ^ 1'b0 ;
  assign n37460 = n4349 & ~n37459 ;
  assign n37461 = n17966 ^ n13825 ^ 1'b0 ;
  assign n37462 = n21152 & ~n37461 ;
  assign n37463 = n18501 & n26366 ;
  assign n37464 = n21384 ^ n12989 ^ 1'b0 ;
  assign n37465 = ~n18833 & n36066 ;
  assign n37466 = ~n9966 & n37465 ;
  assign n37467 = n20532 ^ n13438 ^ 1'b0 ;
  assign n37468 = n32921 ^ x174 ^ 1'b0 ;
  assign n37469 = n37467 & ~n37468 ;
  assign n37470 = n19220 | n28683 ;
  assign n37471 = n37470 ^ n7816 ^ 1'b0 ;
  assign n37472 = n16967 ^ n15422 ^ 1'b0 ;
  assign n37473 = ~n13627 & n37472 ;
  assign n37474 = n37473 ^ n15422 ^ 1'b0 ;
  assign n37475 = ~n2716 & n20791 ;
  assign n37476 = n13761 & ~n21842 ;
  assign n37477 = ( ~n1268 & n5692 ) | ( ~n1268 & n37476 ) | ( n5692 & n37476 ) ;
  assign n37478 = n1725 | n8748 ;
  assign n37479 = n37478 ^ n22292 ^ 1'b0 ;
  assign n37480 = n4537 | n25634 ;
  assign n37481 = n35740 & ~n37480 ;
  assign n37482 = n14980 & ~n18420 ;
  assign n37483 = ( n16177 & n28118 ) | ( n16177 & ~n28769 ) | ( n28118 & ~n28769 ) ;
  assign n37484 = n37483 ^ n5444 ^ 1'b0 ;
  assign n37485 = ~n1968 & n22012 ;
  assign n37486 = n18341 & n23702 ;
  assign n37487 = n6403 & n24960 ;
  assign n37488 = n37487 ^ n13965 ^ 1'b0 ;
  assign n37489 = ( ~n20480 & n29990 ) | ( ~n20480 & n37488 ) | ( n29990 & n37488 ) ;
  assign n37490 = n9954 | n13589 ;
  assign n37491 = ~n3589 & n27950 ;
  assign n37492 = n29329 ^ n12905 ^ 1'b0 ;
  assign n37493 = n16057 ^ n6258 ^ n320 ;
  assign n37494 = n22647 & n27632 ;
  assign n37495 = n2687 | n37494 ;
  assign n37496 = n16332 | n22563 ;
  assign n37497 = n5124 | n8054 ;
  assign n37498 = n37497 ^ n10758 ^ 1'b0 ;
  assign n37499 = n37498 ^ n6698 ^ 1'b0 ;
  assign n37500 = n23456 ^ n18059 ^ n5179 ;
  assign n37501 = n11068 & n37500 ;
  assign n37502 = n37499 & n37501 ;
  assign n37503 = n19907 ^ n14520 ^ 1'b0 ;
  assign n37504 = ~n5642 & n37503 ;
  assign n37505 = n6355 ^ x139 ^ 1'b0 ;
  assign n37506 = n6317 & n37505 ;
  assign n37507 = n13499 & n37506 ;
  assign n37508 = ~n1178 & n37507 ;
  assign n37509 = n1826 & n8358 ;
  assign n37510 = n37509 ^ n536 ^ 1'b0 ;
  assign n37511 = ~n20469 & n37510 ;
  assign n37512 = n37508 & n37511 ;
  assign n37513 = n13809 & n33861 ;
  assign n37514 = n2157 | n23406 ;
  assign n37515 = n31086 | n37514 ;
  assign n37516 = ~n26574 & n36288 ;
  assign n37517 = n37516 ^ n2384 ^ 1'b0 ;
  assign n37518 = n37515 & ~n37517 ;
  assign n37519 = ~n5312 & n12652 ;
  assign n37520 = n37519 ^ n12753 ^ 1'b0 ;
  assign n37521 = n12200 & ~n19476 ;
  assign n37522 = n37521 ^ n9781 ^ 1'b0 ;
  assign n37523 = n23677 ^ n19144 ^ 1'b0 ;
  assign n37524 = n1616 & ~n37523 ;
  assign n37525 = n34044 ^ n13959 ^ 1'b0 ;
  assign n37526 = n445 & n6721 ;
  assign n37527 = n37526 ^ n8089 ^ 1'b0 ;
  assign n37528 = n3221 & ~n7144 ;
  assign n37529 = n32922 & n37528 ;
  assign n37530 = n2760 | n37529 ;
  assign n37531 = n11148 ^ n6048 ^ 1'b0 ;
  assign n37532 = n6653 | n26017 ;
  assign n37533 = n6200 | n34427 ;
  assign n37534 = n37533 ^ n19833 ^ 1'b0 ;
  assign n37535 = n19313 ^ n18508 ^ 1'b0 ;
  assign n37536 = n2210 | n15882 ;
  assign n37537 = n37535 | n37536 ;
  assign n37538 = n24080 ^ n20142 ^ 1'b0 ;
  assign n37539 = n26869 & ~n37538 ;
  assign n37540 = n1515 & n14927 ;
  assign n37541 = n37540 ^ n22618 ^ 1'b0 ;
  assign n37542 = ~n8001 & n20015 ;
  assign n37543 = n6832 | n37542 ;
  assign n37544 = n7832 | n12154 ;
  assign n37545 = n32415 & ~n37544 ;
  assign n37546 = n2946 & n25210 ;
  assign n37547 = ( n3078 & n10465 ) | ( n3078 & ~n30888 ) | ( n10465 & ~n30888 ) ;
  assign n37548 = n10413 | n24493 ;
  assign n37549 = n1740 & ~n8480 ;
  assign n37550 = n2879 & n27850 ;
  assign n37551 = n33288 ^ n2508 ^ 1'b0 ;
  assign n37552 = n37550 & n37551 ;
  assign n37553 = ~n4776 & n37552 ;
  assign n37554 = n37553 ^ n26117 ^ 1'b0 ;
  assign n37555 = ~n14669 & n19974 ;
  assign n37556 = n37555 ^ n7950 ^ 1'b0 ;
  assign n37557 = n37554 | n37556 ;
  assign n37558 = n3606 & n6220 ;
  assign n37559 = n18126 & n37558 ;
  assign n37560 = x226 | n30469 ;
  assign n37561 = n37560 ^ n34651 ^ 1'b0 ;
  assign n37562 = n32442 & ~n36840 ;
  assign n37563 = n37562 ^ n3433 ^ 1'b0 ;
  assign n37564 = n18377 | n25140 ;
  assign n37565 = n979 & ~n10414 ;
  assign n37566 = n3116 ^ n2237 ^ 1'b0 ;
  assign n37567 = n26806 | n34538 ;
  assign n37568 = n8850 ^ n2632 ^ 1'b0 ;
  assign n37569 = n14300 & n37568 ;
  assign n37570 = n37569 ^ n1337 ^ 1'b0 ;
  assign n37571 = x25 & ~n12455 ;
  assign n37572 = n1544 & ~n10892 ;
  assign n37573 = ~n14779 & n37572 ;
  assign n37574 = n31126 | n37573 ;
  assign n37575 = n37574 ^ n29312 ^ 1'b0 ;
  assign n37576 = n9983 & n37575 ;
  assign n37577 = ~n937 & n29648 ;
  assign n37578 = n12470 | n35832 ;
  assign n37579 = ~n18766 & n20503 ;
  assign n37580 = ~n5372 & n20016 ;
  assign n37581 = n37580 ^ n9613 ^ 1'b0 ;
  assign n37582 = n18984 ^ n2466 ^ 1'b0 ;
  assign n37583 = n1890 | n1898 ;
  assign n37584 = n33914 | n37583 ;
  assign n37585 = n7755 & n16640 ;
  assign n37586 = n22414 & ~n23412 ;
  assign n37587 = n37586 ^ n37267 ^ 1'b0 ;
  assign n37588 = n13253 ^ n1815 ^ 1'b0 ;
  assign n37589 = n6886 & ~n8135 ;
  assign n37590 = n23506 ^ n17807 ^ 1'b0 ;
  assign n37591 = n1325 | n37590 ;
  assign n37592 = n9934 & ~n12744 ;
  assign n37593 = n22096 | n32600 ;
  assign n37594 = ~n14774 & n34532 ;
  assign n37595 = n34716 & n37594 ;
  assign n37596 = ~n6729 & n25535 ;
  assign n37597 = n37596 ^ n26898 ^ 1'b0 ;
  assign n37598 = n4069 | n8507 ;
  assign n37599 = n16206 | n37598 ;
  assign n37600 = n37599 ^ n11434 ^ 1'b0 ;
  assign n37601 = n18362 | n27585 ;
  assign n37602 = n37601 ^ n836 ^ 1'b0 ;
  assign n37603 = ~n26228 & n37602 ;
  assign n37604 = n5909 ^ n2664 ^ 1'b0 ;
  assign n37605 = n35224 & n37604 ;
  assign n37606 = ~n32978 & n37605 ;
  assign n37607 = n3171 ^ n1661 ^ 1'b0 ;
  assign n37608 = n37607 ^ n15552 ^ 1'b0 ;
  assign n37609 = n11329 & ~n19710 ;
  assign n37610 = ~n8288 & n37609 ;
  assign n37611 = n37610 ^ n20811 ^ 1'b0 ;
  assign n37612 = ~n6740 & n37611 ;
  assign n37613 = ( n1369 & n13808 ) | ( n1369 & n16150 ) | ( n13808 & n16150 ) ;
  assign n37614 = x97 & n5146 ;
  assign n37615 = n37614 ^ n11886 ^ 1'b0 ;
  assign n37616 = n5261 & ~n37615 ;
  assign n37617 = ~n10381 & n20001 ;
  assign n37618 = ~n8137 & n24978 ;
  assign n37619 = n37618 ^ n16401 ^ 1'b0 ;
  assign n37620 = n37619 ^ n4447 ^ 1'b0 ;
  assign n37621 = n12393 | n14241 ;
  assign n37622 = n915 | n37621 ;
  assign n37623 = n13439 & n19727 ;
  assign n37624 = n37623 ^ n2336 ^ 1'b0 ;
  assign n37625 = n37624 ^ n8921 ^ 1'b0 ;
  assign n37626 = n37625 ^ n5070 ^ 1'b0 ;
  assign n37627 = n8873 | n37626 ;
  assign n37628 = n12305 & ~n20229 ;
  assign n37629 = n19768 & n37068 ;
  assign n37630 = n11455 & n14022 ;
  assign n37631 = n691 & n37630 ;
  assign n37632 = n37631 ^ n18947 ^ 1'b0 ;
  assign n37633 = ~n25928 & n37632 ;
  assign n37634 = n11890 ^ n5083 ^ 1'b0 ;
  assign n37635 = n5619 & n37634 ;
  assign n37636 = n3577 & ~n18299 ;
  assign n37637 = n8536 & ~n37636 ;
  assign n37638 = n3249 & n12141 ;
  assign n37639 = n23282 & n37638 ;
  assign n37640 = n13521 ^ n10377 ^ n2042 ;
  assign n37641 = n4296 & ~n36328 ;
  assign n37642 = ~x252 & n37641 ;
  assign n37643 = n10183 ^ n8061 ^ n1256 ;
  assign n37644 = n37643 ^ n2728 ^ 1'b0 ;
  assign n37645 = n6932 & ~n24446 ;
  assign n37646 = n7179 | n15739 ;
  assign n37647 = ~n13495 & n37646 ;
  assign n37648 = n7609 | n14019 ;
  assign n37649 = n15624 & n23279 ;
  assign n37650 = n2681 & n17370 ;
  assign n37651 = n37650 ^ n7137 ^ 1'b0 ;
  assign n37652 = x226 ^ x177 ^ 1'b0 ;
  assign n37653 = n3432 | n6162 ;
  assign n37654 = n37653 ^ n5466 ^ 1'b0 ;
  assign n37655 = n13533 ^ n3945 ^ n1953 ;
  assign n37656 = n15228 | n37655 ;
  assign n37657 = n37656 ^ n5838 ^ 1'b0 ;
  assign n37658 = n11085 ^ n1188 ^ 1'b0 ;
  assign n37659 = n8957 | n37658 ;
  assign n37660 = n6229 | n37659 ;
  assign n37661 = n11262 | n37660 ;
  assign n37662 = n37661 ^ n18401 ^ 1'b0 ;
  assign n37663 = n17247 & n20787 ;
  assign n37664 = n37663 ^ n18550 ^ 1'b0 ;
  assign n37665 = n3796 ^ n385 ^ 1'b0 ;
  assign n37666 = n25304 & ~n37665 ;
  assign n37667 = x19 & x216 ;
  assign n37668 = n1243 & n37667 ;
  assign n37669 = n37668 ^ n16798 ^ 1'b0 ;
  assign n37670 = n24730 ^ n24060 ^ 1'b0 ;
  assign n37671 = ~n20370 & n37670 ;
  assign n37672 = n18893 ^ n16627 ^ 1'b0 ;
  assign n37673 = n37671 & n37672 ;
  assign n37674 = ~x142 & n692 ;
  assign n37675 = n37674 ^ n25037 ^ 1'b0 ;
  assign n37676 = n27533 ^ n5101 ^ 1'b0 ;
  assign n37677 = ~n11659 & n21799 ;
  assign n37678 = n37677 ^ n23273 ^ 1'b0 ;
  assign n37679 = n4657 & ~n28268 ;
  assign n37680 = n8500 | n15964 ;
  assign n37681 = n26022 | n37680 ;
  assign n37682 = n37679 & ~n37681 ;
  assign n37683 = n3377 & ~n18608 ;
  assign n37684 = n37683 ^ n22917 ^ 1'b0 ;
  assign n37685 = n32077 | n37684 ;
  assign n37686 = n17946 ^ n405 ^ 1'b0 ;
  assign n37687 = n37685 & n37686 ;
  assign n37688 = n16970 ^ n14358 ^ n2495 ;
  assign n37689 = n37688 ^ n14290 ^ 1'b0 ;
  assign n37690 = n37687 & ~n37689 ;
  assign n37691 = ~n825 & n13532 ;
  assign n37692 = n37691 ^ n8538 ^ 1'b0 ;
  assign n37693 = n37692 ^ n2851 ^ 1'b0 ;
  assign n37694 = n5002 & ~n18973 ;
  assign n37695 = n1546 & n37694 ;
  assign n37696 = n20286 ^ n1413 ^ 1'b0 ;
  assign n37697 = ~n37695 & n37696 ;
  assign n37698 = n12904 & n33562 ;
  assign n37699 = n4677 & ~n37698 ;
  assign n37700 = n31272 & n37699 ;
  assign n37703 = n8878 & n28121 ;
  assign n37701 = n6054 | n13382 ;
  assign n37702 = n6558 & n37701 ;
  assign n37704 = n37703 ^ n37702 ^ 1'b0 ;
  assign n37705 = n5067 & ~n9826 ;
  assign n37706 = n37705 ^ n6986 ^ 1'b0 ;
  assign n37707 = n9386 & ~n11954 ;
  assign n37708 = ~n28797 & n37707 ;
  assign n37709 = n37708 ^ n18074 ^ 1'b0 ;
  assign n37710 = n37283 ^ n14300 ^ 1'b0 ;
  assign n37711 = n17068 | n37710 ;
  assign n37712 = n25430 ^ n7241 ^ 1'b0 ;
  assign n37713 = n1450 & ~n37712 ;
  assign n37714 = n13352 & n27655 ;
  assign n37715 = n2949 & n37714 ;
  assign n37716 = n37715 ^ n18235 ^ 1'b0 ;
  assign n37717 = ~n1683 & n27710 ;
  assign n37718 = n15677 & n37717 ;
  assign n37719 = n3057 ^ n2665 ^ 1'b0 ;
  assign n37720 = n9590 & n37719 ;
  assign n37721 = n5988 & n22006 ;
  assign n37722 = x174 & ~n29267 ;
  assign n37723 = n37721 & n37722 ;
  assign n37724 = n20248 & n25694 ;
  assign n37725 = n27521 & ~n36145 ;
  assign n37726 = n10108 & n37725 ;
  assign n37727 = n26237 | n37726 ;
  assign n37728 = n37727 ^ n12242 ^ 1'b0 ;
  assign n37729 = n16624 ^ n4509 ^ 1'b0 ;
  assign n37730 = n15319 & ~n37729 ;
  assign n37731 = n21943 ^ n15323 ^ 1'b0 ;
  assign n37732 = n4811 & ~n37731 ;
  assign y0 = x2 ;
  assign y1 = x5 ;
  assign y2 = x7 ;
  assign y3 = x11 ;
  assign y4 = x13 ;
  assign y5 = x19 ;
  assign y6 = x20 ;
  assign y7 = x24 ;
  assign y8 = x27 ;
  assign y9 = x38 ;
  assign y10 = x42 ;
  assign y11 = x43 ;
  assign y12 = x52 ;
  assign y13 = x56 ;
  assign y14 = x60 ;
  assign y15 = x61 ;
  assign y16 = x62 ;
  assign y17 = x63 ;
  assign y18 = x75 ;
  assign y19 = x81 ;
  assign y20 = x82 ;
  assign y21 = x89 ;
  assign y22 = x92 ;
  assign y23 = x97 ;
  assign y24 = x101 ;
  assign y25 = x107 ;
  assign y26 = x115 ;
  assign y27 = x116 ;
  assign y28 = x124 ;
  assign y29 = x125 ;
  assign y30 = x126 ;
  assign y31 = x128 ;
  assign y32 = x131 ;
  assign y33 = x135 ;
  assign y34 = x136 ;
  assign y35 = x137 ;
  assign y36 = x143 ;
  assign y37 = x144 ;
  assign y38 = x149 ;
  assign y39 = x156 ;
  assign y40 = x167 ;
  assign y41 = x169 ;
  assign y42 = x170 ;
  assign y43 = x176 ;
  assign y44 = x179 ;
  assign y45 = x180 ;
  assign y46 = x188 ;
  assign y47 = x191 ;
  assign y48 = x192 ;
  assign y49 = x195 ;
  assign y50 = x196 ;
  assign y51 = x198 ;
  assign y52 = x202 ;
  assign y53 = x203 ;
  assign y54 = x204 ;
  assign y55 = x214 ;
  assign y56 = x216 ;
  assign y57 = x217 ;
  assign y58 = x219 ;
  assign y59 = x220 ;
  assign y60 = x222 ;
  assign y61 = x225 ;
  assign y62 = x226 ;
  assign y63 = x229 ;
  assign y64 = x231 ;
  assign y65 = x236 ;
  assign y66 = x237 ;
  assign y67 = x241 ;
  assign y68 = x243 ;
  assign y69 = x249 ;
  assign y70 = x254 ;
  assign y71 = n257 ;
  assign y72 = ~n259 ;
  assign y73 = ~n261 ;
  assign y74 = n263 ;
  assign y75 = n265 ;
  assign y76 = ~1'b0 ;
  assign y77 = n267 ;
  assign y78 = n269 ;
  assign y79 = ~n273 ;
  assign y80 = ~n275 ;
  assign y81 = ~n278 ;
  assign y82 = n281 ;
  assign y83 = ~n283 ;
  assign y84 = ~n285 ;
  assign y85 = ~n286 ;
  assign y86 = ~n290 ;
  assign y87 = n292 ;
  assign y88 = ~n294 ;
  assign y89 = n296 ;
  assign y90 = n302 ;
  assign y91 = n305 ;
  assign y92 = n307 ;
  assign y93 = ~n309 ;
  assign y94 = ~n311 ;
  assign y95 = ~n313 ;
  assign y96 = ~n315 ;
  assign y97 = ~n317 ;
  assign y98 = n318 ;
  assign y99 = ~n320 ;
  assign y100 = ~n322 ;
  assign y101 = ~1'b0 ;
  assign y102 = ~n323 ;
  assign y103 = ~n325 ;
  assign y104 = ~n327 ;
  assign y105 = ~n329 ;
  assign y106 = ~n331 ;
  assign y107 = n333 ;
  assign y108 = ~n335 ;
  assign y109 = n337 ;
  assign y110 = n343 ;
  assign y111 = ~n345 ;
  assign y112 = ~n347 ;
  assign y113 = ~n351 ;
  assign y114 = ~n357 ;
  assign y115 = ~n358 ;
  assign y116 = ~n368 ;
  assign y117 = n370 ;
  assign y118 = ~1'b0 ;
  assign y119 = ~1'b0 ;
  assign y120 = ~1'b0 ;
  assign y121 = n372 ;
  assign y122 = n373 ;
  assign y123 = ~n374 ;
  assign y124 = ~1'b0 ;
  assign y125 = ~n376 ;
  assign y126 = n378 ;
  assign y127 = ~n381 ;
  assign y128 = ~1'b0 ;
  assign y129 = ~1'b0 ;
  assign y130 = n387 ;
  assign y131 = n392 ;
  assign y132 = ~1'b0 ;
  assign y133 = ~1'b0 ;
  assign y134 = ~n397 ;
  assign y135 = ~1'b0 ;
  assign y136 = ~1'b0 ;
  assign y137 = ~1'b0 ;
  assign y138 = ~1'b0 ;
  assign y139 = n407 ;
  assign y140 = n409 ;
  assign y141 = ~n421 ;
  assign y142 = n426 ;
  assign y143 = ~n428 ;
  assign y144 = ~n432 ;
  assign y145 = ~n434 ;
  assign y146 = ~n442 ;
  assign y147 = ~1'b0 ;
  assign y148 = n444 ;
  assign y149 = n446 ;
  assign y150 = ~1'b0 ;
  assign y151 = ~1'b0 ;
  assign y152 = ~n448 ;
  assign y153 = ~n456 ;
  assign y154 = ~1'b0 ;
  assign y155 = n461 ;
  assign y156 = 1'b0 ;
  assign y157 = n465 ;
  assign y158 = n467 ;
  assign y159 = ~n468 ;
  assign y160 = ~n472 ;
  assign y161 = x253 ;
  assign y162 = ~1'b0 ;
  assign y163 = ~1'b0 ;
  assign y164 = ~n476 ;
  assign y165 = ~n478 ;
  assign y166 = ~1'b0 ;
  assign y167 = ~n481 ;
  assign y168 = n482 ;
  assign y169 = ~1'b0 ;
  assign y170 = ~1'b0 ;
  assign y171 = ~n493 ;
  assign y172 = n495 ;
  assign y173 = ~n497 ;
  assign y174 = n498 ;
  assign y175 = ~1'b0 ;
  assign y176 = ~n503 ;
  assign y177 = ~n504 ;
  assign y178 = n446 ;
  assign y179 = ~n505 ;
  assign y180 = ~1'b0 ;
  assign y181 = n522 ;
  assign y182 = ~1'b0 ;
  assign y183 = ~n526 ;
  assign y184 = ~1'b0 ;
  assign y185 = n527 ;
  assign y186 = n528 ;
  assign y187 = ~n529 ;
  assign y188 = x127 ;
  assign y189 = ~1'b0 ;
  assign y190 = ~n533 ;
  assign y191 = ~n534 ;
  assign y192 = 1'b0 ;
  assign y193 = ~1'b0 ;
  assign y194 = ~n536 ;
  assign y195 = ~x41 ;
  assign y196 = n538 ;
  assign y197 = ~1'b0 ;
  assign y198 = ~n539 ;
  assign y199 = n546 ;
  assign y200 = n549 ;
  assign y201 = ~n552 ;
  assign y202 = ~1'b0 ;
  assign y203 = n559 ;
  assign y204 = n562 ;
  assign y205 = n570 ;
  assign y206 = ~1'b0 ;
  assign y207 = ~n571 ;
  assign y208 = ~1'b0 ;
  assign y209 = n575 ;
  assign y210 = n579 ;
  assign y211 = ~1'b0 ;
  assign y212 = n583 ;
  assign y213 = n590 ;
  assign y214 = ~1'b0 ;
  assign y215 = ~1'b0 ;
  assign y216 = ~n594 ;
  assign y217 = n595 ;
  assign y218 = ~1'b0 ;
  assign y219 = ~n598 ;
  assign y220 = ~1'b0 ;
  assign y221 = ~1'b0 ;
  assign y222 = x222 ;
  assign y223 = n602 ;
  assign y224 = ~n608 ;
  assign y225 = ~n613 ;
  assign y226 = ~n616 ;
  assign y227 = ~n618 ;
  assign y228 = ~n623 ;
  assign y229 = ~n626 ;
  assign y230 = n629 ;
  assign y231 = ~n296 ;
  assign y232 = ~x22 ;
  assign y233 = ~1'b0 ;
  assign y234 = ~1'b0 ;
  assign y235 = ~n631 ;
  assign y236 = ~1'b0 ;
  assign y237 = n633 ;
  assign y238 = ~n635 ;
  assign y239 = ~1'b0 ;
  assign y240 = n639 ;
  assign y241 = ~n641 ;
  assign y242 = n642 ;
  assign y243 = n643 ;
  assign y244 = ~1'b0 ;
  assign y245 = ~1'b0 ;
  assign y246 = x182 ;
  assign y247 = n644 ;
  assign y248 = n645 ;
  assign y249 = n648 ;
  assign y250 = n655 ;
  assign y251 = n662 ;
  assign y252 = ~n669 ;
  assign y253 = ~n671 ;
  assign y254 = ~n685 ;
  assign y255 = ~1'b0 ;
  assign y256 = ~1'b0 ;
  assign y257 = ~n691 ;
  assign y258 = ~x20 ;
  assign y259 = ~n694 ;
  assign y260 = ~1'b0 ;
  assign y261 = ~n696 ;
  assign y262 = ~1'b0 ;
  assign y263 = ~1'b0 ;
  assign y264 = ~1'b0 ;
  assign y265 = ~n698 ;
  assign y266 = ~n701 ;
  assign y267 = 1'b0 ;
  assign y268 = ~n708 ;
  assign y269 = ~1'b0 ;
  assign y270 = ~n709 ;
  assign y271 = x226 ;
  assign y272 = n710 ;
  assign y273 = ~1'b0 ;
  assign y274 = ~1'b0 ;
  assign y275 = n720 ;
  assign y276 = ~1'b0 ;
  assign y277 = ~1'b0 ;
  assign y278 = n722 ;
  assign y279 = n724 ;
  assign y280 = ~1'b0 ;
  assign y281 = n725 ;
  assign y282 = ~1'b0 ;
  assign y283 = 1'b0 ;
  assign y284 = ~1'b0 ;
  assign y285 = n444 ;
  assign y286 = ~1'b0 ;
  assign y287 = x73 ;
  assign y288 = ~n726 ;
  assign y289 = n728 ;
  assign y290 = ~n729 ;
  assign y291 = n730 ;
  assign y292 = ~1'b0 ;
  assign y293 = ~n748 ;
  assign y294 = ~n749 ;
  assign y295 = n750 ;
  assign y296 = ~1'b0 ;
  assign y297 = ~n752 ;
  assign y298 = ~n753 ;
  assign y299 = ~1'b0 ;
  assign y300 = ~1'b0 ;
  assign y301 = n756 ;
  assign y302 = ~n758 ;
  assign y303 = ~1'b0 ;
  assign y304 = ~x154 ;
  assign y305 = n760 ;
  assign y306 = ~1'b0 ;
  assign y307 = ~n761 ;
  assign y308 = ~1'b0 ;
  assign y309 = n762 ;
  assign y310 = ~1'b0 ;
  assign y311 = ~1'b0 ;
  assign y312 = ~n764 ;
  assign y313 = ~1'b0 ;
  assign y314 = ~1'b0 ;
  assign y315 = ~n770 ;
  assign y316 = ~1'b0 ;
  assign y317 = ~n774 ;
  assign y318 = n778 ;
  assign y319 = ~n780 ;
  assign y320 = ~n781 ;
  assign y321 = ~n784 ;
  assign y322 = ~n766 ;
  assign y323 = ~1'b0 ;
  assign y324 = ~1'b0 ;
  assign y325 = ~n785 ;
  assign y326 = n786 ;
  assign y327 = ~1'b0 ;
  assign y328 = n787 ;
  assign y329 = ~1'b0 ;
  assign y330 = ~1'b0 ;
  assign y331 = ~n790 ;
  assign y332 = ~n796 ;
  assign y333 = ~1'b0 ;
  assign y334 = ~n798 ;
  assign y335 = n800 ;
  assign y336 = x143 ;
  assign y337 = ~1'b0 ;
  assign y338 = ~1'b0 ;
  assign y339 = n801 ;
  assign y340 = ~n803 ;
  assign y341 = 1'b0 ;
  assign y342 = x244 ;
  assign y343 = ~n808 ;
  assign y344 = ~1'b0 ;
  assign y345 = n809 ;
  assign y346 = n817 ;
  assign y347 = ~n821 ;
  assign y348 = x208 ;
  assign y349 = ~n472 ;
  assign y350 = ~n320 ;
  assign y351 = ~1'b0 ;
  assign y352 = n825 ;
  assign y353 = n827 ;
  assign y354 = ~n829 ;
  assign y355 = 1'b0 ;
  assign y356 = ~1'b0 ;
  assign y357 = ~n830 ;
  assign y358 = n833 ;
  assign y359 = n835 ;
  assign y360 = ~n842 ;
  assign y361 = ~n840 ;
  assign y362 = ~n848 ;
  assign y363 = n849 ;
  assign y364 = n853 ;
  assign y365 = n855 ;
  assign y366 = n859 ;
  assign y367 = ~1'b0 ;
  assign y368 = n860 ;
  assign y369 = ~n862 ;
  assign y370 = ~n863 ;
  assign y371 = ~n864 ;
  assign y372 = 1'b0 ;
  assign y373 = ~1'b0 ;
  assign y374 = n867 ;
  assign y375 = ~n871 ;
  assign y376 = ~n874 ;
  assign y377 = ~1'b0 ;
  assign y378 = n876 ;
  assign y379 = n880 ;
  assign y380 = ~n881 ;
  assign y381 = n883 ;
  assign y382 = n886 ;
  assign y383 = ~1'b0 ;
  assign y384 = ~1'b0 ;
  assign y385 = ~1'b0 ;
  assign y386 = n888 ;
  assign y387 = n896 ;
  assign y388 = ~n901 ;
  assign y389 = ~n904 ;
  assign y390 = ~n913 ;
  assign y391 = ~1'b0 ;
  assign y392 = n918 ;
  assign y393 = ~1'b0 ;
  assign y394 = ~n921 ;
  assign y395 = n923 ;
  assign y396 = n924 ;
  assign y397 = n927 ;
  assign y398 = ~1'b0 ;
  assign y399 = n928 ;
  assign y400 = ~n929 ;
  assign y401 = ~n934 ;
  assign y402 = n944 ;
  assign y403 = 1'b0 ;
  assign y404 = ~1'b0 ;
  assign y405 = ~1'b0 ;
  assign y406 = n946 ;
  assign y407 = ~n951 ;
  assign y408 = ~1'b0 ;
  assign y409 = ~n956 ;
  assign y410 = ~1'b0 ;
  assign y411 = x31 ;
  assign y412 = n957 ;
  assign y413 = n958 ;
  assign y414 = n966 ;
  assign y415 = n967 ;
  assign y416 = ~1'b0 ;
  assign y417 = n936 ;
  assign y418 = ~1'b0 ;
  assign y419 = x115 ;
  assign y420 = n969 ;
  assign y421 = ~n971 ;
  assign y422 = n975 ;
  assign y423 = n979 ;
  assign y424 = ~1'b0 ;
  assign y425 = ~n589 ;
  assign y426 = ~n981 ;
  assign y427 = ~n983 ;
  assign y428 = ~n988 ;
  assign y429 = ~1'b0 ;
  assign y430 = ~n989 ;
  assign y431 = n998 ;
  assign y432 = n994 ;
  assign y433 = ~n1007 ;
  assign y434 = ~n1009 ;
  assign y435 = ~n1016 ;
  assign y436 = n1025 ;
  assign y437 = ~1'b0 ;
  assign y438 = ~n1031 ;
  assign y439 = ~1'b0 ;
  assign y440 = n1033 ;
  assign y441 = n1035 ;
  assign y442 = n1037 ;
  assign y443 = n1038 ;
  assign y444 = n1047 ;
  assign y445 = n1050 ;
  assign y446 = ~1'b0 ;
  assign y447 = n1054 ;
  assign y448 = ~1'b0 ;
  assign y449 = n1058 ;
  assign y450 = ~n1061 ;
  assign y451 = ~1'b0 ;
  assign y452 = n1065 ;
  assign y453 = ~n1066 ;
  assign y454 = n1073 ;
  assign y455 = ~n1079 ;
  assign y456 = n1080 ;
  assign y457 = ~n1082 ;
  assign y458 = n1087 ;
  assign y459 = n1089 ;
  assign y460 = ~1'b0 ;
  assign y461 = ~1'b0 ;
  assign y462 = n1096 ;
  assign y463 = ~1'b0 ;
  assign y464 = n1098 ;
  assign y465 = ~1'b0 ;
  assign y466 = ~n1104 ;
  assign y467 = n1105 ;
  assign y468 = ~1'b0 ;
  assign y469 = ~1'b0 ;
  assign y470 = ~1'b0 ;
  assign y471 = ~1'b0 ;
  assign y472 = ~1'b0 ;
  assign y473 = n1106 ;
  assign y474 = ~1'b0 ;
  assign y475 = n1112 ;
  assign y476 = n1114 ;
  assign y477 = ~1'b0 ;
  assign y478 = ~n1118 ;
  assign y479 = n1120 ;
  assign y480 = ~n1126 ;
  assign y481 = ~1'b0 ;
  assign y482 = ~1'b0 ;
  assign y483 = ~n1130 ;
  assign y484 = ~1'b0 ;
  assign y485 = ~1'b0 ;
  assign y486 = n1131 ;
  assign y487 = ~n1135 ;
  assign y488 = n1137 ;
  assign y489 = ~n1141 ;
  assign y490 = n1148 ;
  assign y491 = n1150 ;
  assign y492 = ~1'b0 ;
  assign y493 = ~1'b0 ;
  assign y494 = n1164 ;
  assign y495 = ~1'b0 ;
  assign y496 = n500 ;
  assign y497 = ~1'b0 ;
  assign y498 = ~n1165 ;
  assign y499 = n1167 ;
  assign y500 = ~1'b0 ;
  assign y501 = ~n1169 ;
  assign y502 = ~n1172 ;
  assign y503 = ~x207 ;
  assign y504 = ~1'b0 ;
  assign y505 = ~1'b0 ;
  assign y506 = n1173 ;
  assign y507 = ~n1028 ;
  assign y508 = ~n1182 ;
  assign y509 = ~1'b0 ;
  assign y510 = ~n442 ;
  assign y511 = n1191 ;
  assign y512 = ~1'b0 ;
  assign y513 = n1194 ;
  assign y514 = n1195 ;
  assign y515 = ~1'b0 ;
  assign y516 = ~n1198 ;
  assign y517 = ~1'b0 ;
  assign y518 = n1199 ;
  assign y519 = ~n1202 ;
  assign y520 = n1217 ;
  assign y521 = ~1'b0 ;
  assign y522 = ~1'b0 ;
  assign y523 = ~n1227 ;
  assign y524 = ~n1230 ;
  assign y525 = ~n1234 ;
  assign y526 = ~n1236 ;
  assign y527 = 1'b0 ;
  assign y528 = ~n1239 ;
  assign y529 = ~n1240 ;
  assign y530 = n1247 ;
  assign y531 = ~n1248 ;
  assign y532 = n1249 ;
  assign y533 = n1256 ;
  assign y534 = n1261 ;
  assign y535 = ~1'b0 ;
  assign y536 = n1262 ;
  assign y537 = 1'b0 ;
  assign y538 = n1263 ;
  assign y539 = n1267 ;
  assign y540 = ~n1269 ;
  assign y541 = ~1'b0 ;
  assign y542 = ~n774 ;
  assign y543 = n1277 ;
  assign y544 = ~1'b0 ;
  assign y545 = n1278 ;
  assign y546 = ~n1280 ;
  assign y547 = ~n1285 ;
  assign y548 = n1286 ;
  assign y549 = ~n1290 ;
  assign y550 = x76 ;
  assign y551 = ~n1291 ;
  assign y552 = n1297 ;
  assign y553 = ~n1298 ;
  assign y554 = n1301 ;
  assign y555 = ~n557 ;
  assign y556 = n1302 ;
  assign y557 = ~n1304 ;
  assign y558 = ~1'b0 ;
  assign y559 = ~n1305 ;
  assign y560 = ~1'b0 ;
  assign y561 = ~1'b0 ;
  assign y562 = n1311 ;
  assign y563 = ~n1312 ;
  assign y564 = n1318 ;
  assign y565 = ~1'b0 ;
  assign y566 = ~1'b0 ;
  assign y567 = ~n1327 ;
  assign y568 = n1328 ;
  assign y569 = ~1'b0 ;
  assign y570 = ~1'b0 ;
  assign y571 = ~n1330 ;
  assign y572 = ~n1334 ;
  assign y573 = ~n1335 ;
  assign y574 = ~1'b0 ;
  assign y575 = ~1'b0 ;
  assign y576 = n1336 ;
  assign y577 = ~1'b0 ;
  assign y578 = ~n1337 ;
  assign y579 = n1344 ;
  assign y580 = n1345 ;
  assign y581 = ~n1350 ;
  assign y582 = ~1'b0 ;
  assign y583 = n1351 ;
  assign y584 = ~n1352 ;
  assign y585 = n1269 ;
  assign y586 = ~1'b0 ;
  assign y587 = n1353 ;
  assign y588 = ~n1354 ;
  assign y589 = n1358 ;
  assign y590 = ~1'b0 ;
  assign y591 = n1361 ;
  assign y592 = ~1'b0 ;
  assign y593 = ~n1363 ;
  assign y594 = ~n1372 ;
  assign y595 = ~1'b0 ;
  assign y596 = n1374 ;
  assign y597 = n1378 ;
  assign y598 = ~1'b0 ;
  assign y599 = n1379 ;
  assign y600 = n1380 ;
  assign y601 = ~n1382 ;
  assign y602 = n1389 ;
  assign y603 = ~n1390 ;
  assign y604 = ~1'b0 ;
  assign y605 = ~n1395 ;
  assign y606 = ~1'b0 ;
  assign y607 = ~1'b0 ;
  assign y608 = n1397 ;
  assign y609 = n1400 ;
  assign y610 = ~n1339 ;
  assign y611 = ~n1407 ;
  assign y612 = ~1'b0 ;
  assign y613 = ~n1410 ;
  assign y614 = ~n1414 ;
  assign y615 = n1415 ;
  assign y616 = ~n1421 ;
  assign y617 = ~n1427 ;
  assign y618 = ~1'b0 ;
  assign y619 = n1431 ;
  assign y620 = ~1'b0 ;
  assign y621 = ~1'b0 ;
  assign y622 = n1436 ;
  assign y623 = n1446 ;
  assign y624 = n286 ;
  assign y625 = ~n1449 ;
  assign y626 = ~n1450 ;
  assign y627 = ~1'b0 ;
  assign y628 = ~n1451 ;
  assign y629 = ~n1453 ;
  assign y630 = ~n1455 ;
  assign y631 = ~1'b0 ;
  assign y632 = x155 ;
  assign y633 = n1461 ;
  assign y634 = n1464 ;
  assign y635 = ~1'b0 ;
  assign y636 = ~1'b0 ;
  assign y637 = ~1'b0 ;
  assign y638 = n1468 ;
  assign y639 = ~n1472 ;
  assign y640 = ~n1473 ;
  assign y641 = n1475 ;
  assign y642 = n1477 ;
  assign y643 = n1479 ;
  assign y644 = ~n1480 ;
  assign y645 = ~1'b0 ;
  assign y646 = n1487 ;
  assign y647 = ~1'b0 ;
  assign y648 = ~n1488 ;
  assign y649 = n1489 ;
  assign y650 = ~n1490 ;
  assign y651 = n1492 ;
  assign y652 = ~1'b0 ;
  assign y653 = ~1'b0 ;
  assign y654 = ~1'b0 ;
  assign y655 = ~1'b0 ;
  assign y656 = n1495 ;
  assign y657 = ~1'b0 ;
  assign y658 = n1496 ;
  assign y659 = ~n1503 ;
  assign y660 = ~1'b0 ;
  assign y661 = n1508 ;
  assign y662 = n1511 ;
  assign y663 = n1514 ;
  assign y664 = n1515 ;
  assign y665 = ~n1518 ;
  assign y666 = ~n1522 ;
  assign y667 = ~n1524 ;
  assign y668 = n1525 ;
  assign y669 = ~x93 ;
  assign y670 = ~1'b0 ;
  assign y671 = ~1'b0 ;
  assign y672 = ~n944 ;
  assign y673 = ~n1527 ;
  assign y674 = 1'b0 ;
  assign y675 = ~1'b0 ;
  assign y676 = ~1'b0 ;
  assign y677 = ~n1529 ;
  assign y678 = n345 ;
  assign y679 = ~n1533 ;
  assign y680 = ~n1535 ;
  assign y681 = ~n1538 ;
  assign y682 = ~1'b0 ;
  assign y683 = n1540 ;
  assign y684 = n1549 ;
  assign y685 = ~1'b0 ;
  assign y686 = ~n1553 ;
  assign y687 = n1556 ;
  assign y688 = ~n1557 ;
  assign y689 = ~n1559 ;
  assign y690 = ~1'b0 ;
  assign y691 = ~1'b0 ;
  assign y692 = ~n1560 ;
  assign y693 = ~1'b0 ;
  assign y694 = n1564 ;
  assign y695 = ~n1569 ;
  assign y696 = n1576 ;
  assign y697 = ~1'b0 ;
  assign y698 = n1579 ;
  assign y699 = ~n1580 ;
  assign y700 = n1587 ;
  assign y701 = ~n1588 ;
  assign y702 = n1589 ;
  assign y703 = ~n1591 ;
  assign y704 = ~1'b0 ;
  assign y705 = n1593 ;
  assign y706 = n1594 ;
  assign y707 = ~n1605 ;
  assign y708 = ~1'b0 ;
  assign y709 = ~n1610 ;
  assign y710 = ~n1611 ;
  assign y711 = ~n1613 ;
  assign y712 = ~1'b0 ;
  assign y713 = ~1'b0 ;
  assign y714 = ~1'b0 ;
  assign y715 = ~1'b0 ;
  assign y716 = n1614 ;
  assign y717 = ~1'b0 ;
  assign y718 = n1618 ;
  assign y719 = ~n1619 ;
  assign y720 = ~n1620 ;
  assign y721 = ~1'b0 ;
  assign y722 = n1621 ;
  assign y723 = ~n1626 ;
  assign y724 = ~n1630 ;
  assign y725 = n1635 ;
  assign y726 = n1637 ;
  assign y727 = n1639 ;
  assign y728 = ~1'b0 ;
  assign y729 = ~1'b0 ;
  assign y730 = n1648 ;
  assign y731 = ~n1650 ;
  assign y732 = ~1'b0 ;
  assign y733 = ~n1651 ;
  assign y734 = ~1'b0 ;
  assign y735 = n1654 ;
  assign y736 = n1657 ;
  assign y737 = n1658 ;
  assign y738 = x88 ;
  assign y739 = ~1'b0 ;
  assign y740 = n1663 ;
  assign y741 = ~1'b0 ;
  assign y742 = n1668 ;
  assign y743 = ~1'b0 ;
  assign y744 = 1'b0 ;
  assign y745 = n1671 ;
  assign y746 = ~n1672 ;
  assign y747 = ~n1673 ;
  assign y748 = ~1'b0 ;
  assign y749 = ~1'b0 ;
  assign y750 = n1675 ;
  assign y751 = ~1'b0 ;
  assign y752 = n1512 ;
  assign y753 = n1678 ;
  assign y754 = ~n1680 ;
  assign y755 = ~1'b0 ;
  assign y756 = ~1'b0 ;
  assign y757 = ~1'b0 ;
  assign y758 = n1685 ;
  assign y759 = ~1'b0 ;
  assign y760 = ~n1686 ;
  assign y761 = n1688 ;
  assign y762 = ~n1689 ;
  assign y763 = ~n1690 ;
  assign y764 = ~n1693 ;
  assign y765 = ~n1696 ;
  assign y766 = ~n1698 ;
  assign y767 = ~1'b0 ;
  assign y768 = ~n1703 ;
  assign y769 = n1707 ;
  assign y770 = n1714 ;
  assign y771 = ~1'b0 ;
  assign y772 = n1715 ;
  assign y773 = ~n1718 ;
  assign y774 = n1720 ;
  assign y775 = ~1'b0 ;
  assign y776 = n1724 ;
  assign y777 = ~1'b0 ;
  assign y778 = ~n1725 ;
  assign y779 = n1727 ;
  assign y780 = ~1'b0 ;
  assign y781 = ~1'b0 ;
  assign y782 = ~1'b0 ;
  assign y783 = ~n1729 ;
  assign y784 = n1731 ;
  assign y785 = n1732 ;
  assign y786 = n1735 ;
  assign y787 = ~1'b0 ;
  assign y788 = n1736 ;
  assign y789 = ~1'b0 ;
  assign y790 = ~n1738 ;
  assign y791 = ~1'b0 ;
  assign y792 = ~n1741 ;
  assign y793 = n1743 ;
  assign y794 = ~1'b0 ;
  assign y795 = ~1'b0 ;
  assign y796 = n1744 ;
  assign y797 = ~n1745 ;
  assign y798 = ~1'b0 ;
  assign y799 = ~1'b0 ;
  assign y800 = ~n1746 ;
  assign y801 = ~n1747 ;
  assign y802 = 1'b0 ;
  assign y803 = ~1'b0 ;
  assign y804 = n1749 ;
  assign y805 = ~1'b0 ;
  assign y806 = ~1'b0 ;
  assign y807 = ~1'b0 ;
  assign y808 = ~1'b0 ;
  assign y809 = ~1'b0 ;
  assign y810 = n1758 ;
  assign y811 = ~1'b0 ;
  assign y812 = ~1'b0 ;
  assign y813 = n1762 ;
  assign y814 = n1764 ;
  assign y815 = n1766 ;
  assign y816 = n1770 ;
  assign y817 = ~n1772 ;
  assign y818 = n1779 ;
  assign y819 = ~n1782 ;
  assign y820 = ~n1783 ;
  assign y821 = n1788 ;
  assign y822 = ~1'b0 ;
  assign y823 = n1791 ;
  assign y824 = ~1'b0 ;
  assign y825 = n1792 ;
  assign y826 = ~1'b0 ;
  assign y827 = n1793 ;
  assign y828 = n1797 ;
  assign y829 = ~n1801 ;
  assign y830 = n1803 ;
  assign y831 = 1'b0 ;
  assign y832 = ~n1805 ;
  assign y833 = ~1'b0 ;
  assign y834 = ~1'b0 ;
  assign y835 = n1808 ;
  assign y836 = ~1'b0 ;
  assign y837 = n1809 ;
  assign y838 = ~n894 ;
  assign y839 = n1810 ;
  assign y840 = ~1'b0 ;
  assign y841 = ~1'b0 ;
  assign y842 = ~n1812 ;
  assign y843 = n1815 ;
  assign y844 = n1818 ;
  assign y845 = ~n1820 ;
  assign y846 = ~1'b0 ;
  assign y847 = n1825 ;
  assign y848 = ~1'b0 ;
  assign y849 = ~n1828 ;
  assign y850 = n1832 ;
  assign y851 = ~1'b0 ;
  assign y852 = ~n1834 ;
  assign y853 = ~1'b0 ;
  assign y854 = ~n1835 ;
  assign y855 = ~n1836 ;
  assign y856 = ~n1837 ;
  assign y857 = ~n1840 ;
  assign y858 = n1841 ;
  assign y859 = ~1'b0 ;
  assign y860 = n1846 ;
  assign y861 = ~1'b0 ;
  assign y862 = ~1'b0 ;
  assign y863 = n1849 ;
  assign y864 = ~1'b0 ;
  assign y865 = n1850 ;
  assign y866 = n1854 ;
  assign y867 = n1856 ;
  assign y868 = ~1'b0 ;
  assign y869 = ~1'b0 ;
  assign y870 = ~n1859 ;
  assign y871 = n1861 ;
  assign y872 = ~1'b0 ;
  assign y873 = ~n1863 ;
  assign y874 = n1866 ;
  assign y875 = ~n1867 ;
  assign y876 = ~n1872 ;
  assign y877 = n1873 ;
  assign y878 = ~n1879 ;
  assign y879 = n1885 ;
  assign y880 = ~n1886 ;
  assign y881 = ~x50 ;
  assign y882 = n1892 ;
  assign y883 = ~1'b0 ;
  assign y884 = ~1'b0 ;
  assign y885 = n271 ;
  assign y886 = ~n1893 ;
  assign y887 = n1894 ;
  assign y888 = ~n1897 ;
  assign y889 = ~n1898 ;
  assign y890 = n1900 ;
  assign y891 = ~n325 ;
  assign y892 = x3 ;
  assign y893 = ~1'b0 ;
  assign y894 = ~1'b0 ;
  assign y895 = n1901 ;
  assign y896 = n1909 ;
  assign y897 = n1914 ;
  assign y898 = ~n1683 ;
  assign y899 = ~1'b0 ;
  assign y900 = ~1'b0 ;
  assign y901 = n1916 ;
  assign y902 = n1922 ;
  assign y903 = n1929 ;
  assign y904 = ~1'b0 ;
  assign y905 = n859 ;
  assign y906 = ~n1930 ;
  assign y907 = n1931 ;
  assign y908 = n1932 ;
  assign y909 = ~n1936 ;
  assign y910 = ~1'b0 ;
  assign y911 = 1'b0 ;
  assign y912 = n1883 ;
  assign y913 = ~1'b0 ;
  assign y914 = ~1'b0 ;
  assign y915 = n1937 ;
  assign y916 = ~1'b0 ;
  assign y917 = n1938 ;
  assign y918 = n1941 ;
  assign y919 = n1944 ;
  assign y920 = n1945 ;
  assign y921 = n1947 ;
  assign y922 = ~1'b0 ;
  assign y923 = ~n1949 ;
  assign y924 = n1950 ;
  assign y925 = ~1'b0 ;
  assign y926 = ~1'b0 ;
  assign y927 = ~1'b0 ;
  assign y928 = ~n956 ;
  assign y929 = ~n1951 ;
  assign y930 = ~1'b0 ;
  assign y931 = ~n1952 ;
  assign y932 = n1959 ;
  assign y933 = ~1'b0 ;
  assign y934 = ~1'b0 ;
  assign y935 = ~n1965 ;
  assign y936 = ~1'b0 ;
  assign y937 = ~1'b0 ;
  assign y938 = n1967 ;
  assign y939 = n1969 ;
  assign y940 = ~1'b0 ;
  assign y941 = n1973 ;
  assign y942 = ~1'b0 ;
  assign y943 = n1979 ;
  assign y944 = n1981 ;
  assign y945 = n1793 ;
  assign y946 = ~n1983 ;
  assign y947 = ~n1988 ;
  assign y948 = n1990 ;
  assign y949 = ~1'b0 ;
  assign y950 = ~n1999 ;
  assign y951 = n2001 ;
  assign y952 = ~1'b0 ;
  assign y953 = ~1'b0 ;
  assign y954 = ~n2003 ;
  assign y955 = ~n2004 ;
  assign y956 = ~n2006 ;
  assign y957 = n2008 ;
  assign y958 = n2012 ;
  assign y959 = ~n2019 ;
  assign y960 = ~n2021 ;
  assign y961 = n2035 ;
  assign y962 = ~n2038 ;
  assign y963 = n2044 ;
  assign y964 = n2046 ;
  assign y965 = ~n2047 ;
  assign y966 = ~n2053 ;
  assign y967 = ~n2054 ;
  assign y968 = ~n2055 ;
  assign y969 = n2057 ;
  assign y970 = n2058 ;
  assign y971 = n2060 ;
  assign y972 = ~1'b0 ;
  assign y973 = ~n2061 ;
  assign y974 = n2063 ;
  assign y975 = ~n1181 ;
  assign y976 = ~1'b0 ;
  assign y977 = 1'b0 ;
  assign y978 = ~n2066 ;
  assign y979 = ~1'b0 ;
  assign y980 = ~1'b0 ;
  assign y981 = n2068 ;
  assign y982 = 1'b0 ;
  assign y983 = ~n2070 ;
  assign y984 = ~1'b0 ;
  assign y985 = n2071 ;
  assign y986 = n2073 ;
  assign y987 = ~n2076 ;
  assign y988 = n2078 ;
  assign y989 = ~1'b0 ;
  assign y990 = ~1'b0 ;
  assign y991 = ~1'b0 ;
  assign y992 = ~1'b0 ;
  assign y993 = ~n1239 ;
  assign y994 = n2080 ;
  assign y995 = n2082 ;
  assign y996 = n2083 ;
  assign y997 = ~1'b0 ;
  assign y998 = ~n2087 ;
  assign y999 = ~n2093 ;
  assign y1000 = ~n2098 ;
  assign y1001 = ~1'b0 ;
  assign y1002 = n2109 ;
  assign y1003 = ~1'b0 ;
  assign y1004 = ~n2113 ;
  assign y1005 = ~1'b0 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = ~1'b0 ;
  assign y1008 = ~n2114 ;
  assign y1009 = n2115 ;
  assign y1010 = ~n2116 ;
  assign y1011 = ~n2117 ;
  assign y1012 = ~n2125 ;
  assign y1013 = ~x147 ;
  assign y1014 = n2127 ;
  assign y1015 = n2136 ;
  assign y1016 = ~n2140 ;
  assign y1017 = n2143 ;
  assign y1018 = ~n2149 ;
  assign y1019 = n2150 ;
  assign y1020 = ~1'b0 ;
  assign y1021 = ~1'b0 ;
  assign y1022 = ~1'b0 ;
  assign y1023 = ~1'b0 ;
  assign y1024 = n1784 ;
  assign y1025 = ~1'b0 ;
  assign y1026 = ~1'b0 ;
  assign y1027 = ~n2152 ;
  assign y1028 = ~1'b0 ;
  assign y1029 = n2153 ;
  assign y1030 = n2155 ;
  assign y1031 = n2158 ;
  assign y1032 = ~n2161 ;
  assign y1033 = ~n2162 ;
  assign y1034 = ~1'b0 ;
  assign y1035 = 1'b0 ;
  assign y1036 = ~1'b0 ;
  assign y1037 = ~1'b0 ;
  assign y1038 = ~n2168 ;
  assign y1039 = n2169 ;
  assign y1040 = ~n2173 ;
  assign y1041 = ~x161 ;
  assign y1042 = n2177 ;
  assign y1043 = n2180 ;
  assign y1044 = ~1'b0 ;
  assign y1045 = ~1'b0 ;
  assign y1046 = ~1'b0 ;
  assign y1047 = ~n2181 ;
  assign y1048 = ~n2185 ;
  assign y1049 = ~n2186 ;
  assign y1050 = ~n2187 ;
  assign y1051 = ~1'b0 ;
  assign y1052 = ~1'b0 ;
  assign y1053 = ~1'b0 ;
  assign y1054 = n2188 ;
  assign y1055 = ~x157 ;
  assign y1056 = ~n2191 ;
  assign y1057 = ~1'b0 ;
  assign y1058 = ~1'b0 ;
  assign y1059 = n2197 ;
  assign y1060 = n2203 ;
  assign y1061 = ~n2208 ;
  assign y1062 = ~n2210 ;
  assign y1063 = n2216 ;
  assign y1064 = n571 ;
  assign y1065 = ~1'b0 ;
  assign y1066 = n2217 ;
  assign y1067 = ~n2225 ;
  assign y1068 = ~n2232 ;
  assign y1069 = ~n2243 ;
  assign y1070 = ~1'b0 ;
  assign y1071 = ~n2246 ;
  assign y1072 = ~n2257 ;
  assign y1073 = ~n2259 ;
  assign y1074 = ~n2260 ;
  assign y1075 = ~n2264 ;
  assign y1076 = n2269 ;
  assign y1077 = n2270 ;
  assign y1078 = ~1'b0 ;
  assign y1079 = ~n2272 ;
  assign y1080 = n2273 ;
  assign y1081 = n2185 ;
  assign y1082 = n2274 ;
  assign y1083 = ~1'b0 ;
  assign y1084 = n456 ;
  assign y1085 = ~n647 ;
  assign y1086 = n2275 ;
  assign y1087 = ~1'b0 ;
  assign y1088 = ~1'b0 ;
  assign y1089 = ~1'b0 ;
  assign y1090 = ~n2281 ;
  assign y1091 = ~n2285 ;
  assign y1092 = ~1'b0 ;
  assign y1093 = ~1'b0 ;
  assign y1094 = ~n2286 ;
  assign y1095 = n2292 ;
  assign y1096 = ~n2295 ;
  assign y1097 = ~n2296 ;
  assign y1098 = ~n2301 ;
  assign y1099 = n1345 ;
  assign y1100 = ~n2302 ;
  assign y1101 = ~1'b0 ;
  assign y1102 = ~n2303 ;
  assign y1103 = ~1'b0 ;
  assign y1104 = ~n1859 ;
  assign y1105 = n2304 ;
  assign y1106 = ~1'b0 ;
  assign y1107 = ~n2306 ;
  assign y1108 = ~n2307 ;
  assign y1109 = n2310 ;
  assign y1110 = ~1'b0 ;
  assign y1111 = ~n2311 ;
  assign y1112 = ~n2315 ;
  assign y1113 = ~1'b0 ;
  assign y1114 = ~1'b0 ;
  assign y1115 = ~1'b0 ;
  assign y1116 = 1'b0 ;
  assign y1117 = ~n2325 ;
  assign y1118 = n2326 ;
  assign y1119 = ~n2340 ;
  assign y1120 = ~1'b0 ;
  assign y1121 = n2345 ;
  assign y1122 = ~1'b0 ;
  assign y1123 = ~n2352 ;
  assign y1124 = ~n1883 ;
  assign y1125 = n2356 ;
  assign y1126 = ~n2364 ;
  assign y1127 = ~1'b0 ;
  assign y1128 = n2366 ;
  assign y1129 = n2367 ;
  assign y1130 = n2371 ;
  assign y1131 = n2373 ;
  assign y1132 = n2374 ;
  assign y1133 = n2378 ;
  assign y1134 = n2379 ;
  assign y1135 = ~1'b0 ;
  assign y1136 = ~1'b0 ;
  assign y1137 = ~1'b0 ;
  assign y1138 = n2380 ;
  assign y1139 = ~1'b0 ;
  assign y1140 = ~1'b0 ;
  assign y1141 = ~n2382 ;
  assign y1142 = ~n2384 ;
  assign y1143 = ~1'b0 ;
  assign y1144 = ~1'b0 ;
  assign y1145 = ~n2391 ;
  assign y1146 = ~1'b0 ;
  assign y1147 = n2397 ;
  assign y1148 = ~1'b0 ;
  assign y1149 = x130 ;
  assign y1150 = n2400 ;
  assign y1151 = n2404 ;
  assign y1152 = n2406 ;
  assign y1153 = n2408 ;
  assign y1154 = ~n2409 ;
  assign y1155 = ~n1419 ;
  assign y1156 = n2418 ;
  assign y1157 = n2420 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = ~1'b0 ;
  assign y1160 = ~1'b0 ;
  assign y1161 = ~n2425 ;
  assign y1162 = ~n1877 ;
  assign y1163 = ~n2426 ;
  assign y1164 = ~1'b0 ;
  assign y1165 = ~1'b0 ;
  assign y1166 = ~n2428 ;
  assign y1167 = ~1'b0 ;
  assign y1168 = ~n2435 ;
  assign y1169 = ~n2436 ;
  assign y1170 = n2438 ;
  assign y1171 = ~1'b0 ;
  assign y1172 = ~1'b0 ;
  assign y1173 = ~1'b0 ;
  assign y1174 = n2439 ;
  assign y1175 = n2440 ;
  assign y1176 = n2447 ;
  assign y1177 = ~1'b0 ;
  assign y1178 = ~1'b0 ;
  assign y1179 = n2451 ;
  assign y1180 = ~1'b0 ;
  assign y1181 = ~1'b0 ;
  assign y1182 = ~n2454 ;
  assign y1183 = ~1'b0 ;
  assign y1184 = ~1'b0 ;
  assign y1185 = ~n2457 ;
  assign y1186 = n2459 ;
  assign y1187 = ~1'b0 ;
  assign y1188 = n2463 ;
  assign y1189 = n2465 ;
  assign y1190 = 1'b0 ;
  assign y1191 = n2466 ;
  assign y1192 = ~1'b0 ;
  assign y1193 = ~1'b0 ;
  assign y1194 = ~1'b0 ;
  assign y1195 = n2469 ;
  assign y1196 = ~n2474 ;
  assign y1197 = x174 ;
  assign y1198 = n2480 ;
  assign y1199 = n2482 ;
  assign y1200 = ~n2484 ;
  assign y1201 = n2486 ;
  assign y1202 = ~1'b0 ;
  assign y1203 = n2188 ;
  assign y1204 = 1'b0 ;
  assign y1205 = ~n2487 ;
  assign y1206 = ~n2491 ;
  assign y1207 = n2492 ;
  assign y1208 = n2496 ;
  assign y1209 = n2498 ;
  assign y1210 = ~1'b0 ;
  assign y1211 = ~n2500 ;
  assign y1212 = ~1'b0 ;
  assign y1213 = n2502 ;
  assign y1214 = ~n2503 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = ~n2508 ;
  assign y1217 = ~1'b0 ;
  assign y1218 = ~n2511 ;
  assign y1219 = n1529 ;
  assign y1220 = ~1'b0 ;
  assign y1221 = ~n2515 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = ~n2516 ;
  assign y1224 = n2517 ;
  assign y1225 = n2518 ;
  assign y1226 = ~1'b0 ;
  assign y1227 = ~n2519 ;
  assign y1228 = ~n2523 ;
  assign y1229 = n2526 ;
  assign y1230 = ~n2420 ;
  assign y1231 = n2324 ;
  assign y1232 = n2527 ;
  assign y1233 = n2542 ;
  assign y1234 = ~1'b0 ;
  assign y1235 = n2544 ;
  assign y1236 = ~1'b0 ;
  assign y1237 = ~x6 ;
  assign y1238 = ~1'b0 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = ~n2547 ;
  assign y1241 = ~1'b0 ;
  assign y1242 = n2549 ;
  assign y1243 = ~1'b0 ;
  assign y1244 = ~n2550 ;
  assign y1245 = 1'b0 ;
  assign y1246 = n2554 ;
  assign y1247 = ~1'b0 ;
  assign y1248 = ~n2561 ;
  assign y1249 = n2562 ;
  assign y1250 = n2564 ;
  assign y1251 = ~1'b0 ;
  assign y1252 = ~n2568 ;
  assign y1253 = n2585 ;
  assign y1254 = ~1'b0 ;
  assign y1255 = n2586 ;
  assign y1256 = n2587 ;
  assign y1257 = ~1'b0 ;
  assign y1258 = n2593 ;
  assign y1259 = n1732 ;
  assign y1260 = 1'b0 ;
  assign y1261 = ~1'b0 ;
  assign y1262 = n2602 ;
  assign y1263 = ~1'b0 ;
  assign y1264 = n2607 ;
  assign y1265 = ~1'b0 ;
  assign y1266 = ~n2609 ;
  assign y1267 = n2610 ;
  assign y1268 = ~1'b0 ;
  assign y1269 = n2611 ;
  assign y1270 = 1'b0 ;
  assign y1271 = n2616 ;
  assign y1272 = ~1'b0 ;
  assign y1273 = ~1'b0 ;
  assign y1274 = n2618 ;
  assign y1275 = n2620 ;
  assign y1276 = ~1'b0 ;
  assign y1277 = n2624 ;
  assign y1278 = ~1'b0 ;
  assign y1279 = n2627 ;
  assign y1280 = n2629 ;
  assign y1281 = n2630 ;
  assign y1282 = ~1'b0 ;
  assign y1283 = ~n2634 ;
  assign y1284 = ~n2636 ;
  assign y1285 = ~n2637 ;
  assign y1286 = n2639 ;
  assign y1287 = n2640 ;
  assign y1288 = x65 ;
  assign y1289 = ~n2642 ;
  assign y1290 = ~1'b0 ;
  assign y1291 = ~1'b0 ;
  assign y1292 = ~n2644 ;
  assign y1293 = n2647 ;
  assign y1294 = ~n2650 ;
  assign y1295 = n2653 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~1'b0 ;
  assign y1298 = n2665 ;
  assign y1299 = ~n1646 ;
  assign y1300 = n2667 ;
  assign y1301 = ~1'b0 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = n2669 ;
  assign y1304 = n2671 ;
  assign y1305 = n1738 ;
  assign y1306 = ~1'b0 ;
  assign y1307 = n2675 ;
  assign y1308 = ~n2676 ;
  assign y1309 = ~n1832 ;
  assign y1310 = ~n2677 ;
  assign y1311 = ~n519 ;
  assign y1312 = ~n2426 ;
  assign y1313 = ~n2682 ;
  assign y1314 = ~n2686 ;
  assign y1315 = ~n2689 ;
  assign y1316 = ~n2691 ;
  assign y1317 = n2697 ;
  assign y1318 = n2698 ;
  assign y1319 = ~1'b0 ;
  assign y1320 = ~1'b0 ;
  assign y1321 = ~1'b0 ;
  assign y1322 = ~n2700 ;
  assign y1323 = n2701 ;
  assign y1324 = ~1'b0 ;
  assign y1325 = n2702 ;
  assign y1326 = ~1'b0 ;
  assign y1327 = ~1'b0 ;
  assign y1328 = ~1'b0 ;
  assign y1329 = ~n2706 ;
  assign y1330 = ~1'b0 ;
  assign y1331 = n2707 ;
  assign y1332 = ~n2709 ;
  assign y1333 = ~1'b0 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = ~n2720 ;
  assign y1336 = ~1'b0 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = ~1'b0 ;
  assign y1339 = ~n381 ;
  assign y1340 = n2725 ;
  assign y1341 = ~1'b0 ;
  assign y1342 = ~n2731 ;
  assign y1343 = n2737 ;
  assign y1344 = n2741 ;
  assign y1345 = ~n2743 ;
  assign y1346 = n2744 ;
  assign y1347 = n2746 ;
  assign y1348 = ~n2750 ;
  assign y1349 = ~1'b0 ;
  assign y1350 = 1'b0 ;
  assign y1351 = n2755 ;
  assign y1352 = n2764 ;
  assign y1353 = 1'b0 ;
  assign y1354 = n2766 ;
  assign y1355 = ~n2770 ;
  assign y1356 = ~1'b0 ;
  assign y1357 = ~n2774 ;
  assign y1358 = n2778 ;
  assign y1359 = n2779 ;
  assign y1360 = ~1'b0 ;
  assign y1361 = n2786 ;
  assign y1362 = n2310 ;
  assign y1363 = ~n2787 ;
  assign y1364 = 1'b0 ;
  assign y1365 = ~n2791 ;
  assign y1366 = ~n2793 ;
  assign y1367 = ~1'b0 ;
  assign y1368 = ~1'b0 ;
  assign y1369 = n2798 ;
  assign y1370 = ~n2799 ;
  assign y1371 = ~n2801 ;
  assign y1372 = ~n2803 ;
  assign y1373 = n2812 ;
  assign y1374 = ~1'b0 ;
  assign y1375 = ~1'b0 ;
  assign y1376 = n2820 ;
  assign y1377 = n1521 ;
  assign y1378 = n2822 ;
  assign y1379 = ~n2826 ;
  assign y1380 = ~1'b0 ;
  assign y1381 = ~1'b0 ;
  assign y1382 = n2827 ;
  assign y1383 = n2828 ;
  assign y1384 = n2830 ;
  assign y1385 = ~1'b0 ;
  assign y1386 = ~1'b0 ;
  assign y1387 = ~n2836 ;
  assign y1388 = n2837 ;
  assign y1389 = ~1'b0 ;
  assign y1390 = ~1'b0 ;
  assign y1391 = 1'b0 ;
  assign y1392 = n2838 ;
  assign y1393 = ~1'b0 ;
  assign y1394 = ~1'b0 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = ~1'b0 ;
  assign y1397 = n2465 ;
  assign y1398 = n2839 ;
  assign y1399 = ~n2841 ;
  assign y1400 = ~1'b0 ;
  assign y1401 = ~n2844 ;
  assign y1402 = ~n2845 ;
  assign y1403 = ~1'b0 ;
  assign y1404 = ~n2846 ;
  assign y1405 = ~n1080 ;
  assign y1406 = ~n2849 ;
  assign y1407 = ~1'b0 ;
  assign y1408 = ~1'b0 ;
  assign y1409 = n2851 ;
  assign y1410 = ~1'b0 ;
  assign y1411 = ~1'b0 ;
  assign y1412 = ~n553 ;
  assign y1413 = n2857 ;
  assign y1414 = ~1'b0 ;
  assign y1415 = n2867 ;
  assign y1416 = ~n2868 ;
  assign y1417 = n2870 ;
  assign y1418 = ~n2668 ;
  assign y1419 = ~1'b0 ;
  assign y1420 = ~n1488 ;
  assign y1421 = n2871 ;
  assign y1422 = ~1'b0 ;
  assign y1423 = ~n2872 ;
  assign y1424 = n2875 ;
  assign y1425 = n2878 ;
  assign y1426 = ~1'b0 ;
  assign y1427 = ~n2776 ;
  assign y1428 = ~1'b0 ;
  assign y1429 = 1'b0 ;
  assign y1430 = n2175 ;
  assign y1431 = ~n2887 ;
  assign y1432 = ~1'b0 ;
  assign y1433 = ~1'b0 ;
  assign y1434 = ~n2599 ;
  assign y1435 = ~n2892 ;
  assign y1436 = ~n1337 ;
  assign y1437 = n2897 ;
  assign y1438 = n2900 ;
  assign y1439 = n2901 ;
  assign y1440 = ~n2902 ;
  assign y1441 = ~1'b0 ;
  assign y1442 = ~n2906 ;
  assign y1443 = n1622 ;
  assign y1444 = n2908 ;
  assign y1445 = ~1'b0 ;
  assign y1446 = ~1'b0 ;
  assign y1447 = n2910 ;
  assign y1448 = ~n2911 ;
  assign y1449 = 1'b0 ;
  assign y1450 = ~n2916 ;
  assign y1451 = ~n2922 ;
  assign y1452 = ~1'b0 ;
  assign y1453 = n2932 ;
  assign y1454 = ~n2936 ;
  assign y1455 = ~n2938 ;
  assign y1456 = n2942 ;
  assign y1457 = ~n2951 ;
  assign y1458 = n2955 ;
  assign y1459 = ~1'b0 ;
  assign y1460 = ~n2957 ;
  assign y1461 = n2959 ;
  assign y1462 = n2961 ;
  assign y1463 = ~n2964 ;
  assign y1464 = ~1'b0 ;
  assign y1465 = n2968 ;
  assign y1466 = ~1'b0 ;
  assign y1467 = ~1'b0 ;
  assign y1468 = n2972 ;
  assign y1469 = n2976 ;
  assign y1470 = ~1'b0 ;
  assign y1471 = ~1'b0 ;
  assign y1472 = n2978 ;
  assign y1473 = ~n2849 ;
  assign y1474 = ~n2983 ;
  assign y1475 = n2986 ;
  assign y1476 = n2991 ;
  assign y1477 = ~1'b0 ;
  assign y1478 = ~1'b0 ;
  assign y1479 = ~1'b0 ;
  assign y1480 = ~1'b0 ;
  assign y1481 = ~n3000 ;
  assign y1482 = n3003 ;
  assign y1483 = ~n3013 ;
  assign y1484 = ~n458 ;
  assign y1485 = ~1'b0 ;
  assign y1486 = 1'b0 ;
  assign y1487 = n3014 ;
  assign y1488 = n3015 ;
  assign y1489 = ~1'b0 ;
  assign y1490 = ~1'b0 ;
  assign y1491 = n3016 ;
  assign y1492 = 1'b0 ;
  assign y1493 = ~n1814 ;
  assign y1494 = ~1'b0 ;
  assign y1495 = ~1'b0 ;
  assign y1496 = ~1'b0 ;
  assign y1497 = n3017 ;
  assign y1498 = n1415 ;
  assign y1499 = n1038 ;
  assign y1500 = ~n3022 ;
  assign y1501 = n3026 ;
  assign y1502 = ~n3027 ;
  assign y1503 = n3028 ;
  assign y1504 = n3033 ;
  assign y1505 = ~n3036 ;
  assign y1506 = ~n3039 ;
  assign y1507 = ~n3040 ;
  assign y1508 = ~n3045 ;
  assign y1509 = ~1'b0 ;
  assign y1510 = ~1'b0 ;
  assign y1511 = n3046 ;
  assign y1512 = n3047 ;
  assign y1513 = ~n3049 ;
  assign y1514 = ~n3052 ;
  assign y1515 = n3054 ;
  assign y1516 = ~1'b0 ;
  assign y1517 = ~1'b0 ;
  assign y1518 = ~n3055 ;
  assign y1519 = n3060 ;
  assign y1520 = ~n3064 ;
  assign y1521 = n3068 ;
  assign y1522 = ~n3069 ;
  assign y1523 = ~1'b0 ;
  assign y1524 = ~1'b0 ;
  assign y1525 = n3073 ;
  assign y1526 = ~n3076 ;
  assign y1527 = ~1'b0 ;
  assign y1528 = ~1'b0 ;
  assign y1529 = ~n3080 ;
  assign y1530 = ~n3081 ;
  assign y1531 = ~1'b0 ;
  assign y1532 = n3082 ;
  assign y1533 = n3090 ;
  assign y1534 = 1'b0 ;
  assign y1535 = ~1'b0 ;
  assign y1536 = ~n3095 ;
  assign y1537 = ~n3100 ;
  assign y1538 = n3105 ;
  assign y1539 = ~n3114 ;
  assign y1540 = ~n3115 ;
  assign y1541 = n3116 ;
  assign y1542 = ~n3117 ;
  assign y1543 = n3118 ;
  assign y1544 = ~n3122 ;
  assign y1545 = n1738 ;
  assign y1546 = 1'b0 ;
  assign y1547 = ~1'b0 ;
  assign y1548 = n3124 ;
  assign y1549 = ~n3126 ;
  assign y1550 = n3128 ;
  assign y1551 = ~n3135 ;
  assign y1552 = ~1'b0 ;
  assign y1553 = ~n263 ;
  assign y1554 = ~1'b0 ;
  assign y1555 = ~n3136 ;
  assign y1556 = 1'b0 ;
  assign y1557 = ~1'b0 ;
  assign y1558 = ~1'b0 ;
  assign y1559 = ~n3142 ;
  assign y1560 = n3144 ;
  assign y1561 = n3152 ;
  assign y1562 = ~n1353 ;
  assign y1563 = ~1'b0 ;
  assign y1564 = ~n3153 ;
  assign y1565 = n3154 ;
  assign y1566 = ~n3159 ;
  assign y1567 = ~n3162 ;
  assign y1568 = ~1'b0 ;
  assign y1569 = ~n3165 ;
  assign y1570 = ~1'b0 ;
  assign y1571 = n3166 ;
  assign y1572 = n3167 ;
  assign y1573 = ~1'b0 ;
  assign y1574 = ~n3169 ;
  assign y1575 = ~1'b0 ;
  assign y1576 = n3171 ;
  assign y1577 = ~n3175 ;
  assign y1578 = ~n3180 ;
  assign y1579 = n1164 ;
  assign y1580 = ~n3181 ;
  assign y1581 = ~n3182 ;
  assign y1582 = ~n3184 ;
  assign y1583 = ~1'b0 ;
  assign y1584 = ~1'b0 ;
  assign y1585 = n3189 ;
  assign y1586 = n3193 ;
  assign y1587 = ~n3198 ;
  assign y1588 = n3199 ;
  assign y1589 = ~n3200 ;
  assign y1590 = ~1'b0 ;
  assign y1591 = ~1'b0 ;
  assign y1592 = n3207 ;
  assign y1593 = ~n3213 ;
  assign y1594 = ~1'b0 ;
  assign y1595 = ~n3217 ;
  assign y1596 = ~n3223 ;
  assign y1597 = n2350 ;
  assign y1598 = ~n3224 ;
  assign y1599 = n3227 ;
  assign y1600 = ~1'b0 ;
  assign y1601 = ~n3234 ;
  assign y1602 = ~n3237 ;
  assign y1603 = n3242 ;
  assign y1604 = ~n3243 ;
  assign y1605 = n3245 ;
  assign y1606 = 1'b0 ;
  assign y1607 = n3248 ;
  assign y1608 = n3250 ;
  assign y1609 = n1661 ;
  assign y1610 = n3257 ;
  assign y1611 = 1'b0 ;
  assign y1612 = ~n3258 ;
  assign y1613 = ~n3260 ;
  assign y1614 = ~n3262 ;
  assign y1615 = n3265 ;
  assign y1616 = n3267 ;
  assign y1617 = ~n3274 ;
  assign y1618 = n3275 ;
  assign y1619 = ~1'b0 ;
  assign y1620 = n3278 ;
  assign y1621 = ~n3283 ;
  assign y1622 = ~n3287 ;
  assign y1623 = n3294 ;
  assign y1624 = n3297 ;
  assign y1625 = ~1'b0 ;
  assign y1626 = ~n3298 ;
  assign y1627 = ~n3303 ;
  assign y1628 = ~n3097 ;
  assign y1629 = n3305 ;
  assign y1630 = n3307 ;
  assign y1631 = ~1'b0 ;
  assign y1632 = ~n3310 ;
  assign y1633 = ~1'b0 ;
  assign y1634 = ~n3313 ;
  assign y1635 = ~1'b0 ;
  assign y1636 = n3316 ;
  assign y1637 = ~n3318 ;
  assign y1638 = ~n3321 ;
  assign y1639 = n2633 ;
  assign y1640 = ~1'b0 ;
  assign y1641 = n3322 ;
  assign y1642 = ~1'b0 ;
  assign y1643 = n1628 ;
  assign y1644 = n639 ;
  assign y1645 = n3326 ;
  assign y1646 = ~n3329 ;
  assign y1647 = ~n3332 ;
  assign y1648 = ~n3333 ;
  assign y1649 = ~n3336 ;
  assign y1650 = ~n3337 ;
  assign y1651 = ~n3339 ;
  assign y1652 = ~1'b0 ;
  assign y1653 = ~1'b0 ;
  assign y1654 = ~n700 ;
  assign y1655 = ~n3340 ;
  assign y1656 = ~n3343 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~n3346 ;
  assign y1659 = n3351 ;
  assign y1660 = ~n3353 ;
  assign y1661 = n3356 ;
  assign y1662 = ~n3360 ;
  assign y1663 = n3362 ;
  assign y1664 = ~n3367 ;
  assign y1665 = 1'b0 ;
  assign y1666 = n3378 ;
  assign y1667 = ~1'b0 ;
  assign y1668 = n3379 ;
  assign y1669 = ~n3383 ;
  assign y1670 = ~n3386 ;
  assign y1671 = n3387 ;
  assign y1672 = n3388 ;
  assign y1673 = ~1'b0 ;
  assign y1674 = ~n3083 ;
  assign y1675 = n3390 ;
  assign y1676 = 1'b0 ;
  assign y1677 = ~n3392 ;
  assign y1678 = n3393 ;
  assign y1679 = n3399 ;
  assign y1680 = ~n3403 ;
  assign y1681 = n3407 ;
  assign y1682 = n3408 ;
  assign y1683 = 1'b0 ;
  assign y1684 = n3409 ;
  assign y1685 = n3410 ;
  assign y1686 = n3414 ;
  assign y1687 = ~n3415 ;
  assign y1688 = ~n3416 ;
  assign y1689 = n3417 ;
  assign y1690 = ~n3420 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = ~n3423 ;
  assign y1693 = n1961 ;
  assign y1694 = ~1'b0 ;
  assign y1695 = n3424 ;
  assign y1696 = ~n3430 ;
  assign y1697 = ~1'b0 ;
  assign y1698 = n3431 ;
  assign y1699 = x27 ;
  assign y1700 = ~1'b0 ;
  assign y1701 = ~1'b0 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = 1'b0 ;
  assign y1704 = n3432 ;
  assign y1705 = ~n3434 ;
  assign y1706 = ~x3 ;
  assign y1707 = n2812 ;
  assign y1708 = ~1'b0 ;
  assign y1709 = ~x176 ;
  assign y1710 = ~1'b0 ;
  assign y1711 = ~n3438 ;
  assign y1712 = ~1'b0 ;
  assign y1713 = n3440 ;
  assign y1714 = n3442 ;
  assign y1715 = ~1'b0 ;
  assign y1716 = n3443 ;
  assign y1717 = ~n3446 ;
  assign y1718 = ~1'b0 ;
  assign y1719 = ~n3448 ;
  assign y1720 = ~1'b0 ;
  assign y1721 = n3454 ;
  assign y1722 = n1890 ;
  assign y1723 = ~n3458 ;
  assign y1724 = ~1'b0 ;
  assign y1725 = ~n3461 ;
  assign y1726 = n3463 ;
  assign y1727 = ~1'b0 ;
  assign y1728 = n3467 ;
  assign y1729 = ~1'b0 ;
  assign y1730 = ~1'b0 ;
  assign y1731 = n3469 ;
  assign y1732 = n3476 ;
  assign y1733 = ~1'b0 ;
  assign y1734 = n2143 ;
  assign y1735 = 1'b0 ;
  assign y1736 = ~n3477 ;
  assign y1737 = ~1'b0 ;
  assign y1738 = ~n3479 ;
  assign y1739 = n3481 ;
  assign y1740 = n3484 ;
  assign y1741 = 1'b0 ;
  assign y1742 = n3491 ;
  assign y1743 = ~1'b0 ;
  assign y1744 = ~1'b0 ;
  assign y1745 = ~n3492 ;
  assign y1746 = 1'b0 ;
  assign y1747 = n3496 ;
  assign y1748 = ~1'b0 ;
  assign y1749 = n3499 ;
  assign y1750 = ~n3158 ;
  assign y1751 = n1678 ;
  assign y1752 = ~1'b0 ;
  assign y1753 = ~n3503 ;
  assign y1754 = 1'b0 ;
  assign y1755 = ~1'b0 ;
  assign y1756 = n3431 ;
  assign y1757 = ~1'b0 ;
  assign y1758 = ~n3059 ;
  assign y1759 = ~1'b0 ;
  assign y1760 = ~1'b0 ;
  assign y1761 = ~1'b0 ;
  assign y1762 = n401 ;
  assign y1763 = ~n3505 ;
  assign y1764 = ~n3509 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = ~n3514 ;
  assign y1767 = ~1'b0 ;
  assign y1768 = ~n3458 ;
  assign y1769 = ~n3516 ;
  assign y1770 = ~n3518 ;
  assign y1771 = ~n3521 ;
  assign y1772 = n2655 ;
  assign y1773 = n3526 ;
  assign y1774 = ~n3528 ;
  assign y1775 = ~1'b0 ;
  assign y1776 = n3045 ;
  assign y1777 = ~1'b0 ;
  assign y1778 = ~1'b0 ;
  assign y1779 = ~n3529 ;
  assign y1780 = n3531 ;
  assign y1781 = ~n3532 ;
  assign y1782 = n3533 ;
  assign y1783 = ~n749 ;
  assign y1784 = ~n3536 ;
  assign y1785 = ~n3539 ;
  assign y1786 = n3541 ;
  assign y1787 = ~1'b0 ;
  assign y1788 = n3543 ;
  assign y1789 = ~n3548 ;
  assign y1790 = ~1'b0 ;
  assign y1791 = ~n3549 ;
  assign y1792 = n3555 ;
  assign y1793 = ~1'b0 ;
  assign y1794 = ~1'b0 ;
  assign y1795 = n3556 ;
  assign y1796 = n3558 ;
  assign y1797 = ~1'b0 ;
  assign y1798 = ~n509 ;
  assign y1799 = n3559 ;
  assign y1800 = ~n3561 ;
  assign y1801 = ~1'b0 ;
  assign y1802 = n3563 ;
  assign y1803 = ~n3567 ;
  assign y1804 = ~n3569 ;
  assign y1805 = ~1'b0 ;
  assign y1806 = ~n3575 ;
  assign y1807 = ~1'b0 ;
  assign y1808 = ~1'b0 ;
  assign y1809 = ~1'b0 ;
  assign y1810 = ~n3576 ;
  assign y1811 = ~x98 ;
  assign y1812 = ~n3578 ;
  assign y1813 = ~1'b0 ;
  assign y1814 = ~1'b0 ;
  assign y1815 = ~n3580 ;
  assign y1816 = ~n3582 ;
  assign y1817 = ~n3590 ;
  assign y1818 = ~1'b0 ;
  assign y1819 = ~n3593 ;
  assign y1820 = n3608 ;
  assign y1821 = ~1'b0 ;
  assign y1822 = ~n3613 ;
  assign y1823 = ~n3621 ;
  assign y1824 = ~1'b0 ;
  assign y1825 = ~1'b0 ;
  assign y1826 = ~1'b0 ;
  assign y1827 = ~n3626 ;
  assign y1828 = ~1'b0 ;
  assign y1829 = ~n3629 ;
  assign y1830 = 1'b0 ;
  assign y1831 = n3630 ;
  assign y1832 = ~n3632 ;
  assign y1833 = ~n3635 ;
  assign y1834 = ~n3641 ;
  assign y1835 = ~n519 ;
  assign y1836 = ~n3647 ;
  assign y1837 = ~1'b0 ;
  assign y1838 = n3648 ;
  assign y1839 = x160 ;
  assign y1840 = ~n2949 ;
  assign y1841 = n3651 ;
  assign y1842 = ~n3656 ;
  assign y1843 = ~n3657 ;
  assign y1844 = ~x115 ;
  assign y1845 = ~n3664 ;
  assign y1846 = ~n3667 ;
  assign y1847 = n3670 ;
  assign y1848 = ~1'b0 ;
  assign y1849 = ~1'b0 ;
  assign y1850 = n3672 ;
  assign y1851 = ~n3676 ;
  assign y1852 = ~1'b0 ;
  assign y1853 = ~1'b0 ;
  assign y1854 = ~n3681 ;
  assign y1855 = ~n3685 ;
  assign y1856 = ~n3688 ;
  assign y1857 = ~n3689 ;
  assign y1858 = n3692 ;
  assign y1859 = ~1'b0 ;
  assign y1860 = n836 ;
  assign y1861 = ~1'b0 ;
  assign y1862 = ~1'b0 ;
  assign y1863 = ~1'b0 ;
  assign y1864 = ~n3695 ;
  assign y1865 = ~n631 ;
  assign y1866 = 1'b0 ;
  assign y1867 = n3698 ;
  assign y1868 = n1485 ;
  assign y1869 = n3702 ;
  assign y1870 = ~n3703 ;
  assign y1871 = n3705 ;
  assign y1872 = ~1'b0 ;
  assign y1873 = ~1'b0 ;
  assign y1874 = ~1'b0 ;
  assign y1875 = ~n3709 ;
  assign y1876 = n3710 ;
  assign y1877 = ~1'b0 ;
  assign y1878 = ~n3711 ;
  assign y1879 = 1'b0 ;
  assign y1880 = n3714 ;
  assign y1881 = n1623 ;
  assign y1882 = ~n3715 ;
  assign y1883 = ~n3718 ;
  assign y1884 = n3720 ;
  assign y1885 = ~n3721 ;
  assign y1886 = ~n3723 ;
  assign y1887 = n3725 ;
  assign y1888 = ~n3726 ;
  assign y1889 = ~n3727 ;
  assign y1890 = n3733 ;
  assign y1891 = ~1'b0 ;
  assign y1892 = ~1'b0 ;
  assign y1893 = ~n3739 ;
  assign y1894 = ~1'b0 ;
  assign y1895 = ~n3742 ;
  assign y1896 = ~1'b0 ;
  assign y1897 = n3745 ;
  assign y1898 = ~n3748 ;
  assign y1899 = ~n3749 ;
  assign y1900 = ~n3750 ;
  assign y1901 = ~1'b0 ;
  assign y1902 = ~n3751 ;
  assign y1903 = n3754 ;
  assign y1904 = ~n3755 ;
  assign y1905 = n3756 ;
  assign y1906 = ~n3759 ;
  assign y1907 = n3760 ;
  assign y1908 = ~n3762 ;
  assign y1909 = n3763 ;
  assign y1910 = ~1'b0 ;
  assign y1911 = n3764 ;
  assign y1912 = ~1'b0 ;
  assign y1913 = n3766 ;
  assign y1914 = n3768 ;
  assign y1915 = ~1'b0 ;
  assign y1916 = ~1'b0 ;
  assign y1917 = ~1'b0 ;
  assign y1918 = ~1'b0 ;
  assign y1919 = ~n3770 ;
  assign y1920 = n3772 ;
  assign y1921 = ~n2120 ;
  assign y1922 = 1'b0 ;
  assign y1923 = ~1'b0 ;
  assign y1924 = ~n3773 ;
  assign y1925 = ~n3779 ;
  assign y1926 = n3780 ;
  assign y1927 = ~1'b0 ;
  assign y1928 = ~n3781 ;
  assign y1929 = ~n3784 ;
  assign y1930 = n3786 ;
  assign y1931 = n3791 ;
  assign y1932 = n3792 ;
  assign y1933 = n3794 ;
  assign y1934 = ~1'b0 ;
  assign y1935 = ~n3795 ;
  assign y1936 = n3796 ;
  assign y1937 = n3802 ;
  assign y1938 = ~n3805 ;
  assign y1939 = 1'b0 ;
  assign y1940 = ~n3703 ;
  assign y1941 = n3807 ;
  assign y1942 = ~n3809 ;
  assign y1943 = ~1'b0 ;
  assign y1944 = ~n3810 ;
  assign y1945 = ~1'b0 ;
  assign y1946 = ~n3811 ;
  assign y1947 = ~1'b0 ;
  assign y1948 = n3817 ;
  assign y1949 = 1'b0 ;
  assign y1950 = n3820 ;
  assign y1951 = n3833 ;
  assign y1952 = ~n3834 ;
  assign y1953 = ~n3836 ;
  assign y1954 = ~n3841 ;
  assign y1955 = n3842 ;
  assign y1956 = ~n3845 ;
  assign y1957 = ~1'b0 ;
  assign y1958 = ~1'b0 ;
  assign y1959 = ~1'b0 ;
  assign y1960 = ~n3850 ;
  assign y1961 = ~1'b0 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = n3852 ;
  assign y1964 = ~n3854 ;
  assign y1965 = ~1'b0 ;
  assign y1966 = ~n3856 ;
  assign y1967 = ~n3859 ;
  assign y1968 = ~n3860 ;
  assign y1969 = ~1'b0 ;
  assign y1970 = n3866 ;
  assign y1971 = ~1'b0 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = ~n3870 ;
  assign y1974 = ~1'b0 ;
  assign y1975 = n3872 ;
  assign y1976 = n3875 ;
  assign y1977 = n1361 ;
  assign y1978 = n3878 ;
  assign y1979 = n3879 ;
  assign y1980 = ~1'b0 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = n3883 ;
  assign y1983 = ~1'b0 ;
  assign y1984 = ~n3823 ;
  assign y1985 = ~1'b0 ;
  assign y1986 = ~n3888 ;
  assign y1987 = n3891 ;
  assign y1988 = ~n3893 ;
  assign y1989 = ~n3906 ;
  assign y1990 = n3911 ;
  assign y1991 = n3913 ;
  assign y1992 = ~n1271 ;
  assign y1993 = 1'b0 ;
  assign y1994 = ~1'b0 ;
  assign y1995 = n3914 ;
  assign y1996 = ~1'b0 ;
  assign y1997 = ~n3917 ;
  assign y1998 = ~1'b0 ;
  assign y1999 = ~n3920 ;
  assign y2000 = ~n3922 ;
  assign y2001 = ~1'b0 ;
  assign y2002 = n3925 ;
  assign y2003 = n3936 ;
  assign y2004 = n3938 ;
  assign y2005 = ~n3940 ;
  assign y2006 = ~n3943 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = n3946 ;
  assign y2009 = ~n3948 ;
  assign y2010 = ~n3950 ;
  assign y2011 = ~n3951 ;
  assign y2012 = ~1'b0 ;
  assign y2013 = n3956 ;
  assign y2014 = ~n3960 ;
  assign y2015 = n3964 ;
  assign y2016 = ~1'b0 ;
  assign y2017 = n3965 ;
  assign y2018 = 1'b0 ;
  assign y2019 = n3966 ;
  assign y2020 = ~n3970 ;
  assign y2021 = ~1'b0 ;
  assign y2022 = ~n3971 ;
  assign y2023 = n3974 ;
  assign y2024 = ~1'b0 ;
  assign y2025 = ~1'b0 ;
  assign y2026 = n3976 ;
  assign y2027 = n3982 ;
  assign y2028 = n3984 ;
  assign y2029 = n3988 ;
  assign y2030 = ~n3991 ;
  assign y2031 = ~n3993 ;
  assign y2032 = ~1'b0 ;
  assign y2033 = ~1'b0 ;
  assign y2034 = ~1'b0 ;
  assign y2035 = n3994 ;
  assign y2036 = ~1'b0 ;
  assign y2037 = ~1'b0 ;
  assign y2038 = n3995 ;
  assign y2039 = ~n3996 ;
  assign y2040 = ~1'b0 ;
  assign y2041 = ~n3998 ;
  assign y2042 = n3678 ;
  assign y2043 = ~1'b0 ;
  assign y2044 = ~1'b0 ;
  assign y2045 = ~n4001 ;
  assign y2046 = ~1'b0 ;
  assign y2047 = n3145 ;
  assign y2048 = ~n4002 ;
  assign y2049 = ~1'b0 ;
  assign y2050 = ~n4003 ;
  assign y2051 = ~n4005 ;
  assign y2052 = ~1'b0 ;
  assign y2053 = ~n1264 ;
  assign y2054 = n4008 ;
  assign y2055 = ~1'b0 ;
  assign y2056 = ~n4009 ;
  assign y2057 = ~1'b0 ;
  assign y2058 = ~n4012 ;
  assign y2059 = ~1'b0 ;
  assign y2060 = ~1'b0 ;
  assign y2061 = ~n4013 ;
  assign y2062 = n4014 ;
  assign y2063 = n4016 ;
  assign y2064 = ~1'b0 ;
  assign y2065 = ~1'b0 ;
  assign y2066 = ~n4020 ;
  assign y2067 = ~n4021 ;
  assign y2068 = n4022 ;
  assign y2069 = ~1'b0 ;
  assign y2070 = ~1'b0 ;
  assign y2071 = ~n4024 ;
  assign y2072 = n2970 ;
  assign y2073 = ~1'b0 ;
  assign y2074 = n4027 ;
  assign y2075 = ~1'b0 ;
  assign y2076 = ~1'b0 ;
  assign y2077 = ~n4029 ;
  assign y2078 = ~1'b0 ;
  assign y2079 = ~1'b0 ;
  assign y2080 = n4034 ;
  assign y2081 = ~n4035 ;
  assign y2082 = ~1'b0 ;
  assign y2083 = ~n4037 ;
  assign y2084 = ~1'b0 ;
  assign y2085 = ~1'b0 ;
  assign y2086 = ~n4043 ;
  assign y2087 = ~n4045 ;
  assign y2088 = n2237 ;
  assign y2089 = ~n3953 ;
  assign y2090 = ~n4051 ;
  assign y2091 = ~n4055 ;
  assign y2092 = ~n4059 ;
  assign y2093 = 1'b0 ;
  assign y2094 = ~n4063 ;
  assign y2095 = ~n4066 ;
  assign y2096 = ~1'b0 ;
  assign y2097 = ~1'b0 ;
  assign y2098 = n4067 ;
  assign y2099 = ~n4069 ;
  assign y2100 = 1'b0 ;
  assign y2101 = ~n4074 ;
  assign y2102 = ~1'b0 ;
  assign y2103 = n4076 ;
  assign y2104 = n4077 ;
  assign y2105 = n4079 ;
  assign y2106 = ~n825 ;
  assign y2107 = n994 ;
  assign y2108 = ~1'b0 ;
  assign y2109 = n4080 ;
  assign y2110 = n4081 ;
  assign y2111 = ~n4083 ;
  assign y2112 = n4084 ;
  assign y2113 = ~n4089 ;
  assign y2114 = n4091 ;
  assign y2115 = n4094 ;
  assign y2116 = 1'b0 ;
  assign y2117 = ~1'b0 ;
  assign y2118 = n1605 ;
  assign y2119 = ~1'b0 ;
  assign y2120 = ~n4096 ;
  assign y2121 = ~n4101 ;
  assign y2122 = n4103 ;
  assign y2123 = ~1'b0 ;
  assign y2124 = n4107 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = ~n4108 ;
  assign y2127 = ~1'b0 ;
  assign y2128 = ~n4112 ;
  assign y2129 = ~1'b0 ;
  assign y2130 = ~1'b0 ;
  assign y2131 = ~1'b0 ;
  assign y2132 = ~1'b0 ;
  assign y2133 = ~1'b0 ;
  assign y2134 = ~1'b0 ;
  assign y2135 = n4113 ;
  assign y2136 = ~1'b0 ;
  assign y2137 = ~1'b0 ;
  assign y2138 = n4116 ;
  assign y2139 = ~n4119 ;
  assign y2140 = n4129 ;
  assign y2141 = ~n4132 ;
  assign y2142 = n4136 ;
  assign y2143 = ~n4138 ;
  assign y2144 = ~1'b0 ;
  assign y2145 = ~n4143 ;
  assign y2146 = n4144 ;
  assign y2147 = ~n4147 ;
  assign y2148 = ~n4149 ;
  assign y2149 = ~1'b0 ;
  assign y2150 = ~n4156 ;
  assign y2151 = n4161 ;
  assign y2152 = n4164 ;
  assign y2153 = ~n4168 ;
  assign y2154 = ~n1111 ;
  assign y2155 = n4169 ;
  assign y2156 = ~1'b0 ;
  assign y2157 = ~n4173 ;
  assign y2158 = ~n4176 ;
  assign y2159 = ~n4178 ;
  assign y2160 = n880 ;
  assign y2161 = ~1'b0 ;
  assign y2162 = n4180 ;
  assign y2163 = ~n672 ;
  assign y2164 = ~1'b0 ;
  assign y2165 = ~n4183 ;
  assign y2166 = n2604 ;
  assign y2167 = ~n4188 ;
  assign y2168 = ~n4189 ;
  assign y2169 = ~n4197 ;
  assign y2170 = ~1'b0 ;
  assign y2171 = n4199 ;
  assign y2172 = ~1'b0 ;
  assign y2173 = ~n4201 ;
  assign y2174 = ~1'b0 ;
  assign y2175 = ~n4118 ;
  assign y2176 = ~n4205 ;
  assign y2177 = ~1'b0 ;
  assign y2178 = ~n4118 ;
  assign y2179 = ~n4207 ;
  assign y2180 = n4208 ;
  assign y2181 = ~1'b0 ;
  assign y2182 = ~1'b0 ;
  assign y2183 = ~n4211 ;
  assign y2184 = n4213 ;
  assign y2185 = n4214 ;
  assign y2186 = ~n4217 ;
  assign y2187 = ~1'b0 ;
  assign y2188 = ~1'b0 ;
  assign y2189 = ~1'b0 ;
  assign y2190 = ~n4223 ;
  assign y2191 = n4227 ;
  assign y2192 = n4238 ;
  assign y2193 = n4239 ;
  assign y2194 = n4243 ;
  assign y2195 = n4247 ;
  assign y2196 = n4251 ;
  assign y2197 = ~1'b0 ;
  assign y2198 = n4253 ;
  assign y2199 = ~n4256 ;
  assign y2200 = n4258 ;
  assign y2201 = ~n4260 ;
  assign y2202 = ~1'b0 ;
  assign y2203 = ~1'b0 ;
  assign y2204 = n4270 ;
  assign y2205 = ~x25 ;
  assign y2206 = ~1'b0 ;
  assign y2207 = ~n4274 ;
  assign y2208 = ~1'b0 ;
  assign y2209 = 1'b0 ;
  assign y2210 = ~n4276 ;
  assign y2211 = n4278 ;
  assign y2212 = ~1'b0 ;
  assign y2213 = ~n4281 ;
  assign y2214 = n4284 ;
  assign y2215 = n4287 ;
  assign y2216 = n4291 ;
  assign y2217 = ~1'b0 ;
  assign y2218 = n4296 ;
  assign y2219 = ~1'b0 ;
  assign y2220 = ~n1672 ;
  assign y2221 = n4297 ;
  assign y2222 = ~n4298 ;
  assign y2223 = 1'b0 ;
  assign y2224 = ~n4302 ;
  assign y2225 = n4304 ;
  assign y2226 = ~n4306 ;
  assign y2227 = n4308 ;
  assign y2228 = ~1'b0 ;
  assign y2229 = n4310 ;
  assign y2230 = ~n4314 ;
  assign y2231 = n4315 ;
  assign y2232 = n4316 ;
  assign y2233 = ~1'b0 ;
  assign y2234 = ~1'b0 ;
  assign y2235 = ~1'b0 ;
  assign y2236 = ~n4318 ;
  assign y2237 = n4321 ;
  assign y2238 = n4323 ;
  assign y2239 = n2760 ;
  assign y2240 = ~1'b0 ;
  assign y2241 = ~n4325 ;
  assign y2242 = ~n4327 ;
  assign y2243 = n4329 ;
  assign y2244 = ~n4336 ;
  assign y2245 = n4338 ;
  assign y2246 = ~1'b0 ;
  assign y2247 = ~1'b0 ;
  assign y2248 = ~1'b0 ;
  assign y2249 = n4343 ;
  assign y2250 = 1'b0 ;
  assign y2251 = ~1'b0 ;
  assign y2252 = n4349 ;
  assign y2253 = n4361 ;
  assign y2254 = ~1'b0 ;
  assign y2255 = ~1'b0 ;
  assign y2256 = ~1'b0 ;
  assign y2257 = ~n4366 ;
  assign y2258 = ~n4368 ;
  assign y2259 = ~n4372 ;
  assign y2260 = ~n4373 ;
  assign y2261 = ~1'b0 ;
  assign y2262 = n4376 ;
  assign y2263 = n4378 ;
  assign y2264 = ~1'b0 ;
  assign y2265 = n4380 ;
  assign y2266 = ~1'b0 ;
  assign y2267 = ~n4382 ;
  assign y2268 = x140 ;
  assign y2269 = n4386 ;
  assign y2270 = ~1'b0 ;
  assign y2271 = 1'b0 ;
  assign y2272 = ~n4390 ;
  assign y2273 = n4395 ;
  assign y2274 = ~n1594 ;
  assign y2275 = ~n4396 ;
  assign y2276 = n4398 ;
  assign y2277 = ~1'b0 ;
  assign y2278 = n4399 ;
  assign y2279 = 1'b0 ;
  assign y2280 = n461 ;
  assign y2281 = ~1'b0 ;
  assign y2282 = n4400 ;
  assign y2283 = ~1'b0 ;
  assign y2284 = n4412 ;
  assign y2285 = n4414 ;
  assign y2286 = n4416 ;
  assign y2287 = ~1'b0 ;
  assign y2288 = n4417 ;
  assign y2289 = ~1'b0 ;
  assign y2290 = ~1'b0 ;
  assign y2291 = ~n4418 ;
  assign y2292 = ~n4422 ;
  assign y2293 = ~n4423 ;
  assign y2294 = ~1'b0 ;
  assign y2295 = n4424 ;
  assign y2296 = n3226 ;
  assign y2297 = ~1'b0 ;
  assign y2298 = n4428 ;
  assign y2299 = n4430 ;
  assign y2300 = n4431 ;
  assign y2301 = n4432 ;
  assign y2302 = n4434 ;
  assign y2303 = n4436 ;
  assign y2304 = ~n4438 ;
  assign y2305 = ~n4444 ;
  assign y2306 = n4447 ;
  assign y2307 = ~1'b0 ;
  assign y2308 = ~1'b0 ;
  assign y2309 = n4448 ;
  assign y2310 = ~1'b0 ;
  assign y2311 = ~1'b0 ;
  assign y2312 = ~1'b0 ;
  assign y2313 = n4449 ;
  assign y2314 = n4451 ;
  assign y2315 = n4452 ;
  assign y2316 = ~1'b0 ;
  assign y2317 = ~n4454 ;
  assign y2318 = ~1'b0 ;
  assign y2319 = ~1'b0 ;
  assign y2320 = ~n4455 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = n4460 ;
  assign y2323 = n2561 ;
  assign y2324 = ~1'b0 ;
  assign y2325 = n4465 ;
  assign y2326 = ~n4466 ;
  assign y2327 = n4467 ;
  assign y2328 = 1'b0 ;
  assign y2329 = n4473 ;
  assign y2330 = ~1'b0 ;
  assign y2331 = ~n4475 ;
  assign y2332 = ~n4479 ;
  assign y2333 = ~1'b0 ;
  assign y2334 = ~n4480 ;
  assign y2335 = ~n4484 ;
  assign y2336 = n4487 ;
  assign y2337 = n1475 ;
  assign y2338 = ~n4489 ;
  assign y2339 = ~1'b0 ;
  assign y2340 = n4493 ;
  assign y2341 = n4497 ;
  assign y2342 = n4498 ;
  assign y2343 = ~n4499 ;
  assign y2344 = ~1'b0 ;
  assign y2345 = n4500 ;
  assign y2346 = ~n1656 ;
  assign y2347 = ~1'b0 ;
  assign y2348 = n4501 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = ~1'b0 ;
  assign y2351 = ~n2629 ;
  assign y2352 = n4503 ;
  assign y2353 = ~n4506 ;
  assign y2354 = n4507 ;
  assign y2355 = n4509 ;
  assign y2356 = ~1'b0 ;
  assign y2357 = ~1'b0 ;
  assign y2358 = ~1'b0 ;
  assign y2359 = n966 ;
  assign y2360 = n4510 ;
  assign y2361 = n4516 ;
  assign y2362 = ~n4520 ;
  assign y2363 = ~1'b0 ;
  assign y2364 = 1'b0 ;
  assign y2365 = ~n4526 ;
  assign y2366 = n4529 ;
  assign y2367 = ~1'b0 ;
  assign y2368 = ~1'b0 ;
  assign y2369 = n4537 ;
  assign y2370 = ~1'b0 ;
  assign y2371 = ~n4540 ;
  assign y2372 = n4543 ;
  assign y2373 = ~n4544 ;
  assign y2374 = ~n4546 ;
  assign y2375 = ~n4548 ;
  assign y2376 = ~1'b0 ;
  assign y2377 = n4549 ;
  assign y2378 = n4552 ;
  assign y2379 = n4555 ;
  assign y2380 = n4560 ;
  assign y2381 = n4562 ;
  assign y2382 = ~n3858 ;
  assign y2383 = ~n4565 ;
  assign y2384 = ~1'b0 ;
  assign y2385 = n4566 ;
  assign y2386 = ~n4568 ;
  assign y2387 = ~1'b0 ;
  assign y2388 = ~n4571 ;
  assign y2389 = ~n4573 ;
  assign y2390 = n4574 ;
  assign y2391 = n4577 ;
  assign y2392 = ~1'b0 ;
  assign y2393 = ~1'b0 ;
  assign y2394 = ~1'b0 ;
  assign y2395 = ~n4584 ;
  assign y2396 = ~n4586 ;
  assign y2397 = n4590 ;
  assign y2398 = ~1'b0 ;
  assign y2399 = n4592 ;
  assign y2400 = ~1'b0 ;
  assign y2401 = ~n4595 ;
  assign y2402 = n4596 ;
  assign y2403 = ~1'b0 ;
  assign y2404 = n4601 ;
  assign y2405 = n4562 ;
  assign y2406 = ~1'b0 ;
  assign y2407 = n4582 ;
  assign y2408 = ~n4605 ;
  assign y2409 = ~1'b0 ;
  assign y2410 = ~1'b0 ;
  assign y2411 = ~n4609 ;
  assign y2412 = ~1'b0 ;
  assign y2413 = n4616 ;
  assign y2414 = n4617 ;
  assign y2415 = n4618 ;
  assign y2416 = ~n4620 ;
  assign y2417 = ~n4622 ;
  assign y2418 = ~1'b0 ;
  assign y2419 = ~n4627 ;
  assign y2420 = ~n4637 ;
  assign y2421 = n4641 ;
  assign y2422 = ~n4650 ;
  assign y2423 = ~n4653 ;
  assign y2424 = n4657 ;
  assign y2425 = ~1'b0 ;
  assign y2426 = n651 ;
  assign y2427 = n3995 ;
  assign y2428 = ~n4658 ;
  assign y2429 = ~n4660 ;
  assign y2430 = ~n4661 ;
  assign y2431 = n4664 ;
  assign y2432 = n4668 ;
  assign y2433 = ~n4674 ;
  assign y2434 = ~1'b0 ;
  assign y2435 = ~n4676 ;
  assign y2436 = n4677 ;
  assign y2437 = n4680 ;
  assign y2438 = ~n3676 ;
  assign y2439 = ~1'b0 ;
  assign y2440 = ~1'b0 ;
  assign y2441 = ~1'b0 ;
  assign y2442 = ~1'b0 ;
  assign y2443 = ~1'b0 ;
  assign y2444 = ~n4685 ;
  assign y2445 = ~n4689 ;
  assign y2446 = ~n552 ;
  assign y2447 = 1'b0 ;
  assign y2448 = n4690 ;
  assign y2449 = ~n2495 ;
  assign y2450 = n4693 ;
  assign y2451 = ~n4695 ;
  assign y2452 = n4700 ;
  assign y2453 = x27 ;
  assign y2454 = n4701 ;
  assign y2455 = ~n4703 ;
  assign y2456 = ~1'b0 ;
  assign y2457 = ~1'b0 ;
  assign y2458 = ~1'b0 ;
  assign y2459 = ~n4705 ;
  assign y2460 = ~n4707 ;
  assign y2461 = ~n4708 ;
  assign y2462 = ~n2185 ;
  assign y2463 = ~1'b0 ;
  assign y2464 = n4711 ;
  assign y2465 = n4715 ;
  assign y2466 = ~1'b0 ;
  assign y2467 = ~1'b0 ;
  assign y2468 = 1'b0 ;
  assign y2469 = n4716 ;
  assign y2470 = ~1'b0 ;
  assign y2471 = ~1'b0 ;
  assign y2472 = ~1'b0 ;
  assign y2473 = n4719 ;
  assign y2474 = ~1'b0 ;
  assign y2475 = n1549 ;
  assign y2476 = ~n4724 ;
  assign y2477 = ~n4727 ;
  assign y2478 = n4729 ;
  assign y2479 = ~1'b0 ;
  assign y2480 = ~n4731 ;
  assign y2481 = ~1'b0 ;
  assign y2482 = ~1'b0 ;
  assign y2483 = ~1'b0 ;
  assign y2484 = ~n4733 ;
  assign y2485 = ~n2042 ;
  assign y2486 = n2959 ;
  assign y2487 = n4734 ;
  assign y2488 = n4737 ;
  assign y2489 = ~1'b0 ;
  assign y2490 = ~n4738 ;
  assign y2491 = n4741 ;
  assign y2492 = ~1'b0 ;
  assign y2493 = ~n4172 ;
  assign y2494 = n4745 ;
  assign y2495 = ~n4747 ;
  assign y2496 = n4749 ;
  assign y2497 = n4753 ;
  assign y2498 = ~n4757 ;
  assign y2499 = n1507 ;
  assign y2500 = ~1'b0 ;
  assign y2501 = n4760 ;
  assign y2502 = n4764 ;
  assign y2503 = ~n4766 ;
  assign y2504 = ~1'b0 ;
  assign y2505 = ~1'b0 ;
  assign y2506 = ~1'b0 ;
  assign y2507 = ~n3963 ;
  assign y2508 = ~n4771 ;
  assign y2509 = ~1'b0 ;
  assign y2510 = ~1'b0 ;
  assign y2511 = ~n4773 ;
  assign y2512 = ~n1814 ;
  assign y2513 = ~n4776 ;
  assign y2514 = n4779 ;
  assign y2515 = ~n4780 ;
  assign y2516 = ~1'b0 ;
  assign y2517 = n4782 ;
  assign y2518 = ~n4785 ;
  assign y2519 = n4788 ;
  assign y2520 = ~n1453 ;
  assign y2521 = n4789 ;
  assign y2522 = n4793 ;
  assign y2523 = n897 ;
  assign y2524 = ~n3175 ;
  assign y2525 = n4794 ;
  assign y2526 = ~n4796 ;
  assign y2527 = n4799 ;
  assign y2528 = ~n4804 ;
  assign y2529 = ~n4808 ;
  assign y2530 = ~n4812 ;
  assign y2531 = ~n4815 ;
  assign y2532 = n4816 ;
  assign y2533 = n4400 ;
  assign y2534 = n4819 ;
  assign y2535 = ~n4824 ;
  assign y2536 = ~1'b0 ;
  assign y2537 = ~n4828 ;
  assign y2538 = ~1'b0 ;
  assign y2539 = 1'b0 ;
  assign y2540 = n4831 ;
  assign y2541 = ~1'b0 ;
  assign y2542 = ~1'b0 ;
  assign y2543 = n4834 ;
  assign y2544 = n4835 ;
  assign y2545 = n4836 ;
  assign y2546 = ~1'b0 ;
  assign y2547 = n4838 ;
  assign y2548 = n3748 ;
  assign y2549 = n4841 ;
  assign y2550 = ~1'b0 ;
  assign y2551 = n4845 ;
  assign y2552 = ~n4846 ;
  assign y2553 = ~n4848 ;
  assign y2554 = ~n4849 ;
  assign y2555 = n4851 ;
  assign y2556 = ~n4853 ;
  assign y2557 = n4857 ;
  assign y2558 = n4860 ;
  assign y2559 = n4863 ;
  assign y2560 = n387 ;
  assign y2561 = ~n1181 ;
  assign y2562 = ~1'b0 ;
  assign y2563 = 1'b0 ;
  assign y2564 = ~1'b0 ;
  assign y2565 = ~n4866 ;
  assign y2566 = n4871 ;
  assign y2567 = ~n4734 ;
  assign y2568 = n4872 ;
  assign y2569 = ~n4873 ;
  assign y2570 = ~1'b0 ;
  assign y2571 = ~1'b0 ;
  assign y2572 = ~1'b0 ;
  assign y2573 = ~n4874 ;
  assign y2574 = n4875 ;
  assign y2575 = ~1'b0 ;
  assign y2576 = ~n4877 ;
  assign y2577 = ~n4879 ;
  assign y2578 = n4881 ;
  assign y2579 = ~n4884 ;
  assign y2580 = ~n985 ;
  assign y2581 = n4886 ;
  assign y2582 = n4889 ;
  assign y2583 = ~n4894 ;
  assign y2584 = n4901 ;
  assign y2585 = n4909 ;
  assign y2586 = ~n4910 ;
  assign y2587 = ~1'b0 ;
  assign y2588 = ~n4916 ;
  assign y2589 = ~n4917 ;
  assign y2590 = ~1'b0 ;
  assign y2591 = ~n4923 ;
  assign y2592 = ~n4927 ;
  assign y2593 = ~1'b0 ;
  assign y2594 = n3255 ;
  assign y2595 = ~1'b0 ;
  assign y2596 = ~1'b0 ;
  assign y2597 = ~1'b0 ;
  assign y2598 = n4256 ;
  assign y2599 = ~1'b0 ;
  assign y2600 = n4933 ;
  assign y2601 = n4944 ;
  assign y2602 = ~1'b0 ;
  assign y2603 = n4946 ;
  assign y2604 = n4948 ;
  assign y2605 = n4951 ;
  assign y2606 = ~1'b0 ;
  assign y2607 = n4955 ;
  assign y2608 = n4959 ;
  assign y2609 = ~n4960 ;
  assign y2610 = ~n4961 ;
  assign y2611 = ~n4962 ;
  assign y2612 = ~1'b0 ;
  assign y2613 = ~n4968 ;
  assign y2614 = ~1'b0 ;
  assign y2615 = ~1'b0 ;
  assign y2616 = n4970 ;
  assign y2617 = n4971 ;
  assign y2618 = ~n4974 ;
  assign y2619 = 1'b0 ;
  assign y2620 = ~1'b0 ;
  assign y2621 = ~1'b0 ;
  assign y2622 = 1'b0 ;
  assign y2623 = ~n4979 ;
  assign y2624 = ~n4980 ;
  assign y2625 = n2764 ;
  assign y2626 = ~1'b0 ;
  assign y2627 = ~n1405 ;
  assign y2628 = n4986 ;
  assign y2629 = ~1'b0 ;
  assign y2630 = n4989 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = n4991 ;
  assign y2633 = ~1'b0 ;
  assign y2634 = ~1'b0 ;
  assign y2635 = ~1'b0 ;
  assign y2636 = ~1'b0 ;
  assign y2637 = ~n4993 ;
  assign y2638 = n1444 ;
  assign y2639 = ~1'b0 ;
  assign y2640 = ~n5000 ;
  assign y2641 = ~n4385 ;
  assign y2642 = n5002 ;
  assign y2643 = n5006 ;
  assign y2644 = ~1'b0 ;
  assign y2645 = ~1'b0 ;
  assign y2646 = ~n5012 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = n5013 ;
  assign y2649 = n5014 ;
  assign y2650 = n5017 ;
  assign y2651 = ~n5018 ;
  assign y2652 = n5020 ;
  assign y2653 = n5021 ;
  assign y2654 = n5023 ;
  assign y2655 = ~n5024 ;
  assign y2656 = n5025 ;
  assign y2657 = ~1'b0 ;
  assign y2658 = n5026 ;
  assign y2659 = ~1'b0 ;
  assign y2660 = ~n5029 ;
  assign y2661 = n5036 ;
  assign y2662 = ~1'b0 ;
  assign y2663 = ~1'b0 ;
  assign y2664 = n3210 ;
  assign y2665 = n5042 ;
  assign y2666 = ~n5043 ;
  assign y2667 = ~1'b0 ;
  assign y2668 = n979 ;
  assign y2669 = ~n4300 ;
  assign y2670 = ~1'b0 ;
  assign y2671 = n5047 ;
  assign y2672 = ~1'b0 ;
  assign y2673 = ~n5052 ;
  assign y2674 = ~n3181 ;
  assign y2675 = n5054 ;
  assign y2676 = ~n5062 ;
  assign y2677 = n5064 ;
  assign y2678 = n5066 ;
  assign y2679 = n5067 ;
  assign y2680 = n5068 ;
  assign y2681 = ~1'b0 ;
  assign y2682 = ~n5069 ;
  assign y2683 = ~n3184 ;
  assign y2684 = n5070 ;
  assign y2685 = ~1'b0 ;
  assign y2686 = n1920 ;
  assign y2687 = ~n5071 ;
  assign y2688 = ~1'b0 ;
  assign y2689 = ~1'b0 ;
  assign y2690 = ~1'b0 ;
  assign y2691 = ~1'b0 ;
  assign y2692 = ~n5072 ;
  assign y2693 = n5074 ;
  assign y2694 = ~1'b0 ;
  assign y2695 = n5081 ;
  assign y2696 = n5082 ;
  assign y2697 = x174 ;
  assign y2698 = ~n5085 ;
  assign y2699 = n5088 ;
  assign y2700 = n5089 ;
  assign y2701 = ~1'b0 ;
  assign y2702 = n5094 ;
  assign y2703 = ~1'b0 ;
  assign y2704 = n5099 ;
  assign y2705 = n4857 ;
  assign y2706 = ~n5103 ;
  assign y2707 = n5107 ;
  assign y2708 = ~1'b0 ;
  assign y2709 = ~1'b0 ;
  assign y2710 = ~1'b0 ;
  assign y2711 = ~1'b0 ;
  assign y2712 = ~n5108 ;
  assign y2713 = n5110 ;
  assign y2714 = ~n5111 ;
  assign y2715 = n5112 ;
  assign y2716 = ~n3304 ;
  assign y2717 = ~n5114 ;
  assign y2718 = ~n5116 ;
  assign y2719 = ~n5118 ;
  assign y2720 = ~n5119 ;
  assign y2721 = n5120 ;
  assign y2722 = n5122 ;
  assign y2723 = ~1'b0 ;
  assign y2724 = n5125 ;
  assign y2725 = ~n5126 ;
  assign y2726 = ~n5128 ;
  assign y2727 = ~n3152 ;
  assign y2728 = ~n5129 ;
  assign y2729 = ~n5135 ;
  assign y2730 = ~1'b0 ;
  assign y2731 = ~n5136 ;
  assign y2732 = ~1'b0 ;
  assign y2733 = ~1'b0 ;
  assign y2734 = n5137 ;
  assign y2735 = ~1'b0 ;
  assign y2736 = n5139 ;
  assign y2737 = ~1'b0 ;
  assign y2738 = ~1'b0 ;
  assign y2739 = ~1'b0 ;
  assign y2740 = ~n5143 ;
  assign y2741 = ~n5144 ;
  assign y2742 = ~1'b0 ;
  assign y2743 = ~n5145 ;
  assign y2744 = ~n5148 ;
  assign y2745 = ~n5150 ;
  assign y2746 = ~n5152 ;
  assign y2747 = ~1'b0 ;
  assign y2748 = ~n5155 ;
  assign y2749 = ~n5157 ;
  assign y2750 = ~1'b0 ;
  assign y2751 = n5160 ;
  assign y2752 = 1'b0 ;
  assign y2753 = ~1'b0 ;
  assign y2754 = n5163 ;
  assign y2755 = ~n5166 ;
  assign y2756 = ~n5169 ;
  assign y2757 = ~n5170 ;
  assign y2758 = n5173 ;
  assign y2759 = n5175 ;
  assign y2760 = ~n5176 ;
  assign y2761 = ~n930 ;
  assign y2762 = n5181 ;
  assign y2763 = ~1'b0 ;
  assign y2764 = n5185 ;
  assign y2765 = n5188 ;
  assign y2766 = ~n5189 ;
  assign y2767 = ~n2293 ;
  assign y2768 = ~1'b0 ;
  assign y2769 = n5190 ;
  assign y2770 = ~n5191 ;
  assign y2771 = 1'b0 ;
  assign y2772 = n5192 ;
  assign y2773 = n5195 ;
  assign y2774 = n5196 ;
  assign y2775 = n5198 ;
  assign y2776 = ~n5200 ;
  assign y2777 = n5201 ;
  assign y2778 = ~n628 ;
  assign y2779 = ~1'b0 ;
  assign y2780 = ~1'b0 ;
  assign y2781 = ~n5207 ;
  assign y2782 = n5209 ;
  assign y2783 = ~1'b0 ;
  assign y2784 = ~n5213 ;
  assign y2785 = n5218 ;
  assign y2786 = 1'b0 ;
  assign y2787 = ~n5223 ;
  assign y2788 = ~n5227 ;
  assign y2789 = n5229 ;
  assign y2790 = ~1'b0 ;
  assign y2791 = ~1'b0 ;
  assign y2792 = ~n5232 ;
  assign y2793 = ~n5238 ;
  assign y2794 = n5242 ;
  assign y2795 = ~n5244 ;
  assign y2796 = ~n5246 ;
  assign y2797 = ~1'b0 ;
  assign y2798 = n4608 ;
  assign y2799 = ~1'b0 ;
  assign y2800 = n5252 ;
  assign y2801 = ~n5255 ;
  assign y2802 = ~n2187 ;
  assign y2803 = n5257 ;
  assign y2804 = ~n5262 ;
  assign y2805 = ~1'b0 ;
  assign y2806 = ~1'b0 ;
  assign y2807 = ~n5263 ;
  assign y2808 = n5265 ;
  assign y2809 = ~n5272 ;
  assign y2810 = ~n5277 ;
  assign y2811 = ~n5280 ;
  assign y2812 = ~1'b0 ;
  assign y2813 = ~1'b0 ;
  assign y2814 = n5284 ;
  assign y2815 = n5285 ;
  assign y2816 = ~n5288 ;
  assign y2817 = ~n5290 ;
  assign y2818 = ~1'b0 ;
  assign y2819 = n5292 ;
  assign y2820 = n5298 ;
  assign y2821 = ~n5300 ;
  assign y2822 = n5302 ;
  assign y2823 = ~n5303 ;
  assign y2824 = ~n5304 ;
  assign y2825 = ~n5305 ;
  assign y2826 = ~n5311 ;
  assign y2827 = ~1'b0 ;
  assign y2828 = ~1'b0 ;
  assign y2829 = ~n5312 ;
  assign y2830 = ~n5317 ;
  assign y2831 = ~n5325 ;
  assign y2832 = ~n5328 ;
  assign y2833 = n5330 ;
  assign y2834 = ~n5331 ;
  assign y2835 = n5332 ;
  assign y2836 = ~1'b0 ;
  assign y2837 = ~n3750 ;
  assign y2838 = ~n5336 ;
  assign y2839 = ~1'b0 ;
  assign y2840 = ~1'b0 ;
  assign y2841 = ~1'b0 ;
  assign y2842 = 1'b0 ;
  assign y2843 = ~1'b0 ;
  assign y2844 = ~1'b0 ;
  assign y2845 = ~n5337 ;
  assign y2846 = ~n5338 ;
  assign y2847 = ~1'b0 ;
  assign y2848 = 1'b0 ;
  assign y2849 = n5341 ;
  assign y2850 = 1'b0 ;
  assign y2851 = n3807 ;
  assign y2852 = n4816 ;
  assign y2853 = ~n1126 ;
  assign y2854 = n5344 ;
  assign y2855 = ~n5347 ;
  assign y2856 = n5348 ;
  assign y2857 = ~1'b0 ;
  assign y2858 = ~1'b0 ;
  assign y2859 = n5350 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = ~n5353 ;
  assign y2862 = n5354 ;
  assign y2863 = ~n5357 ;
  assign y2864 = ~1'b0 ;
  assign y2865 = ~1'b0 ;
  assign y2866 = ~1'b0 ;
  assign y2867 = n5358 ;
  assign y2868 = n5364 ;
  assign y2869 = ~1'b0 ;
  assign y2870 = ~n5222 ;
  assign y2871 = n5366 ;
  assign y2872 = n5369 ;
  assign y2873 = n5372 ;
  assign y2874 = ~n5373 ;
  assign y2875 = n5379 ;
  assign y2876 = n5381 ;
  assign y2877 = ~1'b0 ;
  assign y2878 = ~1'b0 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~n5384 ;
  assign y2881 = x228 ;
  assign y2882 = n5386 ;
  assign y2883 = ~n5387 ;
  assign y2884 = n5392 ;
  assign y2885 = ~n5393 ;
  assign y2886 = ~n5396 ;
  assign y2887 = ~1'b0 ;
  assign y2888 = ~n5399 ;
  assign y2889 = ~1'b0 ;
  assign y2890 = ~n5400 ;
  assign y2891 = n5405 ;
  assign y2892 = ~n5408 ;
  assign y2893 = n3443 ;
  assign y2894 = ~n5155 ;
  assign y2895 = ~n5412 ;
  assign y2896 = n5413 ;
  assign y2897 = ~1'b0 ;
  assign y2898 = ~n5415 ;
  assign y2899 = ~n5418 ;
  assign y2900 = ~n5419 ;
  assign y2901 = n5420 ;
  assign y2902 = ~n5422 ;
  assign y2903 = ~1'b0 ;
  assign y2904 = ~1'b0 ;
  assign y2905 = n5423 ;
  assign y2906 = ~n5426 ;
  assign y2907 = n5427 ;
  assign y2908 = ~n5429 ;
  assign y2909 = ~n5431 ;
  assign y2910 = ~n5433 ;
  assign y2911 = ~n5439 ;
  assign y2912 = ~n5443 ;
  assign y2913 = ~1'b0 ;
  assign y2914 = n5447 ;
  assign y2915 = ~n5448 ;
  assign y2916 = ~1'b0 ;
  assign y2917 = ~n5456 ;
  assign y2918 = ~1'b0 ;
  assign y2919 = n5457 ;
  assign y2920 = n5458 ;
  assign y2921 = ~n5460 ;
  assign y2922 = n3879 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = ~n5464 ;
  assign y2925 = ~1'b0 ;
  assign y2926 = ~n5472 ;
  assign y2927 = ~1'b0 ;
  assign y2928 = n5457 ;
  assign y2929 = n5475 ;
  assign y2930 = ~n5476 ;
  assign y2931 = n1405 ;
  assign y2932 = ~n5479 ;
  assign y2933 = ~n5484 ;
  assign y2934 = n5487 ;
  assign y2935 = ~n5505 ;
  assign y2936 = ~1'b0 ;
  assign y2937 = ~1'b0 ;
  assign y2938 = n5507 ;
  assign y2939 = n5508 ;
  assign y2940 = ~n5510 ;
  assign y2941 = ~n4367 ;
  assign y2942 = n5512 ;
  assign y2943 = ~n5514 ;
  assign y2944 = ~1'b0 ;
  assign y2945 = ~1'b0 ;
  assign y2946 = ~n5516 ;
  assign y2947 = ~n5521 ;
  assign y2948 = ~1'b0 ;
  assign y2949 = n5523 ;
  assign y2950 = n5529 ;
  assign y2951 = ~x86 ;
  assign y2952 = n5531 ;
  assign y2953 = ~1'b0 ;
  assign y2954 = ~n5534 ;
  assign y2955 = ~1'b0 ;
  assign y2956 = n5549 ;
  assign y2957 = 1'b0 ;
  assign y2958 = ~1'b0 ;
  assign y2959 = n5551 ;
  assign y2960 = ~n5552 ;
  assign y2961 = ~1'b0 ;
  assign y2962 = ~n5553 ;
  assign y2963 = ~1'b0 ;
  assign y2964 = ~1'b0 ;
  assign y2965 = ~n3776 ;
  assign y2966 = ~1'b0 ;
  assign y2967 = n5555 ;
  assign y2968 = ~1'b0 ;
  assign y2969 = n5557 ;
  assign y2970 = ~n269 ;
  assign y2971 = n5559 ;
  assign y2972 = ~n5560 ;
  assign y2973 = ~1'b0 ;
  assign y2974 = ~1'b0 ;
  assign y2975 = ~1'b0 ;
  assign y2976 = ~1'b0 ;
  assign y2977 = ~1'b0 ;
  assign y2978 = ~n5563 ;
  assign y2979 = n5564 ;
  assign y2980 = ~n5567 ;
  assign y2981 = ~n5571 ;
  assign y2982 = ~n5578 ;
  assign y2983 = n5579 ;
  assign y2984 = n5580 ;
  assign y2985 = ~n5583 ;
  assign y2986 = n5586 ;
  assign y2987 = n5587 ;
  assign y2988 = ~1'b0 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = n5590 ;
  assign y2991 = ~1'b0 ;
  assign y2992 = ~1'b0 ;
  assign y2993 = n5592 ;
  assign y2994 = ~n5595 ;
  assign y2995 = ~n5600 ;
  assign y2996 = ~1'b0 ;
  assign y2997 = n5601 ;
  assign y2998 = ~n5603 ;
  assign y2999 = n5604 ;
  assign y3000 = ~n5606 ;
  assign y3001 = ~n5607 ;
  assign y3002 = ~n5608 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = ~n5612 ;
  assign y3005 = ~1'b0 ;
  assign y3006 = n5618 ;
  assign y3007 = ~1'b0 ;
  assign y3008 = n5619 ;
  assign y3009 = ~n5626 ;
  assign y3010 = ~1'b0 ;
  assign y3011 = ~n5627 ;
  assign y3012 = ~n921 ;
  assign y3013 = ~n5631 ;
  assign y3014 = n5633 ;
  assign y3015 = ~n5634 ;
  assign y3016 = ~1'b0 ;
  assign y3017 = ~1'b0 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = n5639 ;
  assign y3020 = n5398 ;
  assign y3021 = n5643 ;
  assign y3022 = ~1'b0 ;
  assign y3023 = ~1'b0 ;
  assign y3024 = n2035 ;
  assign y3025 = ~1'b0 ;
  assign y3026 = ~1'b0 ;
  assign y3027 = ~n1689 ;
  assign y3028 = ~n5650 ;
  assign y3029 = n5651 ;
  assign y3030 = ~n5654 ;
  assign y3031 = ~n5656 ;
  assign y3032 = 1'b0 ;
  assign y3033 = n5261 ;
  assign y3034 = ~n5658 ;
  assign y3035 = n5659 ;
  assign y3036 = n5660 ;
  assign y3037 = n5662 ;
  assign y3038 = ~n5667 ;
  assign y3039 = ~1'b0 ;
  assign y3040 = ~1'b0 ;
  assign y3041 = n5669 ;
  assign y3042 = n3212 ;
  assign y3043 = n5671 ;
  assign y3044 = ~1'b0 ;
  assign y3045 = n1661 ;
  assign y3046 = n5675 ;
  assign y3047 = ~1'b0 ;
  assign y3048 = ~n5676 ;
  assign y3049 = ~n5682 ;
  assign y3050 = n5688 ;
  assign y3051 = ~1'b0 ;
  assign y3052 = ~n5691 ;
  assign y3053 = n5698 ;
  assign y3054 = ~n5700 ;
  assign y3055 = ~n5702 ;
  assign y3056 = n5706 ;
  assign y3057 = ~n5711 ;
  assign y3058 = ~1'b0 ;
  assign y3059 = n5712 ;
  assign y3060 = n5715 ;
  assign y3061 = ~1'b0 ;
  assign y3062 = n5718 ;
  assign y3063 = ~n5719 ;
  assign y3064 = n5726 ;
  assign y3065 = ~n5728 ;
  assign y3066 = ~n2469 ;
  assign y3067 = ~n5729 ;
  assign y3068 = n5730 ;
  assign y3069 = ~1'b0 ;
  assign y3070 = ~1'b0 ;
  assign y3071 = ~1'b0 ;
  assign y3072 = n5737 ;
  assign y3073 = n5740 ;
  assign y3074 = ~1'b0 ;
  assign y3075 = ~1'b0 ;
  assign y3076 = 1'b0 ;
  assign y3077 = n5742 ;
  assign y3078 = ~n4298 ;
  assign y3079 = ~n5750 ;
  assign y3080 = ~1'b0 ;
  assign y3081 = n5754 ;
  assign y3082 = ~n5755 ;
  assign y3083 = n5758 ;
  assign y3084 = ~1'b0 ;
  assign y3085 = ~n5759 ;
  assign y3086 = ~1'b0 ;
  assign y3087 = ~1'b0 ;
  assign y3088 = ~n788 ;
  assign y3089 = ~n5761 ;
  assign y3090 = n5762 ;
  assign y3091 = ~1'b0 ;
  assign y3092 = ~n5767 ;
  assign y3093 = ~n2910 ;
  assign y3094 = ~1'b0 ;
  assign y3095 = ~n5770 ;
  assign y3096 = ~n5771 ;
  assign y3097 = ~1'b0 ;
  assign y3098 = ~1'b0 ;
  assign y3099 = ~1'b0 ;
  assign y3100 = ~n5775 ;
  assign y3101 = ~n5779 ;
  assign y3102 = ~n5783 ;
  assign y3103 = n5784 ;
  assign y3104 = ~n5790 ;
  assign y3105 = ~n5792 ;
  assign y3106 = ~1'b0 ;
  assign y3107 = ~n5795 ;
  assign y3108 = ~n5796 ;
  assign y3109 = ~n5798 ;
  assign y3110 = n5802 ;
  assign y3111 = ~1'b0 ;
  assign y3112 = ~1'b0 ;
  assign y3113 = ~1'b0 ;
  assign y3114 = ~1'b0 ;
  assign y3115 = n5806 ;
  assign y3116 = n5808 ;
  assign y3117 = n5809 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = ~n1751 ;
  assign y3120 = n5812 ;
  assign y3121 = x161 ;
  assign y3122 = ~1'b0 ;
  assign y3123 = ~n5818 ;
  assign y3124 = ~1'b0 ;
  assign y3125 = ~n2230 ;
  assign y3126 = ~1'b0 ;
  assign y3127 = n5828 ;
  assign y3128 = n5830 ;
  assign y3129 = n5833 ;
  assign y3130 = n5842 ;
  assign y3131 = ~n4579 ;
  assign y3132 = ~n5843 ;
  assign y3133 = 1'b0 ;
  assign y3134 = n5844 ;
  assign y3135 = n5846 ;
  assign y3136 = n5848 ;
  assign y3137 = ~1'b0 ;
  assign y3138 = ~n5851 ;
  assign y3139 = ~1'b0 ;
  assign y3140 = n5852 ;
  assign y3141 = ~1'b0 ;
  assign y3142 = ~n5857 ;
  assign y3143 = n5859 ;
  assign y3144 = ~n5860 ;
  assign y3145 = ~n5861 ;
  assign y3146 = ~n5864 ;
  assign y3147 = ~n5870 ;
  assign y3148 = ~n3153 ;
  assign y3149 = n5872 ;
  assign y3150 = ~n5874 ;
  assign y3151 = ~n5875 ;
  assign y3152 = ~1'b0 ;
  assign y3153 = ~1'b0 ;
  assign y3154 = ~1'b0 ;
  assign y3155 = ~1'b0 ;
  assign y3156 = n5877 ;
  assign y3157 = n5885 ;
  assign y3158 = ~n1286 ;
  assign y3159 = ~n5887 ;
  assign y3160 = ~n5890 ;
  assign y3161 = ~n5891 ;
  assign y3162 = n5892 ;
  assign y3163 = ~n5895 ;
  assign y3164 = ~1'b0 ;
  assign y3165 = n5897 ;
  assign y3166 = n5898 ;
  assign y3167 = ~1'b0 ;
  assign y3168 = ~n5719 ;
  assign y3169 = ~n5904 ;
  assign y3170 = ~n5905 ;
  assign y3171 = ~1'b0 ;
  assign y3172 = ~1'b0 ;
  assign y3173 = n5908 ;
  assign y3174 = n5914 ;
  assign y3175 = ~n5915 ;
  assign y3176 = ~1'b0 ;
  assign y3177 = ~1'b0 ;
  assign y3178 = 1'b0 ;
  assign y3179 = ~1'b0 ;
  assign y3180 = ~n5918 ;
  assign y3181 = ~n5922 ;
  assign y3182 = n5925 ;
  assign y3183 = ~n5926 ;
  assign y3184 = ~n5927 ;
  assign y3185 = n5931 ;
  assign y3186 = n5935 ;
  assign y3187 = n5940 ;
  assign y3188 = ~1'b0 ;
  assign y3189 = ~n5942 ;
  assign y3190 = ~1'b0 ;
  assign y3191 = ~n5943 ;
  assign y3192 = ~1'b0 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = ~1'b0 ;
  assign y3195 = ~1'b0 ;
  assign y3196 = ~1'b0 ;
  assign y3197 = ~1'b0 ;
  assign y3198 = ~n5946 ;
  assign y3199 = n5948 ;
  assign y3200 = ~1'b0 ;
  assign y3201 = ~1'b0 ;
  assign y3202 = n5953 ;
  assign y3203 = ~1'b0 ;
  assign y3204 = ~n5956 ;
  assign y3205 = n5957 ;
  assign y3206 = ~n5958 ;
  assign y3207 = ~n5959 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = ~n5963 ;
  assign y3210 = n5970 ;
  assign y3211 = n5972 ;
  assign y3212 = x12 ;
  assign y3213 = ~1'b0 ;
  assign y3214 = n5973 ;
  assign y3215 = ~1'b0 ;
  assign y3216 = n5974 ;
  assign y3217 = ~n5976 ;
  assign y3218 = ~n5977 ;
  assign y3219 = ~n5983 ;
  assign y3220 = ~n5988 ;
  assign y3221 = ~1'b0 ;
  assign y3222 = n5989 ;
  assign y3223 = ~1'b0 ;
  assign y3224 = n5993 ;
  assign y3225 = n5996 ;
  assign y3226 = ~n6003 ;
  assign y3227 = ~n6005 ;
  assign y3228 = ~n6008 ;
  assign y3229 = ~1'b0 ;
  assign y3230 = ~1'b0 ;
  assign y3231 = n6009 ;
  assign y3232 = ~1'b0 ;
  assign y3233 = ~1'b0 ;
  assign y3234 = n6017 ;
  assign y3235 = n6018 ;
  assign y3236 = n6022 ;
  assign y3237 = ~1'b0 ;
  assign y3238 = ~n6025 ;
  assign y3239 = n6026 ;
  assign y3240 = ~1'b0 ;
  assign y3241 = ~1'b0 ;
  assign y3242 = ~1'b0 ;
  assign y3243 = ~1'b0 ;
  assign y3244 = ~n6031 ;
  assign y3245 = ~n6033 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = ~1'b0 ;
  assign y3248 = n6038 ;
  assign y3249 = n633 ;
  assign y3250 = ~n6043 ;
  assign y3251 = ~1'b0 ;
  assign y3252 = n6049 ;
  assign y3253 = ~n6050 ;
  assign y3254 = ~1'b0 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = n6051 ;
  assign y3257 = n6052 ;
  assign y3258 = 1'b0 ;
  assign y3259 = n6053 ;
  assign y3260 = n6054 ;
  assign y3261 = ~1'b0 ;
  assign y3262 = ~1'b0 ;
  assign y3263 = ~1'b0 ;
  assign y3264 = n6055 ;
  assign y3265 = n6058 ;
  assign y3266 = ~1'b0 ;
  assign y3267 = n6064 ;
  assign y3268 = ~n6067 ;
  assign y3269 = n6070 ;
  assign y3270 = ~n6073 ;
  assign y3271 = ~n6075 ;
  assign y3272 = ~n6078 ;
  assign y3273 = ~n6080 ;
  assign y3274 = n6083 ;
  assign y3275 = ~n6087 ;
  assign y3276 = ~1'b0 ;
  assign y3277 = n6091 ;
  assign y3278 = n6094 ;
  assign y3279 = ~1'b0 ;
  assign y3280 = n6095 ;
  assign y3281 = 1'b0 ;
  assign y3282 = ~1'b0 ;
  assign y3283 = n6096 ;
  assign y3284 = ~1'b0 ;
  assign y3285 = ~1'b0 ;
  assign y3286 = n6097 ;
  assign y3287 = ~1'b0 ;
  assign y3288 = ~n4664 ;
  assign y3289 = ~1'b0 ;
  assign y3290 = ~1'b0 ;
  assign y3291 = 1'b0 ;
  assign y3292 = ~n6098 ;
  assign y3293 = ~1'b0 ;
  assign y3294 = ~1'b0 ;
  assign y3295 = n6100 ;
  assign y3296 = ~1'b0 ;
  assign y3297 = ~n6102 ;
  assign y3298 = x75 ;
  assign y3299 = ~1'b0 ;
  assign y3300 = ~n6104 ;
  assign y3301 = ~1'b0 ;
  assign y3302 = n6110 ;
  assign y3303 = ~1'b0 ;
  assign y3304 = n6114 ;
  assign y3305 = ~n6116 ;
  assign y3306 = ~n6117 ;
  assign y3307 = ~n6118 ;
  assign y3308 = ~1'b0 ;
  assign y3309 = ~n6119 ;
  assign y3310 = ~n6125 ;
  assign y3311 = ~1'b0 ;
  assign y3312 = ~n6131 ;
  assign y3313 = ~n6134 ;
  assign y3314 = ~n6136 ;
  assign y3315 = ~1'b0 ;
  assign y3316 = n6140 ;
  assign y3317 = n1459 ;
  assign y3318 = ~n6143 ;
  assign y3319 = ~n6146 ;
  assign y3320 = n6151 ;
  assign y3321 = ~n6154 ;
  assign y3322 = ~n6156 ;
  assign y3323 = ~n6158 ;
  assign y3324 = ~1'b0 ;
  assign y3325 = ~n6161 ;
  assign y3326 = n6170 ;
  assign y3327 = n6172 ;
  assign y3328 = ~n6179 ;
  assign y3329 = ~n6180 ;
  assign y3330 = 1'b0 ;
  assign y3331 = n6186 ;
  assign y3332 = ~n6187 ;
  assign y3333 = n6190 ;
  assign y3334 = ~n6191 ;
  assign y3335 = ~n6193 ;
  assign y3336 = ~n821 ;
  assign y3337 = ~1'b0 ;
  assign y3338 = ~n6195 ;
  assign y3339 = ~n6196 ;
  assign y3340 = ~n6198 ;
  assign y3341 = n6203 ;
  assign y3342 = ~n6210 ;
  assign y3343 = ~n6213 ;
  assign y3344 = ~1'b0 ;
  assign y3345 = n6217 ;
  assign y3346 = ~1'b0 ;
  assign y3347 = ~n6222 ;
  assign y3348 = ~1'b0 ;
  assign y3349 = ~n6229 ;
  assign y3350 = 1'b0 ;
  assign y3351 = ~1'b0 ;
  assign y3352 = ~n6239 ;
  assign y3353 = ~n6245 ;
  assign y3354 = ~1'b0 ;
  assign y3355 = ~1'b0 ;
  assign y3356 = ~1'b0 ;
  assign y3357 = ~1'b0 ;
  assign y3358 = n6250 ;
  assign y3359 = ~1'b0 ;
  assign y3360 = ~n6252 ;
  assign y3361 = n6253 ;
  assign y3362 = ~n6254 ;
  assign y3363 = n6256 ;
  assign y3364 = ~n6258 ;
  assign y3365 = ~n6259 ;
  assign y3366 = ~n6261 ;
  assign y3367 = ~n6263 ;
  assign y3368 = n6264 ;
  assign y3369 = ~1'b0 ;
  assign y3370 = n6266 ;
  assign y3371 = n4671 ;
  assign y3372 = n6267 ;
  assign y3373 = n6268 ;
  assign y3374 = ~1'b0 ;
  assign y3375 = n6270 ;
  assign y3376 = n6273 ;
  assign y3377 = ~n6274 ;
  assign y3378 = ~n6276 ;
  assign y3379 = ~1'b0 ;
  assign y3380 = ~1'b0 ;
  assign y3381 = ~1'b0 ;
  assign y3382 = ~1'b0 ;
  assign y3383 = ~1'b0 ;
  assign y3384 = ~n6281 ;
  assign y3385 = ~1'b0 ;
  assign y3386 = ~1'b0 ;
  assign y3387 = ~n6286 ;
  assign y3388 = ~1'b0 ;
  assign y3389 = ~1'b0 ;
  assign y3390 = ~1'b0 ;
  assign y3391 = ~1'b0 ;
  assign y3392 = ~n6292 ;
  assign y3393 = ~n6296 ;
  assign y3394 = ~n6297 ;
  assign y3395 = ~n6300 ;
  assign y3396 = ~1'b0 ;
  assign y3397 = ~1'b0 ;
  assign y3398 = n6302 ;
  assign y3399 = n6303 ;
  assign y3400 = n6305 ;
  assign y3401 = ~1'b0 ;
  assign y3402 = ~n6308 ;
  assign y3403 = n5809 ;
  assign y3404 = ~n6312 ;
  assign y3405 = ~1'b0 ;
  assign y3406 = ~n6315 ;
  assign y3407 = n6322 ;
  assign y3408 = ~1'b0 ;
  assign y3409 = n6324 ;
  assign y3410 = n6330 ;
  assign y3411 = ~n6331 ;
  assign y3412 = ~n6333 ;
  assign y3413 = ~n6335 ;
  assign y3414 = ~n6341 ;
  assign y3415 = n1285 ;
  assign y3416 = ~1'b0 ;
  assign y3417 = n6343 ;
  assign y3418 = n6344 ;
  assign y3419 = ~1'b0 ;
  assign y3420 = ~n6348 ;
  assign y3421 = ~1'b0 ;
  assign y3422 = ~1'b0 ;
  assign y3423 = ~1'b0 ;
  assign y3424 = ~n956 ;
  assign y3425 = n6353 ;
  assign y3426 = n6359 ;
  assign y3427 = ~n6362 ;
  assign y3428 = ~n6363 ;
  assign y3429 = n3501 ;
  assign y3430 = ~n6365 ;
  assign y3431 = ~1'b0 ;
  assign y3432 = n6366 ;
  assign y3433 = ~1'b0 ;
  assign y3434 = ~n1704 ;
  assign y3435 = ~1'b0 ;
  assign y3436 = n6368 ;
  assign y3437 = n6371 ;
  assign y3438 = ~1'b0 ;
  assign y3439 = n6378 ;
  assign y3440 = n6379 ;
  assign y3441 = n6382 ;
  assign y3442 = 1'b0 ;
  assign y3443 = ~1'b0 ;
  assign y3444 = n6383 ;
  assign y3445 = ~1'b0 ;
  assign y3446 = n1488 ;
  assign y3447 = n6387 ;
  assign y3448 = ~1'b0 ;
  assign y3449 = ~n6391 ;
  assign y3450 = ~1'b0 ;
  assign y3451 = ~n4549 ;
  assign y3452 = ~n6392 ;
  assign y3453 = ~1'b0 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = ~n6396 ;
  assign y3456 = n6398 ;
  assign y3457 = n3473 ;
  assign y3458 = n6399 ;
  assign y3459 = n6401 ;
  assign y3460 = n6402 ;
  assign y3461 = n6405 ;
  assign y3462 = 1'b0 ;
  assign y3463 = ~n6408 ;
  assign y3464 = ~n6410 ;
  assign y3465 = ~1'b0 ;
  assign y3466 = n6412 ;
  assign y3467 = ~n6418 ;
  assign y3468 = ~1'b0 ;
  assign y3469 = ~1'b0 ;
  assign y3470 = ~1'b0 ;
  assign y3471 = n6419 ;
  assign y3472 = ~n6420 ;
  assign y3473 = ~n6421 ;
  assign y3474 = n6428 ;
  assign y3475 = ~1'b0 ;
  assign y3476 = ~1'b0 ;
  assign y3477 = ~1'b0 ;
  assign y3478 = ~1'b0 ;
  assign y3479 = ~1'b0 ;
  assign y3480 = ~1'b0 ;
  assign y3481 = ~n6430 ;
  assign y3482 = n6431 ;
  assign y3483 = ~n6434 ;
  assign y3484 = n6435 ;
  assign y3485 = x65 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = ~n6439 ;
  assign y3488 = n6446 ;
  assign y3489 = ~n6451 ;
  assign y3490 = ~n6453 ;
  assign y3491 = ~n6460 ;
  assign y3492 = n6461 ;
  assign y3493 = n6468 ;
  assign y3494 = ~n6469 ;
  assign y3495 = 1'b0 ;
  assign y3496 = ~n6471 ;
  assign y3497 = ~1'b0 ;
  assign y3498 = ~1'b0 ;
  assign y3499 = ~1'b0 ;
  assign y3500 = n5891 ;
  assign y3501 = ~1'b0 ;
  assign y3502 = ~1'b0 ;
  assign y3503 = ~1'b0 ;
  assign y3504 = ~n6475 ;
  assign y3505 = ~1'b0 ;
  assign y3506 = n6477 ;
  assign y3507 = ~n6479 ;
  assign y3508 = n6482 ;
  assign y3509 = ~n6484 ;
  assign y3510 = ~1'b0 ;
  assign y3511 = ~n1551 ;
  assign y3512 = ~n6487 ;
  assign y3513 = ~n6491 ;
  assign y3514 = n6493 ;
  assign y3515 = n6494 ;
  assign y3516 = ~n6498 ;
  assign y3517 = ~n6499 ;
  assign y3518 = ~n6502 ;
  assign y3519 = n6505 ;
  assign y3520 = ~n6507 ;
  assign y3521 = ~n6509 ;
  assign y3522 = n6511 ;
  assign y3523 = ~n1644 ;
  assign y3524 = ~n6515 ;
  assign y3525 = n6516 ;
  assign y3526 = n6517 ;
  assign y3527 = 1'b0 ;
  assign y3528 = ~n6519 ;
  assign y3529 = ~1'b0 ;
  assign y3530 = ~1'b0 ;
  assign y3531 = n6522 ;
  assign y3532 = ~n6525 ;
  assign y3533 = ~n6049 ;
  assign y3534 = ~1'b0 ;
  assign y3535 = n6527 ;
  assign y3536 = n6528 ;
  assign y3537 = ~1'b0 ;
  assign y3538 = n6532 ;
  assign y3539 = ~n6534 ;
  assign y3540 = ~1'b0 ;
  assign y3541 = ~1'b0 ;
  assign y3542 = ~n6540 ;
  assign y3543 = n6542 ;
  assign y3544 = n6546 ;
  assign y3545 = ~1'b0 ;
  assign y3546 = ~n6550 ;
  assign y3547 = n6551 ;
  assign y3548 = ~n6553 ;
  assign y3549 = n6555 ;
  assign y3550 = ~n6556 ;
  assign y3551 = ~n6558 ;
  assign y3552 = ~n6560 ;
  assign y3553 = n6562 ;
  assign y3554 = x106 ;
  assign y3555 = ~n6564 ;
  assign y3556 = ~n6572 ;
  assign y3557 = ~1'b0 ;
  assign y3558 = ~1'b0 ;
  assign y3559 = n6576 ;
  assign y3560 = ~1'b0 ;
  assign y3561 = ~1'b0 ;
  assign y3562 = n6578 ;
  assign y3563 = ~1'b0 ;
  assign y3564 = n6583 ;
  assign y3565 = ~n6585 ;
  assign y3566 = ~n6599 ;
  assign y3567 = ~n605 ;
  assign y3568 = ~n6601 ;
  assign y3569 = n6602 ;
  assign y3570 = 1'b0 ;
  assign y3571 = n4395 ;
  assign y3572 = ~1'b0 ;
  assign y3573 = n6603 ;
  assign y3574 = ~1'b0 ;
  assign y3575 = n6614 ;
  assign y3576 = n6619 ;
  assign y3577 = ~n6623 ;
  assign y3578 = n6629 ;
  assign y3579 = ~n6630 ;
  assign y3580 = ~1'b0 ;
  assign y3581 = n6636 ;
  assign y3582 = ~1'b0 ;
  assign y3583 = n6642 ;
  assign y3584 = ~1'b0 ;
  assign y3585 = n6644 ;
  assign y3586 = n6649 ;
  assign y3587 = ~1'b0 ;
  assign y3588 = 1'b0 ;
  assign y3589 = ~n6653 ;
  assign y3590 = ~n6657 ;
  assign y3591 = n6659 ;
  assign y3592 = ~1'b0 ;
  assign y3593 = ~n3065 ;
  assign y3594 = ~n4803 ;
  assign y3595 = ~n6661 ;
  assign y3596 = n1423 ;
  assign y3597 = ~1'b0 ;
  assign y3598 = n3979 ;
  assign y3599 = ~1'b0 ;
  assign y3600 = ~1'b0 ;
  assign y3601 = ~n6662 ;
  assign y3602 = n6665 ;
  assign y3603 = 1'b0 ;
  assign y3604 = n6666 ;
  assign y3605 = ~1'b0 ;
  assign y3606 = ~1'b0 ;
  assign y3607 = ~1'b0 ;
  assign y3608 = n6667 ;
  assign y3609 = ~x160 ;
  assign y3610 = n6668 ;
  assign y3611 = 1'b0 ;
  assign y3612 = ~1'b0 ;
  assign y3613 = ~n6672 ;
  assign y3614 = n6675 ;
  assign y3615 = ~n6682 ;
  assign y3616 = n6686 ;
  assign y3617 = ~1'b0 ;
  assign y3618 = n4730 ;
  assign y3619 = n6687 ;
  assign y3620 = n6689 ;
  assign y3621 = n6694 ;
  assign y3622 = ~1'b0 ;
  assign y3623 = ~1'b0 ;
  assign y3624 = ~x112 ;
  assign y3625 = ~n6698 ;
  assign y3626 = n6700 ;
  assign y3627 = ~n6271 ;
  assign y3628 = 1'b0 ;
  assign y3629 = n6703 ;
  assign y3630 = ~n6707 ;
  assign y3631 = ~n1920 ;
  assign y3632 = n6708 ;
  assign y3633 = ~n6710 ;
  assign y3634 = ~n6712 ;
  assign y3635 = ~n6714 ;
  assign y3636 = 1'b0 ;
  assign y3637 = n6715 ;
  assign y3638 = n6716 ;
  assign y3639 = n6717 ;
  assign y3640 = n6719 ;
  assign y3641 = ~1'b0 ;
  assign y3642 = ~n6727 ;
  assign y3643 = ~1'b0 ;
  assign y3644 = ~1'b0 ;
  assign y3645 = n6738 ;
  assign y3646 = n6742 ;
  assign y3647 = ~1'b0 ;
  assign y3648 = n6743 ;
  assign y3649 = n5703 ;
  assign y3650 = n6745 ;
  assign y3651 = n6747 ;
  assign y3652 = n6748 ;
  assign y3653 = n1395 ;
  assign y3654 = n6750 ;
  assign y3655 = ~1'b0 ;
  assign y3656 = ~n6754 ;
  assign y3657 = ~x86 ;
  assign y3658 = ~1'b0 ;
  assign y3659 = n6757 ;
  assign y3660 = n6759 ;
  assign y3661 = ~1'b0 ;
  assign y3662 = n6761 ;
  assign y3663 = ~n6764 ;
  assign y3664 = n6769 ;
  assign y3665 = ~1'b0 ;
  assign y3666 = ~1'b0 ;
  assign y3667 = ~1'b0 ;
  assign y3668 = ~n6771 ;
  assign y3669 = n6772 ;
  assign y3670 = ~n5031 ;
  assign y3671 = n4824 ;
  assign y3672 = n6780 ;
  assign y3673 = ~1'b0 ;
  assign y3674 = ~1'b0 ;
  assign y3675 = ~n1914 ;
  assign y3676 = n6781 ;
  assign y3677 = n6782 ;
  assign y3678 = n6783 ;
  assign y3679 = 1'b0 ;
  assign y3680 = 1'b0 ;
  assign y3681 = ~n6785 ;
  assign y3682 = n6788 ;
  assign y3683 = ~n6795 ;
  assign y3684 = ~1'b0 ;
  assign y3685 = ~1'b0 ;
  assign y3686 = n6799 ;
  assign y3687 = n6802 ;
  assign y3688 = n6803 ;
  assign y3689 = ~n6805 ;
  assign y3690 = ~1'b0 ;
  assign y3691 = ~n6811 ;
  assign y3692 = 1'b0 ;
  assign y3693 = n6816 ;
  assign y3694 = n6819 ;
  assign y3695 = ~1'b0 ;
  assign y3696 = ~1'b0 ;
  assign y3697 = n3862 ;
  assign y3698 = n6822 ;
  assign y3699 = n6823 ;
  assign y3700 = ~n6824 ;
  assign y3701 = ~n6825 ;
  assign y3702 = ~n6829 ;
  assign y3703 = ~n6838 ;
  assign y3704 = ~1'b0 ;
  assign y3705 = ~1'b0 ;
  assign y3706 = ~1'b0 ;
  assign y3707 = n6050 ;
  assign y3708 = ~1'b0 ;
  assign y3709 = ~n6840 ;
  assign y3710 = ~n6842 ;
  assign y3711 = ~n6845 ;
  assign y3712 = ~n6846 ;
  assign y3713 = n6849 ;
  assign y3714 = ~n3939 ;
  assign y3715 = n415 ;
  assign y3716 = ~n6858 ;
  assign y3717 = n6865 ;
  assign y3718 = ~1'b0 ;
  assign y3719 = n6868 ;
  assign y3720 = n6874 ;
  assign y3721 = ~n6881 ;
  assign y3722 = n6883 ;
  assign y3723 = ~1'b0 ;
  assign y3724 = n6885 ;
  assign y3725 = ~1'b0 ;
  assign y3726 = ~n6888 ;
  assign y3727 = n2310 ;
  assign y3728 = n6893 ;
  assign y3729 = ~n6897 ;
  assign y3730 = n6898 ;
  assign y3731 = ~n6899 ;
  assign y3732 = n6903 ;
  assign y3733 = ~n6904 ;
  assign y3734 = n6924 ;
  assign y3735 = ~1'b0 ;
  assign y3736 = ~1'b0 ;
  assign y3737 = ~n1588 ;
  assign y3738 = ~1'b0 ;
  assign y3739 = ~n6929 ;
  assign y3740 = n6932 ;
  assign y3741 = ~n4166 ;
  assign y3742 = ~n6934 ;
  assign y3743 = n6935 ;
  assign y3744 = ~n6940 ;
  assign y3745 = ~1'b0 ;
  assign y3746 = ~n6941 ;
  assign y3747 = n1854 ;
  assign y3748 = ~1'b0 ;
  assign y3749 = ~n6944 ;
  assign y3750 = 1'b0 ;
  assign y3751 = n6945 ;
  assign y3752 = ~n6948 ;
  assign y3753 = ~1'b0 ;
  assign y3754 = ~1'b0 ;
  assign y3755 = n6951 ;
  assign y3756 = n6956 ;
  assign y3757 = ~n6960 ;
  assign y3758 = ~n6963 ;
  assign y3759 = ~1'b0 ;
  assign y3760 = ~1'b0 ;
  assign y3761 = ~1'b0 ;
  assign y3762 = ~1'b0 ;
  assign y3763 = ~1'b0 ;
  assign y3764 = n6966 ;
  assign y3765 = ~n6969 ;
  assign y3766 = ~n6974 ;
  assign y3767 = 1'b0 ;
  assign y3768 = ~1'b0 ;
  assign y3769 = n6975 ;
  assign y3770 = n6983 ;
  assign y3771 = ~n6988 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = ~n6993 ;
  assign y3774 = ~n6994 ;
  assign y3775 = n7002 ;
  assign y3776 = ~1'b0 ;
  assign y3777 = ~n1369 ;
  assign y3778 = ~1'b0 ;
  assign y3779 = ~1'b0 ;
  assign y3780 = ~n7003 ;
  assign y3781 = ~n7005 ;
  assign y3782 = ~1'b0 ;
  assign y3783 = ~n7010 ;
  assign y3784 = n7013 ;
  assign y3785 = n7014 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = ~n7015 ;
  assign y3788 = ~n7016 ;
  assign y3789 = ~1'b0 ;
  assign y3790 = ~1'b0 ;
  assign y3791 = ~1'b0 ;
  assign y3792 = n7017 ;
  assign y3793 = ~n7021 ;
  assign y3794 = ~n7023 ;
  assign y3795 = ~1'b0 ;
  assign y3796 = ~1'b0 ;
  assign y3797 = ~n7024 ;
  assign y3798 = ~n7025 ;
  assign y3799 = ~n7026 ;
  assign y3800 = n7028 ;
  assign y3801 = ~n7030 ;
  assign y3802 = n7032 ;
  assign y3803 = ~n7036 ;
  assign y3804 = ~1'b0 ;
  assign y3805 = n7037 ;
  assign y3806 = ~1'b0 ;
  assign y3807 = ~1'b0 ;
  assign y3808 = n7039 ;
  assign y3809 = ~n7040 ;
  assign y3810 = ~n407 ;
  assign y3811 = ~n7049 ;
  assign y3812 = ~n7050 ;
  assign y3813 = ~1'b0 ;
  assign y3814 = ~1'b0 ;
  assign y3815 = ~n2071 ;
  assign y3816 = ~1'b0 ;
  assign y3817 = n7051 ;
  assign y3818 = ~1'b0 ;
  assign y3819 = ~1'b0 ;
  assign y3820 = n7052 ;
  assign y3821 = n1810 ;
  assign y3822 = n7055 ;
  assign y3823 = ~n7057 ;
  assign y3824 = ~n7061 ;
  assign y3825 = ~n7062 ;
  assign y3826 = ~1'b0 ;
  assign y3827 = n7066 ;
  assign y3828 = ~n6570 ;
  assign y3829 = ~n7068 ;
  assign y3830 = ~n7069 ;
  assign y3831 = n7070 ;
  assign y3832 = ~n7072 ;
  assign y3833 = 1'b0 ;
  assign y3834 = n1657 ;
  assign y3835 = 1'b0 ;
  assign y3836 = ~n7074 ;
  assign y3837 = ~1'b0 ;
  assign y3838 = ~n7083 ;
  assign y3839 = n7096 ;
  assign y3840 = ~1'b0 ;
  assign y3841 = ~1'b0 ;
  assign y3842 = ~n7100 ;
  assign y3843 = ~1'b0 ;
  assign y3844 = ~1'b0 ;
  assign y3845 = ~n7102 ;
  assign y3846 = ~1'b0 ;
  assign y3847 = n7103 ;
  assign y3848 = ~1'b0 ;
  assign y3849 = ~n7107 ;
  assign y3850 = ~1'b0 ;
  assign y3851 = ~n7108 ;
  assign y3852 = ~1'b0 ;
  assign y3853 = ~n6941 ;
  assign y3854 = ~1'b0 ;
  assign y3855 = ~1'b0 ;
  assign y3856 = ~1'b0 ;
  assign y3857 = ~1'b0 ;
  assign y3858 = ~n7111 ;
  assign y3859 = n807 ;
  assign y3860 = n7120 ;
  assign y3861 = ~n7124 ;
  assign y3862 = n7126 ;
  assign y3863 = ~1'b0 ;
  assign y3864 = ~n2951 ;
  assign y3865 = n7129 ;
  assign y3866 = n7132 ;
  assign y3867 = n7133 ;
  assign y3868 = ~1'b0 ;
  assign y3869 = ~1'b0 ;
  assign y3870 = n7135 ;
  assign y3871 = n7137 ;
  assign y3872 = n7142 ;
  assign y3873 = ~n7149 ;
  assign y3874 = ~n7154 ;
  assign y3875 = ~n7158 ;
  assign y3876 = n7160 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = ~1'b0 ;
  assign y3879 = ~n7161 ;
  assign y3880 = ~1'b0 ;
  assign y3881 = ~1'b0 ;
  assign y3882 = n7162 ;
  assign y3883 = ~n7169 ;
  assign y3884 = ~n7170 ;
  assign y3885 = ~1'b0 ;
  assign y3886 = ~n7171 ;
  assign y3887 = n4932 ;
  assign y3888 = ~n6962 ;
  assign y3889 = ~n7172 ;
  assign y3890 = ~n7173 ;
  assign y3891 = n7177 ;
  assign y3892 = ~n7179 ;
  assign y3893 = n3461 ;
  assign y3894 = 1'b0 ;
  assign y3895 = ~1'b0 ;
  assign y3896 = ~1'b0 ;
  assign y3897 = ~1'b0 ;
  assign y3898 = ~n7189 ;
  assign y3899 = ~n7194 ;
  assign y3900 = n7199 ;
  assign y3901 = ~1'b0 ;
  assign y3902 = ~n7200 ;
  assign y3903 = ~n7204 ;
  assign y3904 = n7207 ;
  assign y3905 = ~n562 ;
  assign y3906 = n7208 ;
  assign y3907 = n7211 ;
  assign y3908 = ~1'b0 ;
  assign y3909 = ~n7215 ;
  assign y3910 = ~n7216 ;
  assign y3911 = n7221 ;
  assign y3912 = ~1'b0 ;
  assign y3913 = n7223 ;
  assign y3914 = n7229 ;
  assign y3915 = ~n7236 ;
  assign y3916 = ~n7237 ;
  assign y3917 = n3073 ;
  assign y3918 = ~n7241 ;
  assign y3919 = ~n7244 ;
  assign y3920 = ~1'b0 ;
  assign y3921 = ~n7251 ;
  assign y3922 = ~n7253 ;
  assign y3923 = ~n7256 ;
  assign y3924 = ~n7257 ;
  assign y3925 = n7258 ;
  assign y3926 = ~n1709 ;
  assign y3927 = n7259 ;
  assign y3928 = ~n7261 ;
  assign y3929 = n7262 ;
  assign y3930 = ~1'b0 ;
  assign y3931 = n7264 ;
  assign y3932 = ~n7265 ;
  assign y3933 = ~1'b0 ;
  assign y3934 = n7268 ;
  assign y3935 = ~1'b0 ;
  assign y3936 = n5686 ;
  assign y3937 = ~n7270 ;
  assign y3938 = ~1'b0 ;
  assign y3939 = ~n7271 ;
  assign y3940 = ~n7275 ;
  assign y3941 = ~1'b0 ;
  assign y3942 = ~1'b0 ;
  assign y3943 = ~1'b0 ;
  assign y3944 = ~1'b0 ;
  assign y3945 = n7280 ;
  assign y3946 = ~1'b0 ;
  assign y3947 = ~n7284 ;
  assign y3948 = n7285 ;
  assign y3949 = n7290 ;
  assign y3950 = ~n7295 ;
  assign y3951 = n7296 ;
  assign y3952 = ~n7299 ;
  assign y3953 = ~n7303 ;
  assign y3954 = ~n7305 ;
  assign y3955 = ~1'b0 ;
  assign y3956 = n7308 ;
  assign y3957 = ~n7314 ;
  assign y3958 = n1368 ;
  assign y3959 = ~1'b0 ;
  assign y3960 = n7317 ;
  assign y3961 = ~n7319 ;
  assign y3962 = ~1'b0 ;
  assign y3963 = ~n7320 ;
  assign y3964 = n7329 ;
  assign y3965 = ~n7331 ;
  assign y3966 = n4265 ;
  assign y3967 = ~1'b0 ;
  assign y3968 = ~n7335 ;
  assign y3969 = ~1'b0 ;
  assign y3970 = n7338 ;
  assign y3971 = n7340 ;
  assign y3972 = ~1'b0 ;
  assign y3973 = ~n7341 ;
  assign y3974 = ~n7343 ;
  assign y3975 = ~1'b0 ;
  assign y3976 = n7350 ;
  assign y3977 = ~1'b0 ;
  assign y3978 = n7353 ;
  assign y3979 = ~n7355 ;
  assign y3980 = ~1'b0 ;
  assign y3981 = n7358 ;
  assign y3982 = ~1'b0 ;
  assign y3983 = ~n3903 ;
  assign y3984 = ~n519 ;
  assign y3985 = ~n7359 ;
  assign y3986 = n7362 ;
  assign y3987 = ~n7365 ;
  assign y3988 = n7366 ;
  assign y3989 = ~1'b0 ;
  assign y3990 = ~n7367 ;
  assign y3991 = ~n7372 ;
  assign y3992 = ~n7373 ;
  assign y3993 = ~1'b0 ;
  assign y3994 = n7378 ;
  assign y3995 = ~1'b0 ;
  assign y3996 = ~n7382 ;
  assign y3997 = ~1'b0 ;
  assign y3998 = ~n7383 ;
  assign y3999 = ~n7384 ;
  assign y4000 = ~1'b0 ;
  assign y4001 = ~n7386 ;
  assign y4002 = ~n7387 ;
  assign y4003 = ~1'b0 ;
  assign y4004 = n7390 ;
  assign y4005 = n7392 ;
  assign y4006 = n7394 ;
  assign y4007 = ~1'b0 ;
  assign y4008 = ~1'b0 ;
  assign y4009 = n7397 ;
  assign y4010 = ~n7401 ;
  assign y4011 = ~1'b0 ;
  assign y4012 = ~1'b0 ;
  assign y4013 = ~n7403 ;
  assign y4014 = n7404 ;
  assign y4015 = ~n7406 ;
  assign y4016 = ~1'b0 ;
  assign y4017 = ~1'b0 ;
  assign y4018 = n7407 ;
  assign y4019 = ~n7410 ;
  assign y4020 = ~1'b0 ;
  assign y4021 = ~1'b0 ;
  assign y4022 = ~1'b0 ;
  assign y4023 = ~1'b0 ;
  assign y4024 = ~n7413 ;
  assign y4025 = n7414 ;
  assign y4026 = ~1'b0 ;
  assign y4027 = 1'b0 ;
  assign y4028 = n7416 ;
  assign y4029 = ~n7420 ;
  assign y4030 = n7429 ;
  assign y4031 = n7430 ;
  assign y4032 = ~1'b0 ;
  assign y4033 = ~n7438 ;
  assign y4034 = n7443 ;
  assign y4035 = n7446 ;
  assign y4036 = ~n7448 ;
  assign y4037 = n7449 ;
  assign y4038 = n7454 ;
  assign y4039 = ~1'b0 ;
  assign y4040 = 1'b0 ;
  assign y4041 = n7457 ;
  assign y4042 = n7459 ;
  assign y4043 = ~n7466 ;
  assign y4044 = n7467 ;
  assign y4045 = n7471 ;
  assign y4046 = n7475 ;
  assign y4047 = ~n7477 ;
  assign y4048 = ~n7481 ;
  assign y4049 = ~n7483 ;
  assign y4050 = ~n7484 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = ~n7485 ;
  assign y4054 = ~1'b0 ;
  assign y4055 = ~1'b0 ;
  assign y4056 = ~1'b0 ;
  assign y4057 = ~n7489 ;
  assign y4058 = ~1'b0 ;
  assign y4059 = n7491 ;
  assign y4060 = n7494 ;
  assign y4061 = ~n7495 ;
  assign y4062 = ~1'b0 ;
  assign y4063 = n7497 ;
  assign y4064 = ~1'b0 ;
  assign y4065 = n7498 ;
  assign y4066 = n7501 ;
  assign y4067 = ~1'b0 ;
  assign y4068 = ~1'b0 ;
  assign y4069 = ~n7513 ;
  assign y4070 = n7515 ;
  assign y4071 = ~1'b0 ;
  assign y4072 = ~1'b0 ;
  assign y4073 = ~n7516 ;
  assign y4074 = ~n7519 ;
  assign y4075 = ~n7527 ;
  assign y4076 = ~1'b0 ;
  assign y4077 = n7531 ;
  assign y4078 = n7533 ;
  assign y4079 = ~n7536 ;
  assign y4080 = n7540 ;
  assign y4081 = ~n7544 ;
  assign y4082 = n7547 ;
  assign y4083 = ~n7549 ;
  assign y4084 = n7550 ;
  assign y4085 = ~n7552 ;
  assign y4086 = n7557 ;
  assign y4087 = ~n7560 ;
  assign y4088 = 1'b0 ;
  assign y4089 = n7562 ;
  assign y4090 = ~n7563 ;
  assign y4091 = ~1'b0 ;
  assign y4092 = ~1'b0 ;
  assign y4093 = ~1'b0 ;
  assign y4094 = n7568 ;
  assign y4095 = ~n7573 ;
  assign y4096 = ~n5826 ;
  assign y4097 = ~n7314 ;
  assign y4098 = ~n7575 ;
  assign y4099 = ~1'b0 ;
  assign y4100 = n7583 ;
  assign y4101 = ~n7584 ;
  assign y4102 = ~n7588 ;
  assign y4103 = n7591 ;
  assign y4104 = ~1'b0 ;
  assign y4105 = ~1'b0 ;
  assign y4106 = ~1'b0 ;
  assign y4107 = n7593 ;
  assign y4108 = ~n7594 ;
  assign y4109 = ~1'b0 ;
  assign y4110 = ~n7595 ;
  assign y4111 = ~n4026 ;
  assign y4112 = ~n5779 ;
  assign y4113 = ~1'b0 ;
  assign y4114 = ~n7601 ;
  assign y4115 = ~n7603 ;
  assign y4116 = ~1'b0 ;
  assign y4117 = ~n7605 ;
  assign y4118 = ~1'b0 ;
  assign y4119 = n305 ;
  assign y4120 = ~n7126 ;
  assign y4121 = n7608 ;
  assign y4122 = ~n7609 ;
  assign y4123 = n7613 ;
  assign y4124 = ~n7618 ;
  assign y4125 = ~1'b0 ;
  assign y4126 = 1'b0 ;
  assign y4127 = ~n7619 ;
  assign y4128 = ~n7622 ;
  assign y4129 = ~n7624 ;
  assign y4130 = ~1'b0 ;
  assign y4131 = ~1'b0 ;
  assign y4132 = n7625 ;
  assign y4133 = n7630 ;
  assign y4134 = n7632 ;
  assign y4135 = n7633 ;
  assign y4136 = ~n7634 ;
  assign y4137 = n7637 ;
  assign y4138 = n7639 ;
  assign y4139 = n7641 ;
  assign y4140 = ~n7642 ;
  assign y4141 = ~n7643 ;
  assign y4142 = ~n6527 ;
  assign y4143 = n7646 ;
  assign y4144 = ~1'b0 ;
  assign y4145 = ~1'b0 ;
  assign y4146 = n7652 ;
  assign y4147 = ~n5381 ;
  assign y4148 = ~n2310 ;
  assign y4149 = n7164 ;
  assign y4150 = ~1'b0 ;
  assign y4151 = ~n7657 ;
  assign y4152 = ~1'b0 ;
  assign y4153 = ~n7660 ;
  assign y4154 = n7661 ;
  assign y4155 = n7668 ;
  assign y4156 = n7670 ;
  assign y4157 = ~n7675 ;
  assign y4158 = n7681 ;
  assign y4159 = n7682 ;
  assign y4160 = ~1'b0 ;
  assign y4161 = ~1'b0 ;
  assign y4162 = ~1'b0 ;
  assign y4163 = n7684 ;
  assign y4164 = ~n7685 ;
  assign y4165 = ~n7688 ;
  assign y4166 = n4274 ;
  assign y4167 = ~1'b0 ;
  assign y4168 = ~n7689 ;
  assign y4169 = ~n7690 ;
  assign y4170 = n7691 ;
  assign y4171 = n7692 ;
  assign y4172 = 1'b0 ;
  assign y4173 = ~x245 ;
  assign y4174 = ~1'b0 ;
  assign y4175 = ~1'b0 ;
  assign y4176 = ~n7694 ;
  assign y4177 = n4395 ;
  assign y4178 = ~n7696 ;
  assign y4179 = ~n7697 ;
  assign y4180 = n7701 ;
  assign y4181 = ~n3480 ;
  assign y4182 = n7703 ;
  assign y4183 = n7704 ;
  assign y4184 = ~n7705 ;
  assign y4185 = n2752 ;
  assign y4186 = n7706 ;
  assign y4187 = n7709 ;
  assign y4188 = ~n7710 ;
  assign y4189 = n7711 ;
  assign y4190 = n7713 ;
  assign y4191 = ~n7717 ;
  assign y4192 = n7726 ;
  assign y4193 = ~1'b0 ;
  assign y4194 = ~1'b0 ;
  assign y4195 = n7729 ;
  assign y4196 = ~n7730 ;
  assign y4197 = n7732 ;
  assign y4198 = n7734 ;
  assign y4199 = ~n6031 ;
  assign y4200 = ~n7736 ;
  assign y4201 = ~1'b0 ;
  assign y4202 = ~n7738 ;
  assign y4203 = n7739 ;
  assign y4204 = ~1'b0 ;
  assign y4205 = n7743 ;
  assign y4206 = n7745 ;
  assign y4207 = n7746 ;
  assign y4208 = n7749 ;
  assign y4209 = 1'b0 ;
  assign y4210 = ~1'b0 ;
  assign y4211 = ~n7750 ;
  assign y4212 = ~n7754 ;
  assign y4213 = ~n7755 ;
  assign y4214 = ~n7756 ;
  assign y4215 = ~1'b0 ;
  assign y4216 = ~n7761 ;
  assign y4217 = ~1'b0 ;
  assign y4218 = ~n7764 ;
  assign y4219 = ~n6198 ;
  assign y4220 = ~1'b0 ;
  assign y4221 = n7769 ;
  assign y4222 = ~1'b0 ;
  assign y4223 = n7777 ;
  assign y4224 = ~n6381 ;
  assign y4225 = ~1'b0 ;
  assign y4226 = ~1'b0 ;
  assign y4227 = n7778 ;
  assign y4228 = ~n5748 ;
  assign y4229 = ~1'b0 ;
  assign y4230 = ~n7781 ;
  assign y4231 = ~n7783 ;
  assign y4232 = ~n7785 ;
  assign y4233 = ~1'b0 ;
  assign y4234 = ~n7787 ;
  assign y4235 = n7788 ;
  assign y4236 = ~n7789 ;
  assign y4237 = ~1'b0 ;
  assign y4238 = ~1'b0 ;
  assign y4239 = ~1'b0 ;
  assign y4240 = n7791 ;
  assign y4241 = 1'b0 ;
  assign y4242 = ~1'b0 ;
  assign y4243 = ~n7792 ;
  assign y4244 = 1'b0 ;
  assign y4245 = n7796 ;
  assign y4246 = ~n7800 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = ~1'b0 ;
  assign y4249 = n7804 ;
  assign y4250 = ~n7807 ;
  assign y4251 = ~1'b0 ;
  assign y4252 = ~n7809 ;
  assign y4253 = n7810 ;
  assign y4254 = ~n7814 ;
  assign y4255 = n7818 ;
  assign y4256 = 1'b0 ;
  assign y4257 = ~n7821 ;
  assign y4258 = ~n7822 ;
  assign y4259 = ~1'b0 ;
  assign y4260 = n7827 ;
  assign y4261 = ~n7828 ;
  assign y4262 = ~n4485 ;
  assign y4263 = ~1'b0 ;
  assign y4264 = n7835 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = n1684 ;
  assign y4267 = ~1'b0 ;
  assign y4268 = ~1'b0 ;
  assign y4269 = ~n7841 ;
  assign y4270 = ~n7846 ;
  assign y4271 = n7847 ;
  assign y4272 = ~1'b0 ;
  assign y4273 = ~n7849 ;
  assign y4274 = ~1'b0 ;
  assign y4275 = ~1'b0 ;
  assign y4276 = ~n7855 ;
  assign y4277 = ~n7858 ;
  assign y4278 = n7870 ;
  assign y4279 = ~1'b0 ;
  assign y4280 = n7880 ;
  assign y4281 = ~1'b0 ;
  assign y4282 = 1'b0 ;
  assign y4283 = ~1'b0 ;
  assign y4284 = n2735 ;
  assign y4285 = ~1'b0 ;
  assign y4286 = ~n7882 ;
  assign y4287 = ~1'b0 ;
  assign y4288 = ~1'b0 ;
  assign y4289 = ~n7883 ;
  assign y4290 = ~1'b0 ;
  assign y4291 = n7885 ;
  assign y4292 = ~n7892 ;
  assign y4293 = n7893 ;
  assign y4294 = n7894 ;
  assign y4295 = ~n7895 ;
  assign y4296 = ~1'b0 ;
  assign y4297 = n7897 ;
  assign y4298 = ~n7899 ;
  assign y4299 = ~1'b0 ;
  assign y4300 = ~1'b0 ;
  assign y4301 = n7901 ;
  assign y4302 = n3714 ;
  assign y4303 = n7905 ;
  assign y4304 = ~1'b0 ;
  assign y4305 = ~1'b0 ;
  assign y4306 = n7908 ;
  assign y4307 = n7912 ;
  assign y4308 = ~n7915 ;
  assign y4309 = n7917 ;
  assign y4310 = n7918 ;
  assign y4311 = n7925 ;
  assign y4312 = 1'b0 ;
  assign y4313 = n7928 ;
  assign y4314 = ~1'b0 ;
  assign y4315 = ~1'b0 ;
  assign y4316 = ~1'b0 ;
  assign y4317 = n7929 ;
  assign y4318 = n7931 ;
  assign y4319 = 1'b0 ;
  assign y4320 = ~n7933 ;
  assign y4321 = ~1'b0 ;
  assign y4322 = n7937 ;
  assign y4323 = ~n7942 ;
  assign y4324 = ~1'b0 ;
  assign y4325 = n7944 ;
  assign y4326 = n7945 ;
  assign y4327 = ~1'b0 ;
  assign y4328 = ~n7947 ;
  assign y4329 = ~1'b0 ;
  assign y4330 = ~1'b0 ;
  assign y4331 = n7949 ;
  assign y4332 = n7950 ;
  assign y4333 = ~1'b0 ;
  assign y4334 = ~1'b0 ;
  assign y4335 = n4118 ;
  assign y4336 = n7953 ;
  assign y4337 = ~n1920 ;
  assign y4338 = n4350 ;
  assign y4339 = 1'b0 ;
  assign y4340 = ~1'b0 ;
  assign y4341 = ~1'b0 ;
  assign y4342 = ~n7954 ;
  assign y4343 = n809 ;
  assign y4344 = ~1'b0 ;
  assign y4345 = ~1'b0 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = ~n7957 ;
  assign y4348 = n7966 ;
  assign y4349 = ~1'b0 ;
  assign y4350 = n7970 ;
  assign y4351 = ~1'b0 ;
  assign y4352 = n7973 ;
  assign y4353 = ~n7974 ;
  assign y4354 = ~n7977 ;
  assign y4355 = ~1'b0 ;
  assign y4356 = ~n2731 ;
  assign y4357 = ~1'b0 ;
  assign y4358 = ~n7981 ;
  assign y4359 = n7988 ;
  assign y4360 = ~n7993 ;
  assign y4361 = n3943 ;
  assign y4362 = ~n7995 ;
  assign y4363 = n7998 ;
  assign y4364 = ~n8001 ;
  assign y4365 = n2798 ;
  assign y4366 = ~n8004 ;
  assign y4367 = ~1'b0 ;
  assign y4368 = ~n8005 ;
  assign y4369 = n8006 ;
  assign y4370 = ~1'b0 ;
  assign y4371 = ~1'b0 ;
  assign y4372 = n8012 ;
  assign y4373 = ~1'b0 ;
  assign y4374 = n8017 ;
  assign y4375 = ~1'b0 ;
  assign y4376 = n8019 ;
  assign y4377 = n8020 ;
  assign y4378 = ~1'b0 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = ~1'b0 ;
  assign y4381 = n8023 ;
  assign y4382 = ~1'b0 ;
  assign y4383 = ~n8024 ;
  assign y4384 = ~1'b0 ;
  assign y4385 = n5091 ;
  assign y4386 = ~n8025 ;
  assign y4387 = n8027 ;
  assign y4388 = ~1'b0 ;
  assign y4389 = ~n8028 ;
  assign y4390 = ~n8035 ;
  assign y4391 = ~n8038 ;
  assign y4392 = ~1'b0 ;
  assign y4393 = ~n7169 ;
  assign y4394 = n8039 ;
  assign y4395 = ~n8041 ;
  assign y4396 = n8045 ;
  assign y4397 = n8048 ;
  assign y4398 = ~n8055 ;
  assign y4399 = ~n8056 ;
  assign y4400 = n8058 ;
  assign y4401 = ~n8059 ;
  assign y4402 = ~n5781 ;
  assign y4403 = n8060 ;
  assign y4404 = ~1'b0 ;
  assign y4405 = n8063 ;
  assign y4406 = ~1'b0 ;
  assign y4407 = ~1'b0 ;
  assign y4408 = n8064 ;
  assign y4409 = ~1'b0 ;
  assign y4410 = ~n8070 ;
  assign y4411 = n8076 ;
  assign y4412 = n8079 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = ~n8081 ;
  assign y4415 = n968 ;
  assign y4416 = ~n8082 ;
  assign y4417 = ~1'b0 ;
  assign y4418 = ~1'b0 ;
  assign y4419 = ~1'b0 ;
  assign y4420 = n8083 ;
  assign y4421 = ~n8084 ;
  assign y4422 = ~n8089 ;
  assign y4423 = ~n8091 ;
  assign y4424 = n8093 ;
  assign y4425 = ~n8095 ;
  assign y4426 = ~1'b0 ;
  assign y4427 = ~1'b0 ;
  assign y4428 = ~n8101 ;
  assign y4429 = ~n5201 ;
  assign y4430 = ~n8104 ;
  assign y4431 = ~1'b0 ;
  assign y4432 = n7567 ;
  assign y4433 = ~1'b0 ;
  assign y4434 = ~n8106 ;
  assign y4435 = ~n8107 ;
  assign y4436 = ~1'b0 ;
  assign y4437 = n8108 ;
  assign y4438 = ~n8111 ;
  assign y4439 = ~n8112 ;
  assign y4440 = ~1'b0 ;
  assign y4441 = ~n8113 ;
  assign y4442 = ~1'b0 ;
  assign y4443 = 1'b0 ;
  assign y4444 = ~n8115 ;
  assign y4445 = ~1'b0 ;
  assign y4446 = ~1'b0 ;
  assign y4447 = ~1'b0 ;
  assign y4448 = ~1'b0 ;
  assign y4449 = n8116 ;
  assign y4450 = n8118 ;
  assign y4451 = n8121 ;
  assign y4452 = ~1'b0 ;
  assign y4453 = ~1'b0 ;
  assign y4454 = ~n8127 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = n562 ;
  assign y4457 = n8128 ;
  assign y4458 = ~n8130 ;
  assign y4459 = ~n8133 ;
  assign y4460 = 1'b0 ;
  assign y4461 = 1'b0 ;
  assign y4462 = ~1'b0 ;
  assign y4463 = n7202 ;
  assign y4464 = n6054 ;
  assign y4465 = n8138 ;
  assign y4466 = ~n8139 ;
  assign y4467 = ~n8144 ;
  assign y4468 = n8145 ;
  assign y4469 = ~n8146 ;
  assign y4470 = ~1'b0 ;
  assign y4471 = n8148 ;
  assign y4472 = ~1'b0 ;
  assign y4473 = ~n8150 ;
  assign y4474 = ~n8151 ;
  assign y4475 = n8155 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = n8161 ;
  assign y4478 = ~n8162 ;
  assign y4479 = ~n7170 ;
  assign y4480 = 1'b0 ;
  assign y4481 = ~1'b0 ;
  assign y4482 = n8168 ;
  assign y4483 = ~1'b0 ;
  assign y4484 = ~n8169 ;
  assign y4485 = ~1'b0 ;
  assign y4486 = n8170 ;
  assign y4487 = ~1'b0 ;
  assign y4488 = n8174 ;
  assign y4489 = ~n8175 ;
  assign y4490 = n8176 ;
  assign y4491 = n8180 ;
  assign y4492 = ~n2315 ;
  assign y4493 = ~n8181 ;
  assign y4494 = ~n8191 ;
  assign y4495 = ~n8195 ;
  assign y4496 = n8196 ;
  assign y4497 = n8202 ;
  assign y4498 = n8203 ;
  assign y4499 = ~n8205 ;
  assign y4500 = n8208 ;
  assign y4501 = n8209 ;
  assign y4502 = ~n8214 ;
  assign y4503 = n8215 ;
  assign y4504 = ~1'b0 ;
  assign y4505 = ~1'b0 ;
  assign y4506 = n8216 ;
  assign y4507 = n8217 ;
  assign y4508 = ~n8221 ;
  assign y4509 = n8226 ;
  assign y4510 = ~n8229 ;
  assign y4511 = ~1'b0 ;
  assign y4512 = ~1'b0 ;
  assign y4513 = ~1'b0 ;
  assign y4514 = ~1'b0 ;
  assign y4515 = ~1'b0 ;
  assign y4516 = ~n8230 ;
  assign y4517 = ~1'b0 ;
  assign y4518 = ~1'b0 ;
  assign y4519 = ~1'b0 ;
  assign y4520 = ~n8231 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n343 ;
  assign y4523 = ~n8232 ;
  assign y4524 = ~n8233 ;
  assign y4525 = n5776 ;
  assign y4526 = ~n8236 ;
  assign y4527 = ~1'b0 ;
  assign y4528 = n8237 ;
  assign y4529 = ~1'b0 ;
  assign y4530 = ~n8241 ;
  assign y4531 = n1610 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = ~1'b0 ;
  assign y4534 = ~1'b0 ;
  assign y4535 = ~n8242 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = ~n3263 ;
  assign y4538 = n2072 ;
  assign y4539 = ~1'b0 ;
  assign y4540 = ~1'b0 ;
  assign y4541 = n8244 ;
  assign y4542 = ~n8246 ;
  assign y4543 = ~n8248 ;
  assign y4544 = ~1'b0 ;
  assign y4545 = ~n8249 ;
  assign y4546 = ~1'b0 ;
  assign y4547 = ~n6647 ;
  assign y4548 = ~1'b0 ;
  assign y4549 = n8250 ;
  assign y4550 = ~n8254 ;
  assign y4551 = n8261 ;
  assign y4552 = ~n8263 ;
  assign y4553 = ~n8273 ;
  assign y4554 = ~n8276 ;
  assign y4555 = n8278 ;
  assign y4556 = n8279 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = n8280 ;
  assign y4559 = ~n8285 ;
  assign y4560 = n8287 ;
  assign y4561 = n8288 ;
  assign y4562 = ~1'b0 ;
  assign y4563 = n8289 ;
  assign y4564 = ~n8291 ;
  assign y4565 = n8293 ;
  assign y4566 = n8294 ;
  assign y4567 = ~1'b0 ;
  assign y4568 = n8295 ;
  assign y4569 = ~1'b0 ;
  assign y4570 = n8297 ;
  assign y4571 = n8299 ;
  assign y4572 = ~n1061 ;
  assign y4573 = ~n8301 ;
  assign y4574 = ~n8305 ;
  assign y4575 = ~n8314 ;
  assign y4576 = n8319 ;
  assign y4577 = ~1'b0 ;
  assign y4578 = ~n8322 ;
  assign y4579 = 1'b0 ;
  assign y4580 = ~1'b0 ;
  assign y4581 = n8329 ;
  assign y4582 = n8331 ;
  assign y4583 = ~n8332 ;
  assign y4584 = ~1'b0 ;
  assign y4585 = n8334 ;
  assign y4586 = ~n8341 ;
  assign y4587 = n8349 ;
  assign y4588 = n8351 ;
  assign y4589 = ~1'b0 ;
  assign y4590 = 1'b0 ;
  assign y4591 = ~n8356 ;
  assign y4592 = ~1'b0 ;
  assign y4593 = n8360 ;
  assign y4594 = ~1'b0 ;
  assign y4595 = ~n8363 ;
  assign y4596 = n8364 ;
  assign y4597 = ~1'b0 ;
  assign y4598 = ~1'b0 ;
  assign y4599 = ~n8365 ;
  assign y4600 = n3181 ;
  assign y4601 = ~1'b0 ;
  assign y4602 = ~n8367 ;
  assign y4603 = ~x28 ;
  assign y4604 = ~n8369 ;
  assign y4605 = ~n8373 ;
  assign y4606 = 1'b0 ;
  assign y4607 = ~1'b0 ;
  assign y4608 = ~1'b0 ;
  assign y4609 = ~n8377 ;
  assign y4610 = ~1'b0 ;
  assign y4611 = ~1'b0 ;
  assign y4612 = ~1'b0 ;
  assign y4613 = ~n8381 ;
  assign y4614 = n8382 ;
  assign y4615 = n3026 ;
  assign y4616 = ~1'b0 ;
  assign y4617 = n8383 ;
  assign y4618 = ~n8384 ;
  assign y4619 = ~n8388 ;
  assign y4620 = ~1'b0 ;
  assign y4621 = ~1'b0 ;
  assign y4622 = ~n3432 ;
  assign y4623 = n8389 ;
  assign y4624 = ~n8401 ;
  assign y4625 = n7864 ;
  assign y4626 = ~1'b0 ;
  assign y4627 = ~n8404 ;
  assign y4628 = ~1'b0 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = n8406 ;
  assign y4631 = ~1'b0 ;
  assign y4632 = ~1'b0 ;
  assign y4633 = ~1'b0 ;
  assign y4634 = ~1'b0 ;
  assign y4635 = 1'b0 ;
  assign y4636 = n8408 ;
  assign y4637 = ~n8410 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = 1'b0 ;
  assign y4640 = n8411 ;
  assign y4641 = ~1'b0 ;
  assign y4642 = ~n8415 ;
  assign y4643 = n8416 ;
  assign y4644 = n7634 ;
  assign y4645 = ~1'b0 ;
  assign y4646 = n8417 ;
  assign y4647 = ~n8427 ;
  assign y4648 = ~1'b0 ;
  assign y4649 = ~n8428 ;
  assign y4650 = ~1'b0 ;
  assign y4651 = ~1'b0 ;
  assign y4652 = n8433 ;
  assign y4653 = ~1'b0 ;
  assign y4654 = ~1'b0 ;
  assign y4655 = ~n3015 ;
  assign y4656 = ~n8436 ;
  assign y4657 = ~1'b0 ;
  assign y4658 = ~n8437 ;
  assign y4659 = ~1'b0 ;
  assign y4660 = ~1'b0 ;
  assign y4661 = n8438 ;
  assign y4662 = ~1'b0 ;
  assign y4663 = n8443 ;
  assign y4664 = ~1'b0 ;
  assign y4665 = ~n8444 ;
  assign y4666 = n8446 ;
  assign y4667 = ~n8137 ;
  assign y4668 = n8448 ;
  assign y4669 = ~n600 ;
  assign y4670 = n8453 ;
  assign y4671 = ~1'b0 ;
  assign y4672 = n8454 ;
  assign y4673 = ~1'b0 ;
  assign y4674 = n8457 ;
  assign y4675 = n8460 ;
  assign y4676 = n8461 ;
  assign y4677 = ~1'b0 ;
  assign y4678 = ~1'b0 ;
  assign y4679 = ~1'b0 ;
  assign y4680 = n4238 ;
  assign y4681 = ~n8462 ;
  assign y4682 = n8463 ;
  assign y4683 = ~1'b0 ;
  assign y4684 = ~1'b0 ;
  assign y4685 = n8464 ;
  assign y4686 = 1'b0 ;
  assign y4687 = ~n8467 ;
  assign y4688 = n8469 ;
  assign y4689 = ~1'b0 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = ~1'b0 ;
  assign y4692 = ~n8470 ;
  assign y4693 = ~1'b0 ;
  assign y4694 = ~n8472 ;
  assign y4695 = ~n8474 ;
  assign y4696 = n8475 ;
  assign y4697 = n1071 ;
  assign y4698 = n8477 ;
  assign y4699 = n8480 ;
  assign y4700 = ~1'b0 ;
  assign y4701 = ~1'b0 ;
  assign y4702 = n8487 ;
  assign y4703 = n8497 ;
  assign y4704 = ~1'b0 ;
  assign y4705 = ~n8500 ;
  assign y4706 = ~n8501 ;
  assign y4707 = ~1'b0 ;
  assign y4708 = ~1'b0 ;
  assign y4709 = ~n8506 ;
  assign y4710 = ~n8507 ;
  assign y4711 = n8508 ;
  assign y4712 = ~n8511 ;
  assign y4713 = n8513 ;
  assign y4714 = ~n8520 ;
  assign y4715 = ~n8522 ;
  assign y4716 = n8524 ;
  assign y4717 = ~n8525 ;
  assign y4718 = ~n8526 ;
  assign y4719 = ~1'b0 ;
  assign y4720 = n8528 ;
  assign y4721 = ~n3243 ;
  assign y4722 = ~1'b0 ;
  assign y4723 = n8536 ;
  assign y4724 = ~1'b0 ;
  assign y4725 = ~1'b0 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = ~1'b0 ;
  assign y4728 = ~n8543 ;
  assign y4729 = ~1'b0 ;
  assign y4730 = n8545 ;
  assign y4731 = n8546 ;
  assign y4732 = ~n8550 ;
  assign y4733 = ~1'b0 ;
  assign y4734 = n8554 ;
  assign y4735 = ~1'b0 ;
  assign y4736 = ~1'b0 ;
  assign y4737 = n8555 ;
  assign y4738 = ~n8559 ;
  assign y4739 = ~n8562 ;
  assign y4740 = ~n8564 ;
  assign y4741 = n8568 ;
  assign y4742 = ~n8572 ;
  assign y4743 = ~n8573 ;
  assign y4744 = ~n8576 ;
  assign y4745 = ~1'b0 ;
  assign y4746 = 1'b0 ;
  assign y4747 = ~n8588 ;
  assign y4748 = ~1'b0 ;
  assign y4749 = ~1'b0 ;
  assign y4750 = ~1'b0 ;
  assign y4751 = ~1'b0 ;
  assign y4752 = ~1'b0 ;
  assign y4753 = ~n8591 ;
  assign y4754 = n8594 ;
  assign y4755 = ~1'b0 ;
  assign y4756 = n8597 ;
  assign y4757 = 1'b0 ;
  assign y4758 = ~n8600 ;
  assign y4759 = ~n8602 ;
  assign y4760 = ~1'b0 ;
  assign y4761 = n8604 ;
  assign y4762 = n8608 ;
  assign y4763 = ~1'b0 ;
  assign y4764 = ~n8609 ;
  assign y4765 = n8613 ;
  assign y4766 = ~n8617 ;
  assign y4767 = 1'b0 ;
  assign y4768 = n8630 ;
  assign y4769 = ~n8631 ;
  assign y4770 = ~n8633 ;
  assign y4771 = ~n8635 ;
  assign y4772 = 1'b0 ;
  assign y4773 = ~1'b0 ;
  assign y4774 = n8640 ;
  assign y4775 = n8642 ;
  assign y4776 = n8645 ;
  assign y4777 = ~n8646 ;
  assign y4778 = ~1'b0 ;
  assign y4779 = n8649 ;
  assign y4780 = ~n8651 ;
  assign y4781 = n8212 ;
  assign y4782 = n8656 ;
  assign y4783 = ~1'b0 ;
  assign y4784 = n8657 ;
  assign y4785 = ~1'b0 ;
  assign y4786 = ~n8659 ;
  assign y4787 = ~1'b0 ;
  assign y4788 = ~n8663 ;
  assign y4789 = 1'b0 ;
  assign y4790 = n1372 ;
  assign y4791 = ~1'b0 ;
  assign y4792 = n8665 ;
  assign y4793 = ~n8667 ;
  assign y4794 = ~n8669 ;
  assign y4795 = ~1'b0 ;
  assign y4796 = ~n8674 ;
  assign y4797 = ~1'b0 ;
  assign y4798 = ~1'b0 ;
  assign y4799 = n8675 ;
  assign y4800 = ~n8677 ;
  assign y4801 = ~1'b0 ;
  assign y4802 = n8679 ;
  assign y4803 = ~n8683 ;
  assign y4804 = n6146 ;
  assign y4805 = n8684 ;
  assign y4806 = ~1'b0 ;
  assign y4807 = n8689 ;
  assign y4808 = ~n8692 ;
  assign y4809 = n8693 ;
  assign y4810 = n8696 ;
  assign y4811 = n8697 ;
  assign y4812 = ~1'b0 ;
  assign y4813 = ~n8698 ;
  assign y4814 = n8700 ;
  assign y4815 = ~1'b0 ;
  assign y4816 = n8702 ;
  assign y4817 = ~n8703 ;
  assign y4818 = n8704 ;
  assign y4819 = ~n8707 ;
  assign y4820 = n8709 ;
  assign y4821 = ~1'b0 ;
  assign y4822 = ~1'b0 ;
  assign y4823 = n8710 ;
  assign y4824 = n8713 ;
  assign y4825 = n8716 ;
  assign y4826 = n2431 ;
  assign y4827 = n8721 ;
  assign y4828 = n926 ;
  assign y4829 = ~n8724 ;
  assign y4830 = n8729 ;
  assign y4831 = ~1'b0 ;
  assign y4832 = ~n8731 ;
  assign y4833 = n8734 ;
  assign y4834 = ~1'b0 ;
  assign y4835 = ~n8735 ;
  assign y4836 = n8740 ;
  assign y4837 = ~1'b0 ;
  assign y4838 = n8743 ;
  assign y4839 = ~1'b0 ;
  assign y4840 = ~1'b0 ;
  assign y4841 = ~1'b0 ;
  assign y4842 = ~n8747 ;
  assign y4843 = ~n8750 ;
  assign y4844 = ~n8752 ;
  assign y4845 = n8759 ;
  assign y4846 = n8761 ;
  assign y4847 = ~n8764 ;
  assign y4848 = n8767 ;
  assign y4849 = n8768 ;
  assign y4850 = ~n8771 ;
  assign y4851 = ~n8774 ;
  assign y4852 = ~n8791 ;
  assign y4853 = ~n8792 ;
  assign y4854 = ~1'b0 ;
  assign y4855 = ~n8793 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = ~n8796 ;
  assign y4858 = ~n8799 ;
  assign y4859 = 1'b0 ;
  assign y4860 = ~1'b0 ;
  assign y4861 = n8804 ;
  assign y4862 = n8809 ;
  assign y4863 = ~n8814 ;
  assign y4864 = ~n8816 ;
  assign y4865 = n8819 ;
  assign y4866 = ~1'b0 ;
  assign y4867 = ~n1920 ;
  assign y4868 = n8820 ;
  assign y4869 = ~1'b0 ;
  assign y4870 = 1'b0 ;
  assign y4871 = ~n8825 ;
  assign y4872 = ~n8830 ;
  assign y4873 = ~1'b0 ;
  assign y4874 = ~n4723 ;
  assign y4875 = n4119 ;
  assign y4876 = ~1'b0 ;
  assign y4877 = ~n8832 ;
  assign y4878 = ~1'b0 ;
  assign y4879 = n8834 ;
  assign y4880 = n8835 ;
  assign y4881 = ~1'b0 ;
  assign y4882 = n8837 ;
  assign y4883 = ~1'b0 ;
  assign y4884 = n3181 ;
  assign y4885 = ~n8841 ;
  assign y4886 = n8842 ;
  assign y4887 = ~1'b0 ;
  assign y4888 = ~n8846 ;
  assign y4889 = ~n8850 ;
  assign y4890 = n6461 ;
  assign y4891 = n8851 ;
  assign y4892 = ~n8855 ;
  assign y4893 = ~1'b0 ;
  assign y4894 = ~n8856 ;
  assign y4895 = ~n8870 ;
  assign y4896 = n8877 ;
  assign y4897 = n8879 ;
  assign y4898 = ~1'b0 ;
  assign y4899 = ~n8881 ;
  assign y4900 = n8888 ;
  assign y4901 = n8889 ;
  assign y4902 = n8892 ;
  assign y4903 = n8893 ;
  assign y4904 = ~1'b0 ;
  assign y4905 = ~1'b0 ;
  assign y4906 = ~n8896 ;
  assign y4907 = n5796 ;
  assign y4908 = ~1'b0 ;
  assign y4909 = 1'b0 ;
  assign y4910 = n8897 ;
  assign y4911 = ~1'b0 ;
  assign y4912 = n8901 ;
  assign y4913 = ~n8905 ;
  assign y4914 = n8907 ;
  assign y4915 = ~1'b0 ;
  assign y4916 = ~n8909 ;
  assign y4917 = ~1'b0 ;
  assign y4918 = ~1'b0 ;
  assign y4919 = 1'b0 ;
  assign y4920 = 1'b0 ;
  assign y4921 = ~n8910 ;
  assign y4922 = ~1'b0 ;
  assign y4923 = n8912 ;
  assign y4924 = ~n8913 ;
  assign y4925 = ~n8916 ;
  assign y4926 = ~1'b0 ;
  assign y4927 = ~1'b0 ;
  assign y4928 = ~1'b0 ;
  assign y4929 = n7032 ;
  assign y4930 = 1'b0 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = ~n8918 ;
  assign y4933 = ~n8919 ;
  assign y4934 = ~1'b0 ;
  assign y4935 = ~1'b0 ;
  assign y4936 = n8923 ;
  assign y4937 = ~1'b0 ;
  assign y4938 = ~1'b0 ;
  assign y4939 = ~n8925 ;
  assign y4940 = ~1'b0 ;
  assign y4941 = ~1'b0 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = ~1'b0 ;
  assign y4944 = ~n8929 ;
  assign y4945 = ~n8932 ;
  assign y4946 = ~1'b0 ;
  assign y4947 = ~1'b0 ;
  assign y4948 = ~1'b0 ;
  assign y4949 = ~n8933 ;
  assign y4950 = ~1'b0 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = n8937 ;
  assign y4953 = n8939 ;
  assign y4954 = ~n8942 ;
  assign y4955 = ~n8945 ;
  assign y4956 = ~1'b0 ;
  assign y4957 = ~1'b0 ;
  assign y4958 = n2860 ;
  assign y4959 = ~n8953 ;
  assign y4960 = n3333 ;
  assign y4961 = ~n8957 ;
  assign y4962 = ~1'b0 ;
  assign y4963 = ~1'b0 ;
  assign y4964 = ~1'b0 ;
  assign y4965 = n8959 ;
  assign y4966 = ~1'b0 ;
  assign y4967 = 1'b0 ;
  assign y4968 = n8960 ;
  assign y4969 = ~n8964 ;
  assign y4970 = ~n8967 ;
  assign y4971 = ~n8972 ;
  assign y4972 = ~1'b0 ;
  assign y4973 = n8976 ;
  assign y4974 = n8989 ;
  assign y4975 = ~1'b0 ;
  assign y4976 = n8990 ;
  assign y4977 = ~1'b0 ;
  assign y4978 = ~1'b0 ;
  assign y4979 = ~1'b0 ;
  assign y4980 = ~1'b0 ;
  assign y4981 = n8993 ;
  assign y4982 = ~1'b0 ;
  assign y4983 = n8750 ;
  assign y4984 = ~n8997 ;
  assign y4985 = n9001 ;
  assign y4986 = ~n9003 ;
  assign y4987 = ~1'b0 ;
  assign y4988 = n9004 ;
  assign y4989 = ~1'b0 ;
  assign y4990 = ~1'b0 ;
  assign y4991 = ~n9005 ;
  assign y4992 = ~1'b0 ;
  assign y4993 = n9010 ;
  assign y4994 = ~n9011 ;
  assign y4995 = n9015 ;
  assign y4996 = n9018 ;
  assign y4997 = ~1'b0 ;
  assign y4998 = n5597 ;
  assign y4999 = ~n9019 ;
  assign y5000 = ~n9026 ;
  assign y5001 = ~n5292 ;
  assign y5002 = n9027 ;
  assign y5003 = n9035 ;
  assign y5004 = 1'b0 ;
  assign y5005 = n9041 ;
  assign y5006 = n9045 ;
  assign y5007 = ~n9049 ;
  assign y5008 = ~1'b0 ;
  assign y5009 = ~1'b0 ;
  assign y5010 = ~1'b0 ;
  assign y5011 = ~1'b0 ;
  assign y5012 = ~n9055 ;
  assign y5013 = n9057 ;
  assign y5014 = ~n9059 ;
  assign y5015 = n9060 ;
  assign y5016 = ~n9061 ;
  assign y5017 = ~n9062 ;
  assign y5018 = ~n9063 ;
  assign y5019 = n9065 ;
  assign y5020 = ~1'b0 ;
  assign y5021 = ~n9072 ;
  assign y5022 = 1'b0 ;
  assign y5023 = ~n9074 ;
  assign y5024 = ~1'b0 ;
  assign y5025 = n9075 ;
  assign y5026 = ~n6423 ;
  assign y5027 = n8706 ;
  assign y5028 = ~1'b0 ;
  assign y5029 = n9076 ;
  assign y5030 = n9078 ;
  assign y5031 = ~n9080 ;
  assign y5032 = n9081 ;
  assign y5033 = ~n9083 ;
  assign y5034 = n9084 ;
  assign y5035 = ~1'b0 ;
  assign y5036 = n9085 ;
  assign y5037 = n9086 ;
  assign y5038 = ~n1630 ;
  assign y5039 = n2901 ;
  assign y5040 = ~1'b0 ;
  assign y5041 = ~1'b0 ;
  assign y5042 = ~n9092 ;
  assign y5043 = ~1'b0 ;
  assign y5044 = ~1'b0 ;
  assign y5045 = ~n9095 ;
  assign y5046 = n9097 ;
  assign y5047 = ~n9099 ;
  assign y5048 = ~n9100 ;
  assign y5049 = ~n4655 ;
  assign y5050 = ~n1727 ;
  assign y5051 = n9101 ;
  assign y5052 = ~1'b0 ;
  assign y5053 = ~1'b0 ;
  assign y5054 = n9103 ;
  assign y5055 = ~n8621 ;
  assign y5056 = ~1'b0 ;
  assign y5057 = ~1'b0 ;
  assign y5058 = n9104 ;
  assign y5059 = ~1'b0 ;
  assign y5060 = ~n9105 ;
  assign y5061 = ~1'b0 ;
  assign y5062 = ~1'b0 ;
  assign y5063 = ~1'b0 ;
  assign y5064 = 1'b0 ;
  assign y5065 = ~1'b0 ;
  assign y5066 = ~1'b0 ;
  assign y5067 = n9108 ;
  assign y5068 = ~1'b0 ;
  assign y5069 = ~n7427 ;
  assign y5070 = n9109 ;
  assign y5071 = ~1'b0 ;
  assign y5072 = n9114 ;
  assign y5073 = n9117 ;
  assign y5074 = ~n9118 ;
  assign y5075 = ~1'b0 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = ~n9125 ;
  assign y5078 = n9126 ;
  assign y5079 = n9128 ;
  assign y5080 = ~n9129 ;
  assign y5081 = ~n9132 ;
  assign y5082 = ~1'b0 ;
  assign y5083 = ~n9139 ;
  assign y5084 = n9141 ;
  assign y5085 = ~n9144 ;
  assign y5086 = ~n9146 ;
  assign y5087 = 1'b0 ;
  assign y5088 = ~1'b0 ;
  assign y5089 = ~n9148 ;
  assign y5090 = ~1'b0 ;
  assign y5091 = ~1'b0 ;
  assign y5092 = ~n3669 ;
  assign y5093 = ~1'b0 ;
  assign y5094 = 1'b0 ;
  assign y5095 = n9152 ;
  assign y5096 = n9153 ;
  assign y5097 = ~1'b0 ;
  assign y5098 = ~1'b0 ;
  assign y5099 = ~n9154 ;
  assign y5100 = ~1'b0 ;
  assign y5101 = n9160 ;
  assign y5102 = ~1'b0 ;
  assign y5103 = ~1'b0 ;
  assign y5104 = ~1'b0 ;
  assign y5105 = ~n8821 ;
  assign y5106 = ~n9167 ;
  assign y5107 = ~n9170 ;
  assign y5108 = n9173 ;
  assign y5109 = ~n9175 ;
  assign y5110 = ~1'b0 ;
  assign y5111 = ~n9176 ;
  assign y5112 = n9181 ;
  assign y5113 = ~n2503 ;
  assign y5114 = ~n9184 ;
  assign y5115 = n9186 ;
  assign y5116 = ~n590 ;
  assign y5117 = ~n9190 ;
  assign y5118 = ~n5225 ;
  assign y5119 = ~1'b0 ;
  assign y5120 = ~1'b0 ;
  assign y5121 = n9194 ;
  assign y5122 = n9195 ;
  assign y5123 = n9196 ;
  assign y5124 = n9197 ;
  assign y5125 = ~1'b0 ;
  assign y5126 = ~1'b0 ;
  assign y5127 = ~1'b0 ;
  assign y5128 = ~1'b0 ;
  assign y5129 = ~1'b0 ;
  assign y5130 = n9203 ;
  assign y5131 = ~1'b0 ;
  assign y5132 = n9205 ;
  assign y5133 = n9207 ;
  assign y5134 = n9211 ;
  assign y5135 = ~n9212 ;
  assign y5136 = ~1'b0 ;
  assign y5137 = ~1'b0 ;
  assign y5138 = ~n7395 ;
  assign y5139 = ~1'b0 ;
  assign y5140 = ~1'b0 ;
  assign y5141 = n9213 ;
  assign y5142 = n9214 ;
  assign y5143 = n9217 ;
  assign y5144 = n9222 ;
  assign y5145 = n9225 ;
  assign y5146 = ~n9227 ;
  assign y5147 = n9231 ;
  assign y5148 = n9232 ;
  assign y5149 = n9233 ;
  assign y5150 = ~1'b0 ;
  assign y5151 = ~n8933 ;
  assign y5152 = 1'b0 ;
  assign y5153 = ~1'b0 ;
  assign y5154 = ~1'b0 ;
  assign y5155 = ~n3454 ;
  assign y5156 = n9238 ;
  assign y5157 = ~1'b0 ;
  assign y5158 = ~n5067 ;
  assign y5159 = ~n9244 ;
  assign y5160 = ~n9248 ;
  assign y5161 = n9250 ;
  assign y5162 = 1'b0 ;
  assign y5163 = ~n9252 ;
  assign y5164 = ~n9263 ;
  assign y5165 = n9264 ;
  assign y5166 = ~n9267 ;
  assign y5167 = n9272 ;
  assign y5168 = ~n9277 ;
  assign y5169 = ~1'b0 ;
  assign y5170 = n4179 ;
  assign y5171 = n9279 ;
  assign y5172 = n9281 ;
  assign y5173 = ~n9287 ;
  assign y5174 = ~1'b0 ;
  assign y5175 = ~n5824 ;
  assign y5176 = ~n5624 ;
  assign y5177 = n9290 ;
  assign y5178 = ~n9291 ;
  assign y5179 = ~n1926 ;
  assign y5180 = ~n9296 ;
  assign y5181 = ~n9300 ;
  assign y5182 = ~1'b0 ;
  assign y5183 = ~1'b0 ;
  assign y5184 = ~n9303 ;
  assign y5185 = ~1'b0 ;
  assign y5186 = ~1'b0 ;
  assign y5187 = ~1'b0 ;
  assign y5188 = n9305 ;
  assign y5189 = n9306 ;
  assign y5190 = n9308 ;
  assign y5191 = n9310 ;
  assign y5192 = n9311 ;
  assign y5193 = ~1'b0 ;
  assign y5194 = ~1'b0 ;
  assign y5195 = ~1'b0 ;
  assign y5196 = ~1'b0 ;
  assign y5197 = n9313 ;
  assign y5198 = 1'b0 ;
  assign y5199 = ~1'b0 ;
  assign y5200 = ~n9314 ;
  assign y5201 = ~n9315 ;
  assign y5202 = n3026 ;
  assign y5203 = n9321 ;
  assign y5204 = n3718 ;
  assign y5205 = ~1'b0 ;
  assign y5206 = ~1'b0 ;
  assign y5207 = ~n9324 ;
  assign y5208 = ~1'b0 ;
  assign y5209 = ~1'b0 ;
  assign y5210 = ~n9326 ;
  assign y5211 = 1'b0 ;
  assign y5212 = ~n9327 ;
  assign y5213 = 1'b0 ;
  assign y5214 = n9335 ;
  assign y5215 = ~1'b0 ;
  assign y5216 = ~1'b0 ;
  assign y5217 = ~n9337 ;
  assign y5218 = ~n965 ;
  assign y5219 = n9341 ;
  assign y5220 = ~n9343 ;
  assign y5221 = ~1'b0 ;
  assign y5222 = ~n9344 ;
  assign y5223 = ~n9349 ;
  assign y5224 = ~1'b0 ;
  assign y5225 = ~n9350 ;
  assign y5226 = ~1'b0 ;
  assign y5227 = n9352 ;
  assign y5228 = n9361 ;
  assign y5229 = ~1'b0 ;
  assign y5230 = ~1'b0 ;
  assign y5231 = ~1'b0 ;
  assign y5232 = ~1'b0 ;
  assign y5233 = ~1'b0 ;
  assign y5234 = ~1'b0 ;
  assign y5235 = n9362 ;
  assign y5236 = ~n9363 ;
  assign y5237 = n2325 ;
  assign y5238 = n9367 ;
  assign y5239 = ~n9368 ;
  assign y5240 = n9369 ;
  assign y5241 = ~n9371 ;
  assign y5242 = ~n9373 ;
  assign y5243 = ~1'b0 ;
  assign y5244 = ~n9374 ;
  assign y5245 = ~n9376 ;
  assign y5246 = ~n9377 ;
  assign y5247 = ~n9378 ;
  assign y5248 = n9381 ;
  assign y5249 = n9382 ;
  assign y5250 = n9386 ;
  assign y5251 = n9388 ;
  assign y5252 = ~1'b0 ;
  assign y5253 = ~n9391 ;
  assign y5254 = ~1'b0 ;
  assign y5255 = 1'b0 ;
  assign y5256 = ~n9393 ;
  assign y5257 = n9394 ;
  assign y5258 = ~1'b0 ;
  assign y5259 = ~1'b0 ;
  assign y5260 = ~1'b0 ;
  assign y5261 = ~n1324 ;
  assign y5262 = ~n9395 ;
  assign y5263 = 1'b0 ;
  assign y5264 = n8672 ;
  assign y5265 = ~n9396 ;
  assign y5266 = n8841 ;
  assign y5267 = n9398 ;
  assign y5268 = n9399 ;
  assign y5269 = n9402 ;
  assign y5270 = n9412 ;
  assign y5271 = ~n9413 ;
  assign y5272 = ~n3798 ;
  assign y5273 = n9415 ;
  assign y5274 = ~1'b0 ;
  assign y5275 = n9417 ;
  assign y5276 = n552 ;
  assign y5277 = ~1'b0 ;
  assign y5278 = ~1'b0 ;
  assign y5279 = n9425 ;
  assign y5280 = n9427 ;
  assign y5281 = ~1'b0 ;
  assign y5282 = ~n9430 ;
  assign y5283 = ~1'b0 ;
  assign y5284 = n9431 ;
  assign y5285 = ~n9432 ;
  assign y5286 = n9438 ;
  assign y5287 = ~1'b0 ;
  assign y5288 = ~1'b0 ;
  assign y5289 = ~n9439 ;
  assign y5290 = n9442 ;
  assign y5291 = ~1'b0 ;
  assign y5292 = n9445 ;
  assign y5293 = ~n9448 ;
  assign y5294 = n9451 ;
  assign y5295 = n9454 ;
  assign y5296 = ~n9465 ;
  assign y5297 = ~n9468 ;
  assign y5298 = ~1'b0 ;
  assign y5299 = ~1'b0 ;
  assign y5300 = ~n8811 ;
  assign y5301 = ~1'b0 ;
  assign y5302 = n9470 ;
  assign y5303 = ~1'b0 ;
  assign y5304 = ~1'b0 ;
  assign y5305 = ~1'b0 ;
  assign y5306 = ~1'b0 ;
  assign y5307 = n9473 ;
  assign y5308 = ~n9475 ;
  assign y5309 = ~1'b0 ;
  assign y5310 = n3940 ;
  assign y5311 = n9479 ;
  assign y5312 = ~1'b0 ;
  assign y5313 = ~1'b0 ;
  assign y5314 = n9482 ;
  assign y5315 = ~1'b0 ;
  assign y5316 = ~n9484 ;
  assign y5317 = ~n9491 ;
  assign y5318 = n9492 ;
  assign y5319 = n9495 ;
  assign y5320 = n9497 ;
  assign y5321 = ~n9498 ;
  assign y5322 = ~n9499 ;
  assign y5323 = ~n9502 ;
  assign y5324 = ~n9514 ;
  assign y5325 = 1'b0 ;
  assign y5326 = n9516 ;
  assign y5327 = n9517 ;
  assign y5328 = n9523 ;
  assign y5329 = ~n9528 ;
  assign y5330 = 1'b0 ;
  assign y5331 = ~n9532 ;
  assign y5332 = n9535 ;
  assign y5333 = ~1'b0 ;
  assign y5334 = n9540 ;
  assign y5335 = ~1'b0 ;
  assign y5336 = ~1'b0 ;
  assign y5337 = ~1'b0 ;
  assign y5338 = n9541 ;
  assign y5339 = n9547 ;
  assign y5340 = ~n9553 ;
  assign y5341 = ~1'b0 ;
  assign y5342 = ~n5110 ;
  assign y5343 = x170 ;
  assign y5344 = ~n2267 ;
  assign y5345 = n9554 ;
  assign y5346 = n9555 ;
  assign y5347 = ~n9556 ;
  assign y5348 = n9559 ;
  assign y5349 = ~1'b0 ;
  assign y5350 = ~1'b0 ;
  assign y5351 = ~x113 ;
  assign y5352 = n9560 ;
  assign y5353 = n9564 ;
  assign y5354 = ~1'b0 ;
  assign y5355 = ~1'b0 ;
  assign y5356 = ~1'b0 ;
  assign y5357 = n9565 ;
  assign y5358 = n9568 ;
  assign y5359 = ~1'b0 ;
  assign y5360 = ~1'b0 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = ~n9571 ;
  assign y5363 = ~1'b0 ;
  assign y5364 = n9576 ;
  assign y5365 = 1'b0 ;
  assign y5366 = n9578 ;
  assign y5367 = n9580 ;
  assign y5368 = ~n9585 ;
  assign y5369 = ~n385 ;
  assign y5370 = n9587 ;
  assign y5371 = n9588 ;
  assign y5372 = x181 ;
  assign y5373 = n5082 ;
  assign y5374 = n9593 ;
  assign y5375 = n9597 ;
  assign y5376 = n9598 ;
  assign y5377 = ~n9600 ;
  assign y5378 = ~1'b0 ;
  assign y5379 = ~1'b0 ;
  assign y5380 = ~x182 ;
  assign y5381 = ~1'b0 ;
  assign y5382 = ~n5670 ;
  assign y5383 = ~1'b0 ;
  assign y5384 = n9606 ;
  assign y5385 = ~n9608 ;
  assign y5386 = n9616 ;
  assign y5387 = ~n9617 ;
  assign y5388 = n9622 ;
  assign y5389 = n9626 ;
  assign y5390 = ~n9627 ;
  assign y5391 = ~1'b0 ;
  assign y5392 = ~n1006 ;
  assign y5393 = n9632 ;
  assign y5394 = ~1'b0 ;
  assign y5395 = ~1'b0 ;
  assign y5396 = n9636 ;
  assign y5397 = ~1'b0 ;
  assign y5398 = ~n9649 ;
  assign y5399 = ~n9655 ;
  assign y5400 = ~1'b0 ;
  assign y5401 = n9661 ;
  assign y5402 = ~n9663 ;
  assign y5403 = ~n9665 ;
  assign y5404 = ~n9677 ;
  assign y5405 = n9684 ;
  assign y5406 = ~n9685 ;
  assign y5407 = ~1'b0 ;
  assign y5408 = ~n9687 ;
  assign y5409 = ~n9690 ;
  assign y5410 = ~n9696 ;
  assign y5411 = ~1'b0 ;
  assign y5412 = n9700 ;
  assign y5413 = ~n9703 ;
  assign y5414 = n9708 ;
  assign y5415 = ~n9710 ;
  assign y5416 = ~n9714 ;
  assign y5417 = ~n9717 ;
  assign y5418 = ~n9720 ;
  assign y5419 = n7749 ;
  assign y5420 = ~1'b0 ;
  assign y5421 = ~1'b0 ;
  assign y5422 = ~n9726 ;
  assign y5423 = n9730 ;
  assign y5424 = n9731 ;
  assign y5425 = ~1'b0 ;
  assign y5426 = ~1'b0 ;
  assign y5427 = ~1'b0 ;
  assign y5428 = ~n7148 ;
  assign y5429 = ~n9732 ;
  assign y5430 = ~1'b0 ;
  assign y5431 = ~1'b0 ;
  assign y5432 = ~n9739 ;
  assign y5433 = ~1'b0 ;
  assign y5434 = ~1'b0 ;
  assign y5435 = n9741 ;
  assign y5436 = ~n9752 ;
  assign y5437 = 1'b0 ;
  assign y5438 = ~1'b0 ;
  assign y5439 = 1'b0 ;
  assign y5440 = ~1'b0 ;
  assign y5441 = ~n9755 ;
  assign y5442 = n9760 ;
  assign y5443 = ~1'b0 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = ~1'b0 ;
  assign y5446 = ~1'b0 ;
  assign y5447 = n9764 ;
  assign y5448 = ~1'b0 ;
  assign y5449 = ~n9766 ;
  assign y5450 = n9771 ;
  assign y5451 = n7475 ;
  assign y5452 = ~1'b0 ;
  assign y5453 = ~n9781 ;
  assign y5454 = n9786 ;
  assign y5455 = ~1'b0 ;
  assign y5456 = ~n9788 ;
  assign y5457 = ~n9789 ;
  assign y5458 = ~n9791 ;
  assign y5459 = ~1'b0 ;
  assign y5460 = 1'b0 ;
  assign y5461 = ~1'b0 ;
  assign y5462 = ~n9793 ;
  assign y5463 = n9794 ;
  assign y5464 = n9795 ;
  assign y5465 = ~n9796 ;
  assign y5466 = ~n9802 ;
  assign y5467 = n9803 ;
  assign y5468 = ~1'b0 ;
  assign y5469 = ~n9806 ;
  assign y5470 = ~n6149 ;
  assign y5471 = ~n9811 ;
  assign y5472 = n9817 ;
  assign y5473 = ~1'b0 ;
  assign y5474 = ~n9819 ;
  assign y5475 = ~1'b0 ;
  assign y5476 = n4814 ;
  assign y5477 = ~1'b0 ;
  assign y5478 = 1'b0 ;
  assign y5479 = ~n9820 ;
  assign y5480 = ~1'b0 ;
  assign y5481 = n9821 ;
  assign y5482 = ~1'b0 ;
  assign y5483 = ~n9827 ;
  assign y5484 = n9831 ;
  assign y5485 = ~1'b0 ;
  assign y5486 = n9834 ;
  assign y5487 = n9793 ;
  assign y5488 = ~n9835 ;
  assign y5489 = n9836 ;
  assign y5490 = ~1'b0 ;
  assign y5491 = n9837 ;
  assign y5492 = ~n9852 ;
  assign y5493 = ~n9854 ;
  assign y5494 = ~1'b0 ;
  assign y5495 = ~n9857 ;
  assign y5496 = ~1'b0 ;
  assign y5497 = ~1'b0 ;
  assign y5498 = 1'b0 ;
  assign y5499 = n1393 ;
  assign y5500 = ~n3485 ;
  assign y5501 = ~1'b0 ;
  assign y5502 = ~1'b0 ;
  assign y5503 = ~n9862 ;
  assign y5504 = ~n9863 ;
  assign y5505 = n9865 ;
  assign y5506 = ~n9866 ;
  assign y5507 = 1'b0 ;
  assign y5508 = n2887 ;
  assign y5509 = n9869 ;
  assign y5510 = ~n9873 ;
  assign y5511 = n9874 ;
  assign y5512 = ~n9876 ;
  assign y5513 = ~n9877 ;
  assign y5514 = ~1'b0 ;
  assign y5515 = ~1'b0 ;
  assign y5516 = ~1'b0 ;
  assign y5517 = ~1'b0 ;
  assign y5518 = n9879 ;
  assign y5519 = ~1'b0 ;
  assign y5520 = ~1'b0 ;
  assign y5521 = n9881 ;
  assign y5522 = ~1'b0 ;
  assign y5523 = ~1'b0 ;
  assign y5524 = ~1'b0 ;
  assign y5525 = ~n5756 ;
  assign y5526 = ~n9888 ;
  assign y5527 = ~n9890 ;
  assign y5528 = ~1'b0 ;
  assign y5529 = ~1'b0 ;
  assign y5530 = 1'b0 ;
  assign y5531 = ~n5875 ;
  assign y5532 = ~1'b0 ;
  assign y5533 = n4664 ;
  assign y5534 = n9891 ;
  assign y5535 = ~n9896 ;
  assign y5536 = ~n9897 ;
  assign y5537 = ~1'b0 ;
  assign y5538 = n9905 ;
  assign y5539 = n9907 ;
  assign y5540 = ~n9909 ;
  assign y5541 = ~n9921 ;
  assign y5542 = n9922 ;
  assign y5543 = ~n9923 ;
  assign y5544 = n9926 ;
  assign y5545 = ~n9928 ;
  assign y5546 = ~1'b0 ;
  assign y5547 = n9933 ;
  assign y5548 = n9934 ;
  assign y5549 = n9937 ;
  assign y5550 = ~n9950 ;
  assign y5551 = n9955 ;
  assign y5552 = ~1'b0 ;
  assign y5553 = ~n9956 ;
  assign y5554 = ~n9963 ;
  assign y5555 = n9964 ;
  assign y5556 = ~1'b0 ;
  assign y5557 = ~1'b0 ;
  assign y5558 = ~1'b0 ;
  assign y5559 = ~n9965 ;
  assign y5560 = ~1'b0 ;
  assign y5561 = n9969 ;
  assign y5562 = ~1'b0 ;
  assign y5563 = ~1'b0 ;
  assign y5564 = n9976 ;
  assign y5565 = n9978 ;
  assign y5566 = n9988 ;
  assign y5567 = ~n9989 ;
  assign y5568 = 1'b0 ;
  assign y5569 = ~1'b0 ;
  assign y5570 = ~n9991 ;
  assign y5571 = ~n9992 ;
  assign y5572 = ~n9993 ;
  assign y5573 = 1'b0 ;
  assign y5574 = ~n3343 ;
  assign y5575 = ~1'b0 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = n9996 ;
  assign y5578 = ~1'b0 ;
  assign y5579 = ~n10002 ;
  assign y5580 = ~n10005 ;
  assign y5581 = ~1'b0 ;
  assign y5582 = ~1'b0 ;
  assign y5583 = ~n10006 ;
  assign y5584 = ~n10008 ;
  assign y5585 = n10016 ;
  assign y5586 = n2725 ;
  assign y5587 = ~1'b0 ;
  assign y5588 = ~1'b0 ;
  assign y5589 = n10017 ;
  assign y5590 = ~1'b0 ;
  assign y5591 = ~n3064 ;
  assign y5592 = ~1'b0 ;
  assign y5593 = n7212 ;
  assign y5594 = ~1'b0 ;
  assign y5595 = n5838 ;
  assign y5596 = ~1'b0 ;
  assign y5597 = ~n10019 ;
  assign y5598 = n10023 ;
  assign y5599 = ~n2210 ;
  assign y5600 = ~1'b0 ;
  assign y5601 = ~n10025 ;
  assign y5602 = ~n10026 ;
  assign y5603 = 1'b0 ;
  assign y5604 = ~n10027 ;
  assign y5605 = ~n10030 ;
  assign y5606 = n6021 ;
  assign y5607 = ~n10033 ;
  assign y5608 = ~n10037 ;
  assign y5609 = n10044 ;
  assign y5610 = ~n10046 ;
  assign y5611 = ~n4118 ;
  assign y5612 = n10048 ;
  assign y5613 = n10051 ;
  assign y5614 = ~n10052 ;
  assign y5615 = n10056 ;
  assign y5616 = ~n10061 ;
  assign y5617 = n10063 ;
  assign y5618 = ~1'b0 ;
  assign y5619 = n10068 ;
  assign y5620 = n10072 ;
  assign y5621 = ~1'b0 ;
  assign y5622 = n10078 ;
  assign y5623 = ~1'b0 ;
  assign y5624 = ~1'b0 ;
  assign y5625 = ~1'b0 ;
  assign y5626 = n10081 ;
  assign y5627 = n10082 ;
  assign y5628 = n10084 ;
  assign y5629 = ~1'b0 ;
  assign y5630 = n5097 ;
  assign y5631 = ~1'b0 ;
  assign y5632 = n10086 ;
  assign y5633 = n10087 ;
  assign y5634 = ~n10095 ;
  assign y5635 = n10098 ;
  assign y5636 = ~1'b0 ;
  assign y5637 = n10101 ;
  assign y5638 = ~1'b0 ;
  assign y5639 = n10102 ;
  assign y5640 = 1'b0 ;
  assign y5641 = n10106 ;
  assign y5642 = ~n10108 ;
  assign y5643 = ~1'b0 ;
  assign y5644 = ~1'b0 ;
  assign y5645 = ~1'b0 ;
  assign y5646 = ~1'b0 ;
  assign y5647 = n10114 ;
  assign y5648 = ~1'b0 ;
  assign y5649 = 1'b0 ;
  assign y5650 = n10120 ;
  assign y5651 = ~n10121 ;
  assign y5652 = n10122 ;
  assign y5653 = 1'b0 ;
  assign y5654 = ~n10124 ;
  assign y5655 = n10133 ;
  assign y5656 = ~n10136 ;
  assign y5657 = n10143 ;
  assign y5658 = n10145 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = ~1'b0 ;
  assign y5661 = ~1'b0 ;
  assign y5662 = n10147 ;
  assign y5663 = ~n3022 ;
  assign y5664 = ~n10150 ;
  assign y5665 = ~n10158 ;
  assign y5666 = ~n10160 ;
  assign y5667 = n10163 ;
  assign y5668 = n10164 ;
  assign y5669 = n10166 ;
  assign y5670 = n10167 ;
  assign y5671 = ~1'b0 ;
  assign y5672 = ~1'b0 ;
  assign y5673 = ~1'b0 ;
  assign y5674 = ~1'b0 ;
  assign y5675 = n10168 ;
  assign y5676 = n10169 ;
  assign y5677 = ~n10171 ;
  assign y5678 = ~n10177 ;
  assign y5679 = n10181 ;
  assign y5680 = ~n10185 ;
  assign y5681 = n10188 ;
  assign y5682 = ~n10189 ;
  assign y5683 = ~n10195 ;
  assign y5684 = ~n10198 ;
  assign y5685 = ~n10201 ;
  assign y5686 = ~1'b0 ;
  assign y5687 = n10203 ;
  assign y5688 = n10205 ;
  assign y5689 = ~1'b0 ;
  assign y5690 = ~1'b0 ;
  assign y5691 = ~n10208 ;
  assign y5692 = ~n10210 ;
  assign y5693 = n10211 ;
  assign y5694 = 1'b0 ;
  assign y5695 = ~1'b0 ;
  assign y5696 = ~1'b0 ;
  assign y5697 = ~1'b0 ;
  assign y5698 = n10218 ;
  assign y5699 = 1'b0 ;
  assign y5700 = ~1'b0 ;
  assign y5701 = ~1'b0 ;
  assign y5702 = ~n10220 ;
  assign y5703 = n10222 ;
  assign y5704 = ~1'b0 ;
  assign y5705 = ~n10225 ;
  assign y5706 = ~1'b0 ;
  assign y5707 = ~n10226 ;
  assign y5708 = ~1'b0 ;
  assign y5709 = ~1'b0 ;
  assign y5710 = ~n10234 ;
  assign y5711 = ~n10237 ;
  assign y5712 = n10238 ;
  assign y5713 = n10239 ;
  assign y5714 = n4720 ;
  assign y5715 = ~1'b0 ;
  assign y5716 = ~n10240 ;
  assign y5717 = n10241 ;
  assign y5718 = ~n9222 ;
  assign y5719 = ~1'b0 ;
  assign y5720 = n10258 ;
  assign y5721 = n10261 ;
  assign y5722 = ~n10262 ;
  assign y5723 = ~1'b0 ;
  assign y5724 = ~n10263 ;
  assign y5725 = ~1'b0 ;
  assign y5726 = n10265 ;
  assign y5727 = ~n10267 ;
  assign y5728 = ~1'b0 ;
  assign y5729 = n10270 ;
  assign y5730 = ~1'b0 ;
  assign y5731 = n10271 ;
  assign y5732 = ~n10273 ;
  assign y5733 = ~n10276 ;
  assign y5734 = ~1'b0 ;
  assign y5735 = ~n10279 ;
  assign y5736 = n10280 ;
  assign y5737 = ~1'b0 ;
  assign y5738 = ~n10281 ;
  assign y5739 = ~1'b0 ;
  assign y5740 = n10283 ;
  assign y5741 = ~n2153 ;
  assign y5742 = n10294 ;
  assign y5743 = n10297 ;
  assign y5744 = ~1'b0 ;
  assign y5745 = n10298 ;
  assign y5746 = n10303 ;
  assign y5747 = ~1'b0 ;
  assign y5748 = ~n820 ;
  assign y5749 = ~n10305 ;
  assign y5750 = ~n6900 ;
  assign y5751 = ~1'b0 ;
  assign y5752 = ~1'b0 ;
  assign y5753 = 1'b0 ;
  assign y5754 = n10308 ;
  assign y5755 = n10311 ;
  assign y5756 = ~n10314 ;
  assign y5757 = ~n10323 ;
  assign y5758 = ~1'b0 ;
  assign y5759 = ~1'b0 ;
  assign y5760 = ~n10325 ;
  assign y5761 = n10332 ;
  assign y5762 = ~n10344 ;
  assign y5763 = n10345 ;
  assign y5764 = ~1'b0 ;
  assign y5765 = n10347 ;
  assign y5766 = n10350 ;
  assign y5767 = n10356 ;
  assign y5768 = ~n10358 ;
  assign y5769 = n5095 ;
  assign y5770 = ~1'b0 ;
  assign y5771 = ~1'b0 ;
  assign y5772 = ~1'b0 ;
  assign y5773 = ~1'b0 ;
  assign y5774 = n10359 ;
  assign y5775 = n9609 ;
  assign y5776 = ~1'b0 ;
  assign y5777 = ~1'b0 ;
  assign y5778 = ~1'b0 ;
  assign y5779 = n10360 ;
  assign y5780 = n10375 ;
  assign y5781 = n10376 ;
  assign y5782 = n10381 ;
  assign y5783 = ~n6703 ;
  assign y5784 = n10382 ;
  assign y5785 = n10383 ;
  assign y5786 = n10389 ;
  assign y5787 = ~n10392 ;
  assign y5788 = ~n10395 ;
  assign y5789 = n10399 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = ~1'b0 ;
  assign y5792 = n10402 ;
  assign y5793 = ~1'b0 ;
  assign y5794 = ~n10406 ;
  assign y5795 = ~1'b0 ;
  assign y5796 = n10408 ;
  assign y5797 = ~n2026 ;
  assign y5798 = n10410 ;
  assign y5799 = n10414 ;
  assign y5800 = ~n10416 ;
  assign y5801 = n10418 ;
  assign y5802 = ~1'b0 ;
  assign y5803 = n10420 ;
  assign y5804 = n10423 ;
  assign y5805 = n10436 ;
  assign y5806 = ~n10443 ;
  assign y5807 = ~1'b0 ;
  assign y5808 = n10445 ;
  assign y5809 = ~1'b0 ;
  assign y5810 = n10451 ;
  assign y5811 = n10452 ;
  assign y5812 = ~1'b0 ;
  assign y5813 = n10454 ;
  assign y5814 = ~1'b0 ;
  assign y5815 = n10457 ;
  assign y5816 = ~n3423 ;
  assign y5817 = ~x95 ;
  assign y5818 = ~n10458 ;
  assign y5819 = 1'b0 ;
  assign y5820 = ~1'b0 ;
  assign y5821 = 1'b0 ;
  assign y5822 = n10462 ;
  assign y5823 = ~n10464 ;
  assign y5824 = n10465 ;
  assign y5825 = ~1'b0 ;
  assign y5826 = ~n10468 ;
  assign y5827 = ~1'b0 ;
  assign y5828 = n10469 ;
  assign y5829 = n10471 ;
  assign y5830 = ~x153 ;
  assign y5831 = ~n3414 ;
  assign y5832 = ~n10472 ;
  assign y5833 = n10473 ;
  assign y5834 = ~1'b0 ;
  assign y5835 = ~n10482 ;
  assign y5836 = ~1'b0 ;
  assign y5837 = ~n10485 ;
  assign y5838 = ~n10490 ;
  assign y5839 = n10492 ;
  assign y5840 = ~n10496 ;
  assign y5841 = n10503 ;
  assign y5842 = n10504 ;
  assign y5843 = 1'b0 ;
  assign y5844 = n10505 ;
  assign y5845 = ~n3622 ;
  assign y5846 = ~1'b0 ;
  assign y5847 = 1'b0 ;
  assign y5848 = ~n10507 ;
  assign y5849 = ~1'b0 ;
  assign y5850 = ~1'b0 ;
  assign y5851 = 1'b0 ;
  assign y5852 = n512 ;
  assign y5853 = ~n10511 ;
  assign y5854 = ~1'b0 ;
  assign y5855 = n10514 ;
  assign y5856 = ~1'b0 ;
  assign y5857 = n10519 ;
  assign y5858 = ~n10522 ;
  assign y5859 = ~1'b0 ;
  assign y5860 = ~n10526 ;
  assign y5861 = n10527 ;
  assign y5862 = n8892 ;
  assign y5863 = ~n10535 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = ~1'b0 ;
  assign y5866 = n10540 ;
  assign y5867 = ~n10545 ;
  assign y5868 = ~1'b0 ;
  assign y5869 = ~n10551 ;
  assign y5870 = ~n10553 ;
  assign y5871 = ~1'b0 ;
  assign y5872 = ~n10556 ;
  assign y5873 = n10557 ;
  assign y5874 = ~1'b0 ;
  assign y5875 = n10558 ;
  assign y5876 = ~n10561 ;
  assign y5877 = ~n10563 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = ~n10573 ;
  assign y5880 = ~1'b0 ;
  assign y5881 = ~1'b0 ;
  assign y5882 = n3862 ;
  assign y5883 = n10576 ;
  assign y5884 = n3177 ;
  assign y5885 = n10577 ;
  assign y5886 = n10583 ;
  assign y5887 = n10584 ;
  assign y5888 = ~1'b0 ;
  assign y5889 = ~1'b0 ;
  assign y5890 = ~1'b0 ;
  assign y5891 = n10587 ;
  assign y5892 = n10588 ;
  assign y5893 = ~1'b0 ;
  assign y5894 = ~n10593 ;
  assign y5895 = ~1'b0 ;
  assign y5896 = ~1'b0 ;
  assign y5897 = ~1'b0 ;
  assign y5898 = ~n10595 ;
  assign y5899 = ~n992 ;
  assign y5900 = ~1'b0 ;
  assign y5901 = ~1'b0 ;
  assign y5902 = ~1'b0 ;
  assign y5903 = n10599 ;
  assign y5904 = ~1'b0 ;
  assign y5905 = ~n10601 ;
  assign y5906 = n10602 ;
  assign y5907 = ~n10604 ;
  assign y5908 = ~n10605 ;
  assign y5909 = n10610 ;
  assign y5910 = ~1'b0 ;
  assign y5911 = n1976 ;
  assign y5912 = n10612 ;
  assign y5913 = ~1'b0 ;
  assign y5914 = ~n3520 ;
  assign y5915 = n10614 ;
  assign y5916 = ~n10616 ;
  assign y5917 = n10617 ;
  assign y5918 = n10622 ;
  assign y5919 = n10623 ;
  assign y5920 = ~n8202 ;
  assign y5921 = ~n10624 ;
  assign y5922 = n10627 ;
  assign y5923 = ~n10629 ;
  assign y5924 = n10632 ;
  assign y5925 = n10642 ;
  assign y5926 = ~1'b0 ;
  assign y5927 = ~1'b0 ;
  assign y5928 = n1451 ;
  assign y5929 = n10643 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = ~1'b0 ;
  assign y5932 = n10646 ;
  assign y5933 = n10649 ;
  assign y5934 = n10653 ;
  assign y5935 = ~1'b0 ;
  assign y5936 = ~n10655 ;
  assign y5937 = ~1'b0 ;
  assign y5938 = n10659 ;
  assign y5939 = ~n10665 ;
  assign y5940 = ~n10666 ;
  assign y5941 = n10669 ;
  assign y5942 = n10672 ;
  assign y5943 = ~1'b0 ;
  assign y5944 = n10674 ;
  assign y5945 = ~1'b0 ;
  assign y5946 = n10679 ;
  assign y5947 = ~1'b0 ;
  assign y5948 = n9312 ;
  assign y5949 = ~n10681 ;
  assign y5950 = ~n10684 ;
  assign y5951 = n10687 ;
  assign y5952 = ~1'b0 ;
  assign y5953 = ~n10690 ;
  assign y5954 = n10692 ;
  assign y5955 = ~n10695 ;
  assign y5956 = ~n458 ;
  assign y5957 = n10697 ;
  assign y5958 = ~1'b0 ;
  assign y5959 = ~1'b0 ;
  assign y5960 = n7659 ;
  assign y5961 = ~1'b0 ;
  assign y5962 = n10698 ;
  assign y5963 = ~1'b0 ;
  assign y5964 = 1'b0 ;
  assign y5965 = n10700 ;
  assign y5966 = n10701 ;
  assign y5967 = ~n10702 ;
  assign y5968 = n10703 ;
  assign y5969 = ~1'b0 ;
  assign y5970 = n10705 ;
  assign y5971 = ~1'b0 ;
  assign y5972 = ~1'b0 ;
  assign y5973 = ~n10708 ;
  assign y5974 = n10709 ;
  assign y5975 = n10712 ;
  assign y5976 = 1'b0 ;
  assign y5977 = ~1'b0 ;
  assign y5978 = n10716 ;
  assign y5979 = ~1'b0 ;
  assign y5980 = 1'b0 ;
  assign y5981 = 1'b0 ;
  assign y5982 = ~1'b0 ;
  assign y5983 = ~1'b0 ;
  assign y5984 = ~n10718 ;
  assign y5985 = n10721 ;
  assign y5986 = ~1'b0 ;
  assign y5987 = ~1'b0 ;
  assign y5988 = n10723 ;
  assign y5989 = ~1'b0 ;
  assign y5990 = 1'b0 ;
  assign y5991 = 1'b0 ;
  assign y5992 = ~1'b0 ;
  assign y5993 = 1'b0 ;
  assign y5994 = ~1'b0 ;
  assign y5995 = n10724 ;
  assign y5996 = n10725 ;
  assign y5997 = ~n10733 ;
  assign y5998 = ~1'b0 ;
  assign y5999 = ~1'b0 ;
  assign y6000 = n10741 ;
  assign y6001 = ~n10742 ;
  assign y6002 = n10748 ;
  assign y6003 = ~n10751 ;
  assign y6004 = ~1'b0 ;
  assign y6005 = n10753 ;
  assign y6006 = ~n10757 ;
  assign y6007 = n10758 ;
  assign y6008 = n10760 ;
  assign y6009 = n10764 ;
  assign y6010 = n10766 ;
  assign y6011 = n10767 ;
  assign y6012 = ~1'b0 ;
  assign y6013 = ~n10768 ;
  assign y6014 = n10770 ;
  assign y6015 = n10771 ;
  assign y6016 = ~1'b0 ;
  assign y6017 = ~n10773 ;
  assign y6018 = n10774 ;
  assign y6019 = ~1'b0 ;
  assign y6020 = ~1'b0 ;
  assign y6021 = ~n10105 ;
  assign y6022 = ~n10776 ;
  assign y6023 = n10777 ;
  assign y6024 = n10778 ;
  assign y6025 = ~n10780 ;
  assign y6026 = n10781 ;
  assign y6027 = ~n10782 ;
  assign y6028 = ~n10783 ;
  assign y6029 = ~1'b0 ;
  assign y6030 = ~n10785 ;
  assign y6031 = ~n10792 ;
  assign y6032 = n10795 ;
  assign y6033 = n10798 ;
  assign y6034 = ~1'b0 ;
  assign y6035 = ~1'b0 ;
  assign y6036 = ~n10803 ;
  assign y6037 = n10809 ;
  assign y6038 = ~n5207 ;
  assign y6039 = ~n10816 ;
  assign y6040 = n10817 ;
  assign y6041 = ~1'b0 ;
  assign y6042 = ~n10818 ;
  assign y6043 = ~n10821 ;
  assign y6044 = ~n10822 ;
  assign y6045 = ~1'b0 ;
  assign y6046 = ~1'b0 ;
  assign y6047 = ~n10824 ;
  assign y6048 = ~n10831 ;
  assign y6049 = n10836 ;
  assign y6050 = ~n5564 ;
  assign y6051 = ~n10838 ;
  assign y6052 = ~1'b0 ;
  assign y6053 = ~1'b0 ;
  assign y6054 = ~n3324 ;
  assign y6055 = n977 ;
  assign y6056 = n10842 ;
  assign y6057 = ~n10843 ;
  assign y6058 = ~1'b0 ;
  assign y6059 = ~n10844 ;
  assign y6060 = ~1'b0 ;
  assign y6061 = ~n10847 ;
  assign y6062 = ~1'b0 ;
  assign y6063 = ~1'b0 ;
  assign y6064 = ~1'b0 ;
  assign y6065 = ~n10851 ;
  assign y6066 = ~1'b0 ;
  assign y6067 = ~n10854 ;
  assign y6068 = ~1'b0 ;
  assign y6069 = ~n4678 ;
  assign y6070 = ~n10855 ;
  assign y6071 = ~n10856 ;
  assign y6072 = ~n1623 ;
  assign y6073 = n10858 ;
  assign y6074 = n10860 ;
  assign y6075 = n10863 ;
  assign y6076 = ~n10864 ;
  assign y6077 = n10867 ;
  assign y6078 = n10871 ;
  assign y6079 = ~1'b0 ;
  assign y6080 = ~1'b0 ;
  assign y6081 = n10873 ;
  assign y6082 = n10878 ;
  assign y6083 = ~n10885 ;
  assign y6084 = ~n10886 ;
  assign y6085 = ~n10888 ;
  assign y6086 = ~1'b0 ;
  assign y6087 = ~1'b0 ;
  assign y6088 = ~n10890 ;
  assign y6089 = n10893 ;
  assign y6090 = ~n1596 ;
  assign y6091 = ~n10895 ;
  assign y6092 = n10898 ;
  assign y6093 = ~n10904 ;
  assign y6094 = ~1'b0 ;
  assign y6095 = n10906 ;
  assign y6096 = ~1'b0 ;
  assign y6097 = ~1'b0 ;
  assign y6098 = ~n10909 ;
  assign y6099 = ~n10911 ;
  assign y6100 = ~n10912 ;
  assign y6101 = ~1'b0 ;
  assign y6102 = ~1'b0 ;
  assign y6103 = ~n10913 ;
  assign y6104 = n10914 ;
  assign y6105 = ~n10915 ;
  assign y6106 = ~n10918 ;
  assign y6107 = ~n10919 ;
  assign y6108 = ~1'b0 ;
  assign y6109 = ~1'b0 ;
  assign y6110 = ~1'b0 ;
  assign y6111 = ~1'b0 ;
  assign y6112 = ~1'b0 ;
  assign y6113 = ~1'b0 ;
  assign y6114 = n10922 ;
  assign y6115 = n10928 ;
  assign y6116 = ~1'b0 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = n10929 ;
  assign y6119 = 1'b0 ;
  assign y6120 = ~1'b0 ;
  assign y6121 = ~n10933 ;
  assign y6122 = n10936 ;
  assign y6123 = ~1'b0 ;
  assign y6124 = ~1'b0 ;
  assign y6125 = n10942 ;
  assign y6126 = 1'b0 ;
  assign y6127 = n10946 ;
  assign y6128 = ~n10948 ;
  assign y6129 = ~1'b0 ;
  assign y6130 = ~n10950 ;
  assign y6131 = ~1'b0 ;
  assign y6132 = n10951 ;
  assign y6133 = n10953 ;
  assign y6134 = ~1'b0 ;
  assign y6135 = ~1'b0 ;
  assign y6136 = ~1'b0 ;
  assign y6137 = ~n10954 ;
  assign y6138 = ~n10955 ;
  assign y6139 = ~n10957 ;
  assign y6140 = ~1'b0 ;
  assign y6141 = ~n10958 ;
  assign y6142 = ~n10960 ;
  assign y6143 = ~1'b0 ;
  assign y6144 = n10962 ;
  assign y6145 = ~1'b0 ;
  assign y6146 = ~n10965 ;
  assign y6147 = ~1'b0 ;
  assign y6148 = ~n10970 ;
  assign y6149 = 1'b0 ;
  assign y6150 = n10979 ;
  assign y6151 = ~1'b0 ;
  assign y6152 = n10980 ;
  assign y6153 = n10981 ;
  assign y6154 = ~1'b0 ;
  assign y6155 = ~n10983 ;
  assign y6156 = n10986 ;
  assign y6157 = ~n10988 ;
  assign y6158 = ~n10991 ;
  assign y6159 = n10994 ;
  assign y6160 = ~1'b0 ;
  assign y6161 = n10996 ;
  assign y6162 = ~1'b0 ;
  assign y6163 = ~x208 ;
  assign y6164 = ~n10999 ;
  assign y6165 = ~n11003 ;
  assign y6166 = 1'b0 ;
  assign y6167 = n11005 ;
  assign y6168 = n11010 ;
  assign y6169 = ~1'b0 ;
  assign y6170 = ~n8592 ;
  assign y6171 = ~1'b0 ;
  assign y6172 = n11016 ;
  assign y6173 = n11032 ;
  assign y6174 = ~1'b0 ;
  assign y6175 = ~1'b0 ;
  assign y6176 = ~1'b0 ;
  assign y6177 = ~n11036 ;
  assign y6178 = n11037 ;
  assign y6179 = ~n11038 ;
  assign y6180 = ~n11040 ;
  assign y6181 = ~n11045 ;
  assign y6182 = n11046 ;
  assign y6183 = ~n11048 ;
  assign y6184 = n11055 ;
  assign y6185 = ~n11058 ;
  assign y6186 = ~n11061 ;
  assign y6187 = 1'b0 ;
  assign y6188 = n11065 ;
  assign y6189 = ~1'b0 ;
  assign y6190 = ~1'b0 ;
  assign y6191 = ~1'b0 ;
  assign y6192 = ~n1514 ;
  assign y6193 = n11066 ;
  assign y6194 = n11068 ;
  assign y6195 = n11071 ;
  assign y6196 = n11073 ;
  assign y6197 = ~1'b0 ;
  assign y6198 = ~n11074 ;
  assign y6199 = n11077 ;
  assign y6200 = ~n11080 ;
  assign y6201 = n11081 ;
  assign y6202 = ~1'b0 ;
  assign y6203 = ~n11082 ;
  assign y6204 = ~1'b0 ;
  assign y6205 = ~n11087 ;
  assign y6206 = ~1'b0 ;
  assign y6207 = n11089 ;
  assign y6208 = n11091 ;
  assign y6209 = ~1'b0 ;
  assign y6210 = n11096 ;
  assign y6211 = ~1'b0 ;
  assign y6212 = 1'b0 ;
  assign y6213 = ~1'b0 ;
  assign y6214 = ~n11099 ;
  assign y6215 = n11104 ;
  assign y6216 = ~1'b0 ;
  assign y6217 = ~1'b0 ;
  assign y6218 = n11108 ;
  assign y6219 = n1562 ;
  assign y6220 = n11109 ;
  assign y6221 = n11113 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = ~1'b0 ;
  assign y6224 = ~n11116 ;
  assign y6225 = ~n11119 ;
  assign y6226 = ~1'b0 ;
  assign y6227 = ~1'b0 ;
  assign y6228 = ~1'b0 ;
  assign y6229 = ~n11120 ;
  assign y6230 = n11123 ;
  assign y6231 = ~n11125 ;
  assign y6232 = n11127 ;
  assign y6233 = ~1'b0 ;
  assign y6234 = ~1'b0 ;
  assign y6235 = ~x31 ;
  assign y6236 = ~n5988 ;
  assign y6237 = n11129 ;
  assign y6238 = n11131 ;
  assign y6239 = ~1'b0 ;
  assign y6240 = n6651 ;
  assign y6241 = ~1'b0 ;
  assign y6242 = n11136 ;
  assign y6243 = n11137 ;
  assign y6244 = ~n11139 ;
  assign y6245 = ~1'b0 ;
  assign y6246 = ~1'b0 ;
  assign y6247 = ~n11143 ;
  assign y6248 = ~n11148 ;
  assign y6249 = ~1'b0 ;
  assign y6250 = n3055 ;
  assign y6251 = n11149 ;
  assign y6252 = n11150 ;
  assign y6253 = ~1'b0 ;
  assign y6254 = ~1'b0 ;
  assign y6255 = n11154 ;
  assign y6256 = n5205 ;
  assign y6257 = n11158 ;
  assign y6258 = n11159 ;
  assign y6259 = ~1'b0 ;
  assign y6260 = 1'b0 ;
  assign y6261 = n11161 ;
  assign y6262 = ~n11162 ;
  assign y6263 = ~1'b0 ;
  assign y6264 = n11165 ;
  assign y6265 = ~1'b0 ;
  assign y6266 = ~1'b0 ;
  assign y6267 = ~n11166 ;
  assign y6268 = ~1'b0 ;
  assign y6269 = n11173 ;
  assign y6270 = n11176 ;
  assign y6271 = n11177 ;
  assign y6272 = n9386 ;
  assign y6273 = 1'b0 ;
  assign y6274 = ~1'b0 ;
  assign y6275 = ~n8506 ;
  assign y6276 = n11184 ;
  assign y6277 = ~n11187 ;
  assign y6278 = ~n11189 ;
  assign y6279 = ~1'b0 ;
  assign y6280 = n11191 ;
  assign y6281 = n11194 ;
  assign y6282 = n11196 ;
  assign y6283 = ~n11197 ;
  assign y6284 = ~1'b0 ;
  assign y6285 = n11199 ;
  assign y6286 = ~1'b0 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = ~1'b0 ;
  assign y6289 = n11205 ;
  assign y6290 = ~n11207 ;
  assign y6291 = n11211 ;
  assign y6292 = ~1'b0 ;
  assign y6293 = ~1'b0 ;
  assign y6294 = ~n11216 ;
  assign y6295 = ~1'b0 ;
  assign y6296 = ~1'b0 ;
  assign y6297 = ~1'b0 ;
  assign y6298 = ~1'b0 ;
  assign y6299 = ~1'b0 ;
  assign y6300 = ~n11219 ;
  assign y6301 = ~n11224 ;
  assign y6302 = n11231 ;
  assign y6303 = ~n11239 ;
  assign y6304 = ~1'b0 ;
  assign y6305 = n11240 ;
  assign y6306 = n11243 ;
  assign y6307 = ~1'b0 ;
  assign y6308 = n11245 ;
  assign y6309 = ~1'b0 ;
  assign y6310 = ~n11246 ;
  assign y6311 = ~n11247 ;
  assign y6312 = ~1'b0 ;
  assign y6313 = n11250 ;
  assign y6314 = n11252 ;
  assign y6315 = x26 ;
  assign y6316 = 1'b0 ;
  assign y6317 = ~n11254 ;
  assign y6318 = ~n11256 ;
  assign y6319 = n11264 ;
  assign y6320 = ~n5305 ;
  assign y6321 = ~1'b0 ;
  assign y6322 = n11268 ;
  assign y6323 = ~n11271 ;
  assign y6324 = ~n11272 ;
  assign y6325 = ~1'b0 ;
  assign y6326 = ~1'b0 ;
  assign y6327 = ~1'b0 ;
  assign y6328 = ~1'b0 ;
  assign y6329 = ~x76 ;
  assign y6330 = n11273 ;
  assign y6331 = ~1'b0 ;
  assign y6332 = 1'b0 ;
  assign y6333 = n11278 ;
  assign y6334 = ~1'b0 ;
  assign y6335 = ~1'b0 ;
  assign y6336 = ~n11282 ;
  assign y6337 = ~1'b0 ;
  assign y6338 = n11287 ;
  assign y6339 = ~1'b0 ;
  assign y6340 = ~1'b0 ;
  assign y6341 = ~n11293 ;
  assign y6342 = 1'b0 ;
  assign y6343 = n11304 ;
  assign y6344 = ~n11308 ;
  assign y6345 = ~n11310 ;
  assign y6346 = n11312 ;
  assign y6347 = ~n11319 ;
  assign y6348 = ~n11322 ;
  assign y6349 = n11323 ;
  assign y6350 = ~n11325 ;
  assign y6351 = ~1'b0 ;
  assign y6352 = ~1'b0 ;
  assign y6353 = ~1'b0 ;
  assign y6354 = ~1'b0 ;
  assign y6355 = ~n11328 ;
  assign y6356 = ~1'b0 ;
  assign y6357 = n11329 ;
  assign y6358 = ~1'b0 ;
  assign y6359 = n11332 ;
  assign y6360 = ~n11333 ;
  assign y6361 = n11335 ;
  assign y6362 = n11339 ;
  assign y6363 = ~n11342 ;
  assign y6364 = ~n11344 ;
  assign y6365 = ~n11345 ;
  assign y6366 = n11346 ;
  assign y6367 = ~1'b0 ;
  assign y6368 = 1'b0 ;
  assign y6369 = ~n11348 ;
  assign y6370 = ~n11350 ;
  assign y6371 = ~n6527 ;
  assign y6372 = ~1'b0 ;
  assign y6373 = ~1'b0 ;
  assign y6374 = ~n11355 ;
  assign y6375 = ~n11359 ;
  assign y6376 = ~n4930 ;
  assign y6377 = ~n11368 ;
  assign y6378 = n11370 ;
  assign y6379 = n6801 ;
  assign y6380 = n11373 ;
  assign y6381 = ~1'b0 ;
  assign y6382 = ~1'b0 ;
  assign y6383 = n11374 ;
  assign y6384 = ~1'b0 ;
  assign y6385 = n11376 ;
  assign y6386 = n11377 ;
  assign y6387 = ~1'b0 ;
  assign y6388 = ~1'b0 ;
  assign y6389 = ~1'b0 ;
  assign y6390 = n11378 ;
  assign y6391 = ~n5991 ;
  assign y6392 = ~1'b0 ;
  assign y6393 = n11380 ;
  assign y6394 = 1'b0 ;
  assign y6395 = ~n11381 ;
  assign y6396 = ~n5290 ;
  assign y6397 = ~n11382 ;
  assign y6398 = ~n11383 ;
  assign y6399 = ~1'b0 ;
  assign y6400 = ~1'b0 ;
  assign y6401 = ~n11388 ;
  assign y6402 = n8773 ;
  assign y6403 = ~n11390 ;
  assign y6404 = n11397 ;
  assign y6405 = ~1'b0 ;
  assign y6406 = ~1'b0 ;
  assign y6407 = n11398 ;
  assign y6408 = ~1'b0 ;
  assign y6409 = n11402 ;
  assign y6410 = 1'b0 ;
  assign y6411 = ~n11403 ;
  assign y6412 = ~n9560 ;
  assign y6413 = ~n11413 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = ~n11415 ;
  assign y6416 = ~1'b0 ;
  assign y6417 = ~n11421 ;
  assign y6418 = ~1'b0 ;
  assign y6419 = 1'b0 ;
  assign y6420 = ~1'b0 ;
  assign y6421 = ~1'b0 ;
  assign y6422 = ~1'b0 ;
  assign y6423 = ~n11427 ;
  assign y6424 = ~1'b0 ;
  assign y6425 = ~1'b0 ;
  assign y6426 = n11428 ;
  assign y6427 = ~1'b0 ;
  assign y6428 = ~n11429 ;
  assign y6429 = ~n6308 ;
  assign y6430 = ~n11432 ;
  assign y6431 = ~1'b0 ;
  assign y6432 = n11438 ;
  assign y6433 = ~n11441 ;
  assign y6434 = ~n2510 ;
  assign y6435 = ~n11442 ;
  assign y6436 = 1'b0 ;
  assign y6437 = n8816 ;
  assign y6438 = ~n11444 ;
  assign y6439 = n11445 ;
  assign y6440 = n11452 ;
  assign y6441 = n11453 ;
  assign y6442 = n11454 ;
  assign y6443 = n11455 ;
  assign y6444 = ~x81 ;
  assign y6445 = ~n11459 ;
  assign y6446 = n11461 ;
  assign y6447 = ~1'b0 ;
  assign y6448 = ~n11462 ;
  assign y6449 = ~1'b0 ;
  assign y6450 = ~1'b0 ;
  assign y6451 = n11463 ;
  assign y6452 = ~1'b0 ;
  assign y6453 = ~1'b0 ;
  assign y6454 = ~1'b0 ;
  assign y6455 = ~1'b0 ;
  assign y6456 = ~n6945 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = ~1'b0 ;
  assign y6459 = ~n11467 ;
  assign y6460 = ~n7832 ;
  assign y6461 = ~1'b0 ;
  assign y6462 = n11473 ;
  assign y6463 = ~1'b0 ;
  assign y6464 = n11474 ;
  assign y6465 = n11478 ;
  assign y6466 = n11479 ;
  assign y6467 = ~n11482 ;
  assign y6468 = ~1'b0 ;
  assign y6469 = n11484 ;
  assign y6470 = ~1'b0 ;
  assign y6471 = ~n11486 ;
  assign y6472 = ~n2145 ;
  assign y6473 = ~n11487 ;
  assign y6474 = n11488 ;
  assign y6475 = ~n11491 ;
  assign y6476 = ~n11492 ;
  assign y6477 = ~1'b0 ;
  assign y6478 = ~1'b0 ;
  assign y6479 = ~1'b0 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = ~n11494 ;
  assign y6482 = ~n11500 ;
  assign y6483 = n11504 ;
  assign y6484 = ~1'b0 ;
  assign y6485 = ~n11506 ;
  assign y6486 = ~n11507 ;
  assign y6487 = n11511 ;
  assign y6488 = ~n11512 ;
  assign y6489 = ~1'b0 ;
  assign y6490 = n9438 ;
  assign y6491 = n796 ;
  assign y6492 = ~1'b0 ;
  assign y6493 = ~1'b0 ;
  assign y6494 = n11517 ;
  assign y6495 = ~n11518 ;
  assign y6496 = ~1'b0 ;
  assign y6497 = ~n11520 ;
  assign y6498 = ~1'b0 ;
  assign y6499 = ~1'b0 ;
  assign y6500 = ~1'b0 ;
  assign y6501 = ~n11522 ;
  assign y6502 = ~1'b0 ;
  assign y6503 = ~n11524 ;
  assign y6504 = ~1'b0 ;
  assign y6505 = ~1'b0 ;
  assign y6506 = ~1'b0 ;
  assign y6507 = ~n11526 ;
  assign y6508 = n11528 ;
  assign y6509 = n11536 ;
  assign y6510 = n11544 ;
  assign y6511 = ~n11563 ;
  assign y6512 = n8387 ;
  assign y6513 = n11566 ;
  assign y6514 = n1111 ;
  assign y6515 = ~n11568 ;
  assign y6516 = ~n11571 ;
  assign y6517 = n3408 ;
  assign y6518 = ~1'b0 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = ~1'b0 ;
  assign y6521 = n11573 ;
  assign y6522 = n11574 ;
  assign y6523 = n11576 ;
  assign y6524 = ~1'b0 ;
  assign y6525 = ~n11577 ;
  assign y6526 = 1'b0 ;
  assign y6527 = ~n11580 ;
  assign y6528 = n11586 ;
  assign y6529 = ~n11595 ;
  assign y6530 = n11596 ;
  assign y6531 = n11599 ;
  assign y6532 = n11604 ;
  assign y6533 = ~n11610 ;
  assign y6534 = ~1'b0 ;
  assign y6535 = ~1'b0 ;
  assign y6536 = ~1'b0 ;
  assign y6537 = n11613 ;
  assign y6538 = ~n11614 ;
  assign y6539 = ~n11615 ;
  assign y6540 = ~1'b0 ;
  assign y6541 = n11621 ;
  assign y6542 = ~n11623 ;
  assign y6543 = n11626 ;
  assign y6544 = ~n11627 ;
  assign y6545 = 1'b0 ;
  assign y6546 = 1'b0 ;
  assign y6547 = ~1'b0 ;
  assign y6548 = ~1'b0 ;
  assign y6549 = ~n11632 ;
  assign y6550 = n11636 ;
  assign y6551 = n11642 ;
  assign y6552 = ~1'b0 ;
  assign y6553 = ~n11649 ;
  assign y6554 = ~1'b0 ;
  assign y6555 = ~1'b0 ;
  assign y6556 = n11651 ;
  assign y6557 = ~1'b0 ;
  assign y6558 = ~n11656 ;
  assign y6559 = ~n11658 ;
  assign y6560 = ~n11659 ;
  assign y6561 = ~n11661 ;
  assign y6562 = n11672 ;
  assign y6563 = n10188 ;
  assign y6564 = ~1'b0 ;
  assign y6565 = ~n11678 ;
  assign y6566 = n11680 ;
  assign y6567 = 1'b0 ;
  assign y6568 = ~1'b0 ;
  assign y6569 = ~n11682 ;
  assign y6570 = ~n11687 ;
  assign y6571 = ~1'b0 ;
  assign y6572 = n11694 ;
  assign y6573 = n11696 ;
  assign y6574 = ~n2425 ;
  assign y6575 = ~n5256 ;
  assign y6576 = ~1'b0 ;
  assign y6577 = ~n11697 ;
  assign y6578 = n11701 ;
  assign y6579 = n2909 ;
  assign y6580 = ~1'b0 ;
  assign y6581 = ~1'b0 ;
  assign y6582 = ~n11702 ;
  assign y6583 = ~1'b0 ;
  assign y6584 = ~n11704 ;
  assign y6585 = n11707 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = n11710 ;
  assign y6588 = ~n11711 ;
  assign y6589 = n11712 ;
  assign y6590 = ~n11714 ;
  assign y6591 = ~n8969 ;
  assign y6592 = n11716 ;
  assign y6593 = ~1'b0 ;
  assign y6594 = n11720 ;
  assign y6595 = n11723 ;
  assign y6596 = ~n11727 ;
  assign y6597 = n11729 ;
  assign y6598 = ~1'b0 ;
  assign y6599 = ~1'b0 ;
  assign y6600 = n11733 ;
  assign y6601 = ~1'b0 ;
  assign y6602 = ~1'b0 ;
  assign y6603 = ~1'b0 ;
  assign y6604 = n11734 ;
  assign y6605 = ~1'b0 ;
  assign y6606 = ~n11738 ;
  assign y6607 = n11740 ;
  assign y6608 = n11743 ;
  assign y6609 = ~n11744 ;
  assign y6610 = ~n11745 ;
  assign y6611 = ~n11746 ;
  assign y6612 = ~1'b0 ;
  assign y6613 = ~n11565 ;
  assign y6614 = ~n11749 ;
  assign y6615 = n11752 ;
  assign y6616 = ~x76 ;
  assign y6617 = n11754 ;
  assign y6618 = n11756 ;
  assign y6619 = n11757 ;
  assign y6620 = ~1'b0 ;
  assign y6621 = n11758 ;
  assign y6622 = ~n11760 ;
  assign y6623 = ~1'b0 ;
  assign y6624 = n11763 ;
  assign y6625 = ~1'b0 ;
  assign y6626 = n11766 ;
  assign y6627 = ~n11770 ;
  assign y6628 = ~n11771 ;
  assign y6629 = n6071 ;
  assign y6630 = n4485 ;
  assign y6631 = n1932 ;
  assign y6632 = n11773 ;
  assign y6633 = n4366 ;
  assign y6634 = ~n11774 ;
  assign y6635 = ~n11775 ;
  assign y6636 = n11777 ;
  assign y6637 = 1'b0 ;
  assign y6638 = n11778 ;
  assign y6639 = ~1'b0 ;
  assign y6640 = n11779 ;
  assign y6641 = n11780 ;
  assign y6642 = ~n11785 ;
  assign y6643 = ~n1580 ;
  assign y6644 = n11787 ;
  assign y6645 = n11789 ;
  assign y6646 = ~1'b0 ;
  assign y6647 = n11790 ;
  assign y6648 = n11793 ;
  assign y6649 = ~n11796 ;
  assign y6650 = n11800 ;
  assign y6651 = ~n11802 ;
  assign y6652 = ~n11804 ;
  assign y6653 = n1977 ;
  assign y6654 = n11808 ;
  assign y6655 = n11810 ;
  assign y6656 = ~1'b0 ;
  assign y6657 = 1'b0 ;
  assign y6658 = n11812 ;
  assign y6659 = ~n11817 ;
  assign y6660 = n11818 ;
  assign y6661 = ~n11819 ;
  assign y6662 = ~1'b0 ;
  assign y6663 = ~1'b0 ;
  assign y6664 = ~n11821 ;
  assign y6665 = ~n11845 ;
  assign y6666 = ~1'b0 ;
  assign y6667 = n11853 ;
  assign y6668 = n11854 ;
  assign y6669 = ~n11855 ;
  assign y6670 = ~1'b0 ;
  assign y6671 = ~n8314 ;
  assign y6672 = ~1'b0 ;
  assign y6673 = ~n11859 ;
  assign y6674 = n11864 ;
  assign y6675 = ~n11865 ;
  assign y6676 = ~1'b0 ;
  assign y6677 = ~n11866 ;
  assign y6678 = ~n11870 ;
  assign y6679 = 1'b0 ;
  assign y6680 = ~n11883 ;
  assign y6681 = ~n11884 ;
  assign y6682 = ~n5471 ;
  assign y6683 = ~n11885 ;
  assign y6684 = ~n11887 ;
  assign y6685 = ~1'b0 ;
  assign y6686 = ~1'b0 ;
  assign y6687 = ~1'b0 ;
  assign y6688 = n11888 ;
  assign y6689 = ~1'b0 ;
  assign y6690 = ~n6736 ;
  assign y6691 = n11890 ;
  assign y6692 = ~1'b0 ;
  assign y6693 = ~n11893 ;
  assign y6694 = n11894 ;
  assign y6695 = 1'b0 ;
  assign y6696 = ~1'b0 ;
  assign y6697 = n11897 ;
  assign y6698 = ~1'b0 ;
  assign y6699 = n11902 ;
  assign y6700 = n11903 ;
  assign y6701 = ~n11908 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = ~1'b0 ;
  assign y6704 = ~1'b0 ;
  assign y6705 = ~1'b0 ;
  assign y6706 = ~n11910 ;
  assign y6707 = n11911 ;
  assign y6708 = ~n11914 ;
  assign y6709 = ~1'b0 ;
  assign y6710 = 1'b0 ;
  assign y6711 = 1'b0 ;
  assign y6712 = n11919 ;
  assign y6713 = ~1'b0 ;
  assign y6714 = n11924 ;
  assign y6715 = ~n11927 ;
  assign y6716 = n11931 ;
  assign y6717 = ~n11932 ;
  assign y6718 = n11934 ;
  assign y6719 = n11935 ;
  assign y6720 = n11938 ;
  assign y6721 = ~n11940 ;
  assign y6722 = ~1'b0 ;
  assign y6723 = n11942 ;
  assign y6724 = n11944 ;
  assign y6725 = n11948 ;
  assign y6726 = n11949 ;
  assign y6727 = n11950 ;
  assign y6728 = ~n6110 ;
  assign y6729 = ~n11951 ;
  assign y6730 = ~1'b0 ;
  assign y6731 = ~n11952 ;
  assign y6732 = n11958 ;
  assign y6733 = ~n11960 ;
  assign y6734 = n11961 ;
  assign y6735 = n11963 ;
  assign y6736 = ~1'b0 ;
  assign y6737 = n11967 ;
  assign y6738 = ~1'b0 ;
  assign y6739 = ~n11968 ;
  assign y6740 = ~n3689 ;
  assign y6741 = ~1'b0 ;
  assign y6742 = n11971 ;
  assign y6743 = 1'b0 ;
  assign y6744 = n11973 ;
  assign y6745 = ~n10229 ;
  assign y6746 = ~n11974 ;
  assign y6747 = ~1'b0 ;
  assign y6748 = ~1'b0 ;
  assign y6749 = n6118 ;
  assign y6750 = ~n11977 ;
  assign y6751 = ~n11979 ;
  assign y6752 = ~n11981 ;
  assign y6753 = ~1'b0 ;
  assign y6754 = ~n11985 ;
  assign y6755 = n11987 ;
  assign y6756 = ~1'b0 ;
  assign y6757 = n11989 ;
  assign y6758 = ~1'b0 ;
  assign y6759 = ~1'b0 ;
  assign y6760 = n11990 ;
  assign y6761 = n11991 ;
  assign y6762 = ~n11992 ;
  assign y6763 = ~n11998 ;
  assign y6764 = n12000 ;
  assign y6765 = ~n12004 ;
  assign y6766 = ~n4079 ;
  assign y6767 = ~n12008 ;
  assign y6768 = ~n12012 ;
  assign y6769 = n12014 ;
  assign y6770 = n12015 ;
  assign y6771 = ~n12018 ;
  assign y6772 = ~n12019 ;
  assign y6773 = ~n12022 ;
  assign y6774 = ~n12023 ;
  assign y6775 = n12024 ;
  assign y6776 = ~n12025 ;
  assign y6777 = 1'b0 ;
  assign y6778 = ~1'b0 ;
  assign y6779 = ~n12026 ;
  assign y6780 = ~n12028 ;
  assign y6781 = n12031 ;
  assign y6782 = ~1'b0 ;
  assign y6783 = ~n12032 ;
  assign y6784 = ~1'b0 ;
  assign y6785 = ~1'b0 ;
  assign y6786 = n12036 ;
  assign y6787 = ~1'b0 ;
  assign y6788 = ~n12040 ;
  assign y6789 = ~1'b0 ;
  assign y6790 = ~n12041 ;
  assign y6791 = ~1'b0 ;
  assign y6792 = ~1'b0 ;
  assign y6793 = n12044 ;
  assign y6794 = n11623 ;
  assign y6795 = ~n12045 ;
  assign y6796 = n12046 ;
  assign y6797 = ~n12052 ;
  assign y6798 = ~1'b0 ;
  assign y6799 = n12054 ;
  assign y6800 = ~1'b0 ;
  assign y6801 = n12055 ;
  assign y6802 = ~n12056 ;
  assign y6803 = n12058 ;
  assign y6804 = n12061 ;
  assign y6805 = n5970 ;
  assign y6806 = ~1'b0 ;
  assign y6807 = ~n12062 ;
  assign y6808 = n12065 ;
  assign y6809 = n12066 ;
  assign y6810 = ~1'b0 ;
  assign y6811 = n12067 ;
  assign y6812 = n2382 ;
  assign y6813 = ~n12069 ;
  assign y6814 = n12071 ;
  assign y6815 = ~1'b0 ;
  assign y6816 = ~1'b0 ;
  assign y6817 = ~n12074 ;
  assign y6818 = n12075 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = ~1'b0 ;
  assign y6821 = n12080 ;
  assign y6822 = ~1'b0 ;
  assign y6823 = n12081 ;
  assign y6824 = n12082 ;
  assign y6825 = 1'b0 ;
  assign y6826 = 1'b0 ;
  assign y6827 = n12086 ;
  assign y6828 = ~n12088 ;
  assign y6829 = ~n12091 ;
  assign y6830 = ~n12094 ;
  assign y6831 = n12114 ;
  assign y6832 = n12115 ;
  assign y6833 = 1'b0 ;
  assign y6834 = ~1'b0 ;
  assign y6835 = n12118 ;
  assign y6836 = n7668 ;
  assign y6837 = ~1'b0 ;
  assign y6838 = n12120 ;
  assign y6839 = ~1'b0 ;
  assign y6840 = ~1'b0 ;
  assign y6841 = ~1'b0 ;
  assign y6842 = ~n12123 ;
  assign y6843 = n12124 ;
  assign y6844 = n12130 ;
  assign y6845 = ~1'b0 ;
  assign y6846 = n12132 ;
  assign y6847 = ~1'b0 ;
  assign y6848 = ~1'b0 ;
  assign y6849 = ~n12137 ;
  assign y6850 = ~1'b0 ;
  assign y6851 = ~n12138 ;
  assign y6852 = n12141 ;
  assign y6853 = ~n12144 ;
  assign y6854 = n12148 ;
  assign y6855 = n12149 ;
  assign y6856 = ~1'b0 ;
  assign y6857 = ~n12151 ;
  assign y6858 = ~n2716 ;
  assign y6859 = ~1'b0 ;
  assign y6860 = ~1'b0 ;
  assign y6861 = 1'b0 ;
  assign y6862 = ~1'b0 ;
  assign y6863 = n12152 ;
  assign y6864 = n12155 ;
  assign y6865 = n12162 ;
  assign y6866 = ~1'b0 ;
  assign y6867 = n12164 ;
  assign y6868 = ~n12167 ;
  assign y6869 = 1'b0 ;
  assign y6870 = ~n12169 ;
  assign y6871 = n12173 ;
  assign y6872 = n12174 ;
  assign y6873 = n12177 ;
  assign y6874 = ~1'b0 ;
  assign y6875 = ~1'b0 ;
  assign y6876 = ~n12178 ;
  assign y6877 = ~n4267 ;
  assign y6878 = n11148 ;
  assign y6879 = ~n12180 ;
  assign y6880 = ~1'b0 ;
  assign y6881 = n12182 ;
  assign y6882 = ~1'b0 ;
  assign y6883 = ~n5903 ;
  assign y6884 = 1'b0 ;
  assign y6885 = n12190 ;
  assign y6886 = ~1'b0 ;
  assign y6887 = n12192 ;
  assign y6888 = n12194 ;
  assign y6889 = 1'b0 ;
  assign y6890 = ~1'b0 ;
  assign y6891 = ~1'b0 ;
  assign y6892 = ~n12196 ;
  assign y6893 = ~n12199 ;
  assign y6894 = ~1'b0 ;
  assign y6895 = n12204 ;
  assign y6896 = ~n12205 ;
  assign y6897 = n12206 ;
  assign y6898 = ~1'b0 ;
  assign y6899 = ~n12208 ;
  assign y6900 = ~1'b0 ;
  assign y6901 = ~n12210 ;
  assign y6902 = ~n10068 ;
  assign y6903 = ~1'b0 ;
  assign y6904 = ~n12211 ;
  assign y6905 = ~1'b0 ;
  assign y6906 = ~1'b0 ;
  assign y6907 = n12213 ;
  assign y6908 = n12214 ;
  assign y6909 = ~n3308 ;
  assign y6910 = ~n12227 ;
  assign y6911 = ~1'b0 ;
  assign y6912 = ~n12237 ;
  assign y6913 = n12238 ;
  assign y6914 = ~1'b0 ;
  assign y6915 = ~n8384 ;
  assign y6916 = n12239 ;
  assign y6917 = n7559 ;
  assign y6918 = n1740 ;
  assign y6919 = ~1'b0 ;
  assign y6920 = ~1'b0 ;
  assign y6921 = ~1'b0 ;
  assign y6922 = ~1'b0 ;
  assign y6923 = n12243 ;
  assign y6924 = 1'b0 ;
  assign y6925 = ~n12248 ;
  assign y6926 = ~n12249 ;
  assign y6927 = n12251 ;
  assign y6928 = ~n12252 ;
  assign y6929 = ~1'b0 ;
  assign y6930 = ~n12253 ;
  assign y6931 = n12256 ;
  assign y6932 = ~1'b0 ;
  assign y6933 = ~1'b0 ;
  assign y6934 = ~n12257 ;
  assign y6935 = ~1'b0 ;
  assign y6936 = ~n12260 ;
  assign y6937 = ~1'b0 ;
  assign y6938 = n12262 ;
  assign y6939 = ~n12263 ;
  assign y6940 = ~1'b0 ;
  assign y6941 = ~1'b0 ;
  assign y6942 = n7271 ;
  assign y6943 = ~n12265 ;
  assign y6944 = ~1'b0 ;
  assign y6945 = 1'b0 ;
  assign y6946 = ~1'b0 ;
  assign y6947 = ~1'b0 ;
  assign y6948 = ~n12266 ;
  assign y6949 = n12268 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = 1'b0 ;
  assign y6952 = n5809 ;
  assign y6953 = ~n12269 ;
  assign y6954 = ~1'b0 ;
  assign y6955 = ~n12270 ;
  assign y6956 = n12272 ;
  assign y6957 = n12285 ;
  assign y6958 = ~1'b0 ;
  assign y6959 = n12288 ;
  assign y6960 = ~1'b0 ;
  assign y6961 = n12292 ;
  assign y6962 = n12293 ;
  assign y6963 = ~n8713 ;
  assign y6964 = n12295 ;
  assign y6965 = ~1'b0 ;
  assign y6966 = n12298 ;
  assign y6967 = n12299 ;
  assign y6968 = ~1'b0 ;
  assign y6969 = n12301 ;
  assign y6970 = ~1'b0 ;
  assign y6971 = ~1'b0 ;
  assign y6972 = ~n9781 ;
  assign y6973 = n12302 ;
  assign y6974 = n12305 ;
  assign y6975 = ~1'b0 ;
  assign y6976 = ~1'b0 ;
  assign y6977 = n10418 ;
  assign y6978 = ~1'b0 ;
  assign y6979 = n12306 ;
  assign y6980 = 1'b0 ;
  assign y6981 = ~n12307 ;
  assign y6982 = 1'b0 ;
  assign y6983 = ~n12309 ;
  assign y6984 = ~n12310 ;
  assign y6985 = n7671 ;
  assign y6986 = 1'b0 ;
  assign y6987 = ~n10150 ;
  assign y6988 = n12311 ;
  assign y6989 = ~n12316 ;
  assign y6990 = ~n12317 ;
  assign y6991 = ~1'b0 ;
  assign y6992 = ~n12326 ;
  assign y6993 = ~n12327 ;
  assign y6994 = ~1'b0 ;
  assign y6995 = ~1'b0 ;
  assign y6996 = n12330 ;
  assign y6997 = ~n12331 ;
  assign y6998 = n9034 ;
  assign y6999 = ~n12332 ;
  assign y7000 = 1'b0 ;
  assign y7001 = ~1'b0 ;
  assign y7002 = ~n12338 ;
  assign y7003 = n12340 ;
  assign y7004 = ~n4238 ;
  assign y7005 = ~n12343 ;
  assign y7006 = ~1'b0 ;
  assign y7007 = n4172 ;
  assign y7008 = ~n12345 ;
  assign y7009 = ~1'b0 ;
  assign y7010 = ~1'b0 ;
  assign y7011 = ~n12346 ;
  assign y7012 = ~1'b0 ;
  assign y7013 = n12352 ;
  assign y7014 = 1'b0 ;
  assign y7015 = n4122 ;
  assign y7016 = n12355 ;
  assign y7017 = n12356 ;
  assign y7018 = ~n12365 ;
  assign y7019 = n12370 ;
  assign y7020 = ~n3255 ;
  assign y7021 = n12374 ;
  assign y7022 = ~1'b0 ;
  assign y7023 = n12377 ;
  assign y7024 = n12380 ;
  assign y7025 = n12381 ;
  assign y7026 = ~1'b0 ;
  assign y7027 = ~1'b0 ;
  assign y7028 = n12383 ;
  assign y7029 = n12387 ;
  assign y7030 = ~n12390 ;
  assign y7031 = ~1'b0 ;
  assign y7032 = ~1'b0 ;
  assign y7033 = ~n12393 ;
  assign y7034 = ~1'b0 ;
  assign y7035 = ~1'b0 ;
  assign y7036 = ~1'b0 ;
  assign y7037 = 1'b0 ;
  assign y7038 = ~1'b0 ;
  assign y7039 = ~1'b0 ;
  assign y7040 = n12394 ;
  assign y7041 = ~n6964 ;
  assign y7042 = ~1'b0 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = 1'b0 ;
  assign y7045 = ~1'b0 ;
  assign y7046 = ~1'b0 ;
  assign y7047 = ~n12396 ;
  assign y7048 = ~1'b0 ;
  assign y7049 = ~1'b0 ;
  assign y7050 = 1'b0 ;
  assign y7051 = ~1'b0 ;
  assign y7052 = ~1'b0 ;
  assign y7053 = n12398 ;
  assign y7054 = ~n12400 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = ~n12404 ;
  assign y7057 = n12408 ;
  assign y7058 = 1'b0 ;
  assign y7059 = ~1'b0 ;
  assign y7060 = ~1'b0 ;
  assign y7061 = ~n12419 ;
  assign y7062 = ~1'b0 ;
  assign y7063 = ~n12421 ;
  assign y7064 = ~1'b0 ;
  assign y7065 = ~1'b0 ;
  assign y7066 = ~1'b0 ;
  assign y7067 = ~1'b0 ;
  assign y7068 = ~n12436 ;
  assign y7069 = n12438 ;
  assign y7070 = n12444 ;
  assign y7071 = n2486 ;
  assign y7072 = ~n12445 ;
  assign y7073 = ~n12447 ;
  assign y7074 = ~1'b0 ;
  assign y7075 = n6025 ;
  assign y7076 = n12448 ;
  assign y7077 = n12452 ;
  assign y7078 = ~1'b0 ;
  assign y7079 = ~1'b0 ;
  assign y7080 = ~1'b0 ;
  assign y7081 = x144 ;
  assign y7082 = ~1'b0 ;
  assign y7083 = ~n12455 ;
  assign y7084 = ~1'b0 ;
  assign y7085 = ~1'b0 ;
  assign y7086 = ~1'b0 ;
  assign y7087 = ~1'b0 ;
  assign y7088 = ~n12456 ;
  assign y7089 = ~1'b0 ;
  assign y7090 = ~1'b0 ;
  assign y7091 = ~n12458 ;
  assign y7092 = ~n12460 ;
  assign y7093 = ~1'b0 ;
  assign y7094 = ~1'b0 ;
  assign y7095 = ~n12461 ;
  assign y7096 = ~1'b0 ;
  assign y7097 = ~n3872 ;
  assign y7098 = ~n12468 ;
  assign y7099 = n12471 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = ~n12473 ;
  assign y7102 = ~n12475 ;
  assign y7103 = n9864 ;
  assign y7104 = n12478 ;
  assign y7105 = ~n2801 ;
  assign y7106 = ~n12154 ;
  assign y7107 = n12479 ;
  assign y7108 = n12492 ;
  assign y7109 = ~1'b0 ;
  assign y7110 = ~1'b0 ;
  assign y7111 = ~1'b0 ;
  assign y7112 = ~n12495 ;
  assign y7113 = n12496 ;
  assign y7114 = ~n12498 ;
  assign y7115 = ~n12500 ;
  assign y7116 = n12502 ;
  assign y7117 = n12505 ;
  assign y7118 = ~1'b0 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = ~n12506 ;
  assign y7121 = ~n12508 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = ~n12512 ;
  assign y7124 = ~n1104 ;
  assign y7125 = ~n12519 ;
  assign y7126 = ~1'b0 ;
  assign y7127 = n12520 ;
  assign y7128 = ~1'b0 ;
  assign y7129 = ~1'b0 ;
  assign y7130 = n12521 ;
  assign y7131 = ~1'b0 ;
  assign y7132 = ~1'b0 ;
  assign y7133 = ~n12522 ;
  assign y7134 = n12524 ;
  assign y7135 = ~n12525 ;
  assign y7136 = n12526 ;
  assign y7137 = ~n9022 ;
  assign y7138 = n12533 ;
  assign y7139 = ~n12536 ;
  assign y7140 = ~n12539 ;
  assign y7141 = ~1'b0 ;
  assign y7142 = n12541 ;
  assign y7143 = ~1'b0 ;
  assign y7144 = ~n12550 ;
  assign y7145 = n12554 ;
  assign y7146 = n12555 ;
  assign y7147 = ~n12556 ;
  assign y7148 = n12561 ;
  assign y7149 = ~n12562 ;
  assign y7150 = n12563 ;
  assign y7151 = n12565 ;
  assign y7152 = ~n12569 ;
  assign y7153 = n12570 ;
  assign y7154 = n12574 ;
  assign y7155 = ~n5676 ;
  assign y7156 = ~1'b0 ;
  assign y7157 = ~1'b0 ;
  assign y7158 = ~n9454 ;
  assign y7159 = ~1'b0 ;
  assign y7160 = ~n12575 ;
  assign y7161 = ~1'b0 ;
  assign y7162 = n12577 ;
  assign y7163 = n12578 ;
  assign y7164 = ~1'b0 ;
  assign y7165 = ~1'b0 ;
  assign y7166 = ~1'b0 ;
  assign y7167 = n12579 ;
  assign y7168 = n12581 ;
  assign y7169 = n12582 ;
  assign y7170 = ~n12584 ;
  assign y7171 = ~1'b0 ;
  assign y7172 = n12585 ;
  assign y7173 = 1'b0 ;
  assign y7174 = ~1'b0 ;
  assign y7175 = n12588 ;
  assign y7176 = n12596 ;
  assign y7177 = ~1'b0 ;
  assign y7178 = ~n12598 ;
  assign y7179 = ~n12600 ;
  assign y7180 = ~1'b0 ;
  assign y7181 = n12605 ;
  assign y7182 = ~1'b0 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = n12610 ;
  assign y7185 = ~1'b0 ;
  assign y7186 = ~1'b0 ;
  assign y7187 = n12611 ;
  assign y7188 = ~n12612 ;
  assign y7189 = ~1'b0 ;
  assign y7190 = n12613 ;
  assign y7191 = n12614 ;
  assign y7192 = n2221 ;
  assign y7193 = ~1'b0 ;
  assign y7194 = x78 ;
  assign y7195 = ~1'b0 ;
  assign y7196 = n8475 ;
  assign y7197 = ~n12615 ;
  assign y7198 = n12617 ;
  assign y7199 = n12618 ;
  assign y7200 = n10164 ;
  assign y7201 = ~1'b0 ;
  assign y7202 = ~1'b0 ;
  assign y7203 = ~n8881 ;
  assign y7204 = ~n12623 ;
  assign y7205 = ~n12627 ;
  assign y7206 = ~1'b0 ;
  assign y7207 = ~n12629 ;
  assign y7208 = n6997 ;
  assign y7209 = 1'b0 ;
  assign y7210 = ~1'b0 ;
  assign y7211 = n12631 ;
  assign y7212 = 1'b0 ;
  assign y7213 = ~1'b0 ;
  assign y7214 = n6207 ;
  assign y7215 = ~1'b0 ;
  assign y7216 = ~n12636 ;
  assign y7217 = n12650 ;
  assign y7218 = n12654 ;
  assign y7219 = ~1'b0 ;
  assign y7220 = ~1'b0 ;
  assign y7221 = n12655 ;
  assign y7222 = ~1'b0 ;
  assign y7223 = n12657 ;
  assign y7224 = ~1'b0 ;
  assign y7225 = ~n12660 ;
  assign y7226 = ~n3286 ;
  assign y7227 = ~1'b0 ;
  assign y7228 = ~n12665 ;
  assign y7229 = n12667 ;
  assign y7230 = ~n12668 ;
  assign y7231 = n4402 ;
  assign y7232 = ~x182 ;
  assign y7233 = n12678 ;
  assign y7234 = 1'b0 ;
  assign y7235 = n12680 ;
  assign y7236 = ~1'b0 ;
  assign y7237 = ~n12682 ;
  assign y7238 = n12684 ;
  assign y7239 = ~n12685 ;
  assign y7240 = n12689 ;
  assign y7241 = ~n12690 ;
  assign y7242 = n12700 ;
  assign y7243 = ~1'b0 ;
  assign y7244 = n12702 ;
  assign y7245 = n12703 ;
  assign y7246 = ~n12704 ;
  assign y7247 = ~n8849 ;
  assign y7248 = 1'b0 ;
  assign y7249 = n12705 ;
  assign y7250 = 1'b0 ;
  assign y7251 = ~n12707 ;
  assign y7252 = n12710 ;
  assign y7253 = ~1'b0 ;
  assign y7254 = ~n12720 ;
  assign y7255 = ~n12723 ;
  assign y7256 = ~n12725 ;
  assign y7257 = n12732 ;
  assign y7258 = ~1'b0 ;
  assign y7259 = n12733 ;
  assign y7260 = ~1'b0 ;
  assign y7261 = ~n12735 ;
  assign y7262 = ~1'b0 ;
  assign y7263 = ~1'b0 ;
  assign y7264 = ~n12736 ;
  assign y7265 = n12737 ;
  assign y7266 = ~1'b0 ;
  assign y7267 = 1'b0 ;
  assign y7268 = n12739 ;
  assign y7269 = ~n12741 ;
  assign y7270 = ~1'b0 ;
  assign y7271 = n12748 ;
  assign y7272 = n607 ;
  assign y7273 = ~n12749 ;
  assign y7274 = n12756 ;
  assign y7275 = ~1'b0 ;
  assign y7276 = n8033 ;
  assign y7277 = ~n12760 ;
  assign y7278 = ~1'b0 ;
  assign y7279 = ~n3390 ;
  assign y7280 = ~n12766 ;
  assign y7281 = ~n12768 ;
  assign y7282 = n12770 ;
  assign y7283 = n4204 ;
  assign y7284 = ~1'b0 ;
  assign y7285 = n12772 ;
  assign y7286 = n12773 ;
  assign y7287 = ~n12775 ;
  assign y7288 = n12780 ;
  assign y7289 = n12781 ;
  assign y7290 = ~1'b0 ;
  assign y7291 = ~1'b0 ;
  assign y7292 = n12783 ;
  assign y7293 = ~n12784 ;
  assign y7294 = n12787 ;
  assign y7295 = ~1'b0 ;
  assign y7296 = ~1'b0 ;
  assign y7297 = n12788 ;
  assign y7298 = n12789 ;
  assign y7299 = n12791 ;
  assign y7300 = n12792 ;
  assign y7301 = ~1'b0 ;
  assign y7302 = ~1'b0 ;
  assign y7303 = n12798 ;
  assign y7304 = ~1'b0 ;
  assign y7305 = n12799 ;
  assign y7306 = n12800 ;
  assign y7307 = n12804 ;
  assign y7308 = n12805 ;
  assign y7309 = ~n12815 ;
  assign y7310 = ~n12818 ;
  assign y7311 = ~1'b0 ;
  assign y7312 = 1'b0 ;
  assign y7313 = ~1'b0 ;
  assign y7314 = ~n7865 ;
  assign y7315 = ~1'b0 ;
  assign y7316 = ~n12820 ;
  assign y7317 = ~n12821 ;
  assign y7318 = ~1'b0 ;
  assign y7319 = n3740 ;
  assign y7320 = ~1'b0 ;
  assign y7321 = n12827 ;
  assign y7322 = n12831 ;
  assign y7323 = ~n12837 ;
  assign y7324 = ~1'b0 ;
  assign y7325 = ~n12839 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = 1'b0 ;
  assign y7328 = ~n12845 ;
  assign y7329 = n12848 ;
  assign y7330 = ~x153 ;
  assign y7331 = n12850 ;
  assign y7332 = ~1'b0 ;
  assign y7333 = n12852 ;
  assign y7334 = ~n12857 ;
  assign y7335 = ~1'b0 ;
  assign y7336 = ~n6178 ;
  assign y7337 = ~n12859 ;
  assign y7338 = n2589 ;
  assign y7339 = n12861 ;
  assign y7340 = ~n12863 ;
  assign y7341 = n12616 ;
  assign y7342 = n12865 ;
  assign y7343 = n12868 ;
  assign y7344 = ~n12872 ;
  assign y7345 = n9652 ;
  assign y7346 = ~1'b0 ;
  assign y7347 = ~1'b0 ;
  assign y7348 = n12874 ;
  assign y7349 = ~n472 ;
  assign y7350 = ~n12877 ;
  assign y7351 = ~n12878 ;
  assign y7352 = ~1'b0 ;
  assign y7353 = ~n12884 ;
  assign y7354 = ~n12885 ;
  assign y7355 = ~1'b0 ;
  assign y7356 = ~1'b0 ;
  assign y7357 = n12891 ;
  assign y7358 = n12892 ;
  assign y7359 = ~1'b0 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = ~1'b0 ;
  assign y7362 = n12896 ;
  assign y7363 = ~n12898 ;
  assign y7364 = ~n12900 ;
  assign y7365 = ~n12903 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = ~1'b0 ;
  assign y7368 = n12905 ;
  assign y7369 = ~n12906 ;
  assign y7370 = n3606 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = ~1'b0 ;
  assign y7373 = n2482 ;
  assign y7374 = ~1'b0 ;
  assign y7375 = ~n12908 ;
  assign y7376 = n12911 ;
  assign y7377 = n12914 ;
  assign y7378 = ~n12915 ;
  assign y7379 = ~1'b0 ;
  assign y7380 = n11704 ;
  assign y7381 = ~n12917 ;
  assign y7382 = ~1'b0 ;
  assign y7383 = n12922 ;
  assign y7384 = n12923 ;
  assign y7385 = ~n12924 ;
  assign y7386 = n12931 ;
  assign y7387 = ~1'b0 ;
  assign y7388 = ~1'b0 ;
  assign y7389 = n12933 ;
  assign y7390 = ~n10715 ;
  assign y7391 = ~1'b0 ;
  assign y7392 = ~1'b0 ;
  assign y7393 = ~1'b0 ;
  assign y7394 = ~1'b0 ;
  assign y7395 = n12934 ;
  assign y7396 = n12941 ;
  assign y7397 = ~1'b0 ;
  assign y7398 = ~1'b0 ;
  assign y7399 = n12949 ;
  assign y7400 = ~n12950 ;
  assign y7401 = ~1'b0 ;
  assign y7402 = ~n2725 ;
  assign y7403 = ~n12952 ;
  assign y7404 = ~1'b0 ;
  assign y7405 = ~n12954 ;
  assign y7406 = ~1'b0 ;
  assign y7407 = n12955 ;
  assign y7408 = ~n12956 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = n12957 ;
  assign y7411 = n12959 ;
  assign y7412 = n12967 ;
  assign y7413 = ~1'b0 ;
  assign y7414 = ~n12969 ;
  assign y7415 = ~1'b0 ;
  assign y7416 = n12973 ;
  assign y7417 = n12974 ;
  assign y7418 = ~1'b0 ;
  assign y7419 = ~1'b0 ;
  assign y7420 = n12979 ;
  assign y7421 = ~1'b0 ;
  assign y7422 = ~n12980 ;
  assign y7423 = 1'b0 ;
  assign y7424 = n12981 ;
  assign y7425 = ~n12983 ;
  assign y7426 = ~n12985 ;
  assign y7427 = ~1'b0 ;
  assign y7428 = ~1'b0 ;
  assign y7429 = n12986 ;
  assign y7430 = n6792 ;
  assign y7431 = ~1'b0 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = ~1'b0 ;
  assign y7434 = ~1'b0 ;
  assign y7435 = ~1'b0 ;
  assign y7436 = ~1'b0 ;
  assign y7437 = ~n12989 ;
  assign y7438 = ~1'b0 ;
  assign y7439 = ~n12995 ;
  assign y7440 = ~n10018 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = ~1'b0 ;
  assign y7443 = n12998 ;
  assign y7444 = ~n13000 ;
  assign y7445 = n13003 ;
  assign y7446 = ~1'b0 ;
  assign y7447 = n13005 ;
  assign y7448 = n13019 ;
  assign y7449 = ~n13020 ;
  assign y7450 = n13022 ;
  assign y7451 = ~n13025 ;
  assign y7452 = ~n13033 ;
  assign y7453 = ~1'b0 ;
  assign y7454 = ~1'b0 ;
  assign y7455 = n13036 ;
  assign y7456 = ~1'b0 ;
  assign y7457 = ~n13042 ;
  assign y7458 = ~n13047 ;
  assign y7459 = ~n13048 ;
  assign y7460 = ~1'b0 ;
  assign y7461 = n13049 ;
  assign y7462 = n8237 ;
  assign y7463 = 1'b0 ;
  assign y7464 = n13053 ;
  assign y7465 = n13057 ;
  assign y7466 = n13064 ;
  assign y7467 = n13069 ;
  assign y7468 = n13070 ;
  assign y7469 = ~n13075 ;
  assign y7470 = ~n13078 ;
  assign y7471 = ~n13080 ;
  assign y7472 = ~1'b0 ;
  assign y7473 = ~1'b0 ;
  assign y7474 = n13081 ;
  assign y7475 = ~1'b0 ;
  assign y7476 = ~1'b0 ;
  assign y7477 = n13086 ;
  assign y7478 = ~1'b0 ;
  assign y7479 = ~n13087 ;
  assign y7480 = 1'b0 ;
  assign y7481 = n13088 ;
  assign y7482 = ~1'b0 ;
  assign y7483 = ~n11486 ;
  assign y7484 = n13089 ;
  assign y7485 = ~n13091 ;
  assign y7486 = ~1'b0 ;
  assign y7487 = ~1'b0 ;
  assign y7488 = n13092 ;
  assign y7489 = n13093 ;
  assign y7490 = n13095 ;
  assign y7491 = n13096 ;
  assign y7492 = ~1'b0 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = ~1'b0 ;
  assign y7495 = n13100 ;
  assign y7496 = n13109 ;
  assign y7497 = ~n9083 ;
  assign y7498 = n13110 ;
  assign y7499 = ~n13111 ;
  assign y7500 = n13118 ;
  assign y7501 = ~1'b0 ;
  assign y7502 = ~1'b0 ;
  assign y7503 = ~n13124 ;
  assign y7504 = ~n13125 ;
  assign y7505 = n13140 ;
  assign y7506 = ~n13142 ;
  assign y7507 = ~1'b0 ;
  assign y7508 = ~1'b0 ;
  assign y7509 = ~1'b0 ;
  assign y7510 = ~1'b0 ;
  assign y7511 = n11207 ;
  assign y7512 = n13144 ;
  assign y7513 = ~1'b0 ;
  assign y7514 = ~n13151 ;
  assign y7515 = ~1'b0 ;
  assign y7516 = ~n13152 ;
  assign y7517 = ~1'b0 ;
  assign y7518 = n13155 ;
  assign y7519 = ~1'b0 ;
  assign y7520 = n13160 ;
  assign y7521 = ~n3678 ;
  assign y7522 = ~1'b0 ;
  assign y7523 = ~1'b0 ;
  assign y7524 = ~n13163 ;
  assign y7525 = ~n13171 ;
  assign y7526 = ~1'b0 ;
  assign y7527 = ~1'b0 ;
  assign y7528 = n13172 ;
  assign y7529 = ~1'b0 ;
  assign y7530 = n13175 ;
  assign y7531 = ~n13177 ;
  assign y7532 = n13178 ;
  assign y7533 = ~1'b0 ;
  assign y7534 = ~n13179 ;
  assign y7535 = ~1'b0 ;
  assign y7536 = ~n13180 ;
  assign y7537 = ~n13182 ;
  assign y7538 = ~1'b0 ;
  assign y7539 = n13184 ;
  assign y7540 = ~n13190 ;
  assign y7541 = ~n13195 ;
  assign y7542 = ~1'b0 ;
  assign y7543 = n13201 ;
  assign y7544 = ~1'b0 ;
  assign y7545 = ~1'b0 ;
  assign y7546 = ~n13203 ;
  assign y7547 = ~1'b0 ;
  assign y7548 = ~n13205 ;
  assign y7549 = ~1'b0 ;
  assign y7550 = ~1'b0 ;
  assign y7551 = ~n13209 ;
  assign y7552 = n13210 ;
  assign y7553 = n13218 ;
  assign y7554 = ~1'b0 ;
  assign y7555 = ~1'b0 ;
  assign y7556 = n13222 ;
  assign y7557 = n13223 ;
  assign y7558 = n13226 ;
  assign y7559 = n13228 ;
  assign y7560 = ~1'b0 ;
  assign y7561 = n13234 ;
  assign y7562 = n13239 ;
  assign y7563 = ~n13241 ;
  assign y7564 = 1'b0 ;
  assign y7565 = n13243 ;
  assign y7566 = ~n13250 ;
  assign y7567 = ~n13258 ;
  assign y7568 = ~n13260 ;
  assign y7569 = ~1'b0 ;
  assign y7570 = ~1'b0 ;
  assign y7571 = ~1'b0 ;
  assign y7572 = ~1'b0 ;
  assign y7573 = n13261 ;
  assign y7574 = n13262 ;
  assign y7575 = ~n13264 ;
  assign y7576 = ~1'b0 ;
  assign y7577 = 1'b0 ;
  assign y7578 = n13266 ;
  assign y7579 = n11329 ;
  assign y7580 = n5262 ;
  assign y7581 = n13268 ;
  assign y7582 = n13270 ;
  assign y7583 = ~n13271 ;
  assign y7584 = ~n13280 ;
  assign y7585 = 1'b0 ;
  assign y7586 = 1'b0 ;
  assign y7587 = n13283 ;
  assign y7588 = ~n13288 ;
  assign y7589 = ~1'b0 ;
  assign y7590 = ~n13294 ;
  assign y7591 = n13295 ;
  assign y7592 = n13296 ;
  assign y7593 = n12159 ;
  assign y7594 = ~1'b0 ;
  assign y7595 = ~1'b0 ;
  assign y7596 = ~n13302 ;
  assign y7597 = ~1'b0 ;
  assign y7598 = ~1'b0 ;
  assign y7599 = ~n13305 ;
  assign y7600 = ~n13306 ;
  assign y7601 = n13310 ;
  assign y7602 = n13311 ;
  assign y7603 = ~1'b0 ;
  assign y7604 = ~n13314 ;
  assign y7605 = n13315 ;
  assign y7606 = ~1'b0 ;
  assign y7607 = ~1'b0 ;
  assign y7608 = ~n13321 ;
  assign y7609 = ~n13323 ;
  assign y7610 = ~n13324 ;
  assign y7611 = ~n13325 ;
  assign y7612 = ~1'b0 ;
  assign y7613 = ~n13326 ;
  assign y7614 = 1'b0 ;
  assign y7615 = n13279 ;
  assign y7616 = ~1'b0 ;
  assign y7617 = n988 ;
  assign y7618 = ~1'b0 ;
  assign y7619 = ~1'b0 ;
  assign y7620 = ~n1514 ;
  assign y7621 = n13327 ;
  assign y7622 = ~n13329 ;
  assign y7623 = ~1'b0 ;
  assign y7624 = n13331 ;
  assign y7625 = 1'b0 ;
  assign y7626 = ~n13341 ;
  assign y7627 = n13346 ;
  assign y7628 = n13348 ;
  assign y7629 = ~1'b0 ;
  assign y7630 = ~1'b0 ;
  assign y7631 = ~n5564 ;
  assign y7632 = n13350 ;
  assign y7633 = ~1'b0 ;
  assign y7634 = ~1'b0 ;
  assign y7635 = ~n13355 ;
  assign y7636 = n13356 ;
  assign y7637 = n13358 ;
  assign y7638 = n13368 ;
  assign y7639 = ~1'b0 ;
  assign y7640 = 1'b0 ;
  assign y7641 = n13369 ;
  assign y7642 = n13370 ;
  assign y7643 = n3599 ;
  assign y7644 = ~n13379 ;
  assign y7645 = ~n13380 ;
  assign y7646 = n13383 ;
  assign y7647 = ~n13385 ;
  assign y7648 = ~n13387 ;
  assign y7649 = ~n13389 ;
  assign y7650 = ~n13391 ;
  assign y7651 = n13394 ;
  assign y7652 = n13396 ;
  assign y7653 = ~1'b0 ;
  assign y7654 = n13397 ;
  assign y7655 = ~1'b0 ;
  assign y7656 = ~n13405 ;
  assign y7657 = n5364 ;
  assign y7658 = ~1'b0 ;
  assign y7659 = ~n13410 ;
  assign y7660 = ~1'b0 ;
  assign y7661 = ~n2293 ;
  assign y7662 = ~1'b0 ;
  assign y7663 = n13411 ;
  assign y7664 = ~1'b0 ;
  assign y7665 = n13413 ;
  assign y7666 = ~1'b0 ;
  assign y7667 = ~n13416 ;
  assign y7668 = ~1'b0 ;
  assign y7669 = ~n13418 ;
  assign y7670 = n13422 ;
  assign y7671 = ~1'b0 ;
  assign y7672 = ~n13430 ;
  assign y7673 = ~n13433 ;
  assign y7674 = ~n13434 ;
  assign y7675 = ~1'b0 ;
  assign y7676 = ~n13437 ;
  assign y7677 = ~1'b0 ;
  assign y7678 = n1435 ;
  assign y7679 = n13443 ;
  assign y7680 = n13446 ;
  assign y7681 = ~1'b0 ;
  assign y7682 = ~n7440 ;
  assign y7683 = ~1'b0 ;
  assign y7684 = ~n13451 ;
  assign y7685 = ~n13452 ;
  assign y7686 = ~n13453 ;
  assign y7687 = ~1'b0 ;
  assign y7688 = ~n13460 ;
  assign y7689 = n13467 ;
  assign y7690 = ~1'b0 ;
  assign y7691 = n13472 ;
  assign y7692 = ~n13473 ;
  assign y7693 = ~n13476 ;
  assign y7694 = n13479 ;
  assign y7695 = ~1'b0 ;
  assign y7696 = ~n13481 ;
  assign y7697 = ~n13485 ;
  assign y7698 = ~n13486 ;
  assign y7699 = n13487 ;
  assign y7700 = n13492 ;
  assign y7701 = ~1'b0 ;
  assign y7702 = 1'b0 ;
  assign y7703 = ~1'b0 ;
  assign y7704 = ~1'b0 ;
  assign y7705 = ~1'b0 ;
  assign y7706 = n13493 ;
  assign y7707 = ~n13495 ;
  assign y7708 = n13499 ;
  assign y7709 = ~1'b0 ;
  assign y7710 = n13500 ;
  assign y7711 = ~1'b0 ;
  assign y7712 = ~1'b0 ;
  assign y7713 = ~1'b0 ;
  assign y7714 = n13501 ;
  assign y7715 = ~n13506 ;
  assign y7716 = ~n13508 ;
  assign y7717 = ~n13511 ;
  assign y7718 = ~n13515 ;
  assign y7719 = ~n13523 ;
  assign y7720 = n13530 ;
  assign y7721 = n6953 ;
  assign y7722 = n13532 ;
  assign y7723 = ~n13535 ;
  assign y7724 = n13538 ;
  assign y7725 = n13540 ;
  assign y7726 = n13543 ;
  assign y7727 = ~n13544 ;
  assign y7728 = ~n13548 ;
  assign y7729 = 1'b0 ;
  assign y7730 = ~n13559 ;
  assign y7731 = n12714 ;
  assign y7732 = n7362 ;
  assign y7733 = ~n13560 ;
  assign y7734 = n13561 ;
  assign y7735 = ~n13562 ;
  assign y7736 = ~1'b0 ;
  assign y7737 = n3879 ;
  assign y7738 = ~1'b0 ;
  assign y7739 = ~n13565 ;
  assign y7740 = ~1'b0 ;
  assign y7741 = ~n13574 ;
  assign y7742 = n13576 ;
  assign y7743 = n13578 ;
  assign y7744 = n4398 ;
  assign y7745 = n12560 ;
  assign y7746 = ~1'b0 ;
  assign y7747 = n13580 ;
  assign y7748 = ~n4230 ;
  assign y7749 = ~1'b0 ;
  assign y7750 = n13590 ;
  assign y7751 = n13595 ;
  assign y7752 = ~1'b0 ;
  assign y7753 = ~1'b0 ;
  assign y7754 = n3376 ;
  assign y7755 = ~n13597 ;
  assign y7756 = ~1'b0 ;
  assign y7757 = ~1'b0 ;
  assign y7758 = n13601 ;
  assign y7759 = ~1'b0 ;
  assign y7760 = n8290 ;
  assign y7761 = ~n13609 ;
  assign y7762 = ~n13610 ;
  assign y7763 = ~n13612 ;
  assign y7764 = ~1'b0 ;
  assign y7765 = n13613 ;
  assign y7766 = 1'b0 ;
  assign y7767 = n13614 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = ~n13616 ;
  assign y7770 = ~1'b0 ;
  assign y7771 = ~1'b0 ;
  assign y7772 = ~n13625 ;
  assign y7773 = ~1'b0 ;
  assign y7774 = ~1'b0 ;
  assign y7775 = n13627 ;
  assign y7776 = ~1'b0 ;
  assign y7777 = ~n13629 ;
  assign y7778 = n13633 ;
  assign y7779 = ~n13638 ;
  assign y7780 = ~1'b0 ;
  assign y7781 = ~n13642 ;
  assign y7782 = ~1'b0 ;
  assign y7783 = ~1'b0 ;
  assign y7784 = ~n13644 ;
  assign y7785 = ~n13653 ;
  assign y7786 = ~n13654 ;
  assign y7787 = ~n13659 ;
  assign y7788 = n13661 ;
  assign y7789 = n13663 ;
  assign y7790 = ~n13665 ;
  assign y7791 = ~n13667 ;
  assign y7792 = ~1'b0 ;
  assign y7793 = ~n13671 ;
  assign y7794 = ~1'b0 ;
  assign y7795 = ~1'b0 ;
  assign y7796 = ~n13676 ;
  assign y7797 = n13677 ;
  assign y7798 = n13681 ;
  assign y7799 = ~n13690 ;
  assign y7800 = ~1'b0 ;
  assign y7801 = ~n1854 ;
  assign y7802 = n13693 ;
  assign y7803 = n13694 ;
  assign y7804 = n13700 ;
  assign y7805 = ~n13703 ;
  assign y7806 = ~n13705 ;
  assign y7807 = ~n3791 ;
  assign y7808 = n13712 ;
  assign y7809 = n13715 ;
  assign y7810 = ~1'b0 ;
  assign y7811 = ~n9786 ;
  assign y7812 = ~1'b0 ;
  assign y7813 = ~n13724 ;
  assign y7814 = ~n13725 ;
  assign y7815 = ~1'b0 ;
  assign y7816 = ~n872 ;
  assign y7817 = ~n13331 ;
  assign y7818 = ~1'b0 ;
  assign y7819 = ~n13729 ;
  assign y7820 = n13733 ;
  assign y7821 = n13735 ;
  assign y7822 = ~n13737 ;
  assign y7823 = ~n13738 ;
  assign y7824 = ~n13742 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = ~n13743 ;
  assign y7827 = ~n13746 ;
  assign y7828 = ~n13747 ;
  assign y7829 = n4920 ;
  assign y7830 = n13749 ;
  assign y7831 = n13750 ;
  assign y7832 = ~n641 ;
  assign y7833 = ~n13752 ;
  assign y7834 = ~n8251 ;
  assign y7835 = ~1'b0 ;
  assign y7836 = ~n7558 ;
  assign y7837 = ~n13763 ;
  assign y7838 = ~n13764 ;
  assign y7839 = ~1'b0 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = ~n13767 ;
  assign y7842 = n13770 ;
  assign y7843 = ~1'b0 ;
  assign y7844 = n13773 ;
  assign y7845 = ~n13775 ;
  assign y7846 = n8956 ;
  assign y7847 = n13785 ;
  assign y7848 = ~1'b0 ;
  assign y7849 = ~1'b0 ;
  assign y7850 = ~n13788 ;
  assign y7851 = n13791 ;
  assign y7852 = ~n13796 ;
  assign y7853 = n4728 ;
  assign y7854 = n13800 ;
  assign y7855 = ~1'b0 ;
  assign y7856 = ~1'b0 ;
  assign y7857 = ~1'b0 ;
  assign y7858 = n13801 ;
  assign y7859 = n13802 ;
  assign y7860 = 1'b0 ;
  assign y7861 = ~1'b0 ;
  assign y7862 = n13804 ;
  assign y7863 = ~n13805 ;
  assign y7864 = ~n13810 ;
  assign y7865 = n13814 ;
  assign y7866 = n13816 ;
  assign y7867 = ~1'b0 ;
  assign y7868 = ~n13817 ;
  assign y7869 = ~n13818 ;
  assign y7870 = ~1'b0 ;
  assign y7871 = ~1'b0 ;
  assign y7872 = n13821 ;
  assign y7873 = ~n13823 ;
  assign y7874 = n13825 ;
  assign y7875 = ~1'b0 ;
  assign y7876 = ~n13826 ;
  assign y7877 = ~1'b0 ;
  assign y7878 = n13827 ;
  assign y7879 = ~n13830 ;
  assign y7880 = ~1'b0 ;
  assign y7881 = ~n13835 ;
  assign y7882 = n13836 ;
  assign y7883 = n13839 ;
  assign y7884 = ~1'b0 ;
  assign y7885 = ~1'b0 ;
  assign y7886 = ~1'b0 ;
  assign y7887 = n13840 ;
  assign y7888 = ~n13842 ;
  assign y7889 = ~1'b0 ;
  assign y7890 = ~1'b0 ;
  assign y7891 = ~1'b0 ;
  assign y7892 = n13845 ;
  assign y7893 = ~1'b0 ;
  assign y7894 = ~n13846 ;
  assign y7895 = n13855 ;
  assign y7896 = 1'b0 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = ~1'b0 ;
  assign y7899 = ~n13856 ;
  assign y7900 = ~n13857 ;
  assign y7901 = ~1'b0 ;
  assign y7902 = n13858 ;
  assign y7903 = n13859 ;
  assign y7904 = ~n13860 ;
  assign y7905 = n13861 ;
  assign y7906 = n4333 ;
  assign y7907 = ~1'b0 ;
  assign y7908 = ~1'b0 ;
  assign y7909 = ~n13865 ;
  assign y7910 = 1'b0 ;
  assign y7911 = ~n6368 ;
  assign y7912 = n13870 ;
  assign y7913 = ~n13876 ;
  assign y7914 = n13879 ;
  assign y7915 = ~n13881 ;
  assign y7916 = ~1'b0 ;
  assign y7917 = n13882 ;
  assign y7918 = ~n13893 ;
  assign y7919 = n13896 ;
  assign y7920 = n13898 ;
  assign y7921 = n13902 ;
  assign y7922 = n12694 ;
  assign y7923 = n13909 ;
  assign y7924 = n7926 ;
  assign y7925 = ~n5106 ;
  assign y7926 = ~n13911 ;
  assign y7927 = ~1'b0 ;
  assign y7928 = ~n13912 ;
  assign y7929 = ~n13913 ;
  assign y7930 = n13914 ;
  assign y7931 = n13919 ;
  assign y7932 = ~n13921 ;
  assign y7933 = n13923 ;
  assign y7934 = ~1'b0 ;
  assign y7935 = ~1'b0 ;
  assign y7936 = ~n13924 ;
  assign y7937 = ~n13925 ;
  assign y7938 = ~1'b0 ;
  assign y7939 = ~n8410 ;
  assign y7940 = ~1'b0 ;
  assign y7941 = ~1'b0 ;
  assign y7942 = ~n13926 ;
  assign y7943 = ~n13931 ;
  assign y7944 = 1'b0 ;
  assign y7945 = n13933 ;
  assign y7946 = ~n13936 ;
  assign y7947 = ~n13938 ;
  assign y7948 = ~1'b0 ;
  assign y7949 = n13939 ;
  assign y7950 = ~1'b0 ;
  assign y7951 = n13941 ;
  assign y7952 = ~1'b0 ;
  assign y7953 = ~1'b0 ;
  assign y7954 = ~1'b0 ;
  assign y7955 = 1'b0 ;
  assign y7956 = ~1'b0 ;
  assign y7957 = ~1'b0 ;
  assign y7958 = n13945 ;
  assign y7959 = n10864 ;
  assign y7960 = ~1'b0 ;
  assign y7961 = ~n11899 ;
  assign y7962 = ~n13950 ;
  assign y7963 = ~1'b0 ;
  assign y7964 = n13951 ;
  assign y7965 = n13952 ;
  assign y7966 = ~1'b0 ;
  assign y7967 = ~n13953 ;
  assign y7968 = ~1'b0 ;
  assign y7969 = ~n13958 ;
  assign y7970 = n13962 ;
  assign y7971 = ~n5105 ;
  assign y7972 = n13963 ;
  assign y7973 = ~1'b0 ;
  assign y7974 = ~1'b0 ;
  assign y7975 = n8045 ;
  assign y7976 = 1'b0 ;
  assign y7977 = n13967 ;
  assign y7978 = n13970 ;
  assign y7979 = ~n13973 ;
  assign y7980 = ~n13976 ;
  assign y7981 = ~n13978 ;
  assign y7982 = ~1'b0 ;
  assign y7983 = n858 ;
  assign y7984 = ~1'b0 ;
  assign y7985 = ~1'b0 ;
  assign y7986 = n13979 ;
  assign y7987 = ~1'b0 ;
  assign y7988 = ~n13980 ;
  assign y7989 = n13985 ;
  assign y7990 = ~n13990 ;
  assign y7991 = ~n13992 ;
  assign y7992 = n14004 ;
  assign y7993 = n14008 ;
  assign y7994 = n14011 ;
  assign y7995 = ~n14015 ;
  assign y7996 = ~1'b0 ;
  assign y7997 = n14017 ;
  assign y7998 = ~1'b0 ;
  assign y7999 = n12922 ;
  assign y8000 = ~n14025 ;
  assign y8001 = ~n14031 ;
  assign y8002 = ~n14033 ;
  assign y8003 = ~n11013 ;
  assign y8004 = ~n14036 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = n7684 ;
  assign y8007 = ~n14038 ;
  assign y8008 = ~1'b0 ;
  assign y8009 = ~1'b0 ;
  assign y8010 = n14040 ;
  assign y8011 = n14041 ;
  assign y8012 = ~n14043 ;
  assign y8013 = ~1'b0 ;
  assign y8014 = ~1'b0 ;
  assign y8015 = ~1'b0 ;
  assign y8016 = ~n14047 ;
  assign y8017 = n14051 ;
  assign y8018 = ~n9636 ;
  assign y8019 = ~n14055 ;
  assign y8020 = ~n14058 ;
  assign y8021 = ~n14061 ;
  assign y8022 = n14063 ;
  assign y8023 = ~1'b0 ;
  assign y8024 = ~n14065 ;
  assign y8025 = n12128 ;
  assign y8026 = n14074 ;
  assign y8027 = ~n14077 ;
  assign y8028 = ~1'b0 ;
  assign y8029 = n14081 ;
  assign y8030 = n14084 ;
  assign y8031 = n14090 ;
  assign y8032 = ~n14091 ;
  assign y8033 = ~n14099 ;
  assign y8034 = n14101 ;
  assign y8035 = ~n5869 ;
  assign y8036 = ~n14103 ;
  assign y8037 = ~n14105 ;
  assign y8038 = ~1'b0 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = 1'b0 ;
  assign y8041 = ~1'b0 ;
  assign y8042 = ~n14110 ;
  assign y8043 = ~n14112 ;
  assign y8044 = ~n14114 ;
  assign y8045 = ~1'b0 ;
  assign y8046 = ~1'b0 ;
  assign y8047 = n14117 ;
  assign y8048 = ~1'b0 ;
  assign y8049 = ~n14119 ;
  assign y8050 = ~1'b0 ;
  assign y8051 = n14121 ;
  assign y8052 = n14122 ;
  assign y8053 = n14125 ;
  assign y8054 = ~n14128 ;
  assign y8055 = n14130 ;
  assign y8056 = n14131 ;
  assign y8057 = ~1'b0 ;
  assign y8058 = ~n14132 ;
  assign y8059 = n14135 ;
  assign y8060 = ~1'b0 ;
  assign y8061 = ~1'b0 ;
  assign y8062 = n14137 ;
  assign y8063 = 1'b0 ;
  assign y8064 = n6413 ;
  assign y8065 = ~n4656 ;
  assign y8066 = ~n14140 ;
  assign y8067 = ~n14155 ;
  assign y8068 = ~1'b0 ;
  assign y8069 = ~n14161 ;
  assign y8070 = ~1'b0 ;
  assign y8071 = n14164 ;
  assign y8072 = ~n14170 ;
  assign y8073 = ~n14173 ;
  assign y8074 = n14177 ;
  assign y8075 = n14180 ;
  assign y8076 = ~n11278 ;
  assign y8077 = ~n14182 ;
  assign y8078 = ~n2546 ;
  assign y8079 = ~1'b0 ;
  assign y8080 = n14184 ;
  assign y8081 = ~1'b0 ;
  assign y8082 = n14185 ;
  assign y8083 = ~n14190 ;
  assign y8084 = n14191 ;
  assign y8085 = ~1'b0 ;
  assign y8086 = ~1'b0 ;
  assign y8087 = n14192 ;
  assign y8088 = ~1'b0 ;
  assign y8089 = 1'b0 ;
  assign y8090 = ~n4927 ;
  assign y8091 = ~1'b0 ;
  assign y8092 = ~n14196 ;
  assign y8093 = ~n14201 ;
  assign y8094 = n14202 ;
  assign y8095 = n14211 ;
  assign y8096 = ~1'b0 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = n14213 ;
  assign y8099 = ~1'b0 ;
  assign y8100 = n14214 ;
  assign y8101 = ~n14216 ;
  assign y8102 = ~1'b0 ;
  assign y8103 = ~n14218 ;
  assign y8104 = ~n14220 ;
  assign y8105 = ~n5433 ;
  assign y8106 = n14221 ;
  assign y8107 = n14223 ;
  assign y8108 = ~n14224 ;
  assign y8109 = n14228 ;
  assign y8110 = ~n14230 ;
  assign y8111 = n14234 ;
  assign y8112 = n14238 ;
  assign y8113 = ~n10844 ;
  assign y8114 = n6182 ;
  assign y8115 = ~n14239 ;
  assign y8116 = n14243 ;
  assign y8117 = ~1'b0 ;
  assign y8118 = ~1'b0 ;
  assign y8119 = ~n14244 ;
  assign y8120 = ~1'b0 ;
  assign y8121 = ~1'b0 ;
  assign y8122 = n14245 ;
  assign y8123 = n14247 ;
  assign y8124 = n14248 ;
  assign y8125 = ~1'b0 ;
  assign y8126 = n14250 ;
  assign y8127 = ~1'b0 ;
  assign y8128 = n14260 ;
  assign y8129 = n14261 ;
  assign y8130 = ~n14263 ;
  assign y8131 = ~n5072 ;
  assign y8132 = n14265 ;
  assign y8133 = n14270 ;
  assign y8134 = ~1'b0 ;
  assign y8135 = n14272 ;
  assign y8136 = ~1'b0 ;
  assign y8137 = n7494 ;
  assign y8138 = ~n14274 ;
  assign y8139 = ~n3167 ;
  assign y8140 = n14275 ;
  assign y8141 = ~n14281 ;
  assign y8142 = 1'b0 ;
  assign y8143 = n14283 ;
  assign y8144 = ~1'b0 ;
  assign y8145 = ~1'b0 ;
  assign y8146 = ~n14287 ;
  assign y8147 = ~1'b0 ;
  assign y8148 = ~n14288 ;
  assign y8149 = ~n14289 ;
  assign y8150 = n14290 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = ~1'b0 ;
  assign y8153 = ~1'b0 ;
  assign y8154 = ~n14292 ;
  assign y8155 = ~n14295 ;
  assign y8156 = ~1'b0 ;
  assign y8157 = ~1'b0 ;
  assign y8158 = ~1'b0 ;
  assign y8159 = ~n14296 ;
  assign y8160 = n14299 ;
  assign y8161 = ~1'b0 ;
  assign y8162 = n14300 ;
  assign y8163 = ~n14301 ;
  assign y8164 = n14302 ;
  assign y8165 = n14304 ;
  assign y8166 = n14305 ;
  assign y8167 = n14306 ;
  assign y8168 = ~1'b0 ;
  assign y8169 = ~n14309 ;
  assign y8170 = ~n14311 ;
  assign y8171 = ~n14313 ;
  assign y8172 = ~1'b0 ;
  assign y8173 = ~n14318 ;
  assign y8174 = ~n14319 ;
  assign y8175 = ~n14320 ;
  assign y8176 = ~1'b0 ;
  assign y8177 = n14321 ;
  assign y8178 = ~1'b0 ;
  assign y8179 = n14327 ;
  assign y8180 = n14329 ;
  assign y8181 = ~1'b0 ;
  assign y8182 = ~1'b0 ;
  assign y8183 = n14331 ;
  assign y8184 = ~1'b0 ;
  assign y8185 = ~n14333 ;
  assign y8186 = ~n14336 ;
  assign y8187 = n14338 ;
  assign y8188 = ~n14339 ;
  assign y8189 = ~1'b0 ;
  assign y8190 = ~n14346 ;
  assign y8191 = n14351 ;
  assign y8192 = ~n14352 ;
  assign y8193 = n5101 ;
  assign y8194 = ~n14354 ;
  assign y8195 = ~n14355 ;
  assign y8196 = ~1'b0 ;
  assign y8197 = ~n5631 ;
  assign y8198 = ~n14361 ;
  assign y8199 = ~n14363 ;
  assign y8200 = ~n14370 ;
  assign y8201 = ~1'b0 ;
  assign y8202 = n14371 ;
  assign y8203 = n14373 ;
  assign y8204 = ~1'b0 ;
  assign y8205 = ~1'b0 ;
  assign y8206 = n14374 ;
  assign y8207 = ~1'b0 ;
  assign y8208 = ~n1766 ;
  assign y8209 = ~1'b0 ;
  assign y8210 = ~1'b0 ;
  assign y8211 = ~n14375 ;
  assign y8212 = ~1'b0 ;
  assign y8213 = ~n14376 ;
  assign y8214 = n14377 ;
  assign y8215 = ~1'b0 ;
  assign y8216 = ~1'b0 ;
  assign y8217 = ~n14387 ;
  assign y8218 = ~1'b0 ;
  assign y8219 = ~1'b0 ;
  assign y8220 = ~n14389 ;
  assign y8221 = n14391 ;
  assign y8222 = ~1'b0 ;
  assign y8223 = n14403 ;
  assign y8224 = ~1'b0 ;
  assign y8225 = 1'b0 ;
  assign y8226 = ~1'b0 ;
  assign y8227 = ~n14404 ;
  assign y8228 = n14405 ;
  assign y8229 = n14406 ;
  assign y8230 = ~n14409 ;
  assign y8231 = n14415 ;
  assign y8232 = ~1'b0 ;
  assign y8233 = ~n3071 ;
  assign y8234 = ~n14417 ;
  assign y8235 = ~n14422 ;
  assign y8236 = ~n14431 ;
  assign y8237 = ~1'b0 ;
  assign y8238 = ~n14432 ;
  assign y8239 = ~n14434 ;
  assign y8240 = ~1'b0 ;
  assign y8241 = n14435 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = ~1'b0 ;
  assign y8244 = ~n14443 ;
  assign y8245 = n14446 ;
  assign y8246 = n14447 ;
  assign y8247 = ~n14451 ;
  assign y8248 = ~n14454 ;
  assign y8249 = ~1'b0 ;
  assign y8250 = ~1'b0 ;
  assign y8251 = ~n14456 ;
  assign y8252 = ~n14459 ;
  assign y8253 = n14463 ;
  assign y8254 = ~n14464 ;
  assign y8255 = n11720 ;
  assign y8256 = ~1'b0 ;
  assign y8257 = n14465 ;
  assign y8258 = ~n14473 ;
  assign y8259 = ~n14476 ;
  assign y8260 = ~1'b0 ;
  assign y8261 = ~n14482 ;
  assign y8262 = ~1'b0 ;
  assign y8263 = ~n14483 ;
  assign y8264 = n14485 ;
  assign y8265 = ~n14488 ;
  assign y8266 = n14491 ;
  assign y8267 = n14493 ;
  assign y8268 = n14496 ;
  assign y8269 = n14497 ;
  assign y8270 = ~1'b0 ;
  assign y8271 = ~n14502 ;
  assign y8272 = ~n14507 ;
  assign y8273 = n14509 ;
  assign y8274 = ~n14511 ;
  assign y8275 = ~n14518 ;
  assign y8276 = ~1'b0 ;
  assign y8277 = ~n14519 ;
  assign y8278 = n14520 ;
  assign y8279 = ~n14522 ;
  assign y8280 = ~1'b0 ;
  assign y8281 = ~1'b0 ;
  assign y8282 = n14523 ;
  assign y8283 = ~n14526 ;
  assign y8284 = ~1'b0 ;
  assign y8285 = ~1'b0 ;
  assign y8286 = n14529 ;
  assign y8287 = ~n4682 ;
  assign y8288 = n7105 ;
  assign y8289 = ~n14530 ;
  assign y8290 = ~1'b0 ;
  assign y8291 = ~n14531 ;
  assign y8292 = ~n14532 ;
  assign y8293 = ~n14534 ;
  assign y8294 = ~1'b0 ;
  assign y8295 = n14535 ;
  assign y8296 = n14536 ;
  assign y8297 = ~1'b0 ;
  assign y8298 = ~1'b0 ;
  assign y8299 = n14539 ;
  assign y8300 = ~n14543 ;
  assign y8301 = ~1'b0 ;
  assign y8302 = n14545 ;
  assign y8303 = n14547 ;
  assign y8304 = ~1'b0 ;
  assign y8305 = ~1'b0 ;
  assign y8306 = n14549 ;
  assign y8307 = ~1'b0 ;
  assign y8308 = n2768 ;
  assign y8309 = ~n14553 ;
  assign y8310 = n7757 ;
  assign y8311 = ~n14554 ;
  assign y8312 = ~n14556 ;
  assign y8313 = ~n10498 ;
  assign y8314 = n14557 ;
  assign y8315 = ~1'b0 ;
  assign y8316 = ~n14559 ;
  assign y8317 = n8081 ;
  assign y8318 = n14560 ;
  assign y8319 = ~n14562 ;
  assign y8320 = ~n14563 ;
  assign y8321 = ~n14565 ;
  assign y8322 = n14567 ;
  assign y8323 = ~1'b0 ;
  assign y8324 = n14576 ;
  assign y8325 = ~1'b0 ;
  assign y8326 = n14581 ;
  assign y8327 = ~n14587 ;
  assign y8328 = ~n14592 ;
  assign y8329 = ~1'b0 ;
  assign y8330 = ~n14593 ;
  assign y8331 = n14594 ;
  assign y8332 = ~n14595 ;
  assign y8333 = n14600 ;
  assign y8334 = n14606 ;
  assign y8335 = ~1'b0 ;
  assign y8336 = n14609 ;
  assign y8337 = n14612 ;
  assign y8338 = n14613 ;
  assign y8339 = n7161 ;
  assign y8340 = ~n14627 ;
  assign y8341 = ~n14628 ;
  assign y8342 = ~n14632 ;
  assign y8343 = n14637 ;
  assign y8344 = 1'b0 ;
  assign y8345 = n8931 ;
  assign y8346 = n14641 ;
  assign y8347 = ~1'b0 ;
  assign y8348 = ~1'b0 ;
  assign y8349 = ~1'b0 ;
  assign y8350 = n14645 ;
  assign y8351 = ~1'b0 ;
  assign y8352 = n14648 ;
  assign y8353 = ~n14649 ;
  assign y8354 = n14650 ;
  assign y8355 = ~1'b0 ;
  assign y8356 = ~1'b0 ;
  assign y8357 = ~n14656 ;
  assign y8358 = ~1'b0 ;
  assign y8359 = ~1'b0 ;
  assign y8360 = ~n14657 ;
  assign y8361 = ~n14659 ;
  assign y8362 = ~n14662 ;
  assign y8363 = n14667 ;
  assign y8364 = ~n14669 ;
  assign y8365 = ~n14670 ;
  assign y8366 = n14672 ;
  assign y8367 = n14676 ;
  assign y8368 = ~1'b0 ;
  assign y8369 = ~n14678 ;
  assign y8370 = ~n14682 ;
  assign y8371 = ~n14683 ;
  assign y8372 = n3336 ;
  assign y8373 = n14690 ;
  assign y8374 = ~1'b0 ;
  assign y8375 = ~1'b0 ;
  assign y8376 = ~n14691 ;
  assign y8377 = ~n14698 ;
  assign y8378 = ~1'b0 ;
  assign y8379 = ~1'b0 ;
  assign y8380 = ~1'b0 ;
  assign y8381 = n14700 ;
  assign y8382 = ~n14705 ;
  assign y8383 = n14332 ;
  assign y8384 = n14708 ;
  assign y8385 = ~1'b0 ;
  assign y8386 = ~n14710 ;
  assign y8387 = n14711 ;
  assign y8388 = 1'b0 ;
  assign y8389 = n14718 ;
  assign y8390 = ~n14754 ;
  assign y8391 = ~n8367 ;
  assign y8392 = ~1'b0 ;
  assign y8393 = ~1'b0 ;
  assign y8394 = n14755 ;
  assign y8395 = ~1'b0 ;
  assign y8396 = ~n14756 ;
  assign y8397 = ~1'b0 ;
  assign y8398 = n12257 ;
  assign y8399 = ~1'b0 ;
  assign y8400 = n14758 ;
  assign y8401 = n14760 ;
  assign y8402 = ~n14762 ;
  assign y8403 = n11785 ;
  assign y8404 = n14773 ;
  assign y8405 = n4787 ;
  assign y8406 = ~1'b0 ;
  assign y8407 = ~1'b0 ;
  assign y8408 = ~n14774 ;
  assign y8409 = ~1'b0 ;
  assign y8410 = ~n14775 ;
  assign y8411 = ~n14777 ;
  assign y8412 = ~1'b0 ;
  assign y8413 = ~n14778 ;
  assign y8414 = n14781 ;
  assign y8415 = ~n14782 ;
  assign y8416 = ~n14783 ;
  assign y8417 = ~n14786 ;
  assign y8418 = ~1'b0 ;
  assign y8419 = ~n14788 ;
  assign y8420 = ~1'b0 ;
  assign y8421 = n14792 ;
  assign y8422 = ~1'b0 ;
  assign y8423 = ~n14797 ;
  assign y8424 = n14799 ;
  assign y8425 = ~n14802 ;
  assign y8426 = n14803 ;
  assign y8427 = ~1'b0 ;
  assign y8428 = ~n14808 ;
  assign y8429 = ~1'b0 ;
  assign y8430 = 1'b0 ;
  assign y8431 = ~1'b0 ;
  assign y8432 = n14809 ;
  assign y8433 = n14810 ;
  assign y8434 = ~n14815 ;
  assign y8435 = ~n14817 ;
  assign y8436 = ~n14819 ;
  assign y8437 = n14821 ;
  assign y8438 = n14826 ;
  assign y8439 = ~n9693 ;
  assign y8440 = ~1'b0 ;
  assign y8441 = ~1'b0 ;
  assign y8442 = ~n14828 ;
  assign y8443 = ~1'b0 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~n14837 ;
  assign y8446 = ~n14839 ;
  assign y8447 = n14846 ;
  assign y8448 = ~1'b0 ;
  assign y8449 = ~1'b0 ;
  assign y8450 = n14847 ;
  assign y8451 = n14854 ;
  assign y8452 = n14856 ;
  assign y8453 = n14858 ;
  assign y8454 = ~n14861 ;
  assign y8455 = ~1'b0 ;
  assign y8456 = n14862 ;
  assign y8457 = ~n14863 ;
  assign y8458 = n14864 ;
  assign y8459 = n14866 ;
  assign y8460 = n14867 ;
  assign y8461 = ~n14871 ;
  assign y8462 = n14873 ;
  assign y8463 = ~1'b0 ;
  assign y8464 = n14875 ;
  assign y8465 = x123 ;
  assign y8466 = ~n14878 ;
  assign y8467 = ~1'b0 ;
  assign y8468 = n14880 ;
  assign y8469 = ~n14881 ;
  assign y8470 = n14883 ;
  assign y8471 = ~n14884 ;
  assign y8472 = ~n14885 ;
  assign y8473 = ~n14887 ;
  assign y8474 = ~n14888 ;
  assign y8475 = ~n14892 ;
  assign y8476 = n14894 ;
  assign y8477 = n14895 ;
  assign y8478 = ~n3748 ;
  assign y8479 = n14897 ;
  assign y8480 = n14898 ;
  assign y8481 = n14900 ;
  assign y8482 = ~n14901 ;
  assign y8483 = n14905 ;
  assign y8484 = ~1'b0 ;
  assign y8485 = ~n2037 ;
  assign y8486 = ~n14910 ;
  assign y8487 = ~1'b0 ;
  assign y8488 = 1'b0 ;
  assign y8489 = n14911 ;
  assign y8490 = ~n14913 ;
  assign y8491 = n14915 ;
  assign y8492 = ~n14921 ;
  assign y8493 = ~n14923 ;
  assign y8494 = ~n14924 ;
  assign y8495 = ~1'b0 ;
  assign y8496 = ~1'b0 ;
  assign y8497 = n14925 ;
  assign y8498 = n14927 ;
  assign y8499 = ~1'b0 ;
  assign y8500 = ~n14930 ;
  assign y8501 = ~n14933 ;
  assign y8502 = ~1'b0 ;
  assign y8503 = ~n14935 ;
  assign y8504 = ~n14941 ;
  assign y8505 = ~1'b0 ;
  assign y8506 = ~1'b0 ;
  assign y8507 = ~n14943 ;
  assign y8508 = n14947 ;
  assign y8509 = ~1'b0 ;
  assign y8510 = n14950 ;
  assign y8511 = ~1'b0 ;
  assign y8512 = n14952 ;
  assign y8513 = ~n14953 ;
  assign y8514 = n14960 ;
  assign y8515 = n14963 ;
  assign y8516 = 1'b0 ;
  assign y8517 = n14968 ;
  assign y8518 = n14969 ;
  assign y8519 = n14972 ;
  assign y8520 = ~1'b0 ;
  assign y8521 = n14974 ;
  assign y8522 = n14977 ;
  assign y8523 = ~n14978 ;
  assign y8524 = ~n14980 ;
  assign y8525 = n14987 ;
  assign y8526 = ~n365 ;
  assign y8527 = ~n14994 ;
  assign y8528 = ~n14997 ;
  assign y8529 = n14999 ;
  assign y8530 = ~1'b0 ;
  assign y8531 = ~n15000 ;
  assign y8532 = ~1'b0 ;
  assign y8533 = ~n15005 ;
  assign y8534 = ~n15007 ;
  assign y8535 = n15008 ;
  assign y8536 = ~1'b0 ;
  assign y8537 = n14757 ;
  assign y8538 = ~1'b0 ;
  assign y8539 = ~n15009 ;
  assign y8540 = n15011 ;
  assign y8541 = ~1'b0 ;
  assign y8542 = ~1'b0 ;
  assign y8543 = ~1'b0 ;
  assign y8544 = ~n15016 ;
  assign y8545 = ~1'b0 ;
  assign y8546 = ~1'b0 ;
  assign y8547 = ~1'b0 ;
  assign y8548 = ~1'b0 ;
  assign y8549 = ~1'b0 ;
  assign y8550 = ~n15021 ;
  assign y8551 = ~n15030 ;
  assign y8552 = ~1'b0 ;
  assign y8553 = ~n7172 ;
  assign y8554 = n2076 ;
  assign y8555 = ~1'b0 ;
  assign y8556 = ~n15031 ;
  assign y8557 = n15035 ;
  assign y8558 = ~n15037 ;
  assign y8559 = n15041 ;
  assign y8560 = ~n9254 ;
  assign y8561 = ~n15043 ;
  assign y8562 = ~1'b0 ;
  assign y8563 = 1'b0 ;
  assign y8564 = ~n15046 ;
  assign y8565 = ~n15047 ;
  assign y8566 = ~n15048 ;
  assign y8567 = ~1'b0 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = ~n15051 ;
  assign y8570 = n15053 ;
  assign y8571 = ~n15056 ;
  assign y8572 = n15058 ;
  assign y8573 = ~n15065 ;
  assign y8574 = ~1'b0 ;
  assign y8575 = ~n15073 ;
  assign y8576 = ~1'b0 ;
  assign y8577 = ~n15075 ;
  assign y8578 = n15078 ;
  assign y8579 = ~n9215 ;
  assign y8580 = ~1'b0 ;
  assign y8581 = ~n15080 ;
  assign y8582 = ~1'b0 ;
  assign y8583 = ~n15091 ;
  assign y8584 = ~n15094 ;
  assign y8585 = ~n15095 ;
  assign y8586 = n15096 ;
  assign y8587 = 1'b0 ;
  assign y8588 = n15098 ;
  assign y8589 = ~1'b0 ;
  assign y8590 = n15103 ;
  assign y8591 = n15104 ;
  assign y8592 = n15108 ;
  assign y8593 = ~1'b0 ;
  assign y8594 = ~n15110 ;
  assign y8595 = ~n15119 ;
  assign y8596 = ~n15121 ;
  assign y8597 = ~1'b0 ;
  assign y8598 = n15122 ;
  assign y8599 = n15126 ;
  assign y8600 = n15128 ;
  assign y8601 = n15130 ;
  assign y8602 = ~n15133 ;
  assign y8603 = n15135 ;
  assign y8604 = n15139 ;
  assign y8605 = ~n15142 ;
  assign y8606 = ~n15148 ;
  assign y8607 = ~1'b0 ;
  assign y8608 = ~n15157 ;
  assign y8609 = n15159 ;
  assign y8610 = ~n15163 ;
  assign y8611 = ~1'b0 ;
  assign y8612 = ~n15165 ;
  assign y8613 = ~1'b0 ;
  assign y8614 = n15167 ;
  assign y8615 = ~n15168 ;
  assign y8616 = ~1'b0 ;
  assign y8617 = n15169 ;
  assign y8618 = ~1'b0 ;
  assign y8619 = ~n15171 ;
  assign y8620 = ~1'b0 ;
  assign y8621 = 1'b0 ;
  assign y8622 = n15172 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = ~1'b0 ;
  assign y8625 = ~1'b0 ;
  assign y8626 = ~1'b0 ;
  assign y8627 = ~n6134 ;
  assign y8628 = n15177 ;
  assign y8629 = n15180 ;
  assign y8630 = n15181 ;
  assign y8631 = ~1'b0 ;
  assign y8632 = ~1'b0 ;
  assign y8633 = ~1'b0 ;
  assign y8634 = n15182 ;
  assign y8635 = n12735 ;
  assign y8636 = ~n15187 ;
  assign y8637 = ~1'b0 ;
  assign y8638 = ~n15192 ;
  assign y8639 = ~1'b0 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = n15194 ;
  assign y8642 = n15196 ;
  assign y8643 = ~n15197 ;
  assign y8644 = ~n15199 ;
  assign y8645 = ~1'b0 ;
  assign y8646 = ~1'b0 ;
  assign y8647 = n4538 ;
  assign y8648 = ~1'b0 ;
  assign y8649 = ~1'b0 ;
  assign y8650 = ~n4718 ;
  assign y8651 = n15201 ;
  assign y8652 = ~n15206 ;
  assign y8653 = n15208 ;
  assign y8654 = ~1'b0 ;
  assign y8655 = 1'b0 ;
  assign y8656 = ~1'b0 ;
  assign y8657 = n15210 ;
  assign y8658 = ~1'b0 ;
  assign y8659 = ~n15217 ;
  assign y8660 = ~n15219 ;
  assign y8661 = ~n15223 ;
  assign y8662 = ~n15227 ;
  assign y8663 = ~n15228 ;
  assign y8664 = ~1'b0 ;
  assign y8665 = ~1'b0 ;
  assign y8666 = ~1'b0 ;
  assign y8667 = n15231 ;
  assign y8668 = ~1'b0 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = 1'b0 ;
  assign y8671 = ~1'b0 ;
  assign y8672 = ~n15235 ;
  assign y8673 = n15236 ;
  assign y8674 = n15237 ;
  assign y8675 = n15239 ;
  assign y8676 = ~n15240 ;
  assign y8677 = n15241 ;
  assign y8678 = ~n9242 ;
  assign y8679 = ~1'b0 ;
  assign y8680 = n15243 ;
  assign y8681 = n15246 ;
  assign y8682 = n15249 ;
  assign y8683 = ~1'b0 ;
  assign y8684 = ~n15250 ;
  assign y8685 = ~n15254 ;
  assign y8686 = n15256 ;
  assign y8687 = ~n15269 ;
  assign y8688 = n15284 ;
  assign y8689 = ~n15294 ;
  assign y8690 = n15297 ;
  assign y8691 = n15300 ;
  assign y8692 = ~n15302 ;
  assign y8693 = n15307 ;
  assign y8694 = ~1'b0 ;
  assign y8695 = ~1'b0 ;
  assign y8696 = ~n15310 ;
  assign y8697 = n15316 ;
  assign y8698 = n15318 ;
  assign y8699 = ~n15320 ;
  assign y8700 = ~1'b0 ;
  assign y8701 = ~1'b0 ;
  assign y8702 = ~n15327 ;
  assign y8703 = ~n15328 ;
  assign y8704 = ~1'b0 ;
  assign y8705 = ~1'b0 ;
  assign y8706 = ~1'b0 ;
  assign y8707 = n15329 ;
  assign y8708 = ~1'b0 ;
  assign y8709 = ~n15330 ;
  assign y8710 = ~n15331 ;
  assign y8711 = ~n15332 ;
  assign y8712 = ~n15335 ;
  assign y8713 = 1'b0 ;
  assign y8714 = n15336 ;
  assign y8715 = n12213 ;
  assign y8716 = n15339 ;
  assign y8717 = 1'b0 ;
  assign y8718 = ~1'b0 ;
  assign y8719 = n15343 ;
  assign y8720 = ~1'b0 ;
  assign y8721 = ~n15346 ;
  assign y8722 = ~1'b0 ;
  assign y8723 = n15348 ;
  assign y8724 = ~n15350 ;
  assign y8725 = ~n15355 ;
  assign y8726 = ~n15007 ;
  assign y8727 = n15357 ;
  assign y8728 = n15361 ;
  assign y8729 = ~1'b0 ;
  assign y8730 = ~n15365 ;
  assign y8731 = ~1'b0 ;
  assign y8732 = n15366 ;
  assign y8733 = n15370 ;
  assign y8734 = n4913 ;
  assign y8735 = ~n15372 ;
  assign y8736 = n15373 ;
  assign y8737 = ~n15376 ;
  assign y8738 = ~1'b0 ;
  assign y8739 = ~n15380 ;
  assign y8740 = ~n15382 ;
  assign y8741 = n15385 ;
  assign y8742 = ~n4568 ;
  assign y8743 = ~1'b0 ;
  assign y8744 = ~1'b0 ;
  assign y8745 = n15386 ;
  assign y8746 = n15387 ;
  assign y8747 = ~n15389 ;
  assign y8748 = n15391 ;
  assign y8749 = ~1'b0 ;
  assign y8750 = n15392 ;
  assign y8751 = n15397 ;
  assign y8752 = ~n15399 ;
  assign y8753 = ~n15400 ;
  assign y8754 = ~1'b0 ;
  assign y8755 = ~1'b0 ;
  assign y8756 = ~n15403 ;
  assign y8757 = ~n15404 ;
  assign y8758 = ~1'b0 ;
  assign y8759 = 1'b0 ;
  assign y8760 = n15408 ;
  assign y8761 = ~n15413 ;
  assign y8762 = ~n15416 ;
  assign y8763 = ~1'b0 ;
  assign y8764 = ~n15417 ;
  assign y8765 = n15419 ;
  assign y8766 = ~1'b0 ;
  assign y8767 = ~n15421 ;
  assign y8768 = ~1'b0 ;
  assign y8769 = ~x142 ;
  assign y8770 = ~1'b0 ;
  assign y8771 = ~1'b0 ;
  assign y8772 = n15422 ;
  assign y8773 = ~1'b0 ;
  assign y8774 = ~n15425 ;
  assign y8775 = ~n15430 ;
  assign y8776 = ~1'b0 ;
  assign y8777 = ~1'b0 ;
  assign y8778 = ~n15432 ;
  assign y8779 = ~n15433 ;
  assign y8780 = ~n15435 ;
  assign y8781 = ~1'b0 ;
  assign y8782 = ~1'b0 ;
  assign y8783 = ~n15436 ;
  assign y8784 = ~n15438 ;
  assign y8785 = n15441 ;
  assign y8786 = ~1'b0 ;
  assign y8787 = ~1'b0 ;
  assign y8788 = n15445 ;
  assign y8789 = n15449 ;
  assign y8790 = ~n15451 ;
  assign y8791 = ~n15454 ;
  assign y8792 = n3143 ;
  assign y8793 = ~1'b0 ;
  assign y8794 = ~1'b0 ;
  assign y8795 = n15460 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = ~n15466 ;
  assign y8798 = ~1'b0 ;
  assign y8799 = ~1'b0 ;
  assign y8800 = ~n15468 ;
  assign y8801 = ~1'b0 ;
  assign y8802 = n15469 ;
  assign y8803 = ~n15470 ;
  assign y8804 = ~n8424 ;
  assign y8805 = ~n15472 ;
  assign y8806 = ~n15474 ;
  assign y8807 = ~n15477 ;
  assign y8808 = n15479 ;
  assign y8809 = n15480 ;
  assign y8810 = n11083 ;
  assign y8811 = ~n15481 ;
  assign y8812 = ~n15491 ;
  assign y8813 = ~n15493 ;
  assign y8814 = ~n15497 ;
  assign y8815 = ~n15501 ;
  assign y8816 = n15503 ;
  assign y8817 = ~n15505 ;
  assign y8818 = ~1'b0 ;
  assign y8819 = ~1'b0 ;
  assign y8820 = ~n15514 ;
  assign y8821 = n15515 ;
  assign y8822 = n15516 ;
  assign y8823 = ~n15519 ;
  assign y8824 = n15521 ;
  assign y8825 = ~n15522 ;
  assign y8826 = n15524 ;
  assign y8827 = ~1'b0 ;
  assign y8828 = n15525 ;
  assign y8829 = ~n15527 ;
  assign y8830 = n15128 ;
  assign y8831 = ~1'b0 ;
  assign y8832 = 1'b0 ;
  assign y8833 = ~n15529 ;
  assign y8834 = ~1'b0 ;
  assign y8835 = n15530 ;
  assign y8836 = ~1'b0 ;
  assign y8837 = n15531 ;
  assign y8838 = n15542 ;
  assign y8839 = n15543 ;
  assign y8840 = ~1'b0 ;
  assign y8841 = ~n15547 ;
  assign y8842 = ~n10473 ;
  assign y8843 = ~n15548 ;
  assign y8844 = ~1'b0 ;
  assign y8845 = ~n15550 ;
  assign y8846 = n15552 ;
  assign y8847 = ~n12837 ;
  assign y8848 = n15554 ;
  assign y8849 = ~n15556 ;
  assign y8850 = ~n15560 ;
  assign y8851 = ~n15561 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = ~n15563 ;
  assign y8854 = n12729 ;
  assign y8855 = ~n15564 ;
  assign y8856 = ~1'b0 ;
  assign y8857 = n15565 ;
  assign y8858 = ~1'b0 ;
  assign y8859 = ~n15569 ;
  assign y8860 = ~n6640 ;
  assign y8861 = ~1'b0 ;
  assign y8862 = n15572 ;
  assign y8863 = ~n15574 ;
  assign y8864 = ~n15576 ;
  assign y8865 = ~n7971 ;
  assign y8866 = ~n15579 ;
  assign y8867 = n15580 ;
  assign y8868 = ~1'b0 ;
  assign y8869 = n15581 ;
  assign y8870 = ~n15582 ;
  assign y8871 = 1'b0 ;
  assign y8872 = ~n15583 ;
  assign y8873 = ~1'b0 ;
  assign y8874 = n15585 ;
  assign y8875 = n15597 ;
  assign y8876 = ~1'b0 ;
  assign y8877 = ~n15601 ;
  assign y8878 = n15602 ;
  assign y8879 = ~n15603 ;
  assign y8880 = n15604 ;
  assign y8881 = n9415 ;
  assign y8882 = n15609 ;
  assign y8883 = ~n15613 ;
  assign y8884 = n15617 ;
  assign y8885 = ~1'b0 ;
  assign y8886 = n15628 ;
  assign y8887 = n15629 ;
  assign y8888 = ~1'b0 ;
  assign y8889 = n15632 ;
  assign y8890 = n15638 ;
  assign y8891 = ~1'b0 ;
  assign y8892 = n15647 ;
  assign y8893 = ~1'b0 ;
  assign y8894 = ~n15650 ;
  assign y8895 = ~n11096 ;
  assign y8896 = n15651 ;
  assign y8897 = n15653 ;
  assign y8898 = ~1'b0 ;
  assign y8899 = ~1'b0 ;
  assign y8900 = ~n15656 ;
  assign y8901 = ~1'b0 ;
  assign y8902 = n15657 ;
  assign y8903 = ~n15660 ;
  assign y8904 = ~n2868 ;
  assign y8905 = n15661 ;
  assign y8906 = ~n15667 ;
  assign y8907 = ~1'b0 ;
  assign y8908 = n15668 ;
  assign y8909 = ~1'b0 ;
  assign y8910 = 1'b0 ;
  assign y8911 = ~n15671 ;
  assign y8912 = ~1'b0 ;
  assign y8913 = ~1'b0 ;
  assign y8914 = ~1'b0 ;
  assign y8915 = ~1'b0 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = n15672 ;
  assign y8918 = ~1'b0 ;
  assign y8919 = ~n15678 ;
  assign y8920 = ~n15680 ;
  assign y8921 = ~1'b0 ;
  assign y8922 = n15681 ;
  assign y8923 = n15684 ;
  assign y8924 = ~1'b0 ;
  assign y8925 = ~1'b0 ;
  assign y8926 = n15685 ;
  assign y8927 = n15689 ;
  assign y8928 = ~1'b0 ;
  assign y8929 = ~1'b0 ;
  assign y8930 = n15693 ;
  assign y8931 = n15695 ;
  assign y8932 = n15696 ;
  assign y8933 = ~n15700 ;
  assign y8934 = n12307 ;
  assign y8935 = ~1'b0 ;
  assign y8936 = ~1'b0 ;
  assign y8937 = ~1'b0 ;
  assign y8938 = ~1'b0 ;
  assign y8939 = ~1'b0 ;
  assign y8940 = ~n15701 ;
  assign y8941 = n635 ;
  assign y8942 = ~n15703 ;
  assign y8943 = ~1'b0 ;
  assign y8944 = n15705 ;
  assign y8945 = n15715 ;
  assign y8946 = x100 ;
  assign y8947 = ~1'b0 ;
  assign y8948 = ~n15717 ;
  assign y8949 = ~n15718 ;
  assign y8950 = n15720 ;
  assign y8951 = n15721 ;
  assign y8952 = ~n15723 ;
  assign y8953 = ~1'b0 ;
  assign y8954 = ~1'b0 ;
  assign y8955 = ~n15726 ;
  assign y8956 = ~n8462 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = n15729 ;
  assign y8959 = ~n15731 ;
  assign y8960 = ~n15734 ;
  assign y8961 = 1'b0 ;
  assign y8962 = n15735 ;
  assign y8963 = n15736 ;
  assign y8964 = ~1'b0 ;
  assign y8965 = n15737 ;
  assign y8966 = ~n15744 ;
  assign y8967 = ~n15749 ;
  assign y8968 = ~n438 ;
  assign y8969 = n15754 ;
  assign y8970 = ~1'b0 ;
  assign y8971 = ~n15756 ;
  assign y8972 = n15757 ;
  assign y8973 = ~1'b0 ;
  assign y8974 = ~1'b0 ;
  assign y8975 = n1587 ;
  assign y8976 = ~1'b0 ;
  assign y8977 = ~n15767 ;
  assign y8978 = ~1'b0 ;
  assign y8979 = n15770 ;
  assign y8980 = n15773 ;
  assign y8981 = n15775 ;
  assign y8982 = ~n15779 ;
  assign y8983 = ~n15781 ;
  assign y8984 = n15783 ;
  assign y8985 = ~n15784 ;
  assign y8986 = n15789 ;
  assign y8987 = ~n15793 ;
  assign y8988 = ~n15794 ;
  assign y8989 = ~n6030 ;
  assign y8990 = ~1'b0 ;
  assign y8991 = ~1'b0 ;
  assign y8992 = ~1'b0 ;
  assign y8993 = 1'b0 ;
  assign y8994 = n15797 ;
  assign y8995 = ~n15799 ;
  assign y8996 = ~1'b0 ;
  assign y8997 = ~n15800 ;
  assign y8998 = ~n15801 ;
  assign y8999 = ~n15804 ;
  assign y9000 = ~1'b0 ;
  assign y9001 = ~1'b0 ;
  assign y9002 = ~1'b0 ;
  assign y9003 = n15807 ;
  assign y9004 = ~n15809 ;
  assign y9005 = n15810 ;
  assign y9006 = ~n15813 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = ~n15814 ;
  assign y9010 = n15817 ;
  assign y9011 = ~n15818 ;
  assign y9012 = n15819 ;
  assign y9013 = ~n15820 ;
  assign y9014 = ~n15822 ;
  assign y9015 = ~1'b0 ;
  assign y9016 = ~n15827 ;
  assign y9017 = ~1'b0 ;
  assign y9018 = ~n15829 ;
  assign y9019 = ~n15831 ;
  assign y9020 = ~n15832 ;
  assign y9021 = ~1'b0 ;
  assign y9022 = ~n15840 ;
  assign y9023 = ~1'b0 ;
  assign y9024 = n15844 ;
  assign y9025 = 1'b0 ;
  assign y9026 = n15847 ;
  assign y9027 = ~1'b0 ;
  assign y9028 = ~1'b0 ;
  assign y9029 = ~1'b0 ;
  assign y9030 = n15851 ;
  assign y9031 = n15852 ;
  assign y9032 = ~1'b0 ;
  assign y9033 = ~1'b0 ;
  assign y9034 = n15853 ;
  assign y9035 = n15854 ;
  assign y9036 = ~1'b0 ;
  assign y9037 = ~n15855 ;
  assign y9038 = ~n15858 ;
  assign y9039 = n15859 ;
  assign y9040 = ~n15860 ;
  assign y9041 = ~n1172 ;
  assign y9042 = n15861 ;
  assign y9043 = n15865 ;
  assign y9044 = n15866 ;
  assign y9045 = n15874 ;
  assign y9046 = ~1'b0 ;
  assign y9047 = ~n15882 ;
  assign y9048 = n15890 ;
  assign y9049 = n15892 ;
  assign y9050 = n15895 ;
  assign y9051 = ~1'b0 ;
  assign y9052 = ~1'b0 ;
  assign y9053 = ~n15901 ;
  assign y9054 = ~n15903 ;
  assign y9055 = ~1'b0 ;
  assign y9056 = ~n15904 ;
  assign y9057 = ~n11973 ;
  assign y9058 = ~1'b0 ;
  assign y9059 = ~n15906 ;
  assign y9060 = n2975 ;
  assign y9061 = ~1'b0 ;
  assign y9062 = 1'b0 ;
  assign y9063 = n15907 ;
  assign y9064 = n15908 ;
  assign y9065 = n4562 ;
  assign y9066 = ~1'b0 ;
  assign y9067 = ~n15909 ;
  assign y9068 = n15910 ;
  assign y9069 = ~n15922 ;
  assign y9070 = ~n15924 ;
  assign y9071 = n15925 ;
  assign y9072 = n15927 ;
  assign y9073 = ~1'b0 ;
  assign y9074 = ~1'b0 ;
  assign y9075 = ~1'b0 ;
  assign y9076 = n13521 ;
  assign y9077 = n15932 ;
  assign y9078 = n15935 ;
  assign y9079 = n15937 ;
  assign y9080 = ~1'b0 ;
  assign y9081 = n15938 ;
  assign y9082 = 1'b0 ;
  assign y9083 = ~1'b0 ;
  assign y9084 = n15939 ;
  assign y9085 = n15943 ;
  assign y9086 = ~1'b0 ;
  assign y9087 = ~n15951 ;
  assign y9088 = ~n15953 ;
  assign y9089 = ~n15955 ;
  assign y9090 = ~1'b0 ;
  assign y9091 = ~n15956 ;
  assign y9092 = ~1'b0 ;
  assign y9093 = ~n15960 ;
  assign y9094 = ~n15964 ;
  assign y9095 = ~n15965 ;
  assign y9096 = ~n15966 ;
  assign y9097 = n15967 ;
  assign y9098 = n9393 ;
  assign y9099 = ~1'b0 ;
  assign y9100 = ~n15969 ;
  assign y9101 = n15971 ;
  assign y9102 = ~1'b0 ;
  assign y9103 = ~1'b0 ;
  assign y9104 = ~1'b0 ;
  assign y9105 = n15973 ;
  assign y9106 = ~n15974 ;
  assign y9107 = 1'b0 ;
  assign y9108 = ~n15975 ;
  assign y9109 = n15978 ;
  assign y9110 = n1016 ;
  assign y9111 = n15980 ;
  assign y9112 = ~1'b0 ;
  assign y9113 = n5203 ;
  assign y9114 = 1'b0 ;
  assign y9115 = n15985 ;
  assign y9116 = ~1'b0 ;
  assign y9117 = n15988 ;
  assign y9118 = n15991 ;
  assign y9119 = 1'b0 ;
  assign y9120 = ~1'b0 ;
  assign y9121 = n15993 ;
  assign y9122 = ~n15997 ;
  assign y9123 = n15998 ;
  assign y9124 = ~n1656 ;
  assign y9125 = n15999 ;
  assign y9126 = ~1'b0 ;
  assign y9127 = n16000 ;
  assign y9128 = ~n16003 ;
  assign y9129 = n16004 ;
  assign y9130 = ~1'b0 ;
  assign y9131 = n16005 ;
  assign y9132 = ~1'b0 ;
  assign y9133 = ~n16014 ;
  assign y9134 = ~1'b0 ;
  assign y9135 = ~1'b0 ;
  assign y9136 = ~1'b0 ;
  assign y9137 = n16015 ;
  assign y9138 = n16016 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = ~1'b0 ;
  assign y9141 = n16018 ;
  assign y9142 = ~1'b0 ;
  assign y9143 = ~n16019 ;
  assign y9144 = ~n5347 ;
  assign y9145 = ~1'b0 ;
  assign y9146 = ~1'b0 ;
  assign y9147 = 1'b0 ;
  assign y9148 = ~n16020 ;
  assign y9149 = ~1'b0 ;
  assign y9150 = ~1'b0 ;
  assign y9151 = n16025 ;
  assign y9152 = ~1'b0 ;
  assign y9153 = n16026 ;
  assign y9154 = ~1'b0 ;
  assign y9155 = n16032 ;
  assign y9156 = n1704 ;
  assign y9157 = n16033 ;
  assign y9158 = ~1'b0 ;
  assign y9159 = ~1'b0 ;
  assign y9160 = ~n16037 ;
  assign y9161 = ~n16038 ;
  assign y9162 = n16039 ;
  assign y9163 = n16041 ;
  assign y9164 = ~1'b0 ;
  assign y9165 = n16042 ;
  assign y9166 = ~1'b0 ;
  assign y9167 = ~n16045 ;
  assign y9168 = ~n10092 ;
  assign y9169 = ~1'b0 ;
  assign y9170 = x106 ;
  assign y9171 = n16048 ;
  assign y9172 = n16052 ;
  assign y9173 = n16054 ;
  assign y9174 = ~1'b0 ;
  assign y9175 = ~n16060 ;
  assign y9176 = n16065 ;
  assign y9177 = n16075 ;
  assign y9178 = ~n16077 ;
  assign y9179 = ~n16079 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = ~n16083 ;
  assign y9182 = ~n16086 ;
  assign y9183 = ~1'b0 ;
  assign y9184 = ~n16089 ;
  assign y9185 = ~1'b0 ;
  assign y9186 = n16092 ;
  assign y9187 = ~n16097 ;
  assign y9188 = n16098 ;
  assign y9189 = n16105 ;
  assign y9190 = ~n16107 ;
  assign y9191 = ~n16109 ;
  assign y9192 = n16114 ;
  assign y9193 = ~n16116 ;
  assign y9194 = ~1'b0 ;
  assign y9195 = ~1'b0 ;
  assign y9196 = n9988 ;
  assign y9197 = ~n16117 ;
  assign y9198 = ~n16119 ;
  assign y9199 = ~n16120 ;
  assign y9200 = ~1'b0 ;
  assign y9201 = n16122 ;
  assign y9202 = n16129 ;
  assign y9203 = ~1'b0 ;
  assign y9204 = ~n16130 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = n16132 ;
  assign y9207 = ~n1145 ;
  assign y9208 = n16135 ;
  assign y9209 = ~n3558 ;
  assign y9210 = 1'b0 ;
  assign y9211 = ~n16139 ;
  assign y9212 = ~1'b0 ;
  assign y9213 = ~n16144 ;
  assign y9214 = ~1'b0 ;
  assign y9215 = ~1'b0 ;
  assign y9216 = n16146 ;
  assign y9217 = n16156 ;
  assign y9218 = n16157 ;
  assign y9219 = ~n16158 ;
  assign y9220 = n16163 ;
  assign y9221 = x106 ;
  assign y9222 = ~n16164 ;
  assign y9223 = ~1'b0 ;
  assign y9224 = ~1'b0 ;
  assign y9225 = ~n16166 ;
  assign y9226 = n16168 ;
  assign y9227 = ~1'b0 ;
  assign y9228 = n16169 ;
  assign y9229 = ~n16170 ;
  assign y9230 = n16171 ;
  assign y9231 = ~1'b0 ;
  assign y9232 = ~1'b0 ;
  assign y9233 = n16172 ;
  assign y9234 = ~n16176 ;
  assign y9235 = n16177 ;
  assign y9236 = ~n16179 ;
  assign y9237 = ~n16181 ;
  assign y9238 = ~n16185 ;
  assign y9239 = n16188 ;
  assign y9240 = ~n16190 ;
  assign y9241 = ~1'b0 ;
  assign y9242 = ~n5641 ;
  assign y9243 = 1'b0 ;
  assign y9244 = ~1'b0 ;
  assign y9245 = ~1'b0 ;
  assign y9246 = ~n16202 ;
  assign y9247 = n16206 ;
  assign y9248 = ~n16209 ;
  assign y9249 = ~n16214 ;
  assign y9250 = ~n16218 ;
  assign y9251 = ~n16219 ;
  assign y9252 = ~n16226 ;
  assign y9253 = ~n16228 ;
  assign y9254 = n16229 ;
  assign y9255 = ~n16232 ;
  assign y9256 = ~1'b0 ;
  assign y9257 = ~1'b0 ;
  assign y9258 = n16234 ;
  assign y9259 = ~n16236 ;
  assign y9260 = ~n16240 ;
  assign y9261 = ~n16241 ;
  assign y9262 = ~1'b0 ;
  assign y9263 = n16242 ;
  assign y9264 = n16245 ;
  assign y9265 = ~n16246 ;
  assign y9266 = ~1'b0 ;
  assign y9267 = n16282 ;
  assign y9268 = ~1'b0 ;
  assign y9269 = n16284 ;
  assign y9270 = n16285 ;
  assign y9271 = ~1'b0 ;
  assign y9272 = n16289 ;
  assign y9273 = ~1'b0 ;
  assign y9274 = ~n16291 ;
  assign y9275 = ~n16295 ;
  assign y9276 = ~1'b0 ;
  assign y9277 = ~1'b0 ;
  assign y9278 = ~n16298 ;
  assign y9279 = n16300 ;
  assign y9280 = ~1'b0 ;
  assign y9281 = n16301 ;
  assign y9282 = n16307 ;
  assign y9283 = ~1'b0 ;
  assign y9284 = n16309 ;
  assign y9285 = ~1'b0 ;
  assign y9286 = ~n16310 ;
  assign y9287 = ~n16313 ;
  assign y9288 = ~n16314 ;
  assign y9289 = n4938 ;
  assign y9290 = ~n16317 ;
  assign y9291 = ~n16318 ;
  assign y9292 = ~n16321 ;
  assign y9293 = ~n16324 ;
  assign y9294 = n10281 ;
  assign y9295 = ~1'b0 ;
  assign y9296 = ~n16328 ;
  assign y9297 = ~n16333 ;
  assign y9298 = ~n16335 ;
  assign y9299 = n16336 ;
  assign y9300 = ~n16339 ;
  assign y9301 = n16342 ;
  assign y9302 = n16343 ;
  assign y9303 = ~1'b0 ;
  assign y9304 = ~n16344 ;
  assign y9305 = ~n16349 ;
  assign y9306 = ~1'b0 ;
  assign y9307 = n16351 ;
  assign y9308 = ~n16353 ;
  assign y9309 = n16355 ;
  assign y9310 = 1'b0 ;
  assign y9311 = n16359 ;
  assign y9312 = ~n16361 ;
  assign y9313 = ~n16362 ;
  assign y9314 = 1'b0 ;
  assign y9315 = ~1'b0 ;
  assign y9316 = ~1'b0 ;
  assign y9317 = ~1'b0 ;
  assign y9318 = n16363 ;
  assign y9319 = n16364 ;
  assign y9320 = ~n16365 ;
  assign y9321 = ~n16368 ;
  assign y9322 = n16373 ;
  assign y9323 = ~1'b0 ;
  assign y9324 = ~1'b0 ;
  assign y9325 = ~1'b0 ;
  assign y9326 = ~1'b0 ;
  assign y9327 = n16375 ;
  assign y9328 = ~n10573 ;
  assign y9329 = ~n16378 ;
  assign y9330 = ~1'b0 ;
  assign y9331 = n16379 ;
  assign y9332 = ~n16386 ;
  assign y9333 = n16389 ;
  assign y9334 = ~1'b0 ;
  assign y9335 = ~1'b0 ;
  assign y9336 = ~n16393 ;
  assign y9337 = n16395 ;
  assign y9338 = n16397 ;
  assign y9339 = ~n16400 ;
  assign y9340 = ~n16407 ;
  assign y9341 = ~n16409 ;
  assign y9342 = ~1'b0 ;
  assign y9343 = ~1'b0 ;
  assign y9344 = ~1'b0 ;
  assign y9345 = ~1'b0 ;
  assign y9346 = ~1'b0 ;
  assign y9347 = n10844 ;
  assign y9348 = ~1'b0 ;
  assign y9349 = ~n16410 ;
  assign y9350 = ~1'b0 ;
  assign y9351 = n16412 ;
  assign y9352 = 1'b0 ;
  assign y9353 = n16415 ;
  assign y9354 = n16417 ;
  assign y9355 = ~1'b0 ;
  assign y9356 = ~1'b0 ;
  assign y9357 = ~n16421 ;
  assign y9358 = ~n16424 ;
  assign y9359 = n14495 ;
  assign y9360 = ~n16427 ;
  assign y9361 = ~1'b0 ;
  assign y9362 = ~1'b0 ;
  assign y9363 = ~1'b0 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = n16434 ;
  assign y9366 = ~n16436 ;
  assign y9367 = ~n16437 ;
  assign y9368 = ~1'b0 ;
  assign y9369 = ~1'b0 ;
  assign y9370 = ~n5575 ;
  assign y9371 = ~1'b0 ;
  assign y9372 = n16440 ;
  assign y9373 = ~n16443 ;
  assign y9374 = ~1'b0 ;
  assign y9375 = n16446 ;
  assign y9376 = ~1'b0 ;
  assign y9377 = ~n16449 ;
  assign y9378 = ~1'b0 ;
  assign y9379 = ~1'b0 ;
  assign y9380 = ~1'b0 ;
  assign y9381 = n16452 ;
  assign y9382 = n16456 ;
  assign y9383 = n3781 ;
  assign y9384 = ~1'b0 ;
  assign y9385 = 1'b0 ;
  assign y9386 = ~n16457 ;
  assign y9387 = n16459 ;
  assign y9388 = n16462 ;
  assign y9389 = n16463 ;
  assign y9390 = ~1'b0 ;
  assign y9391 = ~n16466 ;
  assign y9392 = ~n16468 ;
  assign y9393 = ~1'b0 ;
  assign y9394 = n16469 ;
  assign y9395 = ~1'b0 ;
  assign y9396 = ~n16470 ;
  assign y9397 = ~1'b0 ;
  assign y9398 = n11171 ;
  assign y9399 = n16477 ;
  assign y9400 = ~n16479 ;
  assign y9401 = ~1'b0 ;
  assign y9402 = ~n16483 ;
  assign y9403 = ~n16485 ;
  assign y9404 = ~n15998 ;
  assign y9405 = n16486 ;
  assign y9406 = n16488 ;
  assign y9407 = ~1'b0 ;
  assign y9408 = ~1'b0 ;
  assign y9409 = ~1'b0 ;
  assign y9410 = ~n16490 ;
  assign y9411 = n16492 ;
  assign y9412 = ~1'b0 ;
  assign y9413 = 1'b0 ;
  assign y9414 = ~n16498 ;
  assign y9415 = ~n16500 ;
  assign y9416 = ~1'b0 ;
  assign y9417 = ~1'b0 ;
  assign y9418 = ~n16505 ;
  assign y9419 = n16512 ;
  assign y9420 = ~n11567 ;
  assign y9421 = ~1'b0 ;
  assign y9422 = ~n16515 ;
  assign y9423 = n16516 ;
  assign y9424 = ~n16517 ;
  assign y9425 = ~1'b0 ;
  assign y9426 = ~1'b0 ;
  assign y9427 = ~1'b0 ;
  assign y9428 = ~n16518 ;
  assign y9429 = ~1'b0 ;
  assign y9430 = ~n16519 ;
  assign y9431 = 1'b0 ;
  assign y9432 = ~1'b0 ;
  assign y9433 = ~1'b0 ;
  assign y9434 = ~n16525 ;
  assign y9435 = ~n16533 ;
  assign y9436 = n16545 ;
  assign y9437 = n16548 ;
  assign y9438 = ~1'b0 ;
  assign y9439 = ~1'b0 ;
  assign y9440 = ~n16552 ;
  assign y9441 = 1'b0 ;
  assign y9442 = ~n16553 ;
  assign y9443 = n2459 ;
  assign y9444 = ~n16555 ;
  assign y9445 = n16556 ;
  assign y9446 = ~1'b0 ;
  assign y9447 = ~n16557 ;
  assign y9448 = ~1'b0 ;
  assign y9449 = ~1'b0 ;
  assign y9450 = ~1'b0 ;
  assign y9451 = ~n16560 ;
  assign y9452 = n16562 ;
  assign y9453 = ~1'b0 ;
  assign y9454 = ~n16563 ;
  assign y9455 = ~n16564 ;
  assign y9456 = n7542 ;
  assign y9457 = ~1'b0 ;
  assign y9458 = ~1'b0 ;
  assign y9459 = n16567 ;
  assign y9460 = ~1'b0 ;
  assign y9461 = ~n16569 ;
  assign y9462 = ~1'b0 ;
  assign y9463 = ~n16571 ;
  assign y9464 = ~1'b0 ;
  assign y9465 = ~n16574 ;
  assign y9466 = n16576 ;
  assign y9467 = ~n16578 ;
  assign y9468 = ~n16579 ;
  assign y9469 = n16581 ;
  assign y9470 = ~n16584 ;
  assign y9471 = n16588 ;
  assign y9472 = ~1'b0 ;
  assign y9473 = n16590 ;
  assign y9474 = ~1'b0 ;
  assign y9475 = ~n16593 ;
  assign y9476 = n16596 ;
  assign y9477 = ~n16597 ;
  assign y9478 = ~n16600 ;
  assign y9479 = ~1'b0 ;
  assign y9480 = ~n16602 ;
  assign y9481 = 1'b0 ;
  assign y9482 = ~1'b0 ;
  assign y9483 = ~1'b0 ;
  assign y9484 = n16604 ;
  assign y9485 = ~1'b0 ;
  assign y9486 = ~1'b0 ;
  assign y9487 = n16606 ;
  assign y9488 = ~1'b0 ;
  assign y9489 = ~n16615 ;
  assign y9490 = n16616 ;
  assign y9491 = ~1'b0 ;
  assign y9492 = ~1'b0 ;
  assign y9493 = n16617 ;
  assign y9494 = n16619 ;
  assign y9495 = ~1'b0 ;
  assign y9496 = ~n16629 ;
  assign y9497 = n3473 ;
  assign y9498 = n16632 ;
  assign y9499 = 1'b0 ;
  assign y9500 = n16633 ;
  assign y9501 = ~n16635 ;
  assign y9502 = ~n16636 ;
  assign y9503 = n16637 ;
  assign y9504 = n16640 ;
  assign y9505 = n16642 ;
  assign y9506 = ~1'b0 ;
  assign y9507 = ~n16644 ;
  assign y9508 = ~n16645 ;
  assign y9509 = n16646 ;
  assign y9510 = ~n16648 ;
  assign y9511 = ~n16651 ;
  assign y9512 = ~n16656 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = ~1'b0 ;
  assign y9515 = ~n16657 ;
  assign y9516 = ~1'b0 ;
  assign y9517 = n4955 ;
  assign y9518 = ~1'b0 ;
  assign y9519 = ~n1268 ;
  assign y9520 = ~1'b0 ;
  assign y9521 = ~1'b0 ;
  assign y9522 = n16660 ;
  assign y9523 = n16666 ;
  assign y9524 = ~1'b0 ;
  assign y9525 = n16671 ;
  assign y9526 = n16672 ;
  assign y9527 = ~n16674 ;
  assign y9528 = ~n16676 ;
  assign y9529 = n16680 ;
  assign y9530 = ~1'b0 ;
  assign y9531 = ~1'b0 ;
  assign y9532 = n16683 ;
  assign y9533 = ~n16686 ;
  assign y9534 = n16688 ;
  assign y9535 = ~n16689 ;
  assign y9536 = n16692 ;
  assign y9537 = ~1'b0 ;
  assign y9538 = ~n16694 ;
  assign y9539 = n16695 ;
  assign y9540 = n16698 ;
  assign y9541 = n16699 ;
  assign y9542 = ~1'b0 ;
  assign y9543 = ~n16701 ;
  assign y9544 = ~n16703 ;
  assign y9545 = n16705 ;
  assign y9546 = ~n16711 ;
  assign y9547 = ~1'b0 ;
  assign y9548 = n16712 ;
  assign y9549 = ~n16713 ;
  assign y9550 = n16716 ;
  assign y9551 = ~1'b0 ;
  assign y9552 = ~n16718 ;
  assign y9553 = n16721 ;
  assign y9554 = ~n16724 ;
  assign y9555 = n16725 ;
  assign y9556 = n16726 ;
  assign y9557 = ~1'b0 ;
  assign y9558 = ~1'b0 ;
  assign y9559 = n16727 ;
  assign y9560 = ~1'b0 ;
  assign y9561 = n16730 ;
  assign y9562 = n16736 ;
  assign y9563 = ~n16737 ;
  assign y9564 = n3868 ;
  assign y9565 = ~1'b0 ;
  assign y9566 = n16741 ;
  assign y9567 = n16742 ;
  assign y9568 = n16745 ;
  assign y9569 = ~n16746 ;
  assign y9570 = ~1'b0 ;
  assign y9571 = ~1'b0 ;
  assign y9572 = ~n16749 ;
  assign y9573 = ~n16754 ;
  assign y9574 = ~x57 ;
  assign y9575 = ~1'b0 ;
  assign y9576 = n11869 ;
  assign y9577 = ~n16758 ;
  assign y9578 = n16759 ;
  assign y9579 = ~1'b0 ;
  assign y9580 = ~1'b0 ;
  assign y9581 = n16760 ;
  assign y9582 = ~1'b0 ;
  assign y9583 = ~1'b0 ;
  assign y9584 = 1'b0 ;
  assign y9585 = n3980 ;
  assign y9586 = n16762 ;
  assign y9587 = ~n16764 ;
  assign y9588 = ~n16767 ;
  assign y9589 = ~1'b0 ;
  assign y9590 = ~n16768 ;
  assign y9591 = ~1'b0 ;
  assign y9592 = ~n16770 ;
  assign y9593 = ~n16776 ;
  assign y9594 = ~1'b0 ;
  assign y9595 = ~1'b0 ;
  assign y9596 = 1'b0 ;
  assign y9597 = ~1'b0 ;
  assign y9598 = n16780 ;
  assign y9599 = ~n16783 ;
  assign y9600 = ~n16784 ;
  assign y9601 = ~1'b0 ;
  assign y9602 = ~1'b0 ;
  assign y9603 = 1'b0 ;
  assign y9604 = ~1'b0 ;
  assign y9605 = ~n16788 ;
  assign y9606 = n16789 ;
  assign y9607 = n16792 ;
  assign y9608 = ~n3862 ;
  assign y9609 = ~n16794 ;
  assign y9610 = ~1'b0 ;
  assign y9611 = ~n16799 ;
  assign y9612 = ~1'b0 ;
  assign y9613 = ~n16801 ;
  assign y9614 = ~n16805 ;
  assign y9615 = ~n16811 ;
  assign y9616 = n16814 ;
  assign y9617 = n16819 ;
  assign y9618 = n16821 ;
  assign y9619 = ~1'b0 ;
  assign y9620 = n16824 ;
  assign y9621 = n16826 ;
  assign y9622 = ~1'b0 ;
  assign y9623 = n16827 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = ~1'b0 ;
  assign y9626 = ~1'b0 ;
  assign y9627 = ~n16831 ;
  assign y9628 = n16832 ;
  assign y9629 = n16833 ;
  assign y9630 = n16835 ;
  assign y9631 = ~1'b0 ;
  assign y9632 = ~n12121 ;
  assign y9633 = ~1'b0 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~1'b0 ;
  assign y9636 = ~n16836 ;
  assign y9637 = ~1'b0 ;
  assign y9638 = ~1'b0 ;
  assign y9639 = ~1'b0 ;
  assign y9640 = n11522 ;
  assign y9641 = n16837 ;
  assign y9642 = n16839 ;
  assign y9643 = ~n16841 ;
  assign y9644 = ~1'b0 ;
  assign y9645 = ~1'b0 ;
  assign y9646 = n16842 ;
  assign y9647 = n16843 ;
  assign y9648 = ~n16849 ;
  assign y9649 = ~1'b0 ;
  assign y9650 = ~n16851 ;
  assign y9651 = ~1'b0 ;
  assign y9652 = n16853 ;
  assign y9653 = n16859 ;
  assign y9654 = ~n16860 ;
  assign y9655 = ~n16861 ;
  assign y9656 = n16862 ;
  assign y9657 = ~1'b0 ;
  assign y9658 = n16865 ;
  assign y9659 = n16867 ;
  assign y9660 = ~1'b0 ;
  assign y9661 = n16868 ;
  assign y9662 = n16872 ;
  assign y9663 = ~n16874 ;
  assign y9664 = n16878 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = n16880 ;
  assign y9667 = 1'b0 ;
  assign y9668 = ~1'b0 ;
  assign y9669 = n16882 ;
  assign y9670 = ~n16884 ;
  assign y9671 = ~n16885 ;
  assign y9672 = ~n10309 ;
  assign y9673 = ~1'b0 ;
  assign y9674 = ~1'b0 ;
  assign y9675 = 1'b0 ;
  assign y9676 = ~n7652 ;
  assign y9677 = ~1'b0 ;
  assign y9678 = ~1'b0 ;
  assign y9679 = ~n16887 ;
  assign y9680 = ~1'b0 ;
  assign y9681 = n16891 ;
  assign y9682 = ~n6108 ;
  assign y9683 = ~n16892 ;
  assign y9684 = ~n16893 ;
  assign y9685 = n16896 ;
  assign y9686 = ~1'b0 ;
  assign y9687 = n16897 ;
  assign y9688 = ~n16898 ;
  assign y9689 = ~n16900 ;
  assign y9690 = ~n3768 ;
  assign y9691 = n16902 ;
  assign y9692 = ~1'b0 ;
  assign y9693 = n16903 ;
  assign y9694 = n16910 ;
  assign y9695 = n8454 ;
  assign y9696 = ~1'b0 ;
  assign y9697 = n16920 ;
  assign y9698 = n12427 ;
  assign y9699 = ~1'b0 ;
  assign y9700 = n16923 ;
  assign y9701 = ~n2493 ;
  assign y9702 = ~n6693 ;
  assign y9703 = n16926 ;
  assign y9704 = ~n16929 ;
  assign y9705 = ~n16930 ;
  assign y9706 = ~1'b0 ;
  assign y9707 = ~1'b0 ;
  assign y9708 = 1'b0 ;
  assign y9709 = n16931 ;
  assign y9710 = ~n16938 ;
  assign y9711 = ~n16939 ;
  assign y9712 = ~n16940 ;
  assign y9713 = ~1'b0 ;
  assign y9714 = n16942 ;
  assign y9715 = n16944 ;
  assign y9716 = n16946 ;
  assign y9717 = ~1'b0 ;
  assign y9718 = n16947 ;
  assign y9719 = n16948 ;
  assign y9720 = n16951 ;
  assign y9721 = ~1'b0 ;
  assign y9722 = ~n16953 ;
  assign y9723 = n16954 ;
  assign y9724 = ~n16955 ;
  assign y9725 = ~n16961 ;
  assign y9726 = n16962 ;
  assign y9727 = n16963 ;
  assign y9728 = n6450 ;
  assign y9729 = ~n13226 ;
  assign y9730 = 1'b0 ;
  assign y9731 = ~1'b0 ;
  assign y9732 = n16964 ;
  assign y9733 = n16965 ;
  assign y9734 = n16967 ;
  assign y9735 = ~1'b0 ;
  assign y9736 = ~1'b0 ;
  assign y9737 = ~n16968 ;
  assign y9738 = n16971 ;
  assign y9739 = n16974 ;
  assign y9740 = n16976 ;
  assign y9741 = ~1'b0 ;
  assign y9742 = ~n16984 ;
  assign y9743 = n16985 ;
  assign y9744 = n16986 ;
  assign y9745 = ~1'b0 ;
  assign y9746 = ~n16990 ;
  assign y9747 = ~n16992 ;
  assign y9748 = ~1'b0 ;
  assign y9749 = n16994 ;
  assign y9750 = ~1'b0 ;
  assign y9751 = ~1'b0 ;
  assign y9752 = ~1'b0 ;
  assign y9753 = n16998 ;
  assign y9754 = ~1'b0 ;
  assign y9755 = n16999 ;
  assign y9756 = ~n17000 ;
  assign y9757 = n17002 ;
  assign y9758 = ~1'b0 ;
  assign y9759 = ~n17010 ;
  assign y9760 = ~n17011 ;
  assign y9761 = 1'b0 ;
  assign y9762 = ~n17012 ;
  assign y9763 = ~1'b0 ;
  assign y9764 = ~n17014 ;
  assign y9765 = n17015 ;
  assign y9766 = ~1'b0 ;
  assign y9767 = n17020 ;
  assign y9768 = n7411 ;
  assign y9769 = n17026 ;
  assign y9770 = n6398 ;
  assign y9771 = ~n17028 ;
  assign y9772 = ~n17029 ;
  assign y9773 = ~1'b0 ;
  assign y9774 = n17030 ;
  assign y9775 = ~1'b0 ;
  assign y9776 = n17036 ;
  assign y9777 = n17037 ;
  assign y9778 = n17039 ;
  assign y9779 = ~1'b0 ;
  assign y9780 = ~1'b0 ;
  assign y9781 = ~1'b0 ;
  assign y9782 = n17041 ;
  assign y9783 = ~n17052 ;
  assign y9784 = 1'b0 ;
  assign y9785 = n17053 ;
  assign y9786 = ~n17054 ;
  assign y9787 = n17058 ;
  assign y9788 = n17061 ;
  assign y9789 = ~n17062 ;
  assign y9790 = ~n17064 ;
  assign y9791 = ~1'b0 ;
  assign y9792 = n17066 ;
  assign y9793 = ~n17067 ;
  assign y9794 = ~1'b0 ;
  assign y9795 = ~n17068 ;
  assign y9796 = ~n2463 ;
  assign y9797 = ~1'b0 ;
  assign y9798 = n17069 ;
  assign y9799 = n17070 ;
  assign y9800 = ~n17071 ;
  assign y9801 = ~1'b0 ;
  assign y9802 = ~1'b0 ;
  assign y9803 = n17074 ;
  assign y9804 = n17076 ;
  assign y9805 = ~n17080 ;
  assign y9806 = ~n17084 ;
  assign y9807 = ~1'b0 ;
  assign y9808 = ~n17085 ;
  assign y9809 = n17088 ;
  assign y9810 = n17092 ;
  assign y9811 = ~n17093 ;
  assign y9812 = ~1'b0 ;
  assign y9813 = ~1'b0 ;
  assign y9814 = n17094 ;
  assign y9815 = n17097 ;
  assign y9816 = n17098 ;
  assign y9817 = ~n17100 ;
  assign y9818 = ~n17103 ;
  assign y9819 = n17104 ;
  assign y9820 = ~1'b0 ;
  assign y9821 = ~n17107 ;
  assign y9822 = ~1'b0 ;
  assign y9823 = ~n17108 ;
  assign y9824 = ~n13224 ;
  assign y9825 = ~1'b0 ;
  assign y9826 = ~1'b0 ;
  assign y9827 = ~1'b0 ;
  assign y9828 = n17110 ;
  assign y9829 = ~n17111 ;
  assign y9830 = n11348 ;
  assign y9831 = ~n17116 ;
  assign y9832 = ~1'b0 ;
  assign y9833 = ~1'b0 ;
  assign y9834 = n17119 ;
  assign y9835 = ~n17123 ;
  assign y9836 = ~n17124 ;
  assign y9837 = ~n1704 ;
  assign y9838 = n17132 ;
  assign y9839 = 1'b0 ;
  assign y9840 = ~1'b0 ;
  assign y9841 = ~n17135 ;
  assign y9842 = ~n17136 ;
  assign y9843 = ~1'b0 ;
  assign y9844 = ~1'b0 ;
  assign y9845 = n17137 ;
  assign y9846 = ~n17141 ;
  assign y9847 = ~1'b0 ;
  assign y9848 = ~n17145 ;
  assign y9849 = n1048 ;
  assign y9850 = ~n17146 ;
  assign y9851 = n6953 ;
  assign y9852 = ~n17147 ;
  assign y9853 = n17148 ;
  assign y9854 = ~n17152 ;
  assign y9855 = n3468 ;
  assign y9856 = n17153 ;
  assign y9857 = ~1'b0 ;
  assign y9858 = n17154 ;
  assign y9859 = n647 ;
  assign y9860 = n9238 ;
  assign y9861 = 1'b0 ;
  assign y9862 = ~n17158 ;
  assign y9863 = n17162 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = ~1'b0 ;
  assign y9866 = n17163 ;
  assign y9867 = ~1'b0 ;
  assign y9868 = n17166 ;
  assign y9869 = n17169 ;
  assign y9870 = ~n17171 ;
  assign y9871 = ~n17172 ;
  assign y9872 = n17177 ;
  assign y9873 = ~n17181 ;
  assign y9874 = ~1'b0 ;
  assign y9875 = n17182 ;
  assign y9876 = n17185 ;
  assign y9877 = n17186 ;
  assign y9878 = ~1'b0 ;
  assign y9879 = ~n17188 ;
  assign y9880 = ~1'b0 ;
  assign y9881 = ~1'b0 ;
  assign y9882 = n17189 ;
  assign y9883 = n17190 ;
  assign y9884 = ~1'b0 ;
  assign y9885 = n17192 ;
  assign y9886 = n17196 ;
  assign y9887 = ~1'b0 ;
  assign y9888 = ~1'b0 ;
  assign y9889 = n17198 ;
  assign y9890 = ~n17208 ;
  assign y9891 = ~1'b0 ;
  assign y9892 = ~1'b0 ;
  assign y9893 = n17212 ;
  assign y9894 = n17214 ;
  assign y9895 = ~n17217 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = n17221 ;
  assign y9898 = ~1'b0 ;
  assign y9899 = ~n17222 ;
  assign y9900 = ~1'b0 ;
  assign y9901 = ~n11176 ;
  assign y9902 = ~n17223 ;
  assign y9903 = n17227 ;
  assign y9904 = n17228 ;
  assign y9905 = ~n17230 ;
  assign y9906 = 1'b0 ;
  assign y9907 = ~1'b0 ;
  assign y9908 = ~1'b0 ;
  assign y9909 = ~n17232 ;
  assign y9910 = ~1'b0 ;
  assign y9911 = n17242 ;
  assign y9912 = n17244 ;
  assign y9913 = ~n17246 ;
  assign y9914 = ~n17247 ;
  assign y9915 = ~n17251 ;
  assign y9916 = 1'b0 ;
  assign y9917 = ~n17252 ;
  assign y9918 = ~n17255 ;
  assign y9919 = ~1'b0 ;
  assign y9920 = ~n17257 ;
  assign y9921 = ~n4831 ;
  assign y9922 = 1'b0 ;
  assign y9923 = ~n17262 ;
  assign y9924 = ~n17265 ;
  assign y9925 = n17269 ;
  assign y9926 = ~1'b0 ;
  assign y9927 = n17270 ;
  assign y9928 = ~n17272 ;
  assign y9929 = ~1'b0 ;
  assign y9930 = n17273 ;
  assign y9931 = ~1'b0 ;
  assign y9932 = ~n6563 ;
  assign y9933 = ~1'b0 ;
  assign y9934 = ~1'b0 ;
  assign y9935 = ~n17276 ;
  assign y9936 = ~n17277 ;
  assign y9937 = ~n17282 ;
  assign y9938 = n17286 ;
  assign y9939 = ~1'b0 ;
  assign y9940 = ~n13676 ;
  assign y9941 = n17287 ;
  assign y9942 = ~1'b0 ;
  assign y9943 = ~n17288 ;
  assign y9944 = n17292 ;
  assign y9945 = ~n17293 ;
  assign y9946 = ~1'b0 ;
  assign y9947 = ~1'b0 ;
  assign y9948 = ~1'b0 ;
  assign y9949 = ~1'b0 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = n17294 ;
  assign y9952 = ~n17295 ;
  assign y9953 = n17296 ;
  assign y9954 = ~1'b0 ;
  assign y9955 = 1'b0 ;
  assign y9956 = ~n17297 ;
  assign y9957 = ~1'b0 ;
  assign y9958 = ~n17298 ;
  assign y9959 = ~1'b0 ;
  assign y9960 = 1'b0 ;
  assign y9961 = ~n17303 ;
  assign y9962 = ~1'b0 ;
  assign y9963 = 1'b0 ;
  assign y9964 = n17304 ;
  assign y9965 = n17306 ;
  assign y9966 = ~1'b0 ;
  assign y9967 = ~1'b0 ;
  assign y9968 = ~n17308 ;
  assign y9969 = n17310 ;
  assign y9970 = ~1'b0 ;
  assign y9971 = ~1'b0 ;
  assign y9972 = 1'b0 ;
  assign y9973 = ~n17314 ;
  assign y9974 = ~1'b0 ;
  assign y9975 = n17316 ;
  assign y9976 = ~1'b0 ;
  assign y9977 = ~1'b0 ;
  assign y9978 = ~1'b0 ;
  assign y9979 = ~n17318 ;
  assign y9980 = ~n17320 ;
  assign y9981 = ~1'b0 ;
  assign y9982 = ~n17325 ;
  assign y9983 = n17331 ;
  assign y9984 = 1'b0 ;
  assign y9985 = ~n17344 ;
  assign y9986 = ~n17345 ;
  assign y9987 = ~1'b0 ;
  assign y9988 = n17346 ;
  assign y9989 = ~1'b0 ;
  assign y9990 = ~n17348 ;
  assign y9991 = ~1'b0 ;
  assign y9992 = n17354 ;
  assign y9993 = n17355 ;
  assign y9994 = ~1'b0 ;
  assign y9995 = ~1'b0 ;
  assign y9996 = ~n17357 ;
  assign y9997 = n17360 ;
  assign y9998 = n17362 ;
  assign y9999 = ~n17363 ;
  assign y10000 = ~n14463 ;
  assign y10001 = n17364 ;
  assign y10002 = ~n3747 ;
  assign y10003 = ~n17366 ;
  assign y10004 = ~1'b0 ;
  assign y10005 = ~1'b0 ;
  assign y10006 = ~1'b0 ;
  assign y10007 = n17369 ;
  assign y10008 = n17370 ;
  assign y10009 = n17372 ;
  assign y10010 = n17377 ;
  assign y10011 = n17380 ;
  assign y10012 = ~n17382 ;
  assign y10013 = n17383 ;
  assign y10014 = ~1'b0 ;
  assign y10015 = ~n17390 ;
  assign y10016 = n17391 ;
  assign y10017 = ~n17393 ;
  assign y10018 = ~n17408 ;
  assign y10019 = n17413 ;
  assign y10020 = ~n17414 ;
  assign y10021 = ~1'b0 ;
  assign y10022 = n17415 ;
  assign y10023 = ~1'b0 ;
  assign y10024 = n12805 ;
  assign y10025 = ~1'b0 ;
  assign y10026 = ~n5384 ;
  assign y10027 = ~1'b0 ;
  assign y10028 = ~1'b0 ;
  assign y10029 = ~1'b0 ;
  assign y10030 = ~n17418 ;
  assign y10031 = n17421 ;
  assign y10032 = ~n17422 ;
  assign y10033 = 1'b0 ;
  assign y10034 = ~n17423 ;
  assign y10035 = ~n17424 ;
  assign y10036 = ~1'b0 ;
  assign y10037 = ~1'b0 ;
  assign y10038 = n17425 ;
  assign y10039 = ~1'b0 ;
  assign y10040 = ~n17426 ;
  assign y10041 = n17434 ;
  assign y10042 = ~1'b0 ;
  assign y10043 = n17442 ;
  assign y10044 = ~1'b0 ;
  assign y10045 = ~n17443 ;
  assign y10046 = n17444 ;
  assign y10047 = n17448 ;
  assign y10048 = ~n17457 ;
  assign y10049 = ~1'b0 ;
  assign y10050 = ~n14994 ;
  assign y10051 = n17458 ;
  assign y10052 = n17460 ;
  assign y10053 = ~n17465 ;
  assign y10054 = ~1'b0 ;
  assign y10055 = ~n17469 ;
  assign y10056 = n17470 ;
  assign y10057 = n17473 ;
  assign y10058 = 1'b0 ;
  assign y10059 = ~1'b0 ;
  assign y10060 = ~n17477 ;
  assign y10061 = n17478 ;
  assign y10062 = ~1'b0 ;
  assign y10063 = ~1'b0 ;
  assign y10064 = ~1'b0 ;
  assign y10065 = ~n3705 ;
  assign y10066 = ~1'b0 ;
  assign y10067 = ~1'b0 ;
  assign y10068 = ~1'b0 ;
  assign y10069 = n17480 ;
  assign y10070 = n17482 ;
  assign y10071 = ~1'b0 ;
  assign y10072 = ~1'b0 ;
  assign y10073 = ~n17483 ;
  assign y10074 = ~n17484 ;
  assign y10075 = ~n17487 ;
  assign y10076 = ~n17489 ;
  assign y10077 = n17499 ;
  assign y10078 = n17501 ;
  assign y10079 = ~1'b0 ;
  assign y10080 = n17502 ;
  assign y10081 = n1588 ;
  assign y10082 = ~1'b0 ;
  assign y10083 = n10630 ;
  assign y10084 = ~n17503 ;
  assign y10085 = n17504 ;
  assign y10086 = n17505 ;
  assign y10087 = n17507 ;
  assign y10088 = ~n17508 ;
  assign y10089 = n17510 ;
  assign y10090 = ~n17514 ;
  assign y10091 = n17515 ;
  assign y10092 = ~1'b0 ;
  assign y10093 = ~n17516 ;
  assign y10094 = n4207 ;
  assign y10095 = ~1'b0 ;
  assign y10096 = ~n17521 ;
  assign y10097 = ~1'b0 ;
  assign y10098 = ~1'b0 ;
  assign y10099 = ~n17523 ;
  assign y10100 = ~1'b0 ;
  assign y10101 = ~1'b0 ;
  assign y10102 = ~n17526 ;
  assign y10103 = n13543 ;
  assign y10104 = ~1'b0 ;
  assign y10105 = ~1'b0 ;
  assign y10106 = n17529 ;
  assign y10107 = n17530 ;
  assign y10108 = n17532 ;
  assign y10109 = ~1'b0 ;
  assign y10110 = n17536 ;
  assign y10111 = ~1'b0 ;
  assign y10112 = n17544 ;
  assign y10113 = ~1'b0 ;
  assign y10114 = ~1'b0 ;
  assign y10115 = n17547 ;
  assign y10116 = 1'b0 ;
  assign y10117 = ~1'b0 ;
  assign y10118 = ~1'b0 ;
  assign y10119 = ~n17550 ;
  assign y10120 = n17554 ;
  assign y10121 = n17556 ;
  assign y10122 = n17557 ;
  assign y10123 = ~1'b0 ;
  assign y10124 = ~1'b0 ;
  assign y10125 = n17559 ;
  assign y10126 = ~1'b0 ;
  assign y10127 = n17564 ;
  assign y10128 = n17565 ;
  assign y10129 = n17567 ;
  assign y10130 = 1'b0 ;
  assign y10131 = n17568 ;
  assign y10132 = ~n17569 ;
  assign y10133 = n17572 ;
  assign y10134 = ~1'b0 ;
  assign y10135 = ~n1638 ;
  assign y10136 = ~n17575 ;
  assign y10137 = ~1'b0 ;
  assign y10138 = ~n17577 ;
  assign y10139 = ~1'b0 ;
  assign y10140 = ~n17578 ;
  assign y10141 = n17579 ;
  assign y10142 = n17582 ;
  assign y10143 = n5418 ;
  assign y10144 = ~n11262 ;
  assign y10145 = ~1'b0 ;
  assign y10146 = n17584 ;
  assign y10147 = ~n17596 ;
  assign y10148 = ~n15993 ;
  assign y10149 = n17602 ;
  assign y10150 = n17611 ;
  assign y10151 = ~n17613 ;
  assign y10152 = ~n17615 ;
  assign y10153 = ~1'b0 ;
  assign y10154 = n17620 ;
  assign y10155 = n17621 ;
  assign y10156 = n17626 ;
  assign y10157 = n17627 ;
  assign y10158 = ~n4824 ;
  assign y10159 = ~1'b0 ;
  assign y10160 = ~1'b0 ;
  assign y10161 = n17632 ;
  assign y10162 = n17633 ;
  assign y10163 = ~1'b0 ;
  assign y10164 = n17644 ;
  assign y10165 = 1'b0 ;
  assign y10166 = ~n17651 ;
  assign y10167 = ~1'b0 ;
  assign y10168 = ~1'b0 ;
  assign y10169 = ~1'b0 ;
  assign y10170 = ~n17654 ;
  assign y10171 = ~1'b0 ;
  assign y10172 = ~n17662 ;
  assign y10173 = ~n17663 ;
  assign y10174 = n17667 ;
  assign y10175 = ~1'b0 ;
  assign y10176 = ~1'b0 ;
  assign y10177 = n17669 ;
  assign y10178 = n17670 ;
  assign y10179 = ~1'b0 ;
  assign y10180 = ~1'b0 ;
  assign y10181 = ~n17672 ;
  assign y10182 = n17673 ;
  assign y10183 = n3763 ;
  assign y10184 = n17681 ;
  assign y10185 = n17683 ;
  assign y10186 = n17684 ;
  assign y10187 = ~n17691 ;
  assign y10188 = n5796 ;
  assign y10189 = ~n14528 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = n17693 ;
  assign y10192 = n17694 ;
  assign y10193 = 1'b0 ;
  assign y10194 = ~n17695 ;
  assign y10195 = ~n17696 ;
  assign y10196 = ~1'b0 ;
  assign y10197 = ~1'b0 ;
  assign y10198 = ~n17698 ;
  assign y10199 = ~n17699 ;
  assign y10200 = ~1'b0 ;
  assign y10201 = ~1'b0 ;
  assign y10202 = n13669 ;
  assign y10203 = ~1'b0 ;
  assign y10204 = n17700 ;
  assign y10205 = 1'b0 ;
  assign y10206 = n6861 ;
  assign y10207 = ~n17705 ;
  assign y10208 = ~n17711 ;
  assign y10209 = n17713 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = ~1'b0 ;
  assign y10212 = ~n1656 ;
  assign y10213 = ~n17714 ;
  assign y10214 = n17718 ;
  assign y10215 = n556 ;
  assign y10216 = n17723 ;
  assign y10217 = n5413 ;
  assign y10218 = n17724 ;
  assign y10219 = ~1'b0 ;
  assign y10220 = ~1'b0 ;
  assign y10221 = ~1'b0 ;
  assign y10222 = n17731 ;
  assign y10223 = ~1'b0 ;
  assign y10224 = ~n17734 ;
  assign y10225 = ~n17736 ;
  assign y10226 = ~n12463 ;
  assign y10227 = n7810 ;
  assign y10228 = ~n17739 ;
  assign y10229 = ~n17740 ;
  assign y10230 = n17741 ;
  assign y10231 = n17746 ;
  assign y10232 = n17747 ;
  assign y10233 = ~1'b0 ;
  assign y10234 = n17748 ;
  assign y10235 = n17749 ;
  assign y10236 = ~n17751 ;
  assign y10237 = n17753 ;
  assign y10238 = ~1'b0 ;
  assign y10239 = ~n17758 ;
  assign y10240 = ~n17759 ;
  assign y10241 = n17762 ;
  assign y10242 = n17763 ;
  assign y10243 = ~n17767 ;
  assign y10244 = n17770 ;
  assign y10245 = ~1'b0 ;
  assign y10246 = n3333 ;
  assign y10247 = n17772 ;
  assign y10248 = 1'b0 ;
  assign y10249 = n17774 ;
  assign y10250 = ~n17777 ;
  assign y10251 = n17778 ;
  assign y10252 = ~n6735 ;
  assign y10253 = ~n17781 ;
  assign y10254 = ~1'b0 ;
  assign y10255 = ~n17785 ;
  assign y10256 = ~1'b0 ;
  assign y10257 = 1'b0 ;
  assign y10258 = ~1'b0 ;
  assign y10259 = 1'b0 ;
  assign y10260 = ~1'b0 ;
  assign y10261 = ~n17789 ;
  assign y10262 = n17790 ;
  assign y10263 = ~1'b0 ;
  assign y10264 = n17791 ;
  assign y10265 = n17792 ;
  assign y10266 = ~1'b0 ;
  assign y10267 = ~n17794 ;
  assign y10268 = ~n17796 ;
  assign y10269 = ~1'b0 ;
  assign y10270 = ~n17797 ;
  assign y10271 = ~n17798 ;
  assign y10272 = ~n17800 ;
  assign y10273 = ~n17803 ;
  assign y10274 = ~n17805 ;
  assign y10275 = n17809 ;
  assign y10276 = n17819 ;
  assign y10277 = n17820 ;
  assign y10278 = n17821 ;
  assign y10279 = ~1'b0 ;
  assign y10280 = ~1'b0 ;
  assign y10281 = n17828 ;
  assign y10282 = ~1'b0 ;
  assign y10283 = ~n1920 ;
  assign y10284 = n17830 ;
  assign y10285 = ~1'b0 ;
  assign y10286 = ~n17834 ;
  assign y10287 = ~1'b0 ;
  assign y10288 = ~n17840 ;
  assign y10289 = n17842 ;
  assign y10290 = ~n7466 ;
  assign y10291 = ~n17844 ;
  assign y10292 = ~1'b0 ;
  assign y10293 = ~1'b0 ;
  assign y10294 = ~n17845 ;
  assign y10295 = ~1'b0 ;
  assign y10296 = n17849 ;
  assign y10297 = ~n17854 ;
  assign y10298 = n11258 ;
  assign y10299 = ~1'b0 ;
  assign y10300 = ~1'b0 ;
  assign y10301 = ~n17858 ;
  assign y10302 = ~1'b0 ;
  assign y10303 = n17862 ;
  assign y10304 = n17864 ;
  assign y10305 = ~1'b0 ;
  assign y10306 = ~1'b0 ;
  assign y10307 = ~1'b0 ;
  assign y10308 = n17618 ;
  assign y10309 = ~1'b0 ;
  assign y10310 = 1'b0 ;
  assign y10311 = n17868 ;
  assign y10312 = n17870 ;
  assign y10313 = ~1'b0 ;
  assign y10314 = ~1'b0 ;
  assign y10315 = ~n4493 ;
  assign y10316 = ~n17871 ;
  assign y10317 = ~1'b0 ;
  assign y10318 = ~n17872 ;
  assign y10319 = n17873 ;
  assign y10320 = n17879 ;
  assign y10321 = ~n17882 ;
  assign y10322 = ~n17885 ;
  assign y10323 = ~1'b0 ;
  assign y10324 = ~1'b0 ;
  assign y10325 = n17886 ;
  assign y10326 = ~n4075 ;
  assign y10327 = ~1'b0 ;
  assign y10328 = n17887 ;
  assign y10329 = ~n17889 ;
  assign y10330 = 1'b0 ;
  assign y10331 = ~n17894 ;
  assign y10332 = ~1'b0 ;
  assign y10333 = ~n17895 ;
  assign y10334 = ~n17896 ;
  assign y10335 = ~n17899 ;
  assign y10336 = n17900 ;
  assign y10337 = n17903 ;
  assign y10338 = ~n17906 ;
  assign y10339 = n17907 ;
  assign y10340 = ~n2668 ;
  assign y10341 = n17911 ;
  assign y10342 = ~1'b0 ;
  assign y10343 = ~n14830 ;
  assign y10344 = ~1'b0 ;
  assign y10345 = n17912 ;
  assign y10346 = n11226 ;
  assign y10347 = ~n17914 ;
  assign y10348 = ~n17915 ;
  assign y10349 = n17916 ;
  assign y10350 = n17919 ;
  assign y10351 = n17921 ;
  assign y10352 = ~n17923 ;
  assign y10353 = n17924 ;
  assign y10354 = n17925 ;
  assign y10355 = n17926 ;
  assign y10356 = n17930 ;
  assign y10357 = ~n17933 ;
  assign y10358 = ~1'b0 ;
  assign y10359 = ~1'b0 ;
  assign y10360 = ~n10044 ;
  assign y10361 = ~n17935 ;
  assign y10362 = 1'b0 ;
  assign y10363 = n17937 ;
  assign y10364 = 1'b0 ;
  assign y10365 = ~1'b0 ;
  assign y10366 = ~n17939 ;
  assign y10367 = ~n17941 ;
  assign y10368 = n17942 ;
  assign y10369 = ~n17946 ;
  assign y10370 = ~n17949 ;
  assign y10371 = ~n17950 ;
  assign y10372 = n17952 ;
  assign y10373 = ~1'b0 ;
  assign y10374 = ~n17954 ;
  assign y10375 = ~1'b0 ;
  assign y10376 = 1'b0 ;
  assign y10377 = n17955 ;
  assign y10378 = ~1'b0 ;
  assign y10379 = ~1'b0 ;
  assign y10380 = 1'b0 ;
  assign y10381 = n17957 ;
  assign y10382 = ~1'b0 ;
  assign y10383 = ~1'b0 ;
  assign y10384 = ~n17958 ;
  assign y10385 = ~1'b0 ;
  assign y10386 = n17960 ;
  assign y10387 = n17964 ;
  assign y10388 = ~1'b0 ;
  assign y10389 = ~n6189 ;
  assign y10390 = ~n17965 ;
  assign y10391 = ~n17967 ;
  assign y10392 = ~1'b0 ;
  assign y10393 = ~n17970 ;
  assign y10394 = ~1'b0 ;
  assign y10395 = ~1'b0 ;
  assign y10396 = n17978 ;
  assign y10397 = n17981 ;
  assign y10398 = ~1'b0 ;
  assign y10399 = n17985 ;
  assign y10400 = n17990 ;
  assign y10401 = ~n17991 ;
  assign y10402 = ~1'b0 ;
  assign y10403 = 1'b0 ;
  assign y10404 = n17993 ;
  assign y10405 = n17995 ;
  assign y10406 = ~1'b0 ;
  assign y10407 = ~n18004 ;
  assign y10408 = n2315 ;
  assign y10409 = n18005 ;
  assign y10410 = ~n18006 ;
  assign y10411 = 1'b0 ;
  assign y10412 = ~1'b0 ;
  assign y10413 = ~1'b0 ;
  assign y10414 = n18007 ;
  assign y10415 = ~n18012 ;
  assign y10416 = n18013 ;
  assign y10417 = n18016 ;
  assign y10418 = 1'b0 ;
  assign y10419 = ~n18024 ;
  assign y10420 = ~1'b0 ;
  assign y10421 = n18026 ;
  assign y10422 = n18030 ;
  assign y10423 = ~n18033 ;
  assign y10424 = n18034 ;
  assign y10425 = n18036 ;
  assign y10426 = n1268 ;
  assign y10427 = ~n18039 ;
  assign y10428 = ~n18041 ;
  assign y10429 = ~n18043 ;
  assign y10430 = ~n18048 ;
  assign y10431 = ~1'b0 ;
  assign y10432 = ~1'b0 ;
  assign y10433 = ~n18050 ;
  assign y10434 = ~n18051 ;
  assign y10435 = ~1'b0 ;
  assign y10436 = ~1'b0 ;
  assign y10437 = n17232 ;
  assign y10438 = n18055 ;
  assign y10439 = ~n18057 ;
  assign y10440 = ~1'b0 ;
  assign y10441 = ~n18064 ;
  assign y10442 = n18067 ;
  assign y10443 = ~1'b0 ;
  assign y10444 = ~1'b0 ;
  assign y10445 = n18070 ;
  assign y10446 = n18075 ;
  assign y10447 = n18076 ;
  assign y10448 = ~n18079 ;
  assign y10449 = n18080 ;
  assign y10450 = ~1'b0 ;
  assign y10451 = 1'b0 ;
  assign y10452 = n18082 ;
  assign y10453 = n18089 ;
  assign y10454 = n4321 ;
  assign y10455 = ~1'b0 ;
  assign y10456 = ~1'b0 ;
  assign y10457 = n13523 ;
  assign y10458 = n12345 ;
  assign y10459 = n18096 ;
  assign y10460 = ~n18098 ;
  assign y10461 = ~1'b0 ;
  assign y10462 = ~1'b0 ;
  assign y10463 = 1'b0 ;
  assign y10464 = ~1'b0 ;
  assign y10465 = ~n12095 ;
  assign y10466 = ~n18099 ;
  assign y10467 = n18101 ;
  assign y10468 = n2744 ;
  assign y10469 = ~n18102 ;
  assign y10470 = ~1'b0 ;
  assign y10471 = n18104 ;
  assign y10472 = ~n18105 ;
  assign y10473 = n18106 ;
  assign y10474 = ~1'b0 ;
  assign y10475 = ~1'b0 ;
  assign y10476 = ~n18107 ;
  assign y10477 = ~1'b0 ;
  assign y10478 = n3045 ;
  assign y10479 = n18113 ;
  assign y10480 = ~n18114 ;
  assign y10481 = n18118 ;
  assign y10482 = ~n18121 ;
  assign y10483 = n18122 ;
  assign y10484 = n18123 ;
  assign y10485 = ~n18128 ;
  assign y10486 = ~n18130 ;
  assign y10487 = ~n18131 ;
  assign y10488 = ~n18132 ;
  assign y10489 = ~1'b0 ;
  assign y10490 = ~1'b0 ;
  assign y10491 = ~1'b0 ;
  assign y10492 = ~n18133 ;
  assign y10493 = ~n18138 ;
  assign y10494 = n1298 ;
  assign y10495 = ~1'b0 ;
  assign y10496 = ~n18140 ;
  assign y10497 = ~n7467 ;
  assign y10498 = ~1'b0 ;
  assign y10499 = n18143 ;
  assign y10500 = n18145 ;
  assign y10501 = 1'b0 ;
  assign y10502 = ~1'b0 ;
  assign y10503 = n18147 ;
  assign y10504 = ~1'b0 ;
  assign y10505 = ~n18150 ;
  assign y10506 = ~n18152 ;
  assign y10507 = n18153 ;
  assign y10508 = n8889 ;
  assign y10509 = ~n18154 ;
  assign y10510 = ~n18155 ;
  assign y10511 = ~1'b0 ;
  assign y10512 = n18161 ;
  assign y10513 = ~1'b0 ;
  assign y10514 = ~1'b0 ;
  assign y10515 = ~n18162 ;
  assign y10516 = ~1'b0 ;
  assign y10517 = ~1'b0 ;
  assign y10518 = n18164 ;
  assign y10519 = n18171 ;
  assign y10520 = ~n18175 ;
  assign y10521 = ~1'b0 ;
  assign y10522 = ~n18176 ;
  assign y10523 = ~1'b0 ;
  assign y10524 = ~n18179 ;
  assign y10525 = ~1'b0 ;
  assign y10526 = n18180 ;
  assign y10527 = ~n18182 ;
  assign y10528 = ~n18183 ;
  assign y10529 = ~1'b0 ;
  assign y10530 = ~n18185 ;
  assign y10531 = ~1'b0 ;
  assign y10532 = n18186 ;
  assign y10533 = 1'b0 ;
  assign y10534 = n18190 ;
  assign y10535 = n18198 ;
  assign y10536 = 1'b0 ;
  assign y10537 = ~n18202 ;
  assign y10538 = ~1'b0 ;
  assign y10539 = ~n18208 ;
  assign y10540 = ~n18212 ;
  assign y10541 = n18217 ;
  assign y10542 = ~1'b0 ;
  assign y10543 = ~n18219 ;
  assign y10544 = ~n18222 ;
  assign y10545 = ~n18224 ;
  assign y10546 = n18228 ;
  assign y10547 = ~1'b0 ;
  assign y10548 = ~n18231 ;
  assign y10549 = ~n12616 ;
  assign y10550 = n18235 ;
  assign y10551 = ~1'b0 ;
  assign y10552 = n18237 ;
  assign y10553 = n18239 ;
  assign y10554 = n18240 ;
  assign y10555 = ~n18244 ;
  assign y10556 = ~1'b0 ;
  assign y10557 = ~n18245 ;
  assign y10558 = ~1'b0 ;
  assign y10559 = ~n18246 ;
  assign y10560 = n18247 ;
  assign y10561 = n10259 ;
  assign y10562 = ~n18249 ;
  assign y10563 = ~1'b0 ;
  assign y10564 = ~1'b0 ;
  assign y10565 = ~n17350 ;
  assign y10566 = ~n18251 ;
  assign y10567 = ~n16517 ;
  assign y10568 = n18254 ;
  assign y10569 = n18255 ;
  assign y10570 = ~1'b0 ;
  assign y10571 = ~n18256 ;
  assign y10572 = ~n13286 ;
  assign y10573 = ~n18258 ;
  assign y10574 = ~n18262 ;
  assign y10575 = n18264 ;
  assign y10576 = n18265 ;
  assign y10577 = ~1'b0 ;
  assign y10578 = n18266 ;
  assign y10579 = ~n18274 ;
  assign y10580 = ~1'b0 ;
  assign y10581 = n18275 ;
  assign y10582 = ~n978 ;
  assign y10583 = ~1'b0 ;
  assign y10584 = n18278 ;
  assign y10585 = n18279 ;
  assign y10586 = 1'b0 ;
  assign y10587 = n18280 ;
  assign y10588 = ~1'b0 ;
  assign y10589 = ~n18281 ;
  assign y10590 = n18283 ;
  assign y10591 = n18284 ;
  assign y10592 = n18285 ;
  assign y10593 = 1'b0 ;
  assign y10594 = ~1'b0 ;
  assign y10595 = n18288 ;
  assign y10596 = ~n18289 ;
  assign y10597 = ~n3303 ;
  assign y10598 = ~n18291 ;
  assign y10599 = ~1'b0 ;
  assign y10600 = n18292 ;
  assign y10601 = ~1'b0 ;
  assign y10602 = n18293 ;
  assign y10603 = n18294 ;
  assign y10604 = ~n18295 ;
  assign y10605 = n18300 ;
  assign y10606 = n18311 ;
  assign y10607 = n18312 ;
  assign y10608 = 1'b0 ;
  assign y10609 = ~1'b0 ;
  assign y10610 = ~n18315 ;
  assign y10611 = n18317 ;
  assign y10612 = ~1'b0 ;
  assign y10613 = ~n18319 ;
  assign y10614 = n18326 ;
  assign y10615 = n18327 ;
  assign y10616 = n18330 ;
  assign y10617 = n7266 ;
  assign y10618 = ~1'b0 ;
  assign y10619 = ~1'b0 ;
  assign y10620 = n18331 ;
  assign y10621 = ~1'b0 ;
  assign y10622 = ~1'b0 ;
  assign y10623 = ~n18334 ;
  assign y10624 = ~1'b0 ;
  assign y10625 = ~n18336 ;
  assign y10626 = n18337 ;
  assign y10627 = n405 ;
  assign y10628 = n18340 ;
  assign y10629 = n18342 ;
  assign y10630 = ~n18344 ;
  assign y10631 = n18346 ;
  assign y10632 = ~n18348 ;
  assign y10633 = ~n18351 ;
  assign y10634 = ~1'b0 ;
  assign y10635 = ~1'b0 ;
  assign y10636 = ~n18353 ;
  assign y10637 = ~1'b0 ;
  assign y10638 = ~n18356 ;
  assign y10639 = ~1'b0 ;
  assign y10640 = ~1'b0 ;
  assign y10641 = ~n11252 ;
  assign y10642 = ~n18359 ;
  assign y10643 = ~n4734 ;
  assign y10644 = ~n7685 ;
  assign y10645 = ~n18368 ;
  assign y10646 = ~n18371 ;
  assign y10647 = ~n18375 ;
  assign y10648 = ~n18377 ;
  assign y10649 = ~n18379 ;
  assign y10650 = n18383 ;
  assign y10651 = n18386 ;
  assign y10652 = ~n18388 ;
  assign y10653 = ~n18389 ;
  assign y10654 = ~n2466 ;
  assign y10655 = ~n18390 ;
  assign y10656 = ~n18394 ;
  assign y10657 = ~n18396 ;
  assign y10658 = ~1'b0 ;
  assign y10659 = ~1'b0 ;
  assign y10660 = ~n18397 ;
  assign y10661 = ~n18400 ;
  assign y10662 = n18401 ;
  assign y10663 = ~1'b0 ;
  assign y10664 = ~n18402 ;
  assign y10665 = ~n18404 ;
  assign y10666 = ~n18405 ;
  assign y10667 = 1'b0 ;
  assign y10668 = ~1'b0 ;
  assign y10669 = n18409 ;
  assign y10670 = n18413 ;
  assign y10671 = ~1'b0 ;
  assign y10672 = ~1'b0 ;
  assign y10673 = ~1'b0 ;
  assign y10674 = ~1'b0 ;
  assign y10675 = ~1'b0 ;
  assign y10676 = n18415 ;
  assign y10677 = ~n5101 ;
  assign y10678 = ~n18418 ;
  assign y10679 = ~n18419 ;
  assign y10680 = 1'b0 ;
  assign y10681 = ~n18420 ;
  assign y10682 = ~n11004 ;
  assign y10683 = ~n18425 ;
  assign y10684 = ~n18431 ;
  assign y10685 = ~1'b0 ;
  assign y10686 = n18433 ;
  assign y10687 = ~n18434 ;
  assign y10688 = ~1'b0 ;
  assign y10689 = ~1'b0 ;
  assign y10690 = ~1'b0 ;
  assign y10691 = ~1'b0 ;
  assign y10692 = ~n18438 ;
  assign y10693 = ~1'b0 ;
  assign y10694 = ~n18439 ;
  assign y10695 = ~n18440 ;
  assign y10696 = ~n18442 ;
  assign y10697 = 1'b0 ;
  assign y10698 = ~1'b0 ;
  assign y10699 = ~1'b0 ;
  assign y10700 = n18443 ;
  assign y10701 = n18444 ;
  assign y10702 = ~n18449 ;
  assign y10703 = ~1'b0 ;
  assign y10704 = ~n18453 ;
  assign y10705 = ~n18454 ;
  assign y10706 = ~1'b0 ;
  assign y10707 = ~n18455 ;
  assign y10708 = ~1'b0 ;
  assign y10709 = n18456 ;
  assign y10710 = ~n18458 ;
  assign y10711 = ~n18462 ;
  assign y10712 = ~n18465 ;
  assign y10713 = 1'b0 ;
  assign y10714 = ~n18467 ;
  assign y10715 = ~1'b0 ;
  assign y10716 = 1'b0 ;
  assign y10717 = ~1'b0 ;
  assign y10718 = ~1'b0 ;
  assign y10719 = n18470 ;
  assign y10720 = ~n18471 ;
  assign y10721 = n18473 ;
  assign y10722 = n1969 ;
  assign y10723 = ~1'b0 ;
  assign y10724 = n18474 ;
  assign y10725 = ~1'b0 ;
  assign y10726 = ~1'b0 ;
  assign y10727 = ~1'b0 ;
  assign y10728 = 1'b0 ;
  assign y10729 = ~1'b0 ;
  assign y10730 = n2906 ;
  assign y10731 = ~1'b0 ;
  assign y10732 = ~n18476 ;
  assign y10733 = 1'b0 ;
  assign y10734 = ~1'b0 ;
  assign y10735 = n18481 ;
  assign y10736 = n18482 ;
  assign y10737 = n18484 ;
  assign y10738 = n18485 ;
  assign y10739 = ~n18486 ;
  assign y10740 = n18489 ;
  assign y10741 = n18491 ;
  assign y10742 = ~n18492 ;
  assign y10743 = n18498 ;
  assign y10744 = ~n18500 ;
  assign y10745 = ~1'b0 ;
  assign y10746 = ~1'b0 ;
  assign y10747 = ~1'b0 ;
  assign y10748 = ~n18504 ;
  assign y10749 = n3348 ;
  assign y10750 = ~n18506 ;
  assign y10751 = ~1'b0 ;
  assign y10752 = ~1'b0 ;
  assign y10753 = ~n18512 ;
  assign y10754 = ~1'b0 ;
  assign y10755 = n18513 ;
  assign y10756 = ~n18515 ;
  assign y10757 = ~n18517 ;
  assign y10758 = ~n18520 ;
  assign y10759 = n18521 ;
  assign y10760 = ~1'b0 ;
  assign y10761 = ~n18523 ;
  assign y10762 = n10988 ;
  assign y10763 = ~1'b0 ;
  assign y10764 = ~n4232 ;
  assign y10765 = n18524 ;
  assign y10766 = ~n18529 ;
  assign y10767 = n18530 ;
  assign y10768 = 1'b0 ;
  assign y10769 = ~n18531 ;
  assign y10770 = ~n18535 ;
  assign y10771 = ~1'b0 ;
  assign y10772 = ~1'b0 ;
  assign y10773 = ~n18537 ;
  assign y10774 = ~1'b0 ;
  assign y10775 = ~1'b0 ;
  assign y10776 = ~1'b0 ;
  assign y10777 = n18541 ;
  assign y10778 = ~n18543 ;
  assign y10779 = ~1'b0 ;
  assign y10780 = ~n18545 ;
  assign y10781 = n18552 ;
  assign y10782 = ~1'b0 ;
  assign y10783 = n18553 ;
  assign y10784 = n18554 ;
  assign y10785 = ~n18555 ;
  assign y10786 = ~n13958 ;
  assign y10787 = n18558 ;
  assign y10788 = ~1'b0 ;
  assign y10789 = ~n18561 ;
  assign y10790 = ~1'b0 ;
  assign y10791 = ~n18563 ;
  assign y10792 = 1'b0 ;
  assign y10793 = ~n18566 ;
  assign y10794 = ~n9860 ;
  assign y10795 = n18571 ;
  assign y10796 = n18572 ;
  assign y10797 = n18573 ;
  assign y10798 = ~n18574 ;
  assign y10799 = ~1'b0 ;
  assign y10800 = ~n18580 ;
  assign y10801 = n18582 ;
  assign y10802 = n18584 ;
  assign y10803 = n18585 ;
  assign y10804 = ~1'b0 ;
  assign y10805 = ~n18589 ;
  assign y10806 = n9832 ;
  assign y10807 = ~n18595 ;
  assign y10808 = ~n18597 ;
  assign y10809 = ~n9965 ;
  assign y10810 = ~n18598 ;
  assign y10811 = ~n18599 ;
  assign y10812 = n18603 ;
  assign y10813 = ~n18604 ;
  assign y10814 = ~n18607 ;
  assign y10815 = ~n18611 ;
  assign y10816 = ~n18615 ;
  assign y10817 = n6558 ;
  assign y10818 = ~n18620 ;
  assign y10819 = 1'b0 ;
  assign y10820 = ~1'b0 ;
  assign y10821 = 1'b0 ;
  assign y10822 = ~n18623 ;
  assign y10823 = ~n4493 ;
  assign y10824 = n18626 ;
  assign y10825 = n18630 ;
  assign y10826 = n18634 ;
  assign y10827 = ~1'b0 ;
  assign y10828 = ~n18636 ;
  assign y10829 = ~1'b0 ;
  assign y10830 = ~1'b0 ;
  assign y10831 = ~1'b0 ;
  assign y10832 = ~1'b0 ;
  assign y10833 = n18638 ;
  assign y10834 = ~n18641 ;
  assign y10835 = n18646 ;
  assign y10836 = ~n18648 ;
  assign y10837 = ~1'b0 ;
  assign y10838 = n18649 ;
  assign y10839 = n18651 ;
  assign y10840 = n18661 ;
  assign y10841 = n1608 ;
  assign y10842 = ~1'b0 ;
  assign y10843 = ~n18663 ;
  assign y10844 = ~n11800 ;
  assign y10845 = ~1'b0 ;
  assign y10846 = n18664 ;
  assign y10847 = n18665 ;
  assign y10848 = ~1'b0 ;
  assign y10849 = n18666 ;
  assign y10850 = ~1'b0 ;
  assign y10851 = ~n18671 ;
  assign y10852 = ~1'b0 ;
  assign y10853 = ~1'b0 ;
  assign y10854 = ~n18672 ;
  assign y10855 = ~n18673 ;
  assign y10856 = 1'b0 ;
  assign y10857 = 1'b0 ;
  assign y10858 = ~1'b0 ;
  assign y10859 = ~1'b0 ;
  assign y10860 = ~1'b0 ;
  assign y10861 = n18679 ;
  assign y10862 = ~n13542 ;
  assign y10863 = ~n18682 ;
  assign y10864 = n18684 ;
  assign y10865 = n18685 ;
  assign y10866 = n18686 ;
  assign y10867 = ~n18687 ;
  assign y10868 = n18688 ;
  assign y10869 = ~n18689 ;
  assign y10870 = n18690 ;
  assign y10871 = n18691 ;
  assign y10872 = ~n18693 ;
  assign y10873 = ~1'b0 ;
  assign y10874 = ~n18694 ;
  assign y10875 = n18696 ;
  assign y10876 = n18698 ;
  assign y10877 = n18702 ;
  assign y10878 = n18704 ;
  assign y10879 = ~1'b0 ;
  assign y10880 = n18705 ;
  assign y10881 = n18706 ;
  assign y10882 = ~n18707 ;
  assign y10883 = ~1'b0 ;
  assign y10884 = ~n18711 ;
  assign y10885 = ~1'b0 ;
  assign y10886 = ~n18715 ;
  assign y10887 = ~n1099 ;
  assign y10888 = ~1'b0 ;
  assign y10889 = 1'b0 ;
  assign y10890 = ~1'b0 ;
  assign y10891 = n18717 ;
  assign y10892 = n18721 ;
  assign y10893 = n18729 ;
  assign y10894 = ~1'b0 ;
  assign y10895 = ~1'b0 ;
  assign y10896 = ~n18737 ;
  assign y10897 = n18739 ;
  assign y10898 = ~n18740 ;
  assign y10899 = ~1'b0 ;
  assign y10900 = ~n18742 ;
  assign y10901 = n18744 ;
  assign y10902 = n1404 ;
  assign y10903 = ~n18749 ;
  assign y10904 = n18341 ;
  assign y10905 = ~1'b0 ;
  assign y10906 = ~1'b0 ;
  assign y10907 = n18750 ;
  assign y10908 = ~1'b0 ;
  assign y10909 = n18751 ;
  assign y10910 = n18757 ;
  assign y10911 = n18759 ;
  assign y10912 = ~1'b0 ;
  assign y10913 = n18764 ;
  assign y10914 = ~n18767 ;
  assign y10915 = ~1'b0 ;
  assign y10916 = n18771 ;
  assign y10917 = ~n18772 ;
  assign y10918 = n18778 ;
  assign y10919 = n18779 ;
  assign y10920 = ~n18780 ;
  assign y10921 = ~1'b0 ;
  assign y10922 = n18781 ;
  assign y10923 = ~n18784 ;
  assign y10924 = ~1'b0 ;
  assign y10925 = ~1'b0 ;
  assign y10926 = ~n18786 ;
  assign y10927 = ~1'b0 ;
  assign y10928 = n18787 ;
  assign y10929 = ~1'b0 ;
  assign y10930 = n18788 ;
  assign y10931 = ~n18794 ;
  assign y10932 = ~1'b0 ;
  assign y10933 = ~n18799 ;
  assign y10934 = ~n18800 ;
  assign y10935 = n18802 ;
  assign y10936 = ~n18804 ;
  assign y10937 = ~1'b0 ;
  assign y10938 = n18806 ;
  assign y10939 = ~n18807 ;
  assign y10940 = ~x130 ;
  assign y10941 = ~1'b0 ;
  assign y10942 = n18810 ;
  assign y10943 = ~1'b0 ;
  assign y10944 = ~1'b0 ;
  assign y10945 = n18811 ;
  assign y10946 = n18814 ;
  assign y10947 = n18816 ;
  assign y10948 = n18818 ;
  assign y10949 = ~1'b0 ;
  assign y10950 = n18826 ;
  assign y10951 = ~1'b0 ;
  assign y10952 = ~1'b0 ;
  assign y10953 = n12201 ;
  assign y10954 = n3297 ;
  assign y10955 = n5615 ;
  assign y10956 = ~n18830 ;
  assign y10957 = n18831 ;
  assign y10958 = n17562 ;
  assign y10959 = ~n18355 ;
  assign y10960 = ~1'b0 ;
  assign y10961 = ~n18832 ;
  assign y10962 = ~n18833 ;
  assign y10963 = n18834 ;
  assign y10964 = ~1'b0 ;
  assign y10965 = n18835 ;
  assign y10966 = n18836 ;
  assign y10967 = n18838 ;
  assign y10968 = ~1'b0 ;
  assign y10969 = n18840 ;
  assign y10970 = ~1'b0 ;
  assign y10971 = ~n18842 ;
  assign y10972 = ~1'b0 ;
  assign y10973 = n18848 ;
  assign y10974 = ~n18859 ;
  assign y10975 = ~1'b0 ;
  assign y10976 = ~1'b0 ;
  assign y10977 = n891 ;
  assign y10978 = ~1'b0 ;
  assign y10979 = ~1'b0 ;
  assign y10980 = n18862 ;
  assign y10981 = ~1'b0 ;
  assign y10982 = n18863 ;
  assign y10983 = ~n18864 ;
  assign y10984 = n18865 ;
  assign y10985 = ~n18868 ;
  assign y10986 = ~1'b0 ;
  assign y10987 = ~1'b0 ;
  assign y10988 = ~1'b0 ;
  assign y10989 = ~1'b0 ;
  assign y10990 = n5002 ;
  assign y10991 = ~n18869 ;
  assign y10992 = ~1'b0 ;
  assign y10993 = ~1'b0 ;
  assign y10994 = ~1'b0 ;
  assign y10995 = ~1'b0 ;
  assign y10996 = n18874 ;
  assign y10997 = n18876 ;
  assign y10998 = ~n18877 ;
  assign y10999 = 1'b0 ;
  assign y11000 = n18878 ;
  assign y11001 = n18879 ;
  assign y11002 = n18880 ;
  assign y11003 = ~1'b0 ;
  assign y11004 = n18881 ;
  assign y11005 = ~n11392 ;
  assign y11006 = n18883 ;
  assign y11007 = ~n18885 ;
  assign y11008 = ~n18891 ;
  assign y11009 = n18892 ;
  assign y11010 = ~1'b0 ;
  assign y11011 = ~1'b0 ;
  assign y11012 = ~n18893 ;
  assign y11013 = n7681 ;
  assign y11014 = ~n18898 ;
  assign y11015 = ~n18899 ;
  assign y11016 = ~n18901 ;
  assign y11017 = ~n18904 ;
  assign y11018 = n18908 ;
  assign y11019 = ~n18911 ;
  assign y11020 = ~n18912 ;
  assign y11021 = n2737 ;
  assign y11022 = ~1'b0 ;
  assign y11023 = n5196 ;
  assign y11024 = n18913 ;
  assign y11025 = n18914 ;
  assign y11026 = ~n18919 ;
  assign y11027 = n18922 ;
  assign y11028 = ~1'b0 ;
  assign y11029 = n18924 ;
  assign y11030 = ~n18925 ;
  assign y11031 = ~1'b0 ;
  assign y11032 = ~n18926 ;
  assign y11033 = ~n18930 ;
  assign y11034 = ~1'b0 ;
  assign y11035 = ~n8956 ;
  assign y11036 = 1'b0 ;
  assign y11037 = n18932 ;
  assign y11038 = n18933 ;
  assign y11039 = ~1'b0 ;
  assign y11040 = n18940 ;
  assign y11041 = n18942 ;
  assign y11042 = ~n18947 ;
  assign y11043 = n18949 ;
  assign y11044 = n5411 ;
  assign y11045 = ~1'b0 ;
  assign y11046 = ~n18951 ;
  assign y11047 = n12213 ;
  assign y11048 = n18953 ;
  assign y11049 = ~n18958 ;
  assign y11050 = n18961 ;
  assign y11051 = ~1'b0 ;
  assign y11052 = 1'b0 ;
  assign y11053 = ~1'b0 ;
  assign y11054 = n18971 ;
  assign y11055 = ~n18976 ;
  assign y11056 = ~n7463 ;
  assign y11057 = ~1'b0 ;
  assign y11058 = n18977 ;
  assign y11059 = 1'b0 ;
  assign y11060 = ~1'b0 ;
  assign y11061 = n18978 ;
  assign y11062 = n18981 ;
  assign y11063 = ~1'b0 ;
  assign y11064 = ~x238 ;
  assign y11065 = n18983 ;
  assign y11066 = n18988 ;
  assign y11067 = n18995 ;
  assign y11068 = n7353 ;
  assign y11069 = ~1'b0 ;
  assign y11070 = ~1'b0 ;
  assign y11071 = ~n18999 ;
  assign y11072 = ~n19000 ;
  assign y11073 = ~n19003 ;
  assign y11074 = ~n19006 ;
  assign y11075 = ~1'b0 ;
  assign y11076 = ~n6389 ;
  assign y11077 = 1'b0 ;
  assign y11078 = n19009 ;
  assign y11079 = ~n19012 ;
  assign y11080 = ~n19015 ;
  assign y11081 = n19016 ;
  assign y11082 = ~n19018 ;
  assign y11083 = n19024 ;
  assign y11084 = n3760 ;
  assign y11085 = ~n19025 ;
  assign y11086 = n19026 ;
  assign y11087 = ~n19030 ;
  assign y11088 = n19032 ;
  assign y11089 = ~1'b0 ;
  assign y11090 = n5484 ;
  assign y11091 = ~1'b0 ;
  assign y11092 = n19033 ;
  assign y11093 = n19035 ;
  assign y11094 = ~n19038 ;
  assign y11095 = ~1'b0 ;
  assign y11096 = n19041 ;
  assign y11097 = ~1'b0 ;
  assign y11098 = ~1'b0 ;
  assign y11099 = ~1'b0 ;
  assign y11100 = ~n19043 ;
  assign y11101 = ~n19044 ;
  assign y11102 = ~1'b0 ;
  assign y11103 = n19048 ;
  assign y11104 = ~1'b0 ;
  assign y11105 = ~1'b0 ;
  assign y11106 = ~n19053 ;
  assign y11107 = ~n19055 ;
  assign y11108 = ~n19056 ;
  assign y11109 = ~1'b0 ;
  assign y11110 = ~1'b0 ;
  assign y11111 = ~n19057 ;
  assign y11112 = n19058 ;
  assign y11113 = ~1'b0 ;
  assign y11114 = ~1'b0 ;
  assign y11115 = ~n19060 ;
  assign y11116 = n19061 ;
  assign y11117 = n19062 ;
  assign y11118 = ~n19063 ;
  assign y11119 = n5818 ;
  assign y11120 = ~1'b0 ;
  assign y11121 = n19067 ;
  assign y11122 = ~n19072 ;
  assign y11123 = ~n19074 ;
  assign y11124 = ~n19079 ;
  assign y11125 = n19081 ;
  assign y11126 = ~1'b0 ;
  assign y11127 = ~n19082 ;
  assign y11128 = n5869 ;
  assign y11129 = ~n19083 ;
  assign y11130 = ~1'b0 ;
  assign y11131 = ~1'b0 ;
  assign y11132 = n19092 ;
  assign y11133 = ~1'b0 ;
  assign y11134 = n19095 ;
  assign y11135 = n19097 ;
  assign y11136 = ~n19099 ;
  assign y11137 = n7484 ;
  assign y11138 = n19101 ;
  assign y11139 = ~n19102 ;
  assign y11140 = ~n19104 ;
  assign y11141 = 1'b0 ;
  assign y11142 = n19106 ;
  assign y11143 = ~1'b0 ;
  assign y11144 = n19107 ;
  assign y11145 = ~n19112 ;
  assign y11146 = n19117 ;
  assign y11147 = n19119 ;
  assign y11148 = n19121 ;
  assign y11149 = n5354 ;
  assign y11150 = n19126 ;
  assign y11151 = ~1'b0 ;
  assign y11152 = ~1'b0 ;
  assign y11153 = ~n19131 ;
  assign y11154 = n10078 ;
  assign y11155 = ~1'b0 ;
  assign y11156 = ~n19140 ;
  assign y11157 = ~1'b0 ;
  assign y11158 = n19142 ;
  assign y11159 = 1'b0 ;
  assign y11160 = ~1'b0 ;
  assign y11161 = ~1'b0 ;
  assign y11162 = ~1'b0 ;
  assign y11163 = ~1'b0 ;
  assign y11164 = n19143 ;
  assign y11165 = ~1'b0 ;
  assign y11166 = n19144 ;
  assign y11167 = ~1'b0 ;
  assign y11168 = x180 ;
  assign y11169 = ~1'b0 ;
  assign y11170 = ~1'b0 ;
  assign y11171 = ~n19145 ;
  assign y11172 = ~1'b0 ;
  assign y11173 = ~n19146 ;
  assign y11174 = ~n19169 ;
  assign y11175 = 1'b0 ;
  assign y11176 = ~1'b0 ;
  assign y11177 = ~n10178 ;
  assign y11178 = ~n19170 ;
  assign y11179 = ~n19172 ;
  assign y11180 = ~1'b0 ;
  assign y11181 = n8192 ;
  assign y11182 = ~1'b0 ;
  assign y11183 = ~1'b0 ;
  assign y11184 = n19174 ;
  assign y11185 = n19177 ;
  assign y11186 = n19183 ;
  assign y11187 = n19184 ;
  assign y11188 = 1'b0 ;
  assign y11189 = ~1'b0 ;
  assign y11190 = ~1'b0 ;
  assign y11191 = n19186 ;
  assign y11192 = ~1'b0 ;
  assign y11193 = 1'b0 ;
  assign y11194 = 1'b0 ;
  assign y11195 = n19196 ;
  assign y11196 = ~1'b0 ;
  assign y11197 = ~n19197 ;
  assign y11198 = ~n19198 ;
  assign y11199 = n1754 ;
  assign y11200 = 1'b0 ;
  assign y11201 = ~1'b0 ;
  assign y11202 = ~1'b0 ;
  assign y11203 = ~1'b0 ;
  assign y11204 = ~1'b0 ;
  assign y11205 = ~1'b0 ;
  assign y11206 = n18900 ;
  assign y11207 = ~1'b0 ;
  assign y11208 = ~1'b0 ;
  assign y11209 = ~n19199 ;
  assign y11210 = ~n19204 ;
  assign y11211 = ~1'b0 ;
  assign y11212 = ~n19205 ;
  assign y11213 = n19208 ;
  assign y11214 = 1'b0 ;
  assign y11215 = ~n19211 ;
  assign y11216 = n19213 ;
  assign y11217 = ~n19217 ;
  assign y11218 = ~1'b0 ;
  assign y11219 = ~1'b0 ;
  assign y11220 = ~1'b0 ;
  assign y11221 = n3945 ;
  assign y11222 = ~n19220 ;
  assign y11223 = ~1'b0 ;
  assign y11224 = ~n19222 ;
  assign y11225 = ~1'b0 ;
  assign y11226 = n7937 ;
  assign y11227 = ~n8541 ;
  assign y11228 = ~1'b0 ;
  assign y11229 = 1'b0 ;
  assign y11230 = ~n19224 ;
  assign y11231 = ~1'b0 ;
  assign y11232 = ~1'b0 ;
  assign y11233 = ~n19229 ;
  assign y11234 = n1578 ;
  assign y11235 = ~n19230 ;
  assign y11236 = ~1'b0 ;
  assign y11237 = ~1'b0 ;
  assign y11238 = ~1'b0 ;
  assign y11239 = ~n19231 ;
  assign y11240 = n19232 ;
  assign y11241 = n19233 ;
  assign y11242 = n19234 ;
  assign y11243 = n19235 ;
  assign y11244 = n19236 ;
  assign y11245 = ~n4671 ;
  assign y11246 = 1'b0 ;
  assign y11247 = n19238 ;
  assign y11248 = ~1'b0 ;
  assign y11249 = ~1'b0 ;
  assign y11250 = ~n19239 ;
  assign y11251 = n19245 ;
  assign y11252 = n19249 ;
  assign y11253 = ~1'b0 ;
  assign y11254 = n9374 ;
  assign y11255 = n556 ;
  assign y11256 = ~1'b0 ;
  assign y11257 = ~1'b0 ;
  assign y11258 = n19250 ;
  assign y11259 = ~n19253 ;
  assign y11260 = 1'b0 ;
  assign y11261 = n19255 ;
  assign y11262 = n19262 ;
  assign y11263 = ~n17859 ;
  assign y11264 = n19264 ;
  assign y11265 = ~1'b0 ;
  assign y11266 = ~1'b0 ;
  assign y11267 = n11322 ;
  assign y11268 = n19266 ;
  assign y11269 = n19268 ;
  assign y11270 = ~1'b0 ;
  assign y11271 = ~n19270 ;
  assign y11272 = 1'b0 ;
  assign y11273 = 1'b0 ;
  assign y11274 = n19275 ;
  assign y11275 = n19281 ;
  assign y11276 = ~n19285 ;
  assign y11277 = ~n19286 ;
  assign y11278 = ~n19287 ;
  assign y11279 = ~1'b0 ;
  assign y11280 = ~1'b0 ;
  assign y11281 = ~n19288 ;
  assign y11282 = n5651 ;
  assign y11283 = ~n19291 ;
  assign y11284 = ~n19293 ;
  assign y11285 = ~n19299 ;
  assign y11286 = ~1'b0 ;
  assign y11287 = n19304 ;
  assign y11288 = ~n1692 ;
  assign y11289 = n19305 ;
  assign y11290 = ~n19306 ;
  assign y11291 = ~n19307 ;
  assign y11292 = n19312 ;
  assign y11293 = n19315 ;
  assign y11294 = ~1'b0 ;
  assign y11295 = n19319 ;
  assign y11296 = n19321 ;
  assign y11297 = ~n19322 ;
  assign y11298 = ~n19327 ;
  assign y11299 = ~1'b0 ;
  assign y11300 = ~1'b0 ;
  assign y11301 = ~1'b0 ;
  assign y11302 = n19328 ;
  assign y11303 = ~1'b0 ;
  assign y11304 = n19335 ;
  assign y11305 = ~n19338 ;
  assign y11306 = ~n19341 ;
  assign y11307 = ~1'b0 ;
  assign y11308 = n19344 ;
  assign y11309 = ~1'b0 ;
  assign y11310 = n19351 ;
  assign y11311 = n19356 ;
  assign y11312 = n19358 ;
  assign y11313 = n19360 ;
  assign y11314 = n19362 ;
  assign y11315 = n19368 ;
  assign y11316 = n19370 ;
  assign y11317 = ~n19372 ;
  assign y11318 = ~1'b0 ;
  assign y11319 = ~1'b0 ;
  assign y11320 = ~n19374 ;
  assign y11321 = ~1'b0 ;
  assign y11322 = ~n19383 ;
  assign y11323 = ~1'b0 ;
  assign y11324 = n19385 ;
  assign y11325 = ~n19391 ;
  assign y11326 = ~1'b0 ;
  assign y11327 = n19392 ;
  assign y11328 = n19394 ;
  assign y11329 = n19395 ;
  assign y11330 = ~n19396 ;
  assign y11331 = n19398 ;
  assign y11332 = n19400 ;
  assign y11333 = n19407 ;
  assign y11334 = ~n19409 ;
  assign y11335 = n19410 ;
  assign y11336 = ~n19412 ;
  assign y11337 = ~1'b0 ;
  assign y11338 = ~n19414 ;
  assign y11339 = ~n19416 ;
  assign y11340 = ~n19419 ;
  assign y11341 = n10638 ;
  assign y11342 = n7791 ;
  assign y11343 = ~n19420 ;
  assign y11344 = n19422 ;
  assign y11345 = n19423 ;
  assign y11346 = n19425 ;
  assign y11347 = ~1'b0 ;
  assign y11348 = ~n19427 ;
  assign y11349 = n19434 ;
  assign y11350 = ~1'b0 ;
  assign y11351 = n19435 ;
  assign y11352 = ~n19436 ;
  assign y11353 = ~1'b0 ;
  assign y11354 = ~n19438 ;
  assign y11355 = n11710 ;
  assign y11356 = n19445 ;
  assign y11357 = n19450 ;
  assign y11358 = n19452 ;
  assign y11359 = ~n19457 ;
  assign y11360 = n19459 ;
  assign y11361 = ~n19460 ;
  assign y11362 = ~1'b0 ;
  assign y11363 = ~1'b0 ;
  assign y11364 = n19468 ;
  assign y11365 = ~1'b0 ;
  assign y11366 = n19472 ;
  assign y11367 = n19475 ;
  assign y11368 = n19478 ;
  assign y11369 = n19481 ;
  assign y11370 = ~n19483 ;
  assign y11371 = ~1'b0 ;
  assign y11372 = ~n16954 ;
  assign y11373 = ~1'b0 ;
  assign y11374 = ~n19486 ;
  assign y11375 = n19488 ;
  assign y11376 = ~1'b0 ;
  assign y11377 = ~n19492 ;
  assign y11378 = n5070 ;
  assign y11379 = ~n19494 ;
  assign y11380 = ~1'b0 ;
  assign y11381 = n19501 ;
  assign y11382 = n19502 ;
  assign y11383 = n19504 ;
  assign y11384 = ~n19506 ;
  assign y11385 = ~1'b0 ;
  assign y11386 = ~1'b0 ;
  assign y11387 = ~1'b0 ;
  assign y11388 = n19507 ;
  assign y11389 = 1'b0 ;
  assign y11390 = ~n19509 ;
  assign y11391 = ~n13585 ;
  assign y11392 = ~1'b0 ;
  assign y11393 = ~n19513 ;
  assign y11394 = 1'b0 ;
  assign y11395 = ~n19516 ;
  assign y11396 = ~n2001 ;
  assign y11397 = n19519 ;
  assign y11398 = ~1'b0 ;
  assign y11399 = ~n19520 ;
  assign y11400 = n19521 ;
  assign y11401 = ~1'b0 ;
  assign y11402 = ~n19522 ;
  assign y11403 = ~1'b0 ;
  assign y11404 = ~1'b0 ;
  assign y11405 = ~n19524 ;
  assign y11406 = ~n12520 ;
  assign y11407 = n16751 ;
  assign y11408 = ~n19529 ;
  assign y11409 = ~n19530 ;
  assign y11410 = ~n19531 ;
  assign y11411 = ~1'b0 ;
  assign y11412 = ~n19534 ;
  assign y11413 = n19536 ;
  assign y11414 = ~n19547 ;
  assign y11415 = n19548 ;
  assign y11416 = ~1'b0 ;
  assign y11417 = ~1'b0 ;
  assign y11418 = n10048 ;
  assign y11419 = n19549 ;
  assign y11420 = ~n19551 ;
  assign y11421 = 1'b0 ;
  assign y11422 = ~1'b0 ;
  assign y11423 = ~1'b0 ;
  assign y11424 = n19553 ;
  assign y11425 = n19558 ;
  assign y11426 = ~n19561 ;
  assign y11427 = ~1'b0 ;
  assign y11428 = ~n19567 ;
  assign y11429 = ~n19568 ;
  assign y11430 = n19572 ;
  assign y11431 = ~1'b0 ;
  assign y11432 = ~1'b0 ;
  assign y11433 = ~n19574 ;
  assign y11434 = ~1'b0 ;
  assign y11435 = ~1'b0 ;
  assign y11436 = n16506 ;
  assign y11437 = ~n19577 ;
  assign y11438 = ~1'b0 ;
  assign y11439 = ~1'b0 ;
  assign y11440 = n19578 ;
  assign y11441 = ~1'b0 ;
  assign y11442 = ~1'b0 ;
  assign y11443 = ~n19580 ;
  assign y11444 = ~n19581 ;
  assign y11445 = ~1'b0 ;
  assign y11446 = n19585 ;
  assign y11447 = ~n19588 ;
  assign y11448 = ~n19589 ;
  assign y11449 = ~1'b0 ;
  assign y11450 = ~1'b0 ;
  assign y11451 = n19592 ;
  assign y11452 = ~1'b0 ;
  assign y11453 = ~n19593 ;
  assign y11454 = ~n19595 ;
  assign y11455 = ~n19599 ;
  assign y11456 = ~1'b0 ;
  assign y11457 = ~1'b0 ;
  assign y11458 = ~1'b0 ;
  assign y11459 = n19601 ;
  assign y11460 = ~n19604 ;
  assign y11461 = ~n19614 ;
  assign y11462 = n19615 ;
  assign y11463 = ~1'b0 ;
  assign y11464 = ~1'b0 ;
  assign y11465 = n19617 ;
  assign y11466 = n19619 ;
  assign y11467 = ~1'b0 ;
  assign y11468 = n5091 ;
  assign y11469 = ~1'b0 ;
  assign y11470 = ~1'b0 ;
  assign y11471 = ~1'b0 ;
  assign y11472 = ~1'b0 ;
  assign y11473 = ~1'b0 ;
  assign y11474 = n19620 ;
  assign y11475 = n19622 ;
  assign y11476 = 1'b0 ;
  assign y11477 = ~n19627 ;
  assign y11478 = ~n19630 ;
  assign y11479 = ~n19635 ;
  assign y11480 = ~1'b0 ;
  assign y11481 = n19637 ;
  assign y11482 = ~1'b0 ;
  assign y11483 = ~1'b0 ;
  assign y11484 = n19646 ;
  assign y11485 = ~1'b0 ;
  assign y11486 = ~1'b0 ;
  assign y11487 = ~n19653 ;
  assign y11488 = ~n5290 ;
  assign y11489 = ~n19655 ;
  assign y11490 = ~n19656 ;
  assign y11491 = ~n19665 ;
  assign y11492 = ~n19668 ;
  assign y11493 = ~n19669 ;
  assign y11494 = ~1'b0 ;
  assign y11495 = ~n19673 ;
  assign y11496 = ~1'b0 ;
  assign y11497 = n19675 ;
  assign y11498 = ~1'b0 ;
  assign y11499 = n19678 ;
  assign y11500 = n19679 ;
  assign y11501 = ~n19680 ;
  assign y11502 = ~1'b0 ;
  assign y11503 = ~n19682 ;
  assign y11504 = ~n19687 ;
  assign y11505 = ~1'b0 ;
  assign y11506 = ~n19689 ;
  assign y11507 = n19693 ;
  assign y11508 = ~n19694 ;
  assign y11509 = ~1'b0 ;
  assign y11510 = ~1'b0 ;
  assign y11511 = n19697 ;
  assign y11512 = n19698 ;
  assign y11513 = ~n8309 ;
  assign y11514 = ~n19703 ;
  assign y11515 = ~1'b0 ;
  assign y11516 = ~n19704 ;
  assign y11517 = ~1'b0 ;
  assign y11518 = ~n19707 ;
  assign y11519 = ~n19708 ;
  assign y11520 = ~n19714 ;
  assign y11521 = ~n978 ;
  assign y11522 = ~1'b0 ;
  assign y11523 = n19715 ;
  assign y11524 = ~1'b0 ;
  assign y11525 = n19716 ;
  assign y11526 = ~1'b0 ;
  assign y11527 = ~1'b0 ;
  assign y11528 = ~n19717 ;
  assign y11529 = ~n19720 ;
  assign y11530 = ~n19725 ;
  assign y11531 = n19726 ;
  assign y11532 = ~n19730 ;
  assign y11533 = ~1'b0 ;
  assign y11534 = ~n19731 ;
  assign y11535 = ~1'b0 ;
  assign y11536 = ~1'b0 ;
  assign y11537 = ~1'b0 ;
  assign y11538 = ~n19733 ;
  assign y11539 = ~n19734 ;
  assign y11540 = ~1'b0 ;
  assign y11541 = ~n19740 ;
  assign y11542 = ~1'b0 ;
  assign y11543 = ~n19747 ;
  assign y11544 = n19749 ;
  assign y11545 = ~1'b0 ;
  assign y11546 = n19750 ;
  assign y11547 = ~1'b0 ;
  assign y11548 = ~n19752 ;
  assign y11549 = ~1'b0 ;
  assign y11550 = ~1'b0 ;
  assign y11551 = ~n19753 ;
  assign y11552 = n3988 ;
  assign y11553 = ~n19754 ;
  assign y11554 = ~n19755 ;
  assign y11555 = n19760 ;
  assign y11556 = ~1'b0 ;
  assign y11557 = ~1'b0 ;
  assign y11558 = n19763 ;
  assign y11559 = n19764 ;
  assign y11560 = ~n19766 ;
  assign y11561 = ~n19770 ;
  assign y11562 = n19772 ;
  assign y11563 = ~n19774 ;
  assign y11564 = ~1'b0 ;
  assign y11565 = ~n19779 ;
  assign y11566 = ~1'b0 ;
  assign y11567 = n19791 ;
  assign y11568 = ~1'b0 ;
  assign y11569 = 1'b0 ;
  assign y11570 = ~n19798 ;
  assign y11571 = ~1'b0 ;
  assign y11572 = ~n19800 ;
  assign y11573 = ~n19803 ;
  assign y11574 = n19804 ;
  assign y11575 = n6554 ;
  assign y11576 = ~1'b0 ;
  assign y11577 = n19809 ;
  assign y11578 = ~1'b0 ;
  assign y11579 = ~1'b0 ;
  assign y11580 = ~n19811 ;
  assign y11581 = ~n19813 ;
  assign y11582 = ~n19816 ;
  assign y11583 = ~1'b0 ;
  assign y11584 = ~1'b0 ;
  assign y11585 = ~n11623 ;
  assign y11586 = 1'b0 ;
  assign y11587 = n19822 ;
  assign y11588 = ~n19824 ;
  assign y11589 = ~n19828 ;
  assign y11590 = 1'b0 ;
  assign y11591 = ~1'b0 ;
  assign y11592 = ~1'b0 ;
  assign y11593 = ~n19829 ;
  assign y11594 = n16580 ;
  assign y11595 = ~1'b0 ;
  assign y11596 = n3878 ;
  assign y11597 = n6878 ;
  assign y11598 = n19670 ;
  assign y11599 = 1'b0 ;
  assign y11600 = ~1'b0 ;
  assign y11601 = ~n579 ;
  assign y11602 = n19830 ;
  assign y11603 = ~n19831 ;
  assign y11604 = n19832 ;
  assign y11605 = n19834 ;
  assign y11606 = ~1'b0 ;
  assign y11607 = ~n19839 ;
  assign y11608 = ~1'b0 ;
  assign y11609 = n19845 ;
  assign y11610 = ~n19847 ;
  assign y11611 = ~1'b0 ;
  assign y11612 = ~1'b0 ;
  assign y11613 = n19850 ;
  assign y11614 = n19853 ;
  assign y11615 = 1'b0 ;
  assign y11616 = ~n19856 ;
  assign y11617 = n19857 ;
  assign y11618 = n4438 ;
  assign y11619 = 1'b0 ;
  assign y11620 = ~n19863 ;
  assign y11621 = ~1'b0 ;
  assign y11622 = n7652 ;
  assign y11623 = ~n19865 ;
  assign y11624 = ~n19866 ;
  assign y11625 = ~n19869 ;
  assign y11626 = ~1'b0 ;
  assign y11627 = n19870 ;
  assign y11628 = ~1'b0 ;
  assign y11629 = ~1'b0 ;
  assign y11630 = ~1'b0 ;
  assign y11631 = ~1'b0 ;
  assign y11632 = n19872 ;
  assign y11633 = ~n19873 ;
  assign y11634 = n19878 ;
  assign y11635 = ~n19879 ;
  assign y11636 = ~1'b0 ;
  assign y11637 = n19884 ;
  assign y11638 = ~1'b0 ;
  assign y11639 = n19886 ;
  assign y11640 = ~1'b0 ;
  assign y11641 = n313 ;
  assign y11642 = ~1'b0 ;
  assign y11643 = ~n19887 ;
  assign y11644 = ~n19889 ;
  assign y11645 = ~n19892 ;
  assign y11646 = n19893 ;
  assign y11647 = ~1'b0 ;
  assign y11648 = n10030 ;
  assign y11649 = n19895 ;
  assign y11650 = ~1'b0 ;
  assign y11651 = n19896 ;
  assign y11652 = ~n19897 ;
  assign y11653 = ~n562 ;
  assign y11654 = ~1'b0 ;
  assign y11655 = ~1'b0 ;
  assign y11656 = ~1'b0 ;
  assign y11657 = n19905 ;
  assign y11658 = ~1'b0 ;
  assign y11659 = n19913 ;
  assign y11660 = n19916 ;
  assign y11661 = ~1'b0 ;
  assign y11662 = ~1'b0 ;
  assign y11663 = ~1'b0 ;
  assign y11664 = ~n19917 ;
  assign y11665 = n19919 ;
  assign y11666 = n19921 ;
  assign y11667 = ~1'b0 ;
  assign y11668 = ~n19922 ;
  assign y11669 = ~1'b0 ;
  assign y11670 = n19925 ;
  assign y11671 = n13040 ;
  assign y11672 = n19927 ;
  assign y11673 = ~n19929 ;
  assign y11674 = ~1'b0 ;
  assign y11675 = ~n19931 ;
  assign y11676 = n13800 ;
  assign y11677 = n19933 ;
  assign y11678 = ~n19935 ;
  assign y11679 = ~n5965 ;
  assign y11680 = n19936 ;
  assign y11681 = ~n19939 ;
  assign y11682 = n19940 ;
  assign y11683 = ~n19945 ;
  assign y11684 = ~1'b0 ;
  assign y11685 = ~1'b0 ;
  assign y11686 = 1'b0 ;
  assign y11687 = n19948 ;
  assign y11688 = ~n19446 ;
  assign y11689 = n19951 ;
  assign y11690 = ~1'b0 ;
  assign y11691 = ~1'b0 ;
  assign y11692 = n19953 ;
  assign y11693 = n19956 ;
  assign y11694 = ~1'b0 ;
  assign y11695 = n19959 ;
  assign y11696 = ~1'b0 ;
  assign y11697 = ~n19967 ;
  assign y11698 = n18322 ;
  assign y11699 = n19968 ;
  assign y11700 = ~n19969 ;
  assign y11701 = n19975 ;
  assign y11702 = ~n1302 ;
  assign y11703 = ~n19977 ;
  assign y11704 = ~n19979 ;
  assign y11705 = ~n19982 ;
  assign y11706 = ~n19984 ;
  assign y11707 = ~1'b0 ;
  assign y11708 = n19987 ;
  assign y11709 = ~n19991 ;
  assign y11710 = n19997 ;
  assign y11711 = ~1'b0 ;
  assign y11712 = ~1'b0 ;
  assign y11713 = ~n20003 ;
  assign y11714 = ~n16033 ;
  assign y11715 = ~1'b0 ;
  assign y11716 = ~n20008 ;
  assign y11717 = ~n20011 ;
  assign y11718 = ~1'b0 ;
  assign y11719 = ~1'b0 ;
  assign y11720 = ~n20012 ;
  assign y11721 = ~n20016 ;
  assign y11722 = n20017 ;
  assign y11723 = ~1'b0 ;
  assign y11724 = ~n20021 ;
  assign y11725 = n20023 ;
  assign y11726 = ~1'b0 ;
  assign y11727 = n13505 ;
  assign y11728 = n20025 ;
  assign y11729 = n20027 ;
  assign y11730 = ~1'b0 ;
  assign y11731 = ~1'b0 ;
  assign y11732 = n20028 ;
  assign y11733 = ~n20031 ;
  assign y11734 = ~1'b0 ;
  assign y11735 = ~1'b0 ;
  assign y11736 = ~1'b0 ;
  assign y11737 = ~1'b0 ;
  assign y11738 = n20035 ;
  assign y11739 = n20069 ;
  assign y11740 = ~1'b0 ;
  assign y11741 = n20073 ;
  assign y11742 = ~x81 ;
  assign y11743 = ~1'b0 ;
  assign y11744 = ~n20077 ;
  assign y11745 = ~1'b0 ;
  assign y11746 = ~1'b0 ;
  assign y11747 = n15441 ;
  assign y11748 = ~n20078 ;
  assign y11749 = ~n20079 ;
  assign y11750 = ~n20081 ;
  assign y11751 = ~1'b0 ;
  assign y11752 = ~n20086 ;
  assign y11753 = ~1'b0 ;
  assign y11754 = ~n20089 ;
  assign y11755 = n20090 ;
  assign y11756 = ~1'b0 ;
  assign y11757 = n20091 ;
  assign y11758 = ~n20096 ;
  assign y11759 = ~n20100 ;
  assign y11760 = n20104 ;
  assign y11761 = 1'b0 ;
  assign y11762 = ~1'b0 ;
  assign y11763 = n20106 ;
  assign y11764 = n20108 ;
  assign y11765 = ~1'b0 ;
  assign y11766 = ~1'b0 ;
  assign y11767 = ~1'b0 ;
  assign y11768 = n20118 ;
  assign y11769 = ~1'b0 ;
  assign y11770 = ~n20121 ;
  assign y11771 = n20122 ;
  assign y11772 = n6974 ;
  assign y11773 = ~1'b0 ;
  assign y11774 = n20126 ;
  assign y11775 = n20130 ;
  assign y11776 = ~n20138 ;
  assign y11777 = ~n20139 ;
  assign y11778 = ~1'b0 ;
  assign y11779 = ~n20140 ;
  assign y11780 = ~1'b0 ;
  assign y11781 = 1'b0 ;
  assign y11782 = 1'b0 ;
  assign y11783 = ~1'b0 ;
  assign y11784 = n20144 ;
  assign y11785 = n20147 ;
  assign y11786 = x177 ;
  assign y11787 = ~n20150 ;
  assign y11788 = ~1'b0 ;
  assign y11789 = n6298 ;
  assign y11790 = ~n20151 ;
  assign y11791 = ~1'b0 ;
  assign y11792 = n11310 ;
  assign y11793 = ~n20153 ;
  assign y11794 = 1'b0 ;
  assign y11795 = 1'b0 ;
  assign y11796 = ~1'b0 ;
  assign y11797 = ~n20160 ;
  assign y11798 = ~1'b0 ;
  assign y11799 = ~1'b0 ;
  assign y11800 = ~1'b0 ;
  assign y11801 = ~1'b0 ;
  assign y11802 = n20161 ;
  assign y11803 = n7761 ;
  assign y11804 = ~n20168 ;
  assign y11805 = ~1'b0 ;
  assign y11806 = ~1'b0 ;
  assign y11807 = n20169 ;
  assign y11808 = ~n20170 ;
  assign y11809 = ~1'b0 ;
  assign y11810 = n20172 ;
  assign y11811 = n20174 ;
  assign y11812 = ~1'b0 ;
  assign y11813 = ~1'b0 ;
  assign y11814 = n20176 ;
  assign y11815 = ~n20179 ;
  assign y11816 = ~n741 ;
  assign y11817 = ~n20183 ;
  assign y11818 = ~n20188 ;
  assign y11819 = n20190 ;
  assign y11820 = ~n20193 ;
  assign y11821 = ~n20195 ;
  assign y11822 = ~n20204 ;
  assign y11823 = ~1'b0 ;
  assign y11824 = ~1'b0 ;
  assign y11825 = ~1'b0 ;
  assign y11826 = n20206 ;
  assign y11827 = n20210 ;
  assign y11828 = ~n20215 ;
  assign y11829 = n20218 ;
  assign y11830 = ~1'b0 ;
  assign y11831 = n20222 ;
  assign y11832 = ~n20227 ;
  assign y11833 = ~1'b0 ;
  assign y11834 = n20231 ;
  assign y11835 = ~n20233 ;
  assign y11836 = ~n20234 ;
  assign y11837 = ~1'b0 ;
  assign y11838 = ~n20236 ;
  assign y11839 = ~1'b0 ;
  assign y11840 = n20237 ;
  assign y11841 = ~n20238 ;
  assign y11842 = ~1'b0 ;
  assign y11843 = n20239 ;
  assign y11844 = n20240 ;
  assign y11845 = n13663 ;
  assign y11846 = ~1'b0 ;
  assign y11847 = ~n20247 ;
  assign y11848 = n20248 ;
  assign y11849 = ~n20252 ;
  assign y11850 = ~n20258 ;
  assign y11851 = ~n20259 ;
  assign y11852 = n20261 ;
  assign y11853 = ~1'b0 ;
  assign y11854 = n14601 ;
  assign y11855 = n1717 ;
  assign y11856 = ~1'b0 ;
  assign y11857 = ~1'b0 ;
  assign y11858 = n20265 ;
  assign y11859 = ~1'b0 ;
  assign y11860 = ~n20271 ;
  assign y11861 = n20272 ;
  assign y11862 = ~n20275 ;
  assign y11863 = ~1'b0 ;
  assign y11864 = ~n20276 ;
  assign y11865 = ~1'b0 ;
  assign y11866 = ~n20279 ;
  assign y11867 = n4075 ;
  assign y11868 = n20281 ;
  assign y11869 = 1'b0 ;
  assign y11870 = n20285 ;
  assign y11871 = n20286 ;
  assign y11872 = n20288 ;
  assign y11873 = n20289 ;
  assign y11874 = ~1'b0 ;
  assign y11875 = ~1'b0 ;
  assign y11876 = ~n20290 ;
  assign y11877 = n20291 ;
  assign y11878 = ~1'b0 ;
  assign y11879 = n20292 ;
  assign y11880 = ~1'b0 ;
  assign y11881 = n20294 ;
  assign y11882 = n20295 ;
  assign y11883 = n20301 ;
  assign y11884 = ~1'b0 ;
  assign y11885 = ~1'b0 ;
  assign y11886 = n12855 ;
  assign y11887 = ~1'b0 ;
  assign y11888 = ~1'b0 ;
  assign y11889 = ~n20306 ;
  assign y11890 = ~1'b0 ;
  assign y11891 = n20307 ;
  assign y11892 = n20308 ;
  assign y11893 = ~n12941 ;
  assign y11894 = n20309 ;
  assign y11895 = n20312 ;
  assign y11896 = 1'b0 ;
  assign y11897 = 1'b0 ;
  assign y11898 = n20314 ;
  assign y11899 = n20315 ;
  assign y11900 = ~1'b0 ;
  assign y11901 = ~1'b0 ;
  assign y11902 = ~n20316 ;
  assign y11903 = ~n20318 ;
  assign y11904 = 1'b0 ;
  assign y11905 = n20319 ;
  assign y11906 = ~1'b0 ;
  assign y11907 = ~n20321 ;
  assign y11908 = ~1'b0 ;
  assign y11909 = n20325 ;
  assign y11910 = ~n20327 ;
  assign y11911 = ~1'b0 ;
  assign y11912 = ~n20328 ;
  assign y11913 = ~n20329 ;
  assign y11914 = n20330 ;
  assign y11915 = ~1'b0 ;
  assign y11916 = n20331 ;
  assign y11917 = ~1'b0 ;
  assign y11918 = ~n20334 ;
  assign y11919 = n20335 ;
  assign y11920 = ~1'b0 ;
  assign y11921 = ~1'b0 ;
  assign y11922 = n20336 ;
  assign y11923 = ~1'b0 ;
  assign y11924 = ~n20338 ;
  assign y11925 = n20341 ;
  assign y11926 = ~1'b0 ;
  assign y11927 = ~n20343 ;
  assign y11928 = ~n20345 ;
  assign y11929 = n20346 ;
  assign y11930 = ~1'b0 ;
  assign y11931 = n20348 ;
  assign y11932 = ~1'b0 ;
  assign y11933 = ~1'b0 ;
  assign y11934 = ~1'b0 ;
  assign y11935 = ~1'b0 ;
  assign y11936 = ~1'b0 ;
  assign y11937 = n20349 ;
  assign y11938 = n20350 ;
  assign y11939 = ~n20355 ;
  assign y11940 = n20357 ;
  assign y11941 = n20358 ;
  assign y11942 = n20359 ;
  assign y11943 = ~1'b0 ;
  assign y11944 = ~1'b0 ;
  assign y11945 = ~1'b0 ;
  assign y11946 = n18883 ;
  assign y11947 = ~n20361 ;
  assign y11948 = ~1'b0 ;
  assign y11949 = ~1'b0 ;
  assign y11950 = n20368 ;
  assign y11951 = ~1'b0 ;
  assign y11952 = n6822 ;
  assign y11953 = ~n16810 ;
  assign y11954 = ~1'b0 ;
  assign y11955 = ~n20371 ;
  assign y11956 = ~1'b0 ;
  assign y11957 = 1'b0 ;
  assign y11958 = 1'b0 ;
  assign y11959 = ~n20372 ;
  assign y11960 = ~n20374 ;
  assign y11961 = n20378 ;
  assign y11962 = ~n20380 ;
  assign y11963 = n20382 ;
  assign y11964 = ~1'b0 ;
  assign y11965 = 1'b0 ;
  assign y11966 = ~n20385 ;
  assign y11967 = n20387 ;
  assign y11968 = n20389 ;
  assign y11969 = ~1'b0 ;
  assign y11970 = ~1'b0 ;
  assign y11971 = ~n20391 ;
  assign y11972 = n20392 ;
  assign y11973 = ~n20394 ;
  assign y11974 = n20396 ;
  assign y11975 = ~n20397 ;
  assign y11976 = ~1'b0 ;
  assign y11977 = ~1'b0 ;
  assign y11978 = ~n20399 ;
  assign y11979 = ~1'b0 ;
  assign y11980 = ~n20401 ;
  assign y11981 = ~1'b0 ;
  assign y11982 = ~n20402 ;
  assign y11983 = ~n20406 ;
  assign y11984 = n20408 ;
  assign y11985 = ~1'b0 ;
  assign y11986 = 1'b0 ;
  assign y11987 = 1'b0 ;
  assign y11988 = ~n20411 ;
  assign y11989 = ~1'b0 ;
  assign y11990 = ~1'b0 ;
  assign y11991 = n20416 ;
  assign y11992 = ~n1464 ;
  assign y11993 = ~1'b0 ;
  assign y11994 = ~n20418 ;
  assign y11995 = ~1'b0 ;
  assign y11996 = n3091 ;
  assign y11997 = ~n20420 ;
  assign y11998 = n20422 ;
  assign y11999 = n20423 ;
  assign y12000 = n20425 ;
  assign y12001 = n20426 ;
  assign y12002 = ~1'b0 ;
  assign y12003 = ~1'b0 ;
  assign y12004 = ~1'b0 ;
  assign y12005 = ~1'b0 ;
  assign y12006 = ~n20428 ;
  assign y12007 = 1'b0 ;
  assign y12008 = 1'b0 ;
  assign y12009 = n20433 ;
  assign y12010 = ~1'b0 ;
  assign y12011 = n20434 ;
  assign y12012 = ~n20436 ;
  assign y12013 = n20439 ;
  assign y12014 = n8830 ;
  assign y12015 = ~n20441 ;
  assign y12016 = ~n974 ;
  assign y12017 = ~1'b0 ;
  assign y12018 = ~1'b0 ;
  assign y12019 = ~1'b0 ;
  assign y12020 = n20448 ;
  assign y12021 = ~n20450 ;
  assign y12022 = n20452 ;
  assign y12023 = ~n20453 ;
  assign y12024 = ~n20454 ;
  assign y12025 = n20456 ;
  assign y12026 = n20457 ;
  assign y12027 = n20458 ;
  assign y12028 = ~n20459 ;
  assign y12029 = ~n20460 ;
  assign y12030 = n1260 ;
  assign y12031 = 1'b0 ;
  assign y12032 = n20464 ;
  assign y12033 = n20466 ;
  assign y12034 = n20468 ;
  assign y12035 = n20470 ;
  assign y12036 = ~1'b0 ;
  assign y12037 = n20471 ;
  assign y12038 = ~1'b0 ;
  assign y12039 = n20472 ;
  assign y12040 = n19030 ;
  assign y12041 = ~n20479 ;
  assign y12042 = ~1'b0 ;
  assign y12043 = ~n20480 ;
  assign y12044 = ~1'b0 ;
  assign y12045 = n20482 ;
  assign y12046 = ~n20483 ;
  assign y12047 = ~1'b0 ;
  assign y12048 = ~n20488 ;
  assign y12049 = n1836 ;
  assign y12050 = n20490 ;
  assign y12051 = ~n20493 ;
  assign y12052 = n20494 ;
  assign y12053 = ~1'b0 ;
  assign y12054 = n2991 ;
  assign y12055 = ~n20497 ;
  assign y12056 = ~1'b0 ;
  assign y12057 = n20499 ;
  assign y12058 = ~n20501 ;
  assign y12059 = ~n20503 ;
  assign y12060 = n20508 ;
  assign y12061 = n20511 ;
  assign y12062 = ~1'b0 ;
  assign y12063 = ~n20512 ;
  assign y12064 = n20516 ;
  assign y12065 = ~1'b0 ;
  assign y12066 = ~n20524 ;
  assign y12067 = ~n20525 ;
  assign y12068 = ~1'b0 ;
  assign y12069 = n20529 ;
  assign y12070 = ~1'b0 ;
  assign y12071 = ~n20531 ;
  assign y12072 = ~1'b0 ;
  assign y12073 = n20532 ;
  assign y12074 = n20533 ;
  assign y12075 = ~1'b0 ;
  assign y12076 = ~n20534 ;
  assign y12077 = ~n20551 ;
  assign y12078 = n7042 ;
  assign y12079 = ~n20553 ;
  assign y12080 = ~1'b0 ;
  assign y12081 = ~1'b0 ;
  assign y12082 = ~n20556 ;
  assign y12083 = n20559 ;
  assign y12084 = n20562 ;
  assign y12085 = n3833 ;
  assign y12086 = ~1'b0 ;
  assign y12087 = ~n20565 ;
  assign y12088 = ~n12713 ;
  assign y12089 = ~n20566 ;
  assign y12090 = 1'b0 ;
  assign y12091 = n20568 ;
  assign y12092 = ~1'b0 ;
  assign y12093 = ~n20569 ;
  assign y12094 = ~1'b0 ;
  assign y12095 = ~1'b0 ;
  assign y12096 = n20574 ;
  assign y12097 = n20576 ;
  assign y12098 = ~n20578 ;
  assign y12099 = ~n20580 ;
  assign y12100 = ~n20584 ;
  assign y12101 = ~n20585 ;
  assign y12102 = ~1'b0 ;
  assign y12103 = ~n20588 ;
  assign y12104 = ~1'b0 ;
  assign y12105 = ~1'b0 ;
  assign y12106 = ~1'b0 ;
  assign y12107 = ~n20589 ;
  assign y12108 = n20591 ;
  assign y12109 = n20594 ;
  assign y12110 = n20596 ;
  assign y12111 = n20597 ;
  assign y12112 = ~n20599 ;
  assign y12113 = ~n11083 ;
  assign y12114 = n20602 ;
  assign y12115 = n3509 ;
  assign y12116 = n20607 ;
  assign y12117 = ~1'b0 ;
  assign y12118 = n20608 ;
  assign y12119 = ~n20609 ;
  assign y12120 = ~n13818 ;
  assign y12121 = ~n20611 ;
  assign y12122 = ~n20612 ;
  assign y12123 = ~n20613 ;
  assign y12124 = ~n20617 ;
  assign y12125 = n20619 ;
  assign y12126 = n20622 ;
  assign y12127 = ~1'b0 ;
  assign y12128 = n20623 ;
  assign y12129 = 1'b0 ;
  assign y12130 = ~1'b0 ;
  assign y12131 = ~n20624 ;
  assign y12132 = ~1'b0 ;
  assign y12133 = ~n20628 ;
  assign y12134 = ~n20629 ;
  assign y12135 = ~1'b0 ;
  assign y12136 = n20630 ;
  assign y12137 = n20632 ;
  assign y12138 = n20636 ;
  assign y12139 = ~1'b0 ;
  assign y12140 = ~1'b0 ;
  assign y12141 = n20638 ;
  assign y12142 = n20639 ;
  assign y12143 = ~n20641 ;
  assign y12144 = ~n20642 ;
  assign y12145 = n20646 ;
  assign y12146 = n2744 ;
  assign y12147 = n20648 ;
  assign y12148 = n20649 ;
  assign y12149 = ~1'b0 ;
  assign y12150 = ~1'b0 ;
  assign y12151 = n20655 ;
  assign y12152 = n20657 ;
  assign y12153 = ~n20662 ;
  assign y12154 = n20663 ;
  assign y12155 = n20664 ;
  assign y12156 = ~n20677 ;
  assign y12157 = ~n1463 ;
  assign y12158 = n20679 ;
  assign y12159 = ~n20681 ;
  assign y12160 = n20684 ;
  assign y12161 = n20687 ;
  assign y12162 = ~n20688 ;
  assign y12163 = n20689 ;
  assign y12164 = n4799 ;
  assign y12165 = ~n20691 ;
  assign y12166 = ~1'b0 ;
  assign y12167 = n590 ;
  assign y12168 = ~1'b0 ;
  assign y12169 = ~1'b0 ;
  assign y12170 = n20694 ;
  assign y12171 = 1'b0 ;
  assign y12172 = ~1'b0 ;
  assign y12173 = ~n1050 ;
  assign y12174 = ~n20699 ;
  assign y12175 = ~n13759 ;
  assign y12176 = ~n20700 ;
  assign y12177 = ~1'b0 ;
  assign y12178 = ~1'b0 ;
  assign y12179 = 1'b0 ;
  assign y12180 = ~n20701 ;
  assign y12181 = ~n20702 ;
  assign y12182 = ~1'b0 ;
  assign y12183 = ~1'b0 ;
  assign y12184 = n20703 ;
  assign y12185 = ~1'b0 ;
  assign y12186 = ~1'b0 ;
  assign y12187 = ~n20704 ;
  assign y12188 = ~n20707 ;
  assign y12189 = ~x226 ;
  assign y12190 = n3666 ;
  assign y12191 = ~1'b0 ;
  assign y12192 = ~n20710 ;
  assign y12193 = ~1'b0 ;
  assign y12194 = n20712 ;
  assign y12195 = n20713 ;
  assign y12196 = n20716 ;
  assign y12197 = ~1'b0 ;
  assign y12198 = n20721 ;
  assign y12199 = ~n20731 ;
  assign y12200 = ~1'b0 ;
  assign y12201 = n20733 ;
  assign y12202 = n20734 ;
  assign y12203 = ~n20735 ;
  assign y12204 = 1'b0 ;
  assign y12205 = ~n20740 ;
  assign y12206 = ~1'b0 ;
  assign y12207 = ~n1588 ;
  assign y12208 = ~n20741 ;
  assign y12209 = n20743 ;
  assign y12210 = ~n20745 ;
  assign y12211 = 1'b0 ;
  assign y12212 = ~1'b0 ;
  assign y12213 = ~n20747 ;
  assign y12214 = ~n20748 ;
  assign y12215 = n17188 ;
  assign y12216 = ~1'b0 ;
  assign y12217 = ~n5507 ;
  assign y12218 = ~1'b0 ;
  assign y12219 = ~1'b0 ;
  assign y12220 = ~n20754 ;
  assign y12221 = ~n20755 ;
  assign y12222 = ~n20757 ;
  assign y12223 = ~n540 ;
  assign y12224 = n14863 ;
  assign y12225 = ~1'b0 ;
  assign y12226 = ~n20759 ;
  assign y12227 = ~1'b0 ;
  assign y12228 = ~n20760 ;
  assign y12229 = n3480 ;
  assign y12230 = n20761 ;
  assign y12231 = n20768 ;
  assign y12232 = ~1'b0 ;
  assign y12233 = ~1'b0 ;
  assign y12234 = ~n20769 ;
  assign y12235 = n20772 ;
  assign y12236 = ~n20775 ;
  assign y12237 = ~1'b0 ;
  assign y12238 = n20783 ;
  assign y12239 = n5955 ;
  assign y12240 = ~n20785 ;
  assign y12241 = ~1'b0 ;
  assign y12242 = ~n20786 ;
  assign y12243 = n20787 ;
  assign y12244 = n20788 ;
  assign y12245 = ~n20791 ;
  assign y12246 = ~1'b0 ;
  assign y12247 = n20792 ;
  assign y12248 = ~1'b0 ;
  assign y12249 = ~n20794 ;
  assign y12250 = n20796 ;
  assign y12251 = ~1'b0 ;
  assign y12252 = ~n20799 ;
  assign y12253 = ~n20800 ;
  assign y12254 = ~n20804 ;
  assign y12255 = n20805 ;
  assign y12256 = ~n20806 ;
  assign y12257 = ~n20808 ;
  assign y12258 = n11586 ;
  assign y12259 = ~1'b0 ;
  assign y12260 = ~n20809 ;
  assign y12261 = ~n20813 ;
  assign y12262 = n20815 ;
  assign y12263 = ~1'b0 ;
  assign y12264 = ~1'b0 ;
  assign y12265 = ~n12193 ;
  assign y12266 = ~1'b0 ;
  assign y12267 = ~1'b0 ;
  assign y12268 = ~1'b0 ;
  assign y12269 = n20817 ;
  assign y12270 = ~n20818 ;
  assign y12271 = ~1'b0 ;
  assign y12272 = ~1'b0 ;
  assign y12273 = ~n20822 ;
  assign y12274 = ~n20827 ;
  assign y12275 = ~n20829 ;
  assign y12276 = n20830 ;
  assign y12277 = ~n20834 ;
  assign y12278 = n20838 ;
  assign y12279 = n20839 ;
  assign y12280 = ~n20845 ;
  assign y12281 = ~1'b0 ;
  assign y12282 = ~n20848 ;
  assign y12283 = ~1'b0 ;
  assign y12284 = n20850 ;
  assign y12285 = ~1'b0 ;
  assign y12286 = ~1'b0 ;
  assign y12287 = n20851 ;
  assign y12288 = ~1'b0 ;
  assign y12289 = 1'b0 ;
  assign y12290 = ~1'b0 ;
  assign y12291 = ~1'b0 ;
  assign y12292 = ~n20857 ;
  assign y12293 = n20858 ;
  assign y12294 = 1'b0 ;
  assign y12295 = ~n20863 ;
  assign y12296 = ~1'b0 ;
  assign y12297 = ~n20864 ;
  assign y12298 = ~n20866 ;
  assign y12299 = n20869 ;
  assign y12300 = n20870 ;
  assign y12301 = ~n20874 ;
  assign y12302 = ~1'b0 ;
  assign y12303 = ~1'b0 ;
  assign y12304 = n20876 ;
  assign y12305 = ~1'b0 ;
  assign y12306 = ~1'b0 ;
  assign y12307 = ~1'b0 ;
  assign y12308 = 1'b0 ;
  assign y12309 = ~n20877 ;
  assign y12310 = ~1'b0 ;
  assign y12311 = ~1'b0 ;
  assign y12312 = ~n20883 ;
  assign y12313 = n20884 ;
  assign y12314 = ~1'b0 ;
  assign y12315 = n20885 ;
  assign y12316 = ~1'b0 ;
  assign y12317 = ~1'b0 ;
  assign y12318 = ~1'b0 ;
  assign y12319 = n20888 ;
  assign y12320 = ~n20889 ;
  assign y12321 = 1'b0 ;
  assign y12322 = ~1'b0 ;
  assign y12323 = ~1'b0 ;
  assign y12324 = ~1'b0 ;
  assign y12325 = ~n20891 ;
  assign y12326 = ~n20894 ;
  assign y12327 = ~1'b0 ;
  assign y12328 = n20895 ;
  assign y12329 = ~1'b0 ;
  assign y12330 = ~1'b0 ;
  assign y12331 = n20896 ;
  assign y12332 = ~1'b0 ;
  assign y12333 = ~1'b0 ;
  assign y12334 = ~1'b0 ;
  assign y12335 = ~1'b0 ;
  assign y12336 = ~1'b0 ;
  assign y12337 = ~n20898 ;
  assign y12338 = 1'b0 ;
  assign y12339 = n20900 ;
  assign y12340 = ~n20902 ;
  assign y12341 = ~1'b0 ;
  assign y12342 = ~n20907 ;
  assign y12343 = ~1'b0 ;
  assign y12344 = ~1'b0 ;
  assign y12345 = n20908 ;
  assign y12346 = ~1'b0 ;
  assign y12347 = n20911 ;
  assign y12348 = ~n20914 ;
  assign y12349 = n20919 ;
  assign y12350 = n20920 ;
  assign y12351 = ~1'b0 ;
  assign y12352 = ~1'b0 ;
  assign y12353 = 1'b0 ;
  assign y12354 = ~n20922 ;
  assign y12355 = n20924 ;
  assign y12356 = ~1'b0 ;
  assign y12357 = ~1'b0 ;
  assign y12358 = n20927 ;
  assign y12359 = ~n20929 ;
  assign y12360 = ~1'b0 ;
  assign y12361 = ~1'b0 ;
  assign y12362 = ~n20933 ;
  assign y12363 = ~1'b0 ;
  assign y12364 = ~1'b0 ;
  assign y12365 = 1'b0 ;
  assign y12366 = n20934 ;
  assign y12367 = n20937 ;
  assign y12368 = ~n20938 ;
  assign y12369 = ~n20942 ;
  assign y12370 = n20948 ;
  assign y12371 = n20950 ;
  assign y12372 = ~n20951 ;
  assign y12373 = n20952 ;
  assign y12374 = ~1'b0 ;
  assign y12375 = ~1'b0 ;
  assign y12376 = ~n7337 ;
  assign y12377 = n20957 ;
  assign y12378 = ~n18485 ;
  assign y12379 = n20958 ;
  assign y12380 = ~1'b0 ;
  assign y12381 = ~n20959 ;
  assign y12382 = ~1'b0 ;
  assign y12383 = ~1'b0 ;
  assign y12384 = ~1'b0 ;
  assign y12385 = ~1'b0 ;
  assign y12386 = ~n20964 ;
  assign y12387 = ~1'b0 ;
  assign y12388 = ~n20966 ;
  assign y12389 = n20968 ;
  assign y12390 = ~n20969 ;
  assign y12391 = n20971 ;
  assign y12392 = ~1'b0 ;
  assign y12393 = n20882 ;
  assign y12394 = ~1'b0 ;
  assign y12395 = ~n20973 ;
  assign y12396 = ~1'b0 ;
  assign y12397 = ~n20976 ;
  assign y12398 = 1'b0 ;
  assign y12399 = n20977 ;
  assign y12400 = ~1'b0 ;
  assign y12401 = ~n20979 ;
  assign y12402 = ~1'b0 ;
  assign y12403 = ~n20984 ;
  assign y12404 = 1'b0 ;
  assign y12405 = n5946 ;
  assign y12406 = ~n20987 ;
  assign y12407 = ~1'b0 ;
  assign y12408 = ~n20990 ;
  assign y12409 = ~n4367 ;
  assign y12410 = ~1'b0 ;
  assign y12411 = 1'b0 ;
  assign y12412 = ~n20991 ;
  assign y12413 = ~1'b0 ;
  assign y12414 = ~1'b0 ;
  assign y12415 = n20994 ;
  assign y12416 = n20997 ;
  assign y12417 = ~1'b0 ;
  assign y12418 = n20998 ;
  assign y12419 = n20999 ;
  assign y12420 = ~1'b0 ;
  assign y12421 = ~1'b0 ;
  assign y12422 = ~1'b0 ;
  assign y12423 = ~n21005 ;
  assign y12424 = ~n21006 ;
  assign y12425 = n21008 ;
  assign y12426 = ~1'b0 ;
  assign y12427 = ~1'b0 ;
  assign y12428 = ~1'b0 ;
  assign y12429 = n21010 ;
  assign y12430 = n21013 ;
  assign y12431 = ~1'b0 ;
  assign y12432 = ~n21017 ;
  assign y12433 = ~n21018 ;
  assign y12434 = ~n21020 ;
  assign y12435 = ~1'b0 ;
  assign y12436 = ~1'b0 ;
  assign y12437 = n13585 ;
  assign y12438 = ~1'b0 ;
  assign y12439 = n21025 ;
  assign y12440 = n21029 ;
  assign y12441 = ~1'b0 ;
  assign y12442 = ~1'b0 ;
  assign y12443 = n21031 ;
  assign y12444 = ~n21032 ;
  assign y12445 = ~n21033 ;
  assign y12446 = ~1'b0 ;
  assign y12447 = ~1'b0 ;
  assign y12448 = n21034 ;
  assign y12449 = n21036 ;
  assign y12450 = n21041 ;
  assign y12451 = ~1'b0 ;
  assign y12452 = ~n21044 ;
  assign y12453 = n19888 ;
  assign y12454 = ~n18402 ;
  assign y12455 = ~n21045 ;
  assign y12456 = ~1'b0 ;
  assign y12457 = ~1'b0 ;
  assign y12458 = ~n21049 ;
  assign y12459 = n21050 ;
  assign y12460 = ~n21052 ;
  assign y12461 = n2664 ;
  assign y12462 = ~1'b0 ;
  assign y12463 = ~n21054 ;
  assign y12464 = n21055 ;
  assign y12465 = ~1'b0 ;
  assign y12466 = n19000 ;
  assign y12467 = n21056 ;
  assign y12468 = n1969 ;
  assign y12469 = ~1'b0 ;
  assign y12470 = ~1'b0 ;
  assign y12471 = ~n21057 ;
  assign y12472 = ~1'b0 ;
  assign y12473 = n21061 ;
  assign y12474 = ~1'b0 ;
  assign y12475 = ~1'b0 ;
  assign y12476 = 1'b0 ;
  assign y12477 = n21067 ;
  assign y12478 = ~n21071 ;
  assign y12479 = n21075 ;
  assign y12480 = ~1'b0 ;
  assign y12481 = ~1'b0 ;
  assign y12482 = n21076 ;
  assign y12483 = ~1'b0 ;
  assign y12484 = ~1'b0 ;
  assign y12485 = n21077 ;
  assign y12486 = n21080 ;
  assign y12487 = ~n21082 ;
  assign y12488 = ~1'b0 ;
  assign y12489 = ~n6461 ;
  assign y12490 = n21083 ;
  assign y12491 = n21084 ;
  assign y12492 = ~n21086 ;
  assign y12493 = ~1'b0 ;
  assign y12494 = n10767 ;
  assign y12495 = n21087 ;
  assign y12496 = ~1'b0 ;
  assign y12497 = n3379 ;
  assign y12498 = ~1'b0 ;
  assign y12499 = 1'b0 ;
  assign y12500 = n21088 ;
  assign y12501 = ~n21093 ;
  assign y12502 = ~1'b0 ;
  assign y12503 = n21095 ;
  assign y12504 = ~1'b0 ;
  assign y12505 = ~1'b0 ;
  assign y12506 = n21100 ;
  assign y12507 = ~1'b0 ;
  assign y12508 = ~n21104 ;
  assign y12509 = ~n21105 ;
  assign y12510 = ~n21107 ;
  assign y12511 = n2577 ;
  assign y12512 = n21111 ;
  assign y12513 = ~n21115 ;
  assign y12514 = ~n9951 ;
  assign y12515 = n21117 ;
  assign y12516 = ~1'b0 ;
  assign y12517 = ~1'b0 ;
  assign y12518 = ~n21118 ;
  assign y12519 = n21120 ;
  assign y12520 = ~1'b0 ;
  assign y12521 = ~n21121 ;
  assign y12522 = n21122 ;
  assign y12523 = ~n21127 ;
  assign y12524 = n21128 ;
  assign y12525 = ~n21130 ;
  assign y12526 = n4723 ;
  assign y12527 = n21134 ;
  assign y12528 = ~n21136 ;
  assign y12529 = n1139 ;
  assign y12530 = n21137 ;
  assign y12531 = ~1'b0 ;
  assign y12532 = ~n6031 ;
  assign y12533 = n21139 ;
  assign y12534 = ~1'b0 ;
  assign y12535 = ~1'b0 ;
  assign y12536 = n21142 ;
  assign y12537 = ~1'b0 ;
  assign y12538 = ~1'b0 ;
  assign y12539 = n21144 ;
  assign y12540 = ~1'b0 ;
  assign y12541 = n21155 ;
  assign y12542 = ~n21157 ;
  assign y12543 = ~1'b0 ;
  assign y12544 = ~n21158 ;
  assign y12545 = ~1'b0 ;
  assign y12546 = n10697 ;
  assign y12547 = ~n21160 ;
  assign y12548 = ~n21162 ;
  assign y12549 = ~n5305 ;
  assign y12550 = ~1'b0 ;
  assign y12551 = n18738 ;
  assign y12552 = n21164 ;
  assign y12553 = ~1'b0 ;
  assign y12554 = ~n21165 ;
  assign y12555 = ~1'b0 ;
  assign y12556 = ~n21167 ;
  assign y12557 = ~1'b0 ;
  assign y12558 = ~n21168 ;
  assign y12559 = n21171 ;
  assign y12560 = ~1'b0 ;
  assign y12561 = ~n21121 ;
  assign y12562 = ~1'b0 ;
  assign y12563 = n21173 ;
  assign y12564 = ~1'b0 ;
  assign y12565 = ~n21174 ;
  assign y12566 = ~1'b0 ;
  assign y12567 = ~n21175 ;
  assign y12568 = 1'b0 ;
  assign y12569 = ~1'b0 ;
  assign y12570 = n21177 ;
  assign y12571 = ~n21178 ;
  assign y12572 = n21179 ;
  assign y12573 = ~n21181 ;
  assign y12574 = ~1'b0 ;
  assign y12575 = ~n21184 ;
  assign y12576 = n21185 ;
  assign y12577 = ~n5288 ;
  assign y12578 = n21186 ;
  assign y12579 = ~n21187 ;
  assign y12580 = ~n21188 ;
  assign y12581 = ~n21189 ;
  assign y12582 = ~1'b0 ;
  assign y12583 = n21193 ;
  assign y12584 = ~n21194 ;
  assign y12585 = ~1'b0 ;
  assign y12586 = n21196 ;
  assign y12587 = ~1'b0 ;
  assign y12588 = n21197 ;
  assign y12589 = ~n21198 ;
  assign y12590 = n21202 ;
  assign y12591 = 1'b0 ;
  assign y12592 = n21205 ;
  assign y12593 = ~1'b0 ;
  assign y12594 = ~n21207 ;
  assign y12595 = ~n21209 ;
  assign y12596 = ~n21212 ;
  assign y12597 = ~n21214 ;
  assign y12598 = n21216 ;
  assign y12599 = n21218 ;
  assign y12600 = n21220 ;
  assign y12601 = ~1'b0 ;
  assign y12602 = ~n21228 ;
  assign y12603 = n21231 ;
  assign y12604 = ~n16231 ;
  assign y12605 = ~n21233 ;
  assign y12606 = n21235 ;
  assign y12607 = ~1'b0 ;
  assign y12608 = n21237 ;
  assign y12609 = n21240 ;
  assign y12610 = ~1'b0 ;
  assign y12611 = ~1'b0 ;
  assign y12612 = ~1'b0 ;
  assign y12613 = ~n21241 ;
  assign y12614 = n21244 ;
  assign y12615 = ~1'b0 ;
  assign y12616 = ~1'b0 ;
  assign y12617 = n21248 ;
  assign y12618 = ~n21250 ;
  assign y12619 = ~n6109 ;
  assign y12620 = n21253 ;
  assign y12621 = n21256 ;
  assign y12622 = ~n6215 ;
  assign y12623 = ~1'b0 ;
  assign y12624 = ~1'b0 ;
  assign y12625 = ~n21257 ;
  assign y12626 = n21259 ;
  assign y12627 = ~1'b0 ;
  assign y12628 = ~1'b0 ;
  assign y12629 = ~n21260 ;
  assign y12630 = ~n21261 ;
  assign y12631 = n21264 ;
  assign y12632 = ~n21269 ;
  assign y12633 = ~1'b0 ;
  assign y12634 = n21270 ;
  assign y12635 = ~n21271 ;
  assign y12636 = ~x28 ;
  assign y12637 = ~1'b0 ;
  assign y12638 = ~1'b0 ;
  assign y12639 = ~n21272 ;
  assign y12640 = ~1'b0 ;
  assign y12641 = ~1'b0 ;
  assign y12642 = ~1'b0 ;
  assign y12643 = ~1'b0 ;
  assign y12644 = ~n21273 ;
  assign y12645 = ~1'b0 ;
  assign y12646 = ~n21274 ;
  assign y12647 = n21275 ;
  assign y12648 = ~1'b0 ;
  assign y12649 = ~n21280 ;
  assign y12650 = ~1'b0 ;
  assign y12651 = ~1'b0 ;
  assign y12652 = n21281 ;
  assign y12653 = ~n21284 ;
  assign y12654 = ~n21295 ;
  assign y12655 = n21296 ;
  assign y12656 = n21300 ;
  assign y12657 = ~n21303 ;
  assign y12658 = n21305 ;
  assign y12659 = ~1'b0 ;
  assign y12660 = n21307 ;
  assign y12661 = n21309 ;
  assign y12662 = ~1'b0 ;
  assign y12663 = ~1'b0 ;
  assign y12664 = ~1'b0 ;
  assign y12665 = ~n21313 ;
  assign y12666 = ~n20631 ;
  assign y12667 = ~1'b0 ;
  assign y12668 = ~n21314 ;
  assign y12669 = ~n7285 ;
  assign y12670 = ~n21317 ;
  assign y12671 = ~n1710 ;
  assign y12672 = ~1'b0 ;
  assign y12673 = n21320 ;
  assign y12674 = 1'b0 ;
  assign y12675 = n9768 ;
  assign y12676 = ~n21323 ;
  assign y12677 = ~1'b0 ;
  assign y12678 = ~n21331 ;
  assign y12679 = ~n21332 ;
  assign y12680 = ~1'b0 ;
  assign y12681 = ~n21333 ;
  assign y12682 = ~n6401 ;
  assign y12683 = ~n21336 ;
  assign y12684 = ~1'b0 ;
  assign y12685 = 1'b0 ;
  assign y12686 = ~n21340 ;
  assign y12687 = n21343 ;
  assign y12688 = n21344 ;
  assign y12689 = n21346 ;
  assign y12690 = n21348 ;
  assign y12691 = ~n21349 ;
  assign y12692 = ~1'b0 ;
  assign y12693 = n21350 ;
  assign y12694 = ~n21354 ;
  assign y12695 = ~n21358 ;
  assign y12696 = ~n21359 ;
  assign y12697 = ~n21365 ;
  assign y12698 = ~n21370 ;
  assign y12699 = n21371 ;
  assign y12700 = ~n21373 ;
  assign y12701 = ~1'b0 ;
  assign y12702 = n21374 ;
  assign y12703 = ~n21381 ;
  assign y12704 = ~1'b0 ;
  assign y12705 = n21382 ;
  assign y12706 = n21383 ;
  assign y12707 = n6057 ;
  assign y12708 = n4527 ;
  assign y12709 = ~1'b0 ;
  assign y12710 = n2143 ;
  assign y12711 = n21385 ;
  assign y12712 = ~n21393 ;
  assign y12713 = ~n21395 ;
  assign y12714 = ~1'b0 ;
  assign y12715 = n1691 ;
  assign y12716 = ~n21398 ;
  assign y12717 = ~1'b0 ;
  assign y12718 = ~1'b0 ;
  assign y12719 = n21399 ;
  assign y12720 = ~n21401 ;
  assign y12721 = ~n21402 ;
  assign y12722 = ~1'b0 ;
  assign y12723 = ~n21414 ;
  assign y12724 = n21417 ;
  assign y12725 = 1'b0 ;
  assign y12726 = ~n21418 ;
  assign y12727 = ~1'b0 ;
  assign y12728 = ~n21421 ;
  assign y12729 = n21423 ;
  assign y12730 = n21425 ;
  assign y12731 = n21426 ;
  assign y12732 = n21427 ;
  assign y12733 = ~1'b0 ;
  assign y12734 = ~1'b0 ;
  assign y12735 = ~n20841 ;
  assign y12736 = ~n7662 ;
  assign y12737 = ~1'b0 ;
  assign y12738 = ~n21429 ;
  assign y12739 = ~1'b0 ;
  assign y12740 = n21432 ;
  assign y12741 = ~1'b0 ;
  assign y12742 = ~n21434 ;
  assign y12743 = n9061 ;
  assign y12744 = ~n21435 ;
  assign y12745 = ~1'b0 ;
  assign y12746 = ~n21436 ;
  assign y12747 = ~n21438 ;
  assign y12748 = n9978 ;
  assign y12749 = ~1'b0 ;
  assign y12750 = ~1'b0 ;
  assign y12751 = ~n21440 ;
  assign y12752 = ~1'b0 ;
  assign y12753 = 1'b0 ;
  assign y12754 = 1'b0 ;
  assign y12755 = ~n21442 ;
  assign y12756 = ~n21443 ;
  assign y12757 = ~n21445 ;
  assign y12758 = ~n11944 ;
  assign y12759 = n1573 ;
  assign y12760 = n21447 ;
  assign y12761 = ~1'b0 ;
  assign y12762 = 1'b0 ;
  assign y12763 = ~x221 ;
  assign y12764 = n21448 ;
  assign y12765 = n21449 ;
  assign y12766 = ~n21451 ;
  assign y12767 = n21452 ;
  assign y12768 = ~n21457 ;
  assign y12769 = ~1'b0 ;
  assign y12770 = ~1'b0 ;
  assign y12771 = ~n21458 ;
  assign y12772 = ~1'b0 ;
  assign y12773 = ~1'b0 ;
  assign y12774 = ~n21459 ;
  assign y12775 = ~n4118 ;
  assign y12776 = n21460 ;
  assign y12777 = ~1'b0 ;
  assign y12778 = ~n21466 ;
  assign y12779 = ~1'b0 ;
  assign y12780 = n21468 ;
  assign y12781 = n21469 ;
  assign y12782 = n21470 ;
  assign y12783 = n21472 ;
  assign y12784 = ~n21475 ;
  assign y12785 = ~1'b0 ;
  assign y12786 = ~n18459 ;
  assign y12787 = ~n21478 ;
  assign y12788 = n21488 ;
  assign y12789 = ~n21489 ;
  assign y12790 = ~1'b0 ;
  assign y12791 = ~n21490 ;
  assign y12792 = ~n21493 ;
  assign y12793 = ~1'b0 ;
  assign y12794 = ~n21494 ;
  assign y12795 = ~1'b0 ;
  assign y12796 = ~n21496 ;
  assign y12797 = n12329 ;
  assign y12798 = ~1'b0 ;
  assign y12799 = ~1'b0 ;
  assign y12800 = n21497 ;
  assign y12801 = ~1'b0 ;
  assign y12802 = n21499 ;
  assign y12803 = ~n21500 ;
  assign y12804 = 1'b0 ;
  assign y12805 = ~1'b0 ;
  assign y12806 = ~1'b0 ;
  assign y12807 = n13596 ;
  assign y12808 = n21501 ;
  assign y12809 = ~n21502 ;
  assign y12810 = ~1'b0 ;
  assign y12811 = ~1'b0 ;
  assign y12812 = n21503 ;
  assign y12813 = ~1'b0 ;
  assign y12814 = n21506 ;
  assign y12815 = ~n1273 ;
  assign y12816 = ~1'b0 ;
  assign y12817 = ~n21507 ;
  assign y12818 = n1825 ;
  assign y12819 = ~1'b0 ;
  assign y12820 = ~1'b0 ;
  assign y12821 = n21508 ;
  assign y12822 = n21513 ;
  assign y12823 = ~1'b0 ;
  assign y12824 = ~n21516 ;
  assign y12825 = ~1'b0 ;
  assign y12826 = ~n21518 ;
  assign y12827 = ~n21524 ;
  assign y12828 = ~n21525 ;
  assign y12829 = ~1'b0 ;
  assign y12830 = ~1'b0 ;
  assign y12831 = 1'b0 ;
  assign y12832 = ~n21530 ;
  assign y12833 = 1'b0 ;
  assign y12834 = ~n17073 ;
  assign y12835 = ~n21532 ;
  assign y12836 = ~n15521 ;
  assign y12837 = ~1'b0 ;
  assign y12838 = n21533 ;
  assign y12839 = ~1'b0 ;
  assign y12840 = n21534 ;
  assign y12841 = n21539 ;
  assign y12842 = ~1'b0 ;
  assign y12843 = n21541 ;
  assign y12844 = n21543 ;
  assign y12845 = ~n21544 ;
  assign y12846 = ~1'b0 ;
  assign y12847 = n21547 ;
  assign y12848 = n21549 ;
  assign y12849 = ~n21553 ;
  assign y12850 = ~1'b0 ;
  assign y12851 = ~n21555 ;
  assign y12852 = ~1'b0 ;
  assign y12853 = ~n21556 ;
  assign y12854 = n21560 ;
  assign y12855 = n3127 ;
  assign y12856 = ~n21566 ;
  assign y12857 = ~1'b0 ;
  assign y12858 = n21568 ;
  assign y12859 = ~n21570 ;
  assign y12860 = n21574 ;
  assign y12861 = ~1'b0 ;
  assign y12862 = ~n21575 ;
  assign y12863 = n21578 ;
  assign y12864 = ~n21583 ;
  assign y12865 = ~n21591 ;
  assign y12866 = n12801 ;
  assign y12867 = ~1'b0 ;
  assign y12868 = ~1'b0 ;
  assign y12869 = ~n21592 ;
  assign y12870 = ~1'b0 ;
  assign y12871 = n21593 ;
  assign y12872 = ~1'b0 ;
  assign y12873 = ~1'b0 ;
  assign y12874 = n21599 ;
  assign y12875 = ~n21601 ;
  assign y12876 = n21606 ;
  assign y12877 = n21607 ;
  assign y12878 = n21610 ;
  assign y12879 = 1'b0 ;
  assign y12880 = n21612 ;
  assign y12881 = ~1'b0 ;
  assign y12882 = n21614 ;
  assign y12883 = ~n21615 ;
  assign y12884 = n4513 ;
  assign y12885 = n21618 ;
  assign y12886 = ~n21623 ;
  assign y12887 = ~n4868 ;
  assign y12888 = ~n21626 ;
  assign y12889 = n21628 ;
  assign y12890 = ~n21631 ;
  assign y12891 = ~n21632 ;
  assign y12892 = ~n21640 ;
  assign y12893 = ~n15993 ;
  assign y12894 = ~n19771 ;
  assign y12895 = 1'b0 ;
  assign y12896 = ~n21646 ;
  assign y12897 = ~n21648 ;
  assign y12898 = ~1'b0 ;
  assign y12899 = ~1'b0 ;
  assign y12900 = n15401 ;
  assign y12901 = n21652 ;
  assign y12902 = ~1'b0 ;
  assign y12903 = n2210 ;
  assign y12904 = n21654 ;
  assign y12905 = ~1'b0 ;
  assign y12906 = n21656 ;
  assign y12907 = n21658 ;
  assign y12908 = n21662 ;
  assign y12909 = ~1'b0 ;
  assign y12910 = ~1'b0 ;
  assign y12911 = ~n21663 ;
  assign y12912 = ~1'b0 ;
  assign y12913 = ~1'b0 ;
  assign y12914 = ~1'b0 ;
  assign y12915 = 1'b0 ;
  assign y12916 = ~n21665 ;
  assign y12917 = ~n21666 ;
  assign y12918 = ~n21667 ;
  assign y12919 = ~1'b0 ;
  assign y12920 = ~1'b0 ;
  assign y12921 = n21668 ;
  assign y12922 = ~1'b0 ;
  assign y12923 = n11585 ;
  assign y12924 = ~n21670 ;
  assign y12925 = ~n14995 ;
  assign y12926 = ~n21671 ;
  assign y12927 = ~1'b0 ;
  assign y12928 = ~n4075 ;
  assign y12929 = n16008 ;
  assign y12930 = n21673 ;
  assign y12931 = ~n21675 ;
  assign y12932 = ~n21678 ;
  assign y12933 = n1651 ;
  assign y12934 = ~1'b0 ;
  assign y12935 = 1'b0 ;
  assign y12936 = ~1'b0 ;
  assign y12937 = n1402 ;
  assign y12938 = n21680 ;
  assign y12939 = ~1'b0 ;
  assign y12940 = n21681 ;
  assign y12941 = n21682 ;
  assign y12942 = ~1'b0 ;
  assign y12943 = n21690 ;
  assign y12944 = ~n21696 ;
  assign y12945 = ~1'b0 ;
  assign y12946 = n21697 ;
  assign y12947 = ~n9128 ;
  assign y12948 = ~n21700 ;
  assign y12949 = ~n21704 ;
  assign y12950 = ~1'b0 ;
  assign y12951 = n8041 ;
  assign y12952 = ~n21706 ;
  assign y12953 = ~1'b0 ;
  assign y12954 = ~1'b0 ;
  assign y12955 = ~n361 ;
  assign y12956 = ~n21710 ;
  assign y12957 = ~n21716 ;
  assign y12958 = ~1'b0 ;
  assign y12959 = ~1'b0 ;
  assign y12960 = ~1'b0 ;
  assign y12961 = ~n8774 ;
  assign y12962 = ~1'b0 ;
  assign y12963 = ~1'b0 ;
  assign y12964 = ~n21718 ;
  assign y12965 = 1'b0 ;
  assign y12966 = ~1'b0 ;
  assign y12967 = ~n21723 ;
  assign y12968 = ~n21724 ;
  assign y12969 = ~1'b0 ;
  assign y12970 = ~n21725 ;
  assign y12971 = ~1'b0 ;
  assign y12972 = ~1'b0 ;
  assign y12973 = ~1'b0 ;
  assign y12974 = ~n21727 ;
  assign y12975 = n21728 ;
  assign y12976 = ~1'b0 ;
  assign y12977 = ~1'b0 ;
  assign y12978 = n988 ;
  assign y12979 = ~1'b0 ;
  assign y12980 = ~n21729 ;
  assign y12981 = n21730 ;
  assign y12982 = 1'b0 ;
  assign y12983 = n21731 ;
  assign y12984 = ~1'b0 ;
  assign y12985 = ~1'b0 ;
  assign y12986 = ~1'b0 ;
  assign y12987 = ~n21736 ;
  assign y12988 = ~1'b0 ;
  assign y12989 = ~1'b0 ;
  assign y12990 = ~n21738 ;
  assign y12991 = n21739 ;
  assign y12992 = ~1'b0 ;
  assign y12993 = ~1'b0 ;
  assign y12994 = n21740 ;
  assign y12995 = ~1'b0 ;
  assign y12996 = ~1'b0 ;
  assign y12997 = 1'b0 ;
  assign y12998 = ~1'b0 ;
  assign y12999 = n21741 ;
  assign y13000 = ~n21743 ;
  assign y13001 = 1'b0 ;
  assign y13002 = ~1'b0 ;
  assign y13003 = n21744 ;
  assign y13004 = ~n21745 ;
  assign y13005 = ~1'b0 ;
  assign y13006 = ~1'b0 ;
  assign y13007 = n19309 ;
  assign y13008 = n21746 ;
  assign y13009 = ~n11486 ;
  assign y13010 = n21748 ;
  assign y13011 = ~n21750 ;
  assign y13012 = n21751 ;
  assign y13013 = n21753 ;
  assign y13014 = ~n21754 ;
  assign y13015 = ~1'b0 ;
  assign y13016 = ~n21758 ;
  assign y13017 = ~1'b0 ;
  assign y13018 = n21759 ;
  assign y13019 = ~n21761 ;
  assign y13020 = 1'b0 ;
  assign y13021 = n21763 ;
  assign y13022 = n21766 ;
  assign y13023 = ~n21769 ;
  assign y13024 = n21771 ;
  assign y13025 = n21773 ;
  assign y13026 = n3407 ;
  assign y13027 = ~n21774 ;
  assign y13028 = n21775 ;
  assign y13029 = ~1'b0 ;
  assign y13030 = ~n21776 ;
  assign y13031 = ~1'b0 ;
  assign y13032 = ~n21779 ;
  assign y13033 = ~n21780 ;
  assign y13034 = ~n21785 ;
  assign y13035 = ~n21786 ;
  assign y13036 = ~n21788 ;
  assign y13037 = ~1'b0 ;
  assign y13038 = n21790 ;
  assign y13039 = 1'b0 ;
  assign y13040 = n21798 ;
  assign y13041 = n10273 ;
  assign y13042 = 1'b0 ;
  assign y13043 = ~1'b0 ;
  assign y13044 = ~1'b0 ;
  assign y13045 = ~n21802 ;
  assign y13046 = ~n21803 ;
  assign y13047 = n21805 ;
  assign y13048 = ~n9439 ;
  assign y13049 = 1'b0 ;
  assign y13050 = ~1'b0 ;
  assign y13051 = ~1'b0 ;
  assign y13052 = ~n21807 ;
  assign y13053 = n5613 ;
  assign y13054 = ~n21812 ;
  assign y13055 = ~n21816 ;
  assign y13056 = ~1'b0 ;
  assign y13057 = 1'b0 ;
  assign y13058 = n21818 ;
  assign y13059 = ~1'b0 ;
  assign y13060 = ~n21819 ;
  assign y13061 = ~n21820 ;
  assign y13062 = ~n21823 ;
  assign y13063 = ~1'b0 ;
  assign y13064 = n21829 ;
  assign y13065 = ~n21832 ;
  assign y13066 = n21833 ;
  assign y13067 = ~n21837 ;
  assign y13068 = n3581 ;
  assign y13069 = n21839 ;
  assign y13070 = ~1'b0 ;
  assign y13071 = ~1'b0 ;
  assign y13072 = n21843 ;
  assign y13073 = ~n21844 ;
  assign y13074 = ~n21847 ;
  assign y13075 = ~1'b0 ;
  assign y13076 = ~n21849 ;
  assign y13077 = n21854 ;
  assign y13078 = ~n21856 ;
  assign y13079 = ~1'b0 ;
  assign y13080 = n21857 ;
  assign y13081 = ~n21858 ;
  assign y13082 = n21859 ;
  assign y13083 = ~1'b0 ;
  assign y13084 = ~n21862 ;
  assign y13085 = ~1'b0 ;
  assign y13086 = n21863 ;
  assign y13087 = ~n14474 ;
  assign y13088 = n21864 ;
  assign y13089 = ~1'b0 ;
  assign y13090 = ~n21865 ;
  assign y13091 = n21869 ;
  assign y13092 = ~n21871 ;
  assign y13093 = n21873 ;
  assign y13094 = ~1'b0 ;
  assign y13095 = n21874 ;
  assign y13096 = n21876 ;
  assign y13097 = n21877 ;
  assign y13098 = ~1'b0 ;
  assign y13099 = ~1'b0 ;
  assign y13100 = ~1'b0 ;
  assign y13101 = 1'b0 ;
  assign y13102 = ~n21879 ;
  assign y13103 = n12713 ;
  assign y13104 = ~n21881 ;
  assign y13105 = ~n21882 ;
  assign y13106 = 1'b0 ;
  assign y13107 = ~n21885 ;
  assign y13108 = 1'b0 ;
  assign y13109 = ~n21887 ;
  assign y13110 = ~n21889 ;
  assign y13111 = ~1'b0 ;
  assign y13112 = ~n21891 ;
  assign y13113 = ~1'b0 ;
  assign y13114 = ~1'b0 ;
  assign y13115 = ~n21893 ;
  assign y13116 = n21895 ;
  assign y13117 = ~1'b0 ;
  assign y13118 = ~n21899 ;
  assign y13119 = n21901 ;
  assign y13120 = ~n7387 ;
  assign y13121 = n21903 ;
  assign y13122 = ~1'b0 ;
  assign y13123 = ~n21905 ;
  assign y13124 = ~n21907 ;
  assign y13125 = n21908 ;
  assign y13126 = ~1'b0 ;
  assign y13127 = n21910 ;
  assign y13128 = ~1'b0 ;
  assign y13129 = ~1'b0 ;
  assign y13130 = ~n21911 ;
  assign y13131 = ~1'b0 ;
  assign y13132 = ~n21913 ;
  assign y13133 = ~n21915 ;
  assign y13134 = n21917 ;
  assign y13135 = ~1'b0 ;
  assign y13136 = n21918 ;
  assign y13137 = ~1'b0 ;
  assign y13138 = ~n21921 ;
  assign y13139 = ~1'b0 ;
  assign y13140 = n21923 ;
  assign y13141 = n21924 ;
  assign y13142 = n21927 ;
  assign y13143 = n21928 ;
  assign y13144 = ~1'b0 ;
  assign y13145 = ~1'b0 ;
  assign y13146 = n21931 ;
  assign y13147 = n21935 ;
  assign y13148 = ~1'b0 ;
  assign y13149 = ~1'b0 ;
  assign y13150 = n11034 ;
  assign y13151 = ~1'b0 ;
  assign y13152 = ~1'b0 ;
  assign y13153 = ~n21943 ;
  assign y13154 = ~1'b0 ;
  assign y13155 = n21944 ;
  assign y13156 = n21946 ;
  assign y13157 = ~1'b0 ;
  assign y13158 = n4059 ;
  assign y13159 = ~1'b0 ;
  assign y13160 = ~n21948 ;
  assign y13161 = n21954 ;
  assign y13162 = ~n21955 ;
  assign y13163 = ~1'b0 ;
  assign y13164 = ~1'b0 ;
  assign y13165 = n21961 ;
  assign y13166 = 1'b0 ;
  assign y13167 = ~1'b0 ;
  assign y13168 = ~1'b0 ;
  assign y13169 = ~1'b0 ;
  assign y13170 = n14980 ;
  assign y13171 = ~1'b0 ;
  assign y13172 = 1'b0 ;
  assign y13173 = ~1'b0 ;
  assign y13174 = n21962 ;
  assign y13175 = 1'b0 ;
  assign y13176 = ~n21971 ;
  assign y13177 = ~1'b0 ;
  assign y13178 = ~n12427 ;
  assign y13179 = ~n21972 ;
  assign y13180 = ~1'b0 ;
  assign y13181 = ~1'b0 ;
  assign y13182 = 1'b0 ;
  assign y13183 = ~1'b0 ;
  assign y13184 = ~1'b0 ;
  assign y13185 = n18159 ;
  assign y13186 = n21976 ;
  assign y13187 = ~1'b0 ;
  assign y13188 = ~n21978 ;
  assign y13189 = n21980 ;
  assign y13190 = ~1'b0 ;
  assign y13191 = n6781 ;
  assign y13192 = ~1'b0 ;
  assign y13193 = ~1'b0 ;
  assign y13194 = ~n21981 ;
  assign y13195 = ~n10599 ;
  assign y13196 = ~n21983 ;
  assign y13197 = ~n21988 ;
  assign y13198 = ~1'b0 ;
  assign y13199 = n21992 ;
  assign y13200 = ~n22003 ;
  assign y13201 = n22004 ;
  assign y13202 = 1'b0 ;
  assign y13203 = ~1'b0 ;
  assign y13204 = n2561 ;
  assign y13205 = ~n22005 ;
  assign y13206 = ~1'b0 ;
  assign y13207 = ~1'b0 ;
  assign y13208 = ~n22011 ;
  assign y13209 = n22012 ;
  assign y13210 = ~1'b0 ;
  assign y13211 = n22014 ;
  assign y13212 = ~1'b0 ;
  assign y13213 = 1'b0 ;
  assign y13214 = n22018 ;
  assign y13215 = n22020 ;
  assign y13216 = ~n22022 ;
  assign y13217 = ~n22029 ;
  assign y13218 = ~n22030 ;
  assign y13219 = n22031 ;
  assign y13220 = ~n22032 ;
  assign y13221 = n22033 ;
  assign y13222 = n22034 ;
  assign y13223 = ~1'b0 ;
  assign y13224 = n22037 ;
  assign y13225 = n22050 ;
  assign y13226 = ~n22051 ;
  assign y13227 = ~1'b0 ;
  assign y13228 = ~1'b0 ;
  assign y13229 = n22052 ;
  assign y13230 = n22053 ;
  assign y13231 = ~n22059 ;
  assign y13232 = ~n22060 ;
  assign y13233 = n15580 ;
  assign y13234 = ~1'b0 ;
  assign y13235 = n22062 ;
  assign y13236 = ~1'b0 ;
  assign y13237 = ~1'b0 ;
  assign y13238 = ~n22067 ;
  assign y13239 = ~1'b0 ;
  assign y13240 = ~1'b0 ;
  assign y13241 = ~n22070 ;
  assign y13242 = ~1'b0 ;
  assign y13243 = ~n19211 ;
  assign y13244 = n22071 ;
  assign y13245 = ~1'b0 ;
  assign y13246 = ~n22074 ;
  assign y13247 = ~n22079 ;
  assign y13248 = ~1'b0 ;
  assign y13249 = n22081 ;
  assign y13250 = ~1'b0 ;
  assign y13251 = n22083 ;
  assign y13252 = ~n22084 ;
  assign y13253 = ~1'b0 ;
  assign y13254 = n22085 ;
  assign y13255 = ~n1239 ;
  assign y13256 = n22091 ;
  assign y13257 = n17305 ;
  assign y13258 = ~n22094 ;
  assign y13259 = n22098 ;
  assign y13260 = ~n22099 ;
  assign y13261 = ~1'b0 ;
  assign y13262 = n22101 ;
  assign y13263 = n22102 ;
  assign y13264 = ~n22108 ;
  assign y13265 = ~n22110 ;
  assign y13266 = ~1'b0 ;
  assign y13267 = ~1'b0 ;
  assign y13268 = ~1'b0 ;
  assign y13269 = ~n22115 ;
  assign y13270 = n22116 ;
  assign y13271 = n22118 ;
  assign y13272 = ~n22119 ;
  assign y13273 = ~1'b0 ;
  assign y13274 = ~1'b0 ;
  assign y13275 = n22120 ;
  assign y13276 = ~1'b0 ;
  assign y13277 = ~n7883 ;
  assign y13278 = ~1'b0 ;
  assign y13279 = n22122 ;
  assign y13280 = n22125 ;
  assign y13281 = n22127 ;
  assign y13282 = ~1'b0 ;
  assign y13283 = ~n22134 ;
  assign y13284 = n22139 ;
  assign y13285 = ~n22141 ;
  assign y13286 = ~1'b0 ;
  assign y13287 = ~1'b0 ;
  assign y13288 = ~n7558 ;
  assign y13289 = ~1'b0 ;
  assign y13290 = n22143 ;
  assign y13291 = n22144 ;
  assign y13292 = ~1'b0 ;
  assign y13293 = n21358 ;
  assign y13294 = n22145 ;
  assign y13295 = ~1'b0 ;
  assign y13296 = ~1'b0 ;
  assign y13297 = ~1'b0 ;
  assign y13298 = ~n22148 ;
  assign y13299 = ~n22150 ;
  assign y13300 = ~n22154 ;
  assign y13301 = ~1'b0 ;
  assign y13302 = n22155 ;
  assign y13303 = ~1'b0 ;
  assign y13304 = ~1'b0 ;
  assign y13305 = ~n22164 ;
  assign y13306 = n22170 ;
  assign y13307 = n22173 ;
  assign y13308 = ~n22176 ;
  assign y13309 = ~n22181 ;
  assign y13310 = ~n22182 ;
  assign y13311 = ~n22183 ;
  assign y13312 = n22185 ;
  assign y13313 = ~n22189 ;
  assign y13314 = ~n22201 ;
  assign y13315 = ~1'b0 ;
  assign y13316 = n22203 ;
  assign y13317 = ~n22205 ;
  assign y13318 = ~n22208 ;
  assign y13319 = n3069 ;
  assign y13320 = n22210 ;
  assign y13321 = ~n22216 ;
  assign y13322 = ~n22217 ;
  assign y13323 = n22219 ;
  assign y13324 = ~n22220 ;
  assign y13325 = n22221 ;
  assign y13326 = n22224 ;
  assign y13327 = ~1'b0 ;
  assign y13328 = ~n22227 ;
  assign y13329 = ~n22228 ;
  assign y13330 = 1'b0 ;
  assign y13331 = n22230 ;
  assign y13332 = ~1'b0 ;
  assign y13333 = ~1'b0 ;
  assign y13334 = ~1'b0 ;
  assign y13335 = ~n22231 ;
  assign y13336 = ~n22232 ;
  assign y13337 = ~n22234 ;
  assign y13338 = n22235 ;
  assign y13339 = ~n22238 ;
  assign y13340 = ~1'b0 ;
  assign y13341 = n22239 ;
  assign y13342 = ~1'b0 ;
  assign y13343 = ~1'b0 ;
  assign y13344 = ~n22241 ;
  assign y13345 = ~n22243 ;
  assign y13346 = n22248 ;
  assign y13347 = ~n22254 ;
  assign y13348 = ~n22257 ;
  assign y13349 = ~n22258 ;
  assign y13350 = n22260 ;
  assign y13351 = ~n22263 ;
  assign y13352 = ~1'b0 ;
  assign y13353 = ~n937 ;
  assign y13354 = n22265 ;
  assign y13355 = ~n22269 ;
  assign y13356 = ~1'b0 ;
  assign y13357 = ~1'b0 ;
  assign y13358 = ~1'b0 ;
  assign y13359 = ~1'b0 ;
  assign y13360 = ~1'b0 ;
  assign y13361 = n22270 ;
  assign y13362 = ~n22271 ;
  assign y13363 = ~n22274 ;
  assign y13364 = n22277 ;
  assign y13365 = n22280 ;
  assign y13366 = ~1'b0 ;
  assign y13367 = ~n22290 ;
  assign y13368 = ~n22291 ;
  assign y13369 = ~1'b0 ;
  assign y13370 = ~1'b0 ;
  assign y13371 = ~1'b0 ;
  assign y13372 = ~n22293 ;
  assign y13373 = n22304 ;
  assign y13374 = ~n22305 ;
  assign y13375 = ~n22306 ;
  assign y13376 = n22308 ;
  assign y13377 = ~n22315 ;
  assign y13378 = ~1'b0 ;
  assign y13379 = ~1'b0 ;
  assign y13380 = ~1'b0 ;
  assign y13381 = n22316 ;
  assign y13382 = ~n22320 ;
  assign y13383 = ~n22322 ;
  assign y13384 = ~1'b0 ;
  assign y13385 = ~1'b0 ;
  assign y13386 = n22325 ;
  assign y13387 = n22326 ;
  assign y13388 = 1'b0 ;
  assign y13389 = ~n22331 ;
  assign y13390 = ~1'b0 ;
  assign y13391 = ~1'b0 ;
  assign y13392 = ~n22332 ;
  assign y13393 = n22333 ;
  assign y13394 = n22335 ;
  assign y13395 = ~1'b0 ;
  assign y13396 = ~n22338 ;
  assign y13397 = ~1'b0 ;
  assign y13398 = n22340 ;
  assign y13399 = ~n22341 ;
  assign y13400 = ~1'b0 ;
  assign y13401 = n22345 ;
  assign y13402 = ~n22349 ;
  assign y13403 = ~n22356 ;
  assign y13404 = ~n22358 ;
  assign y13405 = 1'b0 ;
  assign y13406 = ~1'b0 ;
  assign y13407 = ~1'b0 ;
  assign y13408 = ~n22360 ;
  assign y13409 = ~1'b0 ;
  assign y13410 = n22363 ;
  assign y13411 = ~1'b0 ;
  assign y13412 = n22365 ;
  assign y13413 = ~1'b0 ;
  assign y13414 = ~1'b0 ;
  assign y13415 = ~1'b0 ;
  assign y13416 = 1'b0 ;
  assign y13417 = ~n22369 ;
  assign y13418 = n22372 ;
  assign y13419 = ~n22373 ;
  assign y13420 = ~n22377 ;
  assign y13421 = ~n22382 ;
  assign y13422 = n22384 ;
  assign y13423 = ~1'b0 ;
  assign y13424 = ~1'b0 ;
  assign y13425 = ~n22389 ;
  assign y13426 = n22390 ;
  assign y13427 = n22391 ;
  assign y13428 = 1'b0 ;
  assign y13429 = ~1'b0 ;
  assign y13430 = ~1'b0 ;
  assign y13431 = ~1'b0 ;
  assign y13432 = ~1'b0 ;
  assign y13433 = ~n10797 ;
  assign y13434 = ~1'b0 ;
  assign y13435 = 1'b0 ;
  assign y13436 = ~n22393 ;
  assign y13437 = ~1'b0 ;
  assign y13438 = ~n2106 ;
  assign y13439 = n22400 ;
  assign y13440 = ~n22406 ;
  assign y13441 = ~1'b0 ;
  assign y13442 = 1'b0 ;
  assign y13443 = ~1'b0 ;
  assign y13444 = ~n22411 ;
  assign y13445 = ~1'b0 ;
  assign y13446 = ~1'b0 ;
  assign y13447 = ~1'b0 ;
  assign y13448 = ~1'b0 ;
  assign y13449 = n22412 ;
  assign y13450 = ~1'b0 ;
  assign y13451 = 1'b0 ;
  assign y13452 = ~1'b0 ;
  assign y13453 = n22414 ;
  assign y13454 = ~n22415 ;
  assign y13455 = ~n22419 ;
  assign y13456 = ~1'b0 ;
  assign y13457 = 1'b0 ;
  assign y13458 = ~1'b0 ;
  assign y13459 = ~1'b0 ;
  assign y13460 = n22421 ;
  assign y13461 = ~n22427 ;
  assign y13462 = ~1'b0 ;
  assign y13463 = n22429 ;
  assign y13464 = ~n22432 ;
  assign y13465 = n7885 ;
  assign y13466 = ~1'b0 ;
  assign y13467 = n3695 ;
  assign y13468 = ~1'b0 ;
  assign y13469 = ~1'b0 ;
  assign y13470 = ~1'b0 ;
  assign y13471 = ~n22437 ;
  assign y13472 = n22439 ;
  assign y13473 = n22440 ;
  assign y13474 = ~n4094 ;
  assign y13475 = ~n22441 ;
  assign y13476 = 1'b0 ;
  assign y13477 = n9589 ;
  assign y13478 = n22446 ;
  assign y13479 = ~1'b0 ;
  assign y13480 = ~n22453 ;
  assign y13481 = ~n22454 ;
  assign y13482 = ~n22456 ;
  assign y13483 = ~n22457 ;
  assign y13484 = n12913 ;
  assign y13485 = ~1'b0 ;
  assign y13486 = ~1'b0 ;
  assign y13487 = n22458 ;
  assign y13488 = ~n22460 ;
  assign y13489 = ~1'b0 ;
  assign y13490 = ~n22461 ;
  assign y13491 = ~1'b0 ;
  assign y13492 = ~n22462 ;
  assign y13493 = n22463 ;
  assign y13494 = ~1'b0 ;
  assign y13495 = ~1'b0 ;
  assign y13496 = ~n22466 ;
  assign y13497 = ~1'b0 ;
  assign y13498 = ~n22468 ;
  assign y13499 = ~n22469 ;
  assign y13500 = n22470 ;
  assign y13501 = ~n22472 ;
  assign y13502 = n3476 ;
  assign y13503 = n22476 ;
  assign y13504 = ~1'b0 ;
  assign y13505 = ~1'b0 ;
  assign y13506 = ~n22479 ;
  assign y13507 = n22484 ;
  assign y13508 = ~1'b0 ;
  assign y13509 = ~1'b0 ;
  assign y13510 = n22487 ;
  assign y13511 = n22491 ;
  assign y13512 = ~n22492 ;
  assign y13513 = n22494 ;
  assign y13514 = ~1'b0 ;
  assign y13515 = n22495 ;
  assign y13516 = ~1'b0 ;
  assign y13517 = ~1'b0 ;
  assign y13518 = n22496 ;
  assign y13519 = ~n22499 ;
  assign y13520 = ~1'b0 ;
  assign y13521 = ~n22502 ;
  assign y13522 = ~n22504 ;
  assign y13523 = ~1'b0 ;
  assign y13524 = ~1'b0 ;
  assign y13525 = ~n22506 ;
  assign y13526 = ~n22507 ;
  assign y13527 = ~1'b0 ;
  assign y13528 = ~n22513 ;
  assign y13529 = ~n22517 ;
  assign y13530 = ~n22518 ;
  assign y13531 = n22519 ;
  assign y13532 = ~n22520 ;
  assign y13533 = ~n15721 ;
  assign y13534 = ~1'b0 ;
  assign y13535 = ~1'b0 ;
  assign y13536 = ~n22523 ;
  assign y13537 = n22524 ;
  assign y13538 = ~1'b0 ;
  assign y13539 = ~n22525 ;
  assign y13540 = ~1'b0 ;
  assign y13541 = n22528 ;
  assign y13542 = ~n22531 ;
  assign y13543 = n22534 ;
  assign y13544 = ~n22537 ;
  assign y13545 = ~1'b0 ;
  assign y13546 = ~n22539 ;
  assign y13547 = ~1'b0 ;
  assign y13548 = n22541 ;
  assign y13549 = ~1'b0 ;
  assign y13550 = ~n7650 ;
  assign y13551 = n22542 ;
  assign y13552 = ~n22546 ;
  assign y13553 = 1'b0 ;
  assign y13554 = n22550 ;
  assign y13555 = ~n22554 ;
  assign y13556 = ~n22555 ;
  assign y13557 = ~1'b0 ;
  assign y13558 = ~1'b0 ;
  assign y13559 = 1'b0 ;
  assign y13560 = ~n22558 ;
  assign y13561 = 1'b0 ;
  assign y13562 = ~n22560 ;
  assign y13563 = ~1'b0 ;
  assign y13564 = ~1'b0 ;
  assign y13565 = ~1'b0 ;
  assign y13566 = n22288 ;
  assign y13567 = n22561 ;
  assign y13568 = n22565 ;
  assign y13569 = ~1'b0 ;
  assign y13570 = n22570 ;
  assign y13571 = n22573 ;
  assign y13572 = n22575 ;
  assign y13573 = ~n22579 ;
  assign y13574 = ~n22583 ;
  assign y13575 = ~1'b0 ;
  assign y13576 = ~1'b0 ;
  assign y13577 = 1'b0 ;
  assign y13578 = n22584 ;
  assign y13579 = ~1'b0 ;
  assign y13580 = n22588 ;
  assign y13581 = ~n22598 ;
  assign y13582 = ~1'b0 ;
  assign y13583 = n11810 ;
  assign y13584 = n22599 ;
  assign y13585 = ~1'b0 ;
  assign y13586 = ~1'b0 ;
  assign y13587 = n22601 ;
  assign y13588 = ~n22605 ;
  assign y13589 = n22607 ;
  assign y13590 = n21395 ;
  assign y13591 = ~n22610 ;
  assign y13592 = ~1'b0 ;
  assign y13593 = ~n22611 ;
  assign y13594 = n22614 ;
  assign y13595 = n22616 ;
  assign y13596 = n22617 ;
  assign y13597 = ~n22618 ;
  assign y13598 = ~1'b0 ;
  assign y13599 = n22623 ;
  assign y13600 = n22624 ;
  assign y13601 = n22625 ;
  assign y13602 = n22628 ;
  assign y13603 = ~n22629 ;
  assign y13604 = n22632 ;
  assign y13605 = ~1'b0 ;
  assign y13606 = ~1'b0 ;
  assign y13607 = ~1'b0 ;
  assign y13608 = ~n22633 ;
  assign y13609 = n22637 ;
  assign y13610 = ~1'b0 ;
  assign y13611 = ~n16208 ;
  assign y13612 = ~n22639 ;
  assign y13613 = ~1'b0 ;
  assign y13614 = n22644 ;
  assign y13615 = ~n7373 ;
  assign y13616 = ~n22645 ;
  assign y13617 = ~1'b0 ;
  assign y13618 = ~1'b0 ;
  assign y13619 = ~n22646 ;
  assign y13620 = n4227 ;
  assign y13621 = ~1'b0 ;
  assign y13622 = ~1'b0 ;
  assign y13623 = ~1'b0 ;
  assign y13624 = ~n22647 ;
  assign y13625 = ~n22650 ;
  assign y13626 = ~1'b0 ;
  assign y13627 = n22652 ;
  assign y13628 = n22654 ;
  assign y13629 = n22655 ;
  assign y13630 = n22659 ;
  assign y13631 = n18387 ;
  assign y13632 = ~1'b0 ;
  assign y13633 = ~n22661 ;
  assign y13634 = ~n22665 ;
  assign y13635 = ~1'b0 ;
  assign y13636 = ~1'b0 ;
  assign y13637 = ~n3187 ;
  assign y13638 = n5891 ;
  assign y13639 = ~n399 ;
  assign y13640 = ~1'b0 ;
  assign y13641 = ~1'b0 ;
  assign y13642 = ~1'b0 ;
  assign y13643 = ~n22674 ;
  assign y13644 = ~1'b0 ;
  assign y13645 = ~n22678 ;
  assign y13646 = n22686 ;
  assign y13647 = n22688 ;
  assign y13648 = n22690 ;
  assign y13649 = n22693 ;
  assign y13650 = ~1'b0 ;
  assign y13651 = ~n22694 ;
  assign y13652 = ~n22697 ;
  assign y13653 = ~1'b0 ;
  assign y13654 = n22700 ;
  assign y13655 = ~1'b0 ;
  assign y13656 = ~n22701 ;
  assign y13657 = 1'b0 ;
  assign y13658 = n22704 ;
  assign y13659 = ~1'b0 ;
  assign y13660 = ~n22705 ;
  assign y13661 = n22706 ;
  assign y13662 = 1'b0 ;
  assign y13663 = n3337 ;
  assign y13664 = n22709 ;
  assign y13665 = ~1'b0 ;
  assign y13666 = n22713 ;
  assign y13667 = ~1'b0 ;
  assign y13668 = n22714 ;
  assign y13669 = ~1'b0 ;
  assign y13670 = n22717 ;
  assign y13671 = ~n22718 ;
  assign y13672 = n22720 ;
  assign y13673 = n22721 ;
  assign y13674 = ~1'b0 ;
  assign y13675 = ~1'b0 ;
  assign y13676 = ~n22723 ;
  assign y13677 = ~n22726 ;
  assign y13678 = ~n22731 ;
  assign y13679 = ~n22735 ;
  assign y13680 = ~1'b0 ;
  assign y13681 = n22736 ;
  assign y13682 = ~1'b0 ;
  assign y13683 = ~1'b0 ;
  assign y13684 = ~1'b0 ;
  assign y13685 = n22738 ;
  assign y13686 = ~n1985 ;
  assign y13687 = ~n22741 ;
  assign y13688 = ~n22743 ;
  assign y13689 = ~1'b0 ;
  assign y13690 = n22744 ;
  assign y13691 = ~1'b0 ;
  assign y13692 = n4217 ;
  assign y13693 = ~1'b0 ;
  assign y13694 = ~n10672 ;
  assign y13695 = n22749 ;
  assign y13696 = ~1'b0 ;
  assign y13697 = ~n22753 ;
  assign y13698 = ~n22758 ;
  assign y13699 = n22759 ;
  assign y13700 = n22762 ;
  assign y13701 = n22769 ;
  assign y13702 = ~n22770 ;
  assign y13703 = ~1'b0 ;
  assign y13704 = ~1'b0 ;
  assign y13705 = ~n22771 ;
  assign y13706 = ~1'b0 ;
  assign y13707 = 1'b0 ;
  assign y13708 = ~n22772 ;
  assign y13709 = n22778 ;
  assign y13710 = n10462 ;
  assign y13711 = n22779 ;
  assign y13712 = n22780 ;
  assign y13713 = ~n22782 ;
  assign y13714 = ~n21449 ;
  assign y13715 = ~n22783 ;
  assign y13716 = ~n22784 ;
  assign y13717 = ~1'b0 ;
  assign y13718 = ~1'b0 ;
  assign y13719 = n1773 ;
  assign y13720 = ~1'b0 ;
  assign y13721 = ~1'b0 ;
  assign y13722 = ~1'b0 ;
  assign y13723 = n22786 ;
  assign y13724 = ~1'b0 ;
  assign y13725 = n22787 ;
  assign y13726 = ~1'b0 ;
  assign y13727 = ~1'b0 ;
  assign y13728 = ~n22793 ;
  assign y13729 = ~1'b0 ;
  assign y13730 = ~n22795 ;
  assign y13731 = ~1'b0 ;
  assign y13732 = n22796 ;
  assign y13733 = ~1'b0 ;
  assign y13734 = ~1'b0 ;
  assign y13735 = n22797 ;
  assign y13736 = ~n22800 ;
  assign y13737 = n22802 ;
  assign y13738 = 1'b0 ;
  assign y13739 = ~n22803 ;
  assign y13740 = n22804 ;
  assign y13741 = 1'b0 ;
  assign y13742 = ~1'b0 ;
  assign y13743 = n22807 ;
  assign y13744 = n22808 ;
  assign y13745 = ~1'b0 ;
  assign y13746 = ~n22809 ;
  assign y13747 = n22811 ;
  assign y13748 = ~1'b0 ;
  assign y13749 = ~1'b0 ;
  assign y13750 = ~n22814 ;
  assign y13751 = ~n22815 ;
  assign y13752 = n22821 ;
  assign y13753 = n22825 ;
  assign y13754 = ~n22827 ;
  assign y13755 = ~1'b0 ;
  assign y13756 = ~1'b0 ;
  assign y13757 = n22833 ;
  assign y13758 = ~n22834 ;
  assign y13759 = ~1'b0 ;
  assign y13760 = ~1'b0 ;
  assign y13761 = ~1'b0 ;
  assign y13762 = ~1'b0 ;
  assign y13763 = ~1'b0 ;
  assign y13764 = n22840 ;
  assign y13765 = n1421 ;
  assign y13766 = n4538 ;
  assign y13767 = ~n22841 ;
  assign y13768 = ~n22844 ;
  assign y13769 = n22845 ;
  assign y13770 = ~n22847 ;
  assign y13771 = ~n22852 ;
  assign y13772 = n14945 ;
  assign y13773 = ~n22867 ;
  assign y13774 = ~1'b0 ;
  assign y13775 = ~1'b0 ;
  assign y13776 = 1'b0 ;
  assign y13777 = n22868 ;
  assign y13778 = n22869 ;
  assign y13779 = ~1'b0 ;
  assign y13780 = n7504 ;
  assign y13781 = ~1'b0 ;
  assign y13782 = ~1'b0 ;
  assign y13783 = n22870 ;
  assign y13784 = ~n22872 ;
  assign y13785 = ~n22877 ;
  assign y13786 = ~1'b0 ;
  assign y13787 = ~1'b0 ;
  assign y13788 = ~1'b0 ;
  assign y13789 = ~1'b0 ;
  assign y13790 = n22880 ;
  assign y13791 = ~1'b0 ;
  assign y13792 = ~n22881 ;
  assign y13793 = 1'b0 ;
  assign y13794 = ~1'b0 ;
  assign y13795 = ~1'b0 ;
  assign y13796 = n22882 ;
  assign y13797 = ~1'b0 ;
  assign y13798 = ~n22886 ;
  assign y13799 = ~n22889 ;
  assign y13800 = ~1'b0 ;
  assign y13801 = ~n22893 ;
  assign y13802 = n22894 ;
  assign y13803 = ~n22897 ;
  assign y13804 = n22900 ;
  assign y13805 = n22901 ;
  assign y13806 = ~1'b0 ;
  assign y13807 = ~n22903 ;
  assign y13808 = ~n22905 ;
  assign y13809 = ~n22906 ;
  assign y13810 = n22907 ;
  assign y13811 = n22912 ;
  assign y13812 = n22915 ;
  assign y13813 = ~n22921 ;
  assign y13814 = n22922 ;
  assign y13815 = 1'b0 ;
  assign y13816 = ~n22923 ;
  assign y13817 = n2187 ;
  assign y13818 = ~n22927 ;
  assign y13819 = n1455 ;
  assign y13820 = n22928 ;
  assign y13821 = ~1'b0 ;
  assign y13822 = 1'b0 ;
  assign y13823 = ~n16157 ;
  assign y13824 = ~n22929 ;
  assign y13825 = ~n12094 ;
  assign y13826 = n1066 ;
  assign y13827 = ~n22930 ;
  assign y13828 = ~1'b0 ;
  assign y13829 = ~n22936 ;
  assign y13830 = n22937 ;
  assign y13831 = n22938 ;
  assign y13832 = ~n22939 ;
  assign y13833 = 1'b0 ;
  assign y13834 = ~1'b0 ;
  assign y13835 = ~n22940 ;
  assign y13836 = n22944 ;
  assign y13837 = ~1'b0 ;
  assign y13838 = n22945 ;
  assign y13839 = ~n22950 ;
  assign y13840 = 1'b0 ;
  assign y13841 = n22952 ;
  assign y13842 = ~1'b0 ;
  assign y13843 = n4848 ;
  assign y13844 = ~1'b0 ;
  assign y13845 = n22954 ;
  assign y13846 = ~n22955 ;
  assign y13847 = n22957 ;
  assign y13848 = ~n22959 ;
  assign y13849 = ~1'b0 ;
  assign y13850 = n22960 ;
  assign y13851 = ~1'b0 ;
  assign y13852 = ~n7673 ;
  assign y13853 = ~1'b0 ;
  assign y13854 = ~n22963 ;
  assign y13855 = ~n22965 ;
  assign y13856 = ~1'b0 ;
  assign y13857 = ~n22967 ;
  assign y13858 = ~n22970 ;
  assign y13859 = n22973 ;
  assign y13860 = ~1'b0 ;
  assign y13861 = n22975 ;
  assign y13862 = ~1'b0 ;
  assign y13863 = n22978 ;
  assign y13864 = n22981 ;
  assign y13865 = n22983 ;
  assign y13866 = ~1'b0 ;
  assign y13867 = ~n22984 ;
  assign y13868 = ~1'b0 ;
  assign y13869 = ~n22994 ;
  assign y13870 = ~n22995 ;
  assign y13871 = ~1'b0 ;
  assign y13872 = n22996 ;
  assign y13873 = ~n22997 ;
  assign y13874 = n23001 ;
  assign y13875 = ~1'b0 ;
  assign y13876 = n23003 ;
  assign y13877 = ~1'b0 ;
  assign y13878 = ~n23005 ;
  assign y13879 = n23010 ;
  assign y13880 = ~n23011 ;
  assign y13881 = ~n23013 ;
  assign y13882 = ~1'b0 ;
  assign y13883 = ~n23014 ;
  assign y13884 = ~n23018 ;
  assign y13885 = ~n23020 ;
  assign y13886 = n23022 ;
  assign y13887 = ~n23023 ;
  assign y13888 = n23024 ;
  assign y13889 = ~1'b0 ;
  assign y13890 = ~1'b0 ;
  assign y13891 = ~1'b0 ;
  assign y13892 = ~1'b0 ;
  assign y13893 = ~n23025 ;
  assign y13894 = ~n23034 ;
  assign y13895 = n23037 ;
  assign y13896 = ~1'b0 ;
  assign y13897 = n23038 ;
  assign y13898 = ~n23041 ;
  assign y13899 = 1'b0 ;
  assign y13900 = n12848 ;
  assign y13901 = ~1'b0 ;
  assign y13902 = n23044 ;
  assign y13903 = ~n23045 ;
  assign y13904 = n23050 ;
  assign y13905 = ~n23053 ;
  assign y13906 = ~1'b0 ;
  assign y13907 = ~1'b0 ;
  assign y13908 = ~n23055 ;
  assign y13909 = n23057 ;
  assign y13910 = ~n23059 ;
  assign y13911 = ~1'b0 ;
  assign y13912 = ~1'b0 ;
  assign y13913 = ~1'b0 ;
  assign y13914 = ~n23060 ;
  assign y13915 = n23062 ;
  assign y13916 = ~n23063 ;
  assign y13917 = ~n23064 ;
  assign y13918 = ~n23067 ;
  assign y13919 = ~n23069 ;
  assign y13920 = ~1'b0 ;
  assign y13921 = ~n23070 ;
  assign y13922 = ~1'b0 ;
  assign y13923 = ~1'b0 ;
  assign y13924 = n23071 ;
  assign y13925 = n9493 ;
  assign y13926 = ~1'b0 ;
  assign y13927 = ~n4352 ;
  assign y13928 = ~n23074 ;
  assign y13929 = ~1'b0 ;
  assign y13930 = n23076 ;
  assign y13931 = ~n23077 ;
  assign y13932 = ~1'b0 ;
  assign y13933 = ~n14000 ;
  assign y13934 = ~1'b0 ;
  assign y13935 = ~1'b0 ;
  assign y13936 = ~1'b0 ;
  assign y13937 = n23078 ;
  assign y13938 = ~n23083 ;
  assign y13939 = n23094 ;
  assign y13940 = ~n23095 ;
  assign y13941 = ~1'b0 ;
  assign y13942 = ~n23097 ;
  assign y13943 = n23098 ;
  assign y13944 = ~1'b0 ;
  assign y13945 = ~n23103 ;
  assign y13946 = n23105 ;
  assign y13947 = ~1'b0 ;
  assign y13948 = ~1'b0 ;
  assign y13949 = n23106 ;
  assign y13950 = ~n23107 ;
  assign y13951 = ~n23121 ;
  assign y13952 = n23122 ;
  assign y13953 = n23124 ;
  assign y13954 = n23129 ;
  assign y13955 = ~1'b0 ;
  assign y13956 = ~n4075 ;
  assign y13957 = ~1'b0 ;
  assign y13958 = ~1'b0 ;
  assign y13959 = ~1'b0 ;
  assign y13960 = n23130 ;
  assign y13961 = ~n14578 ;
  assign y13962 = ~n23133 ;
  assign y13963 = ~1'b0 ;
  assign y13964 = ~n23136 ;
  assign y13965 = n23138 ;
  assign y13966 = ~n23139 ;
  assign y13967 = n23141 ;
  assign y13968 = ~n23143 ;
  assign y13969 = n23146 ;
  assign y13970 = ~1'b0 ;
  assign y13971 = ~1'b0 ;
  assign y13972 = ~1'b0 ;
  assign y13973 = n23148 ;
  assign y13974 = ~n23153 ;
  assign y13975 = 1'b0 ;
  assign y13976 = ~1'b0 ;
  assign y13977 = ~1'b0 ;
  assign y13978 = ~1'b0 ;
  assign y13979 = ~n23154 ;
  assign y13980 = ~1'b0 ;
  assign y13981 = n23155 ;
  assign y13982 = n23161 ;
  assign y13983 = ~n22760 ;
  assign y13984 = ~n23164 ;
  assign y13985 = ~n23165 ;
  assign y13986 = ~1'b0 ;
  assign y13987 = ~1'b0 ;
  assign y13988 = ~n23184 ;
  assign y13989 = ~1'b0 ;
  assign y13990 = n23185 ;
  assign y13991 = ~1'b0 ;
  assign y13992 = n5368 ;
  assign y13993 = ~n23187 ;
  assign y13994 = n22361 ;
  assign y13995 = ~1'b0 ;
  assign y13996 = ~1'b0 ;
  assign y13997 = ~n1815 ;
  assign y13998 = ~1'b0 ;
  assign y13999 = n22288 ;
  assign y14000 = ~1'b0 ;
  assign y14001 = 1'b0 ;
  assign y14002 = ~1'b0 ;
  assign y14003 = ~n23191 ;
  assign y14004 = n23192 ;
  assign y14005 = n23195 ;
  assign y14006 = ~1'b0 ;
  assign y14007 = ~n23200 ;
  assign y14008 = ~n23201 ;
  assign y14009 = ~1'b0 ;
  assign y14010 = n4363 ;
  assign y14011 = n23202 ;
  assign y14012 = ~1'b0 ;
  assign y14013 = n23207 ;
  assign y14014 = n23213 ;
  assign y14015 = ~1'b0 ;
  assign y14016 = n23216 ;
  assign y14017 = ~1'b0 ;
  assign y14018 = n23217 ;
  assign y14019 = n23219 ;
  assign y14020 = ~1'b0 ;
  assign y14021 = ~n23224 ;
  assign y14022 = ~1'b0 ;
  assign y14023 = ~n23225 ;
  assign y14024 = ~n23230 ;
  assign y14025 = n23232 ;
  assign y14026 = n23234 ;
  assign y14027 = n23235 ;
  assign y14028 = 1'b0 ;
  assign y14029 = ~n23236 ;
  assign y14030 = 1'b0 ;
  assign y14031 = n23237 ;
  assign y14032 = ~1'b0 ;
  assign y14033 = ~n12613 ;
  assign y14034 = ~n23241 ;
  assign y14035 = ~n23242 ;
  assign y14036 = ~n23247 ;
  assign y14037 = ~1'b0 ;
  assign y14038 = ~1'b0 ;
  assign y14039 = ~1'b0 ;
  assign y14040 = n23248 ;
  assign y14041 = ~1'b0 ;
  assign y14042 = ~n23249 ;
  assign y14043 = ~1'b0 ;
  assign y14044 = n3140 ;
  assign y14045 = 1'b0 ;
  assign y14046 = ~n23252 ;
  assign y14047 = ~n23256 ;
  assign y14048 = n23258 ;
  assign y14049 = n23262 ;
  assign y14050 = ~n23263 ;
  assign y14051 = ~1'b0 ;
  assign y14052 = n23264 ;
  assign y14053 = ~1'b0 ;
  assign y14054 = n23267 ;
  assign y14055 = 1'b0 ;
  assign y14056 = ~n23269 ;
  assign y14057 = ~n23270 ;
  assign y14058 = ~n23274 ;
  assign y14059 = n23277 ;
  assign y14060 = ~n23284 ;
  assign y14061 = ~n23285 ;
  assign y14062 = n23286 ;
  assign y14063 = n23288 ;
  assign y14064 = ~n23289 ;
  assign y14065 = n23291 ;
  assign y14066 = ~n23293 ;
  assign y14067 = n23295 ;
  assign y14068 = ~n23299 ;
  assign y14069 = 1'b0 ;
  assign y14070 = ~n23303 ;
  assign y14071 = n23305 ;
  assign y14072 = n23308 ;
  assign y14073 = ~1'b0 ;
  assign y14074 = ~n23311 ;
  assign y14075 = 1'b0 ;
  assign y14076 = ~1'b0 ;
  assign y14077 = ~n23312 ;
  assign y14078 = ~1'b0 ;
  assign y14079 = ~n23316 ;
  assign y14080 = n23319 ;
  assign y14081 = ~n23324 ;
  assign y14082 = ~n23327 ;
  assign y14083 = ~n23329 ;
  assign y14084 = n23331 ;
  assign y14085 = ~n11494 ;
  assign y14086 = ~1'b0 ;
  assign y14087 = ~n23333 ;
  assign y14088 = ~1'b0 ;
  assign y14089 = n23334 ;
  assign y14090 = ~n23337 ;
  assign y14091 = ~n7902 ;
  assign y14092 = ~n23339 ;
  assign y14093 = ~n23343 ;
  assign y14094 = n23344 ;
  assign y14095 = ~n23346 ;
  assign y14096 = ~1'b0 ;
  assign y14097 = ~1'b0 ;
  assign y14098 = n7997 ;
  assign y14099 = n23350 ;
  assign y14100 = ~n23352 ;
  assign y14101 = ~1'b0 ;
  assign y14102 = n23353 ;
  assign y14103 = n23357 ;
  assign y14104 = n23358 ;
  assign y14105 = n16818 ;
  assign y14106 = ~1'b0 ;
  assign y14107 = n23362 ;
  assign y14108 = ~n23364 ;
  assign y14109 = 1'b0 ;
  assign y14110 = ~1'b0 ;
  assign y14111 = ~1'b0 ;
  assign y14112 = ~1'b0 ;
  assign y14113 = ~1'b0 ;
  assign y14114 = n23366 ;
  assign y14115 = n23369 ;
  assign y14116 = 1'b0 ;
  assign y14117 = ~n23373 ;
  assign y14118 = x88 ;
  assign y14119 = ~n23374 ;
  assign y14120 = ~1'b0 ;
  assign y14121 = n23376 ;
  assign y14122 = ~n23380 ;
  assign y14123 = ~1'b0 ;
  assign y14124 = 1'b0 ;
  assign y14125 = ~1'b0 ;
  assign y14126 = n23389 ;
  assign y14127 = ~1'b0 ;
  assign y14128 = ~1'b0 ;
  assign y14129 = 1'b0 ;
  assign y14130 = ~1'b0 ;
  assign y14131 = n23393 ;
  assign y14132 = n23398 ;
  assign y14133 = n7358 ;
  assign y14134 = ~1'b0 ;
  assign y14135 = ~n23399 ;
  assign y14136 = n23400 ;
  assign y14137 = ~1'b0 ;
  assign y14138 = n23405 ;
  assign y14139 = ~1'b0 ;
  assign y14140 = ~n23409 ;
  assign y14141 = ~1'b0 ;
  assign y14142 = ~1'b0 ;
  assign y14143 = 1'b0 ;
  assign y14144 = ~n23410 ;
  assign y14145 = ~1'b0 ;
  assign y14146 = ~n14308 ;
  assign y14147 = n23413 ;
  assign y14148 = ~n23414 ;
  assign y14149 = ~1'b0 ;
  assign y14150 = x92 ;
  assign y14151 = ~n23415 ;
  assign y14152 = ~n23422 ;
  assign y14153 = 1'b0 ;
  assign y14154 = ~n6840 ;
  assign y14155 = ~n23427 ;
  assign y14156 = ~n23428 ;
  assign y14157 = n23429 ;
  assign y14158 = n1510 ;
  assign y14159 = n23431 ;
  assign y14160 = ~n6333 ;
  assign y14161 = ~1'b0 ;
  assign y14162 = ~1'b0 ;
  assign y14163 = ~1'b0 ;
  assign y14164 = ~n23432 ;
  assign y14165 = n23433 ;
  assign y14166 = n23437 ;
  assign y14167 = ~n23438 ;
  assign y14168 = ~1'b0 ;
  assign y14169 = n9721 ;
  assign y14170 = ~n23440 ;
  assign y14171 = ~n18869 ;
  assign y14172 = n23442 ;
  assign y14173 = ~1'b0 ;
  assign y14174 = n4549 ;
  assign y14175 = ~1'b0 ;
  assign y14176 = ~n23444 ;
  assign y14177 = ~1'b0 ;
  assign y14178 = n583 ;
  assign y14179 = ~n23453 ;
  assign y14180 = n23459 ;
  assign y14181 = 1'b0 ;
  assign y14182 = ~n20491 ;
  assign y14183 = n23461 ;
  assign y14184 = ~n23462 ;
  assign y14185 = ~1'b0 ;
  assign y14186 = ~n23465 ;
  assign y14187 = ~n23005 ;
  assign y14188 = n23467 ;
  assign y14189 = ~1'b0 ;
  assign y14190 = ~1'b0 ;
  assign y14191 = n23469 ;
  assign y14192 = n9327 ;
  assign y14193 = ~n23471 ;
  assign y14194 = ~1'b0 ;
  assign y14195 = n23472 ;
  assign y14196 = n23475 ;
  assign y14197 = ~1'b0 ;
  assign y14198 = 1'b0 ;
  assign y14199 = n23477 ;
  assign y14200 = ~1'b0 ;
  assign y14201 = n23479 ;
  assign y14202 = ~n23485 ;
  assign y14203 = 1'b0 ;
  assign y14204 = n6152 ;
  assign y14205 = n23486 ;
  assign y14206 = ~1'b0 ;
  assign y14207 = n23487 ;
  assign y14208 = ~1'b0 ;
  assign y14209 = ~n23489 ;
  assign y14210 = ~1'b0 ;
  assign y14211 = n23495 ;
  assign y14212 = ~n23498 ;
  assign y14213 = ~n23499 ;
  assign y14214 = ~1'b0 ;
  assign y14215 = ~1'b0 ;
  assign y14216 = ~1'b0 ;
  assign y14217 = ~n23500 ;
  assign y14218 = ~1'b0 ;
  assign y14219 = n23503 ;
  assign y14220 = ~1'b0 ;
  assign y14221 = ~n14675 ;
  assign y14222 = ~1'b0 ;
  assign y14223 = n2503 ;
  assign y14224 = n23505 ;
  assign y14225 = ~1'b0 ;
  assign y14226 = ~n23513 ;
  assign y14227 = ~1'b0 ;
  assign y14228 = n23514 ;
  assign y14229 = ~n23517 ;
  assign y14230 = ~n23521 ;
  assign y14231 = ~n23528 ;
  assign y14232 = ~n23529 ;
  assign y14233 = ~n23530 ;
  assign y14234 = ~n23533 ;
  assign y14235 = n23534 ;
  assign y14236 = ~1'b0 ;
  assign y14237 = ~n23536 ;
  assign y14238 = ~n23540 ;
  assign y14239 = ~n23541 ;
  assign y14240 = ~1'b0 ;
  assign y14241 = ~1'b0 ;
  assign y14242 = n23542 ;
  assign y14243 = ~n23543 ;
  assign y14244 = n23545 ;
  assign y14245 = ~1'b0 ;
  assign y14246 = n23546 ;
  assign y14247 = ~n23547 ;
  assign y14248 = n23549 ;
  assign y14249 = ~n23553 ;
  assign y14250 = ~1'b0 ;
  assign y14251 = n23556 ;
  assign y14252 = n23557 ;
  assign y14253 = ~1'b0 ;
  assign y14254 = n23558 ;
  assign y14255 = ~n23561 ;
  assign y14256 = n23566 ;
  assign y14257 = ~n11264 ;
  assign y14258 = n23567 ;
  assign y14259 = ~1'b0 ;
  assign y14260 = ~n23571 ;
  assign y14261 = ~n23572 ;
  assign y14262 = n23574 ;
  assign y14263 = ~n23575 ;
  assign y14264 = n23578 ;
  assign y14265 = ~n23582 ;
  assign y14266 = ~n23584 ;
  assign y14267 = ~n8095 ;
  assign y14268 = ~n15569 ;
  assign y14269 = 1'b0 ;
  assign y14270 = ~n23596 ;
  assign y14271 = ~1'b0 ;
  assign y14272 = n9029 ;
  assign y14273 = 1'b0 ;
  assign y14274 = n23597 ;
  assign y14275 = n23602 ;
  assign y14276 = n23603 ;
  assign y14277 = ~1'b0 ;
  assign y14278 = ~1'b0 ;
  assign y14279 = n23604 ;
  assign y14280 = ~n23607 ;
  assign y14281 = n23608 ;
  assign y14282 = ~1'b0 ;
  assign y14283 = n23612 ;
  assign y14284 = n23613 ;
  assign y14285 = n23614 ;
  assign y14286 = ~n23617 ;
  assign y14287 = n23619 ;
  assign y14288 = n23620 ;
  assign y14289 = n23626 ;
  assign y14290 = n23635 ;
  assign y14291 = n23639 ;
  assign y14292 = n23642 ;
  assign y14293 = n4333 ;
  assign y14294 = n23644 ;
  assign y14295 = ~1'b0 ;
  assign y14296 = ~1'b0 ;
  assign y14297 = ~1'b0 ;
  assign y14298 = n23645 ;
  assign y14299 = ~1'b0 ;
  assign y14300 = ~1'b0 ;
  assign y14301 = ~n5146 ;
  assign y14302 = ~n23646 ;
  assign y14303 = n23650 ;
  assign y14304 = n23656 ;
  assign y14305 = n23660 ;
  assign y14306 = ~1'b0 ;
  assign y14307 = ~n23661 ;
  assign y14308 = n23662 ;
  assign y14309 = ~1'b0 ;
  assign y14310 = ~n15953 ;
  assign y14311 = ~n23664 ;
  assign y14312 = n23665 ;
  assign y14313 = n23666 ;
  assign y14314 = n23674 ;
  assign y14315 = ~n23679 ;
  assign y14316 = ~1'b0 ;
  assign y14317 = ~1'b0 ;
  assign y14318 = ~1'b0 ;
  assign y14319 = ~1'b0 ;
  assign y14320 = ~n23682 ;
  assign y14321 = ~n23684 ;
  assign y14322 = n23685 ;
  assign y14323 = ~1'b0 ;
  assign y14324 = ~1'b0 ;
  assign y14325 = ~1'b0 ;
  assign y14326 = ~n23688 ;
  assign y14327 = ~n23689 ;
  assign y14328 = n23690 ;
  assign y14329 = n23691 ;
  assign y14330 = n23693 ;
  assign y14331 = ~1'b0 ;
  assign y14332 = n23698 ;
  assign y14333 = ~n23702 ;
  assign y14334 = ~n23706 ;
  assign y14335 = n23707 ;
  assign y14336 = ~1'b0 ;
  assign y14337 = ~n23711 ;
  assign y14338 = n1541 ;
  assign y14339 = ~1'b0 ;
  assign y14340 = ~n23712 ;
  assign y14341 = ~n23713 ;
  assign y14342 = ~n23714 ;
  assign y14343 = ~1'b0 ;
  assign y14344 = ~n23716 ;
  assign y14345 = ~1'b0 ;
  assign y14346 = n23717 ;
  assign y14347 = n23718 ;
  assign y14348 = n23724 ;
  assign y14349 = ~1'b0 ;
  assign y14350 = ~1'b0 ;
  assign y14351 = 1'b0 ;
  assign y14352 = ~1'b0 ;
  assign y14353 = ~1'b0 ;
  assign y14354 = ~1'b0 ;
  assign y14355 = ~1'b0 ;
  assign y14356 = ~1'b0 ;
  assign y14357 = ~1'b0 ;
  assign y14358 = 1'b0 ;
  assign y14359 = n4824 ;
  assign y14360 = ~n23728 ;
  assign y14361 = n23731 ;
  assign y14362 = ~1'b0 ;
  assign y14363 = n23735 ;
  assign y14364 = n23737 ;
  assign y14365 = ~1'b0 ;
  assign y14366 = n23739 ;
  assign y14367 = ~n23741 ;
  assign y14368 = 1'b0 ;
  assign y14369 = ~1'b0 ;
  assign y14370 = ~1'b0 ;
  assign y14371 = ~1'b0 ;
  assign y14372 = ~1'b0 ;
  assign y14373 = n23743 ;
  assign y14374 = n23747 ;
  assign y14375 = ~1'b0 ;
  assign y14376 = ~n23757 ;
  assign y14377 = ~1'b0 ;
  assign y14378 = n23758 ;
  assign y14379 = ~1'b0 ;
  assign y14380 = ~1'b0 ;
  assign y14381 = ~n23759 ;
  assign y14382 = ~1'b0 ;
  assign y14383 = n23761 ;
  assign y14384 = n23766 ;
  assign y14385 = n23767 ;
  assign y14386 = n23772 ;
  assign y14387 = n23773 ;
  assign y14388 = ~1'b0 ;
  assign y14389 = ~1'b0 ;
  assign y14390 = n23777 ;
  assign y14391 = ~n23779 ;
  assign y14392 = n23784 ;
  assign y14393 = n22263 ;
  assign y14394 = ~n23786 ;
  assign y14395 = ~1'b0 ;
  assign y14396 = ~1'b0 ;
  assign y14397 = ~1'b0 ;
  assign y14398 = ~n23788 ;
  assign y14399 = ~n5462 ;
  assign y14400 = ~n23789 ;
  assign y14401 = ~1'b0 ;
  assign y14402 = n23791 ;
  assign y14403 = ~n23796 ;
  assign y14404 = n6217 ;
  assign y14405 = ~n23799 ;
  assign y14406 = n23801 ;
  assign y14407 = ~n23804 ;
  assign y14408 = n23808 ;
  assign y14409 = n7482 ;
  assign y14410 = ~1'b0 ;
  assign y14411 = ~1'b0 ;
  assign y14412 = ~1'b0 ;
  assign y14413 = ~1'b0 ;
  assign y14414 = ~1'b0 ;
  assign y14415 = ~n23816 ;
  assign y14416 = ~n23820 ;
  assign y14417 = ~1'b0 ;
  assign y14418 = ~1'b0 ;
  assign y14419 = ~1'b0 ;
  assign y14420 = 1'b0 ;
  assign y14421 = ~1'b0 ;
  assign y14422 = ~n23824 ;
  assign y14423 = ~1'b0 ;
  assign y14424 = ~1'b0 ;
  assign y14425 = ~1'b0 ;
  assign y14426 = ~1'b0 ;
  assign y14427 = n23827 ;
  assign y14428 = n23829 ;
  assign y14429 = n23831 ;
  assign y14430 = ~n1890 ;
  assign y14431 = ~n23833 ;
  assign y14432 = n23838 ;
  assign y14433 = ~1'b0 ;
  assign y14434 = n23839 ;
  assign y14435 = n23842 ;
  assign y14436 = n23844 ;
  assign y14437 = ~n23848 ;
  assign y14438 = ~1'b0 ;
  assign y14439 = ~1'b0 ;
  assign y14440 = ~n23853 ;
  assign y14441 = ~n23861 ;
  assign y14442 = ~1'b0 ;
  assign y14443 = 1'b0 ;
  assign y14444 = ~1'b0 ;
  assign y14445 = ~n23862 ;
  assign y14446 = n23864 ;
  assign y14447 = ~1'b0 ;
  assign y14448 = ~n23866 ;
  assign y14449 = ~n23870 ;
  assign y14450 = ~1'b0 ;
  assign y14451 = ~n23874 ;
  assign y14452 = ~n23878 ;
  assign y14453 = ~1'b0 ;
  assign y14454 = ~n2491 ;
  assign y14455 = ~n11683 ;
  assign y14456 = ~n23880 ;
  assign y14457 = n23882 ;
  assign y14458 = n23888 ;
  assign y14459 = ~n23894 ;
  assign y14460 = ~1'b0 ;
  assign y14461 = n23896 ;
  assign y14462 = n23899 ;
  assign y14463 = ~n23902 ;
  assign y14464 = n23906 ;
  assign y14465 = ~1'b0 ;
  assign y14466 = n23908 ;
  assign y14467 = n23912 ;
  assign y14468 = n23920 ;
  assign y14469 = ~n23921 ;
  assign y14470 = n23924 ;
  assign y14471 = ~n23927 ;
  assign y14472 = ~1'b0 ;
  assign y14473 = ~n23930 ;
  assign y14474 = ~n23931 ;
  assign y14475 = ~n23932 ;
  assign y14476 = n19762 ;
  assign y14477 = n14897 ;
  assign y14478 = ~n19814 ;
  assign y14479 = n23935 ;
  assign y14480 = ~n23937 ;
  assign y14481 = n23938 ;
  assign y14482 = n23940 ;
  assign y14483 = n23943 ;
  assign y14484 = n23946 ;
  assign y14485 = n23947 ;
  assign y14486 = ~1'b0 ;
  assign y14487 = n9527 ;
  assign y14488 = ~n23954 ;
  assign y14489 = ~1'b0 ;
  assign y14490 = n23955 ;
  assign y14491 = ~1'b0 ;
  assign y14492 = ~1'b0 ;
  assign y14493 = 1'b0 ;
  assign y14494 = ~n23958 ;
  assign y14495 = 1'b0 ;
  assign y14496 = n23959 ;
  assign y14497 = ~n23963 ;
  assign y14498 = n23967 ;
  assign y14499 = ~n23972 ;
  assign y14500 = ~1'b0 ;
  assign y14501 = ~n23973 ;
  assign y14502 = n23974 ;
  assign y14503 = n23975 ;
  assign y14504 = n4065 ;
  assign y14505 = n23980 ;
  assign y14506 = n7961 ;
  assign y14507 = ~1'b0 ;
  assign y14508 = ~n7671 ;
  assign y14509 = n23982 ;
  assign y14510 = ~1'b0 ;
  assign y14511 = n23986 ;
  assign y14512 = ~1'b0 ;
  assign y14513 = n23987 ;
  assign y14514 = 1'b0 ;
  assign y14515 = ~n23988 ;
  assign y14516 = ~1'b0 ;
  assign y14517 = ~1'b0 ;
  assign y14518 = n23993 ;
  assign y14519 = ~1'b0 ;
  assign y14520 = ~1'b0 ;
  assign y14521 = ~n23999 ;
  assign y14522 = ~1'b0 ;
  assign y14523 = ~n24009 ;
  assign y14524 = ~n24011 ;
  assign y14525 = n24013 ;
  assign y14526 = n24014 ;
  assign y14527 = ~n24020 ;
  assign y14528 = ~n24027 ;
  assign y14529 = ~n24030 ;
  assign y14530 = n6401 ;
  assign y14531 = n6740 ;
  assign y14532 = ~n8631 ;
  assign y14533 = ~n24033 ;
  assign y14534 = ~1'b0 ;
  assign y14535 = ~1'b0 ;
  assign y14536 = n24035 ;
  assign y14537 = ~1'b0 ;
  assign y14538 = ~n24036 ;
  assign y14539 = ~n24039 ;
  assign y14540 = ~n24040 ;
  assign y14541 = ~n20769 ;
  assign y14542 = ~n24043 ;
  assign y14543 = ~1'b0 ;
  assign y14544 = ~1'b0 ;
  assign y14545 = ~n24046 ;
  assign y14546 = ~n24047 ;
  assign y14547 = n24048 ;
  assign y14548 = ~n24051 ;
  assign y14549 = ~1'b0 ;
  assign y14550 = ~1'b0 ;
  assign y14551 = n4675 ;
  assign y14552 = ~1'b0 ;
  assign y14553 = ~n24054 ;
  assign y14554 = ~n24059 ;
  assign y14555 = ~n7609 ;
  assign y14556 = ~n24067 ;
  assign y14557 = ~1'b0 ;
  assign y14558 = ~1'b0 ;
  assign y14559 = n24071 ;
  assign y14560 = n16075 ;
  assign y14561 = ~n24073 ;
  assign y14562 = ~n24075 ;
  assign y14563 = n24080 ;
  assign y14564 = ~1'b0 ;
  assign y14565 = ~1'b0 ;
  assign y14566 = ~1'b0 ;
  assign y14567 = ~1'b0 ;
  assign y14568 = n24084 ;
  assign y14569 = ~1'b0 ;
  assign y14570 = ~n24086 ;
  assign y14571 = n24087 ;
  assign y14572 = ~1'b0 ;
  assign y14573 = ~n24090 ;
  assign y14574 = ~1'b0 ;
  assign y14575 = n24093 ;
  assign y14576 = ~n24097 ;
  assign y14577 = ~n24098 ;
  assign y14578 = ~1'b0 ;
  assign y14579 = ~1'b0 ;
  assign y14580 = n24101 ;
  assign y14581 = n6625 ;
  assign y14582 = ~n24105 ;
  assign y14583 = n24106 ;
  assign y14584 = ~1'b0 ;
  assign y14585 = ~1'b0 ;
  assign y14586 = n24108 ;
  assign y14587 = n24110 ;
  assign y14588 = n24111 ;
  assign y14589 = ~1'b0 ;
  assign y14590 = n24113 ;
  assign y14591 = n24114 ;
  assign y14592 = ~1'b0 ;
  assign y14593 = ~1'b0 ;
  assign y14594 = ~n10116 ;
  assign y14595 = ~1'b0 ;
  assign y14596 = n24115 ;
  assign y14597 = ~1'b0 ;
  assign y14598 = 1'b0 ;
  assign y14599 = n24117 ;
  assign y14600 = ~n24122 ;
  assign y14601 = ~n4738 ;
  assign y14602 = n24126 ;
  assign y14603 = ~n24127 ;
  assign y14604 = 1'b0 ;
  assign y14605 = ~n24129 ;
  assign y14606 = n24130 ;
  assign y14607 = n24136 ;
  assign y14608 = ~n24137 ;
  assign y14609 = ~n24139 ;
  assign y14610 = ~n24140 ;
  assign y14611 = 1'b0 ;
  assign y14612 = n24143 ;
  assign y14613 = ~n24145 ;
  assign y14614 = ~n24147 ;
  assign y14615 = ~n24148 ;
  assign y14616 = ~n24152 ;
  assign y14617 = n24153 ;
  assign y14618 = ~1'b0 ;
  assign y14619 = ~n24167 ;
  assign y14620 = n24171 ;
  assign y14621 = ~n24174 ;
  assign y14622 = 1'b0 ;
  assign y14623 = ~1'b0 ;
  assign y14624 = n24178 ;
  assign y14625 = ~1'b0 ;
  assign y14626 = ~1'b0 ;
  assign y14627 = ~1'b0 ;
  assign y14628 = n24179 ;
  assign y14629 = ~n24181 ;
  assign y14630 = ~n24184 ;
  assign y14631 = n24187 ;
  assign y14632 = ~1'b0 ;
  assign y14633 = ~n24189 ;
  assign y14634 = n24190 ;
  assign y14635 = ~1'b0 ;
  assign y14636 = ~n24191 ;
  assign y14637 = 1'b0 ;
  assign y14638 = n24195 ;
  assign y14639 = ~n24197 ;
  assign y14640 = n24198 ;
  assign y14641 = ~n24204 ;
  assign y14642 = ~n24206 ;
  assign y14643 = n24207 ;
  assign y14644 = ~1'b0 ;
  assign y14645 = ~1'b0 ;
  assign y14646 = n24213 ;
  assign y14647 = ~1'b0 ;
  assign y14648 = ~n24215 ;
  assign y14649 = ~n24216 ;
  assign y14650 = ~1'b0 ;
  assign y14651 = ~n24217 ;
  assign y14652 = n18648 ;
  assign y14653 = ~n24218 ;
  assign y14654 = ~1'b0 ;
  assign y14655 = ~1'b0 ;
  assign y14656 = ~1'b0 ;
  assign y14657 = n24219 ;
  assign y14658 = n24224 ;
  assign y14659 = ~1'b0 ;
  assign y14660 = ~n24226 ;
  assign y14661 = ~n13763 ;
  assign y14662 = n24228 ;
  assign y14663 = ~1'b0 ;
  assign y14664 = ~1'b0 ;
  assign y14665 = n3746 ;
  assign y14666 = n24229 ;
  assign y14667 = ~1'b0 ;
  assign y14668 = ~n20283 ;
  assign y14669 = ~1'b0 ;
  assign y14670 = n24231 ;
  assign y14671 = n24232 ;
  assign y14672 = ~1'b0 ;
  assign y14673 = ~1'b0 ;
  assign y14674 = ~n16892 ;
  assign y14675 = ~1'b0 ;
  assign y14676 = n24235 ;
  assign y14677 = ~1'b0 ;
  assign y14678 = ~1'b0 ;
  assign y14679 = ~n24237 ;
  assign y14680 = 1'b0 ;
  assign y14681 = ~1'b0 ;
  assign y14682 = ~n24238 ;
  assign y14683 = ~1'b0 ;
  assign y14684 = ~n24240 ;
  assign y14685 = 1'b0 ;
  assign y14686 = ~1'b0 ;
  assign y14687 = ~n24241 ;
  assign y14688 = ~n24242 ;
  assign y14689 = n24243 ;
  assign y14690 = n24244 ;
  assign y14691 = ~n24249 ;
  assign y14692 = n19503 ;
  assign y14693 = ~n24253 ;
  assign y14694 = ~1'b0 ;
  assign y14695 = ~1'b0 ;
  assign y14696 = n24258 ;
  assign y14697 = n24260 ;
  assign y14698 = ~1'b0 ;
  assign y14699 = n24262 ;
  assign y14700 = ~1'b0 ;
  assign y14701 = n24265 ;
  assign y14702 = ~n24272 ;
  assign y14703 = ~n24273 ;
  assign y14704 = ~1'b0 ;
  assign y14705 = n24274 ;
  assign y14706 = ~1'b0 ;
  assign y14707 = ~n24275 ;
  assign y14708 = ~n24277 ;
  assign y14709 = ~1'b0 ;
  assign y14710 = n24278 ;
  assign y14711 = ~1'b0 ;
  assign y14712 = ~n24279 ;
  assign y14713 = ~1'b0 ;
  assign y14714 = n24280 ;
  assign y14715 = n24284 ;
  assign y14716 = ~1'b0 ;
  assign y14717 = ~n24285 ;
  assign y14718 = ~n4279 ;
  assign y14719 = ~1'b0 ;
  assign y14720 = ~n24286 ;
  assign y14721 = n24288 ;
  assign y14722 = n5079 ;
  assign y14723 = n24294 ;
  assign y14724 = n24296 ;
  assign y14725 = ~1'b0 ;
  assign y14726 = n24298 ;
  assign y14727 = ~n24300 ;
  assign y14728 = ~n24304 ;
  assign y14729 = ~n24306 ;
  assign y14730 = ~1'b0 ;
  assign y14731 = ~n24310 ;
  assign y14732 = ~1'b0 ;
  assign y14733 = ~n24311 ;
  assign y14734 = ~1'b0 ;
  assign y14735 = n24312 ;
  assign y14736 = ~n24314 ;
  assign y14737 = ~n24316 ;
  assign y14738 = ~n24317 ;
  assign y14739 = ~n24318 ;
  assign y14740 = ~1'b0 ;
  assign y14741 = n24320 ;
  assign y14742 = ~1'b0 ;
  assign y14743 = ~n24325 ;
  assign y14744 = ~1'b0 ;
  assign y14745 = n24329 ;
  assign y14746 = ~n7741 ;
  assign y14747 = ~1'b0 ;
  assign y14748 = ~n24331 ;
  assign y14749 = ~1'b0 ;
  assign y14750 = ~n24333 ;
  assign y14751 = n24337 ;
  assign y14752 = n24338 ;
  assign y14753 = n24340 ;
  assign y14754 = ~1'b0 ;
  assign y14755 = ~1'b0 ;
  assign y14756 = n24341 ;
  assign y14757 = ~1'b0 ;
  assign y14758 = n24342 ;
  assign y14759 = n24343 ;
  assign y14760 = ~n24345 ;
  assign y14761 = ~n24351 ;
  assign y14762 = ~n21387 ;
  assign y14763 = ~n24352 ;
  assign y14764 = ~1'b0 ;
  assign y14765 = ~1'b0 ;
  assign y14766 = ~1'b0 ;
  assign y14767 = n18759 ;
  assign y14768 = n24353 ;
  assign y14769 = ~1'b0 ;
  assign y14770 = ~1'b0 ;
  assign y14771 = ~n24355 ;
  assign y14772 = ~1'b0 ;
  assign y14773 = n24357 ;
  assign y14774 = 1'b0 ;
  assign y14775 = n24359 ;
  assign y14776 = ~1'b0 ;
  assign y14777 = n24363 ;
  assign y14778 = ~1'b0 ;
  assign y14779 = ~1'b0 ;
  assign y14780 = ~1'b0 ;
  assign y14781 = n24367 ;
  assign y14782 = ~1'b0 ;
  assign y14783 = ~1'b0 ;
  assign y14784 = ~n24368 ;
  assign y14785 = ~n24373 ;
  assign y14786 = ~1'b0 ;
  assign y14787 = ~n24376 ;
  assign y14788 = ~1'b0 ;
  assign y14789 = ~n24378 ;
  assign y14790 = 1'b0 ;
  assign y14791 = n24380 ;
  assign y14792 = ~n24382 ;
  assign y14793 = ~n22906 ;
  assign y14794 = ~n9264 ;
  assign y14795 = ~1'b0 ;
  assign y14796 = ~n24384 ;
  assign y14797 = ~n24385 ;
  assign y14798 = ~1'b0 ;
  assign y14799 = n3230 ;
  assign y14800 = ~n24389 ;
  assign y14801 = n24390 ;
  assign y14802 = ~1'b0 ;
  assign y14803 = n24391 ;
  assign y14804 = ~1'b0 ;
  assign y14805 = 1'b0 ;
  assign y14806 = ~1'b0 ;
  assign y14807 = n24394 ;
  assign y14808 = ~n3714 ;
  assign y14809 = ~n24397 ;
  assign y14810 = n24398 ;
  assign y14811 = ~n24402 ;
  assign y14812 = ~n10682 ;
  assign y14813 = ~1'b0 ;
  assign y14814 = n24405 ;
  assign y14815 = ~1'b0 ;
  assign y14816 = ~n24410 ;
  assign y14817 = n24412 ;
  assign y14818 = ~n24417 ;
  assign y14819 = n5615 ;
  assign y14820 = ~1'b0 ;
  assign y14821 = ~1'b0 ;
  assign y14822 = n24418 ;
  assign y14823 = n24421 ;
  assign y14824 = n24422 ;
  assign y14825 = ~n17586 ;
  assign y14826 = ~1'b0 ;
  assign y14827 = ~1'b0 ;
  assign y14828 = n24423 ;
  assign y14829 = n24425 ;
  assign y14830 = ~n24427 ;
  assign y14831 = ~n24430 ;
  assign y14832 = ~n3703 ;
  assign y14833 = n6570 ;
  assign y14834 = ~1'b0 ;
  assign y14835 = ~1'b0 ;
  assign y14836 = ~n24432 ;
  assign y14837 = ~1'b0 ;
  assign y14838 = ~1'b0 ;
  assign y14839 = ~1'b0 ;
  assign y14840 = ~n24435 ;
  assign y14841 = n24439 ;
  assign y14842 = 1'b0 ;
  assign y14843 = 1'b0 ;
  assign y14844 = ~n9248 ;
  assign y14845 = ~1'b0 ;
  assign y14846 = n24441 ;
  assign y14847 = n24442 ;
  assign y14848 = n24448 ;
  assign y14849 = ~n1605 ;
  assign y14850 = n24449 ;
  assign y14851 = ~n24452 ;
  assign y14852 = ~n24453 ;
  assign y14853 = n24458 ;
  assign y14854 = n19697 ;
  assign y14855 = ~1'b0 ;
  assign y14856 = n24462 ;
  assign y14857 = ~n24464 ;
  assign y14858 = ~1'b0 ;
  assign y14859 = ~1'b0 ;
  assign y14860 = ~1'b0 ;
  assign y14861 = ~1'b0 ;
  assign y14862 = ~n24465 ;
  assign y14863 = ~1'b0 ;
  assign y14864 = ~1'b0 ;
  assign y14865 = ~n24468 ;
  assign y14866 = n24469 ;
  assign y14867 = n24474 ;
  assign y14868 = n24476 ;
  assign y14869 = ~n24479 ;
  assign y14870 = n1404 ;
  assign y14871 = n24481 ;
  assign y14872 = n24484 ;
  assign y14873 = n24490 ;
  assign y14874 = n24494 ;
  assign y14875 = ~n4241 ;
  assign y14876 = ~n24498 ;
  assign y14877 = ~1'b0 ;
  assign y14878 = ~1'b0 ;
  assign y14879 = ~n24499 ;
  assign y14880 = ~n18600 ;
  assign y14881 = ~1'b0 ;
  assign y14882 = n24501 ;
  assign y14883 = ~n13370 ;
  assign y14884 = ~1'b0 ;
  assign y14885 = n24502 ;
  assign y14886 = 1'b0 ;
  assign y14887 = ~n24504 ;
  assign y14888 = ~n7867 ;
  assign y14889 = ~n24507 ;
  assign y14890 = ~1'b0 ;
  assign y14891 = n24508 ;
  assign y14892 = ~1'b0 ;
  assign y14893 = ~1'b0 ;
  assign y14894 = n24511 ;
  assign y14895 = ~n24513 ;
  assign y14896 = ~n24516 ;
  assign y14897 = ~n1102 ;
  assign y14898 = ~n24517 ;
  assign y14899 = ~1'b0 ;
  assign y14900 = ~n24518 ;
  assign y14901 = ~n24520 ;
  assign y14902 = ~n8978 ;
  assign y14903 = n24522 ;
  assign y14904 = ~1'b0 ;
  assign y14905 = ~n24523 ;
  assign y14906 = ~n24526 ;
  assign y14907 = 1'b0 ;
  assign y14908 = ~1'b0 ;
  assign y14909 = n24528 ;
  assign y14910 = ~1'b0 ;
  assign y14911 = ~n24529 ;
  assign y14912 = ~n24533 ;
  assign y14913 = n24534 ;
  assign y14914 = ~1'b0 ;
  assign y14915 = n24537 ;
  assign y14916 = ~1'b0 ;
  assign y14917 = ~n24539 ;
  assign y14918 = ~n24540 ;
  assign y14919 = ~1'b0 ;
  assign y14920 = ~1'b0 ;
  assign y14921 = n24541 ;
  assign y14922 = 1'b0 ;
  assign y14923 = ~n24543 ;
  assign y14924 = n10185 ;
  assign y14925 = ~1'b0 ;
  assign y14926 = n959 ;
  assign y14927 = n24545 ;
  assign y14928 = n24546 ;
  assign y14929 = ~1'b0 ;
  assign y14930 = ~n24547 ;
  assign y14931 = ~n24549 ;
  assign y14932 = ~1'b0 ;
  assign y14933 = n24550 ;
  assign y14934 = n24551 ;
  assign y14935 = n24559 ;
  assign y14936 = ~1'b0 ;
  assign y14937 = n24560 ;
  assign y14938 = ~1'b0 ;
  assign y14939 = ~1'b0 ;
  assign y14940 = ~1'b0 ;
  assign y14941 = n24563 ;
  assign y14942 = n24568 ;
  assign y14943 = ~n24569 ;
  assign y14944 = ~n24570 ;
  assign y14945 = ~n24571 ;
  assign y14946 = ~n24574 ;
  assign y14947 = ~n24603 ;
  assign y14948 = ~1'b0 ;
  assign y14949 = n24610 ;
  assign y14950 = ~1'b0 ;
  assign y14951 = ~n24613 ;
  assign y14952 = 1'b0 ;
  assign y14953 = 1'b0 ;
  assign y14954 = n2572 ;
  assign y14955 = ~n24618 ;
  assign y14956 = ~n24624 ;
  assign y14957 = n24626 ;
  assign y14958 = n24627 ;
  assign y14959 = ~1'b0 ;
  assign y14960 = ~n24628 ;
  assign y14961 = ~1'b0 ;
  assign y14962 = n24630 ;
  assign y14963 = ~n24631 ;
  assign y14964 = ~n24633 ;
  assign y14965 = n24635 ;
  assign y14966 = ~1'b0 ;
  assign y14967 = ~1'b0 ;
  assign y14968 = ~n24638 ;
  assign y14969 = ~1'b0 ;
  assign y14970 = n24640 ;
  assign y14971 = n24642 ;
  assign y14972 = ~n24649 ;
  assign y14973 = ~1'b0 ;
  assign y14974 = ~n24652 ;
  assign y14975 = n24660 ;
  assign y14976 = n24664 ;
  assign y14977 = n24667 ;
  assign y14978 = ~1'b0 ;
  assign y14979 = ~n7257 ;
  assign y14980 = ~1'b0 ;
  assign y14981 = ~n24669 ;
  assign y14982 = n19508 ;
  assign y14983 = ~n24670 ;
  assign y14984 = ~1'b0 ;
  assign y14985 = ~n24676 ;
  assign y14986 = ~n24677 ;
  assign y14987 = ~n24681 ;
  assign y14988 = ~1'b0 ;
  assign y14989 = ~1'b0 ;
  assign y14990 = ~1'b0 ;
  assign y14991 = ~n24683 ;
  assign y14992 = ~n2449 ;
  assign y14993 = ~1'b0 ;
  assign y14994 = n23593 ;
  assign y14995 = ~n24688 ;
  assign y14996 = ~n24691 ;
  assign y14997 = 1'b0 ;
  assign y14998 = ~1'b0 ;
  assign y14999 = n24693 ;
  assign y15000 = ~n24700 ;
  assign y15001 = ~n24703 ;
  assign y15002 = ~n24704 ;
  assign y15003 = ~n24706 ;
  assign y15004 = ~n24707 ;
  assign y15005 = ~n24708 ;
  assign y15006 = n24713 ;
  assign y15007 = ~n24714 ;
  assign y15008 = n24716 ;
  assign y15009 = ~n24719 ;
  assign y15010 = ~1'b0 ;
  assign y15011 = n24721 ;
  assign y15012 = n24726 ;
  assign y15013 = ~n24730 ;
  assign y15014 = ~n24732 ;
  assign y15015 = n24733 ;
  assign y15016 = ~n24735 ;
  assign y15017 = n24736 ;
  assign y15018 = ~n24737 ;
  assign y15019 = ~1'b0 ;
  assign y15020 = ~1'b0 ;
  assign y15021 = n24780 ;
  assign y15022 = 1'b0 ;
  assign y15023 = n24783 ;
  assign y15024 = n24787 ;
  assign y15025 = ~n24789 ;
  assign y15026 = n24791 ;
  assign y15027 = n24794 ;
  assign y15028 = ~1'b0 ;
  assign y15029 = ~1'b0 ;
  assign y15030 = n4968 ;
  assign y15031 = n24797 ;
  assign y15032 = n24799 ;
  assign y15033 = n24801 ;
  assign y15034 = ~n24802 ;
  assign y15035 = n24803 ;
  assign y15036 = ~n5534 ;
  assign y15037 = n24805 ;
  assign y15038 = ~n24809 ;
  assign y15039 = ~1'b0 ;
  assign y15040 = n24810 ;
  assign y15041 = ~1'b0 ;
  assign y15042 = ~n6617 ;
  assign y15043 = ~1'b0 ;
  assign y15044 = n4785 ;
  assign y15045 = ~1'b0 ;
  assign y15046 = ~n24811 ;
  assign y15047 = ~1'b0 ;
  assign y15048 = 1'b0 ;
  assign y15049 = ~n24812 ;
  assign y15050 = ~n12635 ;
  assign y15051 = n24814 ;
  assign y15052 = ~1'b0 ;
  assign y15053 = n24817 ;
  assign y15054 = n16635 ;
  assign y15055 = n24818 ;
  assign y15056 = n24824 ;
  assign y15057 = ~1'b0 ;
  assign y15058 = 1'b0 ;
  assign y15059 = n24825 ;
  assign y15060 = ~1'b0 ;
  assign y15061 = ~n24826 ;
  assign y15062 = ~1'b0 ;
  assign y15063 = ~1'b0 ;
  assign y15064 = ~n24828 ;
  assign y15065 = ~1'b0 ;
  assign y15066 = n24831 ;
  assign y15067 = n24832 ;
  assign y15068 = n24836 ;
  assign y15069 = ~1'b0 ;
  assign y15070 = n24839 ;
  assign y15071 = ~n24842 ;
  assign y15072 = ~n24846 ;
  assign y15073 = ~n24850 ;
  assign y15074 = ~1'b0 ;
  assign y15075 = ~1'b0 ;
  assign y15076 = n24852 ;
  assign y15077 = n24853 ;
  assign y15078 = n24854 ;
  assign y15079 = ~n24864 ;
  assign y15080 = n24865 ;
  assign y15081 = n24869 ;
  assign y15082 = ~n24873 ;
  assign y15083 = n24874 ;
  assign y15084 = ~1'b0 ;
  assign y15085 = ~n24875 ;
  assign y15086 = n24878 ;
  assign y15087 = ~1'b0 ;
  assign y15088 = ~1'b0 ;
  assign y15089 = n24880 ;
  assign y15090 = n6944 ;
  assign y15091 = ~1'b0 ;
  assign y15092 = ~1'b0 ;
  assign y15093 = ~1'b0 ;
  assign y15094 = ~1'b0 ;
  assign y15095 = n24882 ;
  assign y15096 = 1'b0 ;
  assign y15097 = n24883 ;
  assign y15098 = n19697 ;
  assign y15099 = ~n24886 ;
  assign y15100 = ~n24887 ;
  assign y15101 = ~1'b0 ;
  assign y15102 = ~n822 ;
  assign y15103 = n24888 ;
  assign y15104 = ~n24892 ;
  assign y15105 = n24901 ;
  assign y15106 = n16371 ;
  assign y15107 = n21955 ;
  assign y15108 = ~n24917 ;
  assign y15109 = ~1'b0 ;
  assign y15110 = ~1'b0 ;
  assign y15111 = n24919 ;
  assign y15112 = ~1'b0 ;
  assign y15113 = ~1'b0 ;
  assign y15114 = ~n24921 ;
  assign y15115 = ~1'b0 ;
  assign y15116 = n24922 ;
  assign y15117 = ~n24923 ;
  assign y15118 = ~n24924 ;
  assign y15119 = ~1'b0 ;
  assign y15120 = ~n17039 ;
  assign y15121 = ~n24928 ;
  assign y15122 = ~1'b0 ;
  assign y15123 = ~1'b0 ;
  assign y15124 = ~n17773 ;
  assign y15125 = ~1'b0 ;
  assign y15126 = ~n24930 ;
  assign y15127 = ~1'b0 ;
  assign y15128 = ~n24931 ;
  assign y15129 = ~1'b0 ;
  assign y15130 = n24932 ;
  assign y15131 = ~n24934 ;
  assign y15132 = ~1'b0 ;
  assign y15133 = n24937 ;
  assign y15134 = ~n24938 ;
  assign y15135 = ~n15161 ;
  assign y15136 = ~1'b0 ;
  assign y15137 = ~n24939 ;
  assign y15138 = 1'b0 ;
  assign y15139 = n24941 ;
  assign y15140 = ~1'b0 ;
  assign y15141 = ~1'b0 ;
  assign y15142 = ~n24942 ;
  assign y15143 = n24945 ;
  assign y15144 = ~1'b0 ;
  assign y15145 = ~n24949 ;
  assign y15146 = ~1'b0 ;
  assign y15147 = n24950 ;
  assign y15148 = ~n24951 ;
  assign y15149 = ~1'b0 ;
  assign y15150 = n24952 ;
  assign y15151 = ~1'b0 ;
  assign y15152 = ~1'b0 ;
  assign y15153 = n21076 ;
  assign y15154 = n24958 ;
  assign y15155 = n24959 ;
  assign y15156 = n24961 ;
  assign y15157 = ~1'b0 ;
  assign y15158 = ~1'b0 ;
  assign y15159 = ~n4536 ;
  assign y15160 = ~1'b0 ;
  assign y15161 = 1'b0 ;
  assign y15162 = n24962 ;
  assign y15163 = ~n24964 ;
  assign y15164 = ~1'b0 ;
  assign y15165 = n24967 ;
  assign y15166 = ~n24969 ;
  assign y15167 = ~n24973 ;
  assign y15168 = ~n24977 ;
  assign y15169 = n24982 ;
  assign y15170 = ~n24987 ;
  assign y15171 = ~n24988 ;
  assign y15172 = ~n11421 ;
  assign y15173 = ~1'b0 ;
  assign y15174 = n22907 ;
  assign y15175 = ~n24989 ;
  assign y15176 = ~1'b0 ;
  assign y15177 = ~1'b0 ;
  assign y15178 = 1'b0 ;
  assign y15179 = n24991 ;
  assign y15180 = 1'b0 ;
  assign y15181 = 1'b0 ;
  assign y15182 = 1'b0 ;
  assign y15183 = ~1'b0 ;
  assign y15184 = n24994 ;
  assign y15185 = ~n24997 ;
  assign y15186 = ~n24998 ;
  assign y15187 = n25004 ;
  assign y15188 = n25006 ;
  assign y15189 = ~1'b0 ;
  assign y15190 = ~n25010 ;
  assign y15191 = n25012 ;
  assign y15192 = ~n25013 ;
  assign y15193 = ~n25016 ;
  assign y15194 = ~n25017 ;
  assign y15195 = ~n12461 ;
  assign y15196 = ~n25018 ;
  assign y15197 = ~n25020 ;
  assign y15198 = ~n25024 ;
  assign y15199 = n25025 ;
  assign y15200 = ~1'b0 ;
  assign y15201 = n25026 ;
  assign y15202 = n25028 ;
  assign y15203 = ~n25029 ;
  assign y15204 = ~n25032 ;
  assign y15205 = ~1'b0 ;
  assign y15206 = ~n16379 ;
  assign y15207 = ~1'b0 ;
  assign y15208 = n25034 ;
  assign y15209 = ~n25039 ;
  assign y15210 = ~n25042 ;
  assign y15211 = ~1'b0 ;
  assign y15212 = ~n6985 ;
  assign y15213 = n25043 ;
  assign y15214 = ~n25045 ;
  assign y15215 = ~1'b0 ;
  assign y15216 = n13072 ;
  assign y15217 = ~n25046 ;
  assign y15218 = n25048 ;
  assign y15219 = ~1'b0 ;
  assign y15220 = ~n25050 ;
  assign y15221 = n25053 ;
  assign y15222 = ~n25056 ;
  assign y15223 = ~n25058 ;
  assign y15224 = n25060 ;
  assign y15225 = ~1'b0 ;
  assign y15226 = ~n25062 ;
  assign y15227 = ~1'b0 ;
  assign y15228 = n25063 ;
  assign y15229 = ~1'b0 ;
  assign y15230 = ~1'b0 ;
  assign y15231 = ~n25064 ;
  assign y15232 = ~1'b0 ;
  assign y15233 = ~n25069 ;
  assign y15234 = 1'b0 ;
  assign y15235 = ~n25070 ;
  assign y15236 = ~n25071 ;
  assign y15237 = n25073 ;
  assign y15238 = ~1'b0 ;
  assign y15239 = n25082 ;
  assign y15240 = 1'b0 ;
  assign y15241 = ~1'b0 ;
  assign y15242 = ~1'b0 ;
  assign y15243 = ~n25083 ;
  assign y15244 = n4336 ;
  assign y15245 = ~1'b0 ;
  assign y15246 = ~n25085 ;
  assign y15247 = ~n25088 ;
  assign y15248 = n4276 ;
  assign y15249 = n25089 ;
  assign y15250 = n25091 ;
  assign y15251 = ~n25097 ;
  assign y15252 = n25099 ;
  assign y15253 = ~1'b0 ;
  assign y15254 = ~n25100 ;
  assign y15255 = ~n25102 ;
  assign y15256 = ~n25103 ;
  assign y15257 = ~1'b0 ;
  assign y15258 = 1'b0 ;
  assign y15259 = ~1'b0 ;
  assign y15260 = ~n25105 ;
  assign y15261 = ~1'b0 ;
  assign y15262 = ~n25106 ;
  assign y15263 = n5523 ;
  assign y15264 = ~1'b0 ;
  assign y15265 = ~1'b0 ;
  assign y15266 = ~1'b0 ;
  assign y15267 = ~1'b0 ;
  assign y15268 = ~1'b0 ;
  assign y15269 = n25107 ;
  assign y15270 = n25116 ;
  assign y15271 = ~1'b0 ;
  assign y15272 = n25117 ;
  assign y15273 = ~n25118 ;
  assign y15274 = n25119 ;
  assign y15275 = n25120 ;
  assign y15276 = 1'b0 ;
  assign y15277 = ~n25123 ;
  assign y15278 = n25124 ;
  assign y15279 = ~1'b0 ;
  assign y15280 = n25126 ;
  assign y15281 = ~n25133 ;
  assign y15282 = ~n25135 ;
  assign y15283 = ~n25136 ;
  assign y15284 = n25138 ;
  assign y15285 = ~1'b0 ;
  assign y15286 = ~1'b0 ;
  assign y15287 = ~1'b0 ;
  assign y15288 = ~1'b0 ;
  assign y15289 = ~n25139 ;
  assign y15290 = ~1'b0 ;
  assign y15291 = ~1'b0 ;
  assign y15292 = ~n25141 ;
  assign y15293 = n25143 ;
  assign y15294 = ~n25144 ;
  assign y15295 = ~n25146 ;
  assign y15296 = ~n24990 ;
  assign y15297 = n25147 ;
  assign y15298 = n19670 ;
  assign y15299 = n14101 ;
  assign y15300 = ~n25149 ;
  assign y15301 = ~1'b0 ;
  assign y15302 = ~1'b0 ;
  assign y15303 = ~n25150 ;
  assign y15304 = ~1'b0 ;
  assign y15305 = ~1'b0 ;
  assign y15306 = ~1'b0 ;
  assign y15307 = ~n25152 ;
  assign y15308 = n25153 ;
  assign y15309 = n25157 ;
  assign y15310 = ~1'b0 ;
  assign y15311 = n25159 ;
  assign y15312 = ~n25160 ;
  assign y15313 = ~1'b0 ;
  assign y15314 = n25161 ;
  assign y15315 = n25163 ;
  assign y15316 = ~n25166 ;
  assign y15317 = ~n25170 ;
  assign y15318 = n25171 ;
  assign y15319 = ~n25172 ;
  assign y15320 = n25174 ;
  assign y15321 = ~n25175 ;
  assign y15322 = n25176 ;
  assign y15323 = ~1'b0 ;
  assign y15324 = 1'b0 ;
  assign y15325 = n19215 ;
  assign y15326 = ~n25179 ;
  assign y15327 = ~1'b0 ;
  assign y15328 = ~1'b0 ;
  assign y15329 = ~n25186 ;
  assign y15330 = ~n25189 ;
  assign y15331 = n8525 ;
  assign y15332 = ~n18467 ;
  assign y15333 = ~n25191 ;
  assign y15334 = ~1'b0 ;
  assign y15335 = ~n25194 ;
  assign y15336 = ~n15698 ;
  assign y15337 = ~n25197 ;
  assign y15338 = ~n9253 ;
  assign y15339 = ~n25200 ;
  assign y15340 = n25202 ;
  assign y15341 = ~1'b0 ;
  assign y15342 = ~1'b0 ;
  assign y15343 = ~1'b0 ;
  assign y15344 = n25203 ;
  assign y15345 = ~1'b0 ;
  assign y15346 = n9639 ;
  assign y15347 = ~1'b0 ;
  assign y15348 = ~1'b0 ;
  assign y15349 = ~1'b0 ;
  assign y15350 = ~n25205 ;
  assign y15351 = n25208 ;
  assign y15352 = ~n17254 ;
  assign y15353 = n25210 ;
  assign y15354 = ~n25211 ;
  assign y15355 = ~n25212 ;
  assign y15356 = ~n24459 ;
  assign y15357 = ~1'b0 ;
  assign y15358 = ~n25216 ;
  assign y15359 = ~n17947 ;
  assign y15360 = ~1'b0 ;
  assign y15361 = ~n25220 ;
  assign y15362 = ~1'b0 ;
  assign y15363 = ~1'b0 ;
  assign y15364 = 1'b0 ;
  assign y15365 = ~n20031 ;
  assign y15366 = ~n25221 ;
  assign y15367 = n25223 ;
  assign y15368 = ~1'b0 ;
  assign y15369 = ~n25225 ;
  assign y15370 = ~n956 ;
  assign y15371 = ~1'b0 ;
  assign y15372 = ~1'b0 ;
  assign y15373 = ~1'b0 ;
  assign y15374 = n10617 ;
  assign y15375 = ~1'b0 ;
  assign y15376 = n25226 ;
  assign y15377 = ~1'b0 ;
  assign y15378 = n25228 ;
  assign y15379 = ~n25230 ;
  assign y15380 = n25233 ;
  assign y15381 = ~1'b0 ;
  assign y15382 = ~n25236 ;
  assign y15383 = ~n25239 ;
  assign y15384 = ~1'b0 ;
  assign y15385 = ~1'b0 ;
  assign y15386 = n25240 ;
  assign y15387 = ~n25241 ;
  assign y15388 = n25246 ;
  assign y15389 = 1'b0 ;
  assign y15390 = ~n25247 ;
  assign y15391 = n25254 ;
  assign y15392 = ~1'b0 ;
  assign y15393 = ~1'b0 ;
  assign y15394 = n25256 ;
  assign y15395 = ~n25259 ;
  assign y15396 = n25261 ;
  assign y15397 = ~n25263 ;
  assign y15398 = ~1'b0 ;
  assign y15399 = ~n25268 ;
  assign y15400 = ~n25276 ;
  assign y15401 = ~1'b0 ;
  assign y15402 = ~1'b0 ;
  assign y15403 = ~n25281 ;
  assign y15404 = n25282 ;
  assign y15405 = n25285 ;
  assign y15406 = ~n25286 ;
  assign y15407 = ~n25291 ;
  assign y15408 = ~1'b0 ;
  assign y15409 = ~n25298 ;
  assign y15410 = ~1'b0 ;
  assign y15411 = ~1'b0 ;
  assign y15412 = n25299 ;
  assign y15413 = ~n25306 ;
  assign y15414 = n25307 ;
  assign y15415 = ~n25308 ;
  assign y15416 = ~n25309 ;
  assign y15417 = ~1'b0 ;
  assign y15418 = n25310 ;
  assign y15419 = n25317 ;
  assign y15420 = n25331 ;
  assign y15421 = ~n25340 ;
  assign y15422 = n25343 ;
  assign y15423 = n25347 ;
  assign y15424 = ~1'b0 ;
  assign y15425 = ~n25349 ;
  assign y15426 = ~1'b0 ;
  assign y15427 = ~n25353 ;
  assign y15428 = ~1'b0 ;
  assign y15429 = ~1'b0 ;
  assign y15430 = n25355 ;
  assign y15431 = ~1'b0 ;
  assign y15432 = ~n25358 ;
  assign y15433 = n16200 ;
  assign y15434 = n25359 ;
  assign y15435 = n25361 ;
  assign y15436 = n25362 ;
  assign y15437 = ~n25369 ;
  assign y15438 = ~n20499 ;
  assign y15439 = ~n25374 ;
  assign y15440 = n25375 ;
  assign y15441 = ~n25376 ;
  assign y15442 = ~n25377 ;
  assign y15443 = ~1'b0 ;
  assign y15444 = ~n6708 ;
  assign y15445 = n25379 ;
  assign y15446 = n25382 ;
  assign y15447 = ~n25383 ;
  assign y15448 = ~n25386 ;
  assign y15449 = ~n25387 ;
  assign y15450 = n25391 ;
  assign y15451 = n25397 ;
  assign y15452 = n25398 ;
  assign y15453 = ~n25400 ;
  assign y15454 = n25403 ;
  assign y15455 = n25406 ;
  assign y15456 = ~1'b0 ;
  assign y15457 = n25410 ;
  assign y15458 = ~n25411 ;
  assign y15459 = ~n25412 ;
  assign y15460 = n25418 ;
  assign y15461 = ~n25419 ;
  assign y15462 = n25421 ;
  assign y15463 = n17294 ;
  assign y15464 = n25422 ;
  assign y15465 = ~1'b0 ;
  assign y15466 = ~1'b0 ;
  assign y15467 = ~n25423 ;
  assign y15468 = n25424 ;
  assign y15469 = ~1'b0 ;
  assign y15470 = n25427 ;
  assign y15471 = ~1'b0 ;
  assign y15472 = n25430 ;
  assign y15473 = ~n25431 ;
  assign y15474 = ~1'b0 ;
  assign y15475 = ~1'b0 ;
  assign y15476 = n25439 ;
  assign y15477 = ~1'b0 ;
  assign y15478 = n25441 ;
  assign y15479 = ~n25442 ;
  assign y15480 = n25447 ;
  assign y15481 = ~1'b0 ;
  assign y15482 = ~n25448 ;
  assign y15483 = n25449 ;
  assign y15484 = ~n25451 ;
  assign y15485 = 1'b0 ;
  assign y15486 = ~1'b0 ;
  assign y15487 = n25453 ;
  assign y15488 = ~1'b0 ;
  assign y15489 = ~n25454 ;
  assign y15490 = ~1'b0 ;
  assign y15491 = n25459 ;
  assign y15492 = n25461 ;
  assign y15493 = ~n715 ;
  assign y15494 = ~n25462 ;
  assign y15495 = ~n25463 ;
  assign y15496 = ~1'b0 ;
  assign y15497 = ~1'b0 ;
  assign y15498 = ~1'b0 ;
  assign y15499 = ~1'b0 ;
  assign y15500 = n25466 ;
  assign y15501 = ~n25469 ;
  assign y15502 = ~1'b0 ;
  assign y15503 = n25470 ;
  assign y15504 = 1'b0 ;
  assign y15505 = ~1'b0 ;
  assign y15506 = ~n25492 ;
  assign y15507 = n25494 ;
  assign y15508 = n25496 ;
  assign y15509 = n25500 ;
  assign y15510 = ~1'b0 ;
  assign y15511 = ~n25504 ;
  assign y15512 = ~n25507 ;
  assign y15513 = ~n25510 ;
  assign y15514 = n25514 ;
  assign y15515 = 1'b0 ;
  assign y15516 = ~n25517 ;
  assign y15517 = ~1'b0 ;
  assign y15518 = ~1'b0 ;
  assign y15519 = ~1'b0 ;
  assign y15520 = ~n25524 ;
  assign y15521 = n25525 ;
  assign y15522 = 1'b0 ;
  assign y15523 = ~n25526 ;
  assign y15524 = ~1'b0 ;
  assign y15525 = ~n25530 ;
  assign y15526 = n25533 ;
  assign y15527 = ~1'b0 ;
  assign y15528 = ~1'b0 ;
  assign y15529 = ~n25535 ;
  assign y15530 = n25536 ;
  assign y15531 = ~n25537 ;
  assign y15532 = ~n25541 ;
  assign y15533 = n25546 ;
  assign y15534 = n25548 ;
  assign y15535 = n25553 ;
  assign y15536 = 1'b0 ;
  assign y15537 = n25554 ;
  assign y15538 = n25555 ;
  assign y15539 = ~1'b0 ;
  assign y15540 = n25558 ;
  assign y15541 = n25560 ;
  assign y15542 = ~1'b0 ;
  assign y15543 = n25561 ;
  assign y15544 = ~n25562 ;
  assign y15545 = n4618 ;
  assign y15546 = n25566 ;
  assign y15547 = ~1'b0 ;
  assign y15548 = ~n14897 ;
  assign y15549 = ~1'b0 ;
  assign y15550 = ~n25567 ;
  assign y15551 = ~n25568 ;
  assign y15552 = n25571 ;
  assign y15553 = 1'b0 ;
  assign y15554 = ~1'b0 ;
  assign y15555 = n25572 ;
  assign y15556 = n25574 ;
  assign y15557 = ~1'b0 ;
  assign y15558 = ~1'b0 ;
  assign y15559 = ~n25575 ;
  assign y15560 = n25581 ;
  assign y15561 = ~1'b0 ;
  assign y15562 = ~1'b0 ;
  assign y15563 = n25582 ;
  assign y15564 = ~n25588 ;
  assign y15565 = ~1'b0 ;
  assign y15566 = ~1'b0 ;
  assign y15567 = ~n25591 ;
  assign y15568 = ~1'b0 ;
  assign y15569 = ~n25595 ;
  assign y15570 = ~n25596 ;
  assign y15571 = ~n25599 ;
  assign y15572 = n25603 ;
  assign y15573 = n25606 ;
  assign y15574 = n25610 ;
  assign y15575 = ~n25612 ;
  assign y15576 = ~n25614 ;
  assign y15577 = 1'b0 ;
  assign y15578 = ~n25615 ;
  assign y15579 = ~1'b0 ;
  assign y15580 = ~n25616 ;
  assign y15581 = n6966 ;
  assign y15582 = n25617 ;
  assign y15583 = n25619 ;
  assign y15584 = ~n25622 ;
  assign y15585 = ~1'b0 ;
  assign y15586 = ~1'b0 ;
  assign y15587 = ~1'b0 ;
  assign y15588 = ~1'b0 ;
  assign y15589 = ~1'b0 ;
  assign y15590 = ~1'b0 ;
  assign y15591 = n25625 ;
  assign y15592 = n25627 ;
  assign y15593 = n25633 ;
  assign y15594 = ~1'b0 ;
  assign y15595 = ~n25634 ;
  assign y15596 = ~n25636 ;
  assign y15597 = ~1'b0 ;
  assign y15598 = ~n25639 ;
  assign y15599 = ~n25642 ;
  assign y15600 = ~1'b0 ;
  assign y15601 = ~n25643 ;
  assign y15602 = n25645 ;
  assign y15603 = ~1'b0 ;
  assign y15604 = ~1'b0 ;
  assign y15605 = ~1'b0 ;
  assign y15606 = n25646 ;
  assign y15607 = n25650 ;
  assign y15608 = n25651 ;
  assign y15609 = n25657 ;
  assign y15610 = ~1'b0 ;
  assign y15611 = n5664 ;
  assign y15612 = ~1'b0 ;
  assign y15613 = ~n25661 ;
  assign y15614 = ~n25663 ;
  assign y15615 = 1'b0 ;
  assign y15616 = 1'b0 ;
  assign y15617 = ~n25669 ;
  assign y15618 = ~1'b0 ;
  assign y15619 = ~n25671 ;
  assign y15620 = ~n25672 ;
  assign y15621 = ~n25675 ;
  assign y15622 = ~n25677 ;
  assign y15623 = ~1'b0 ;
  assign y15624 = ~n25681 ;
  assign y15625 = n25686 ;
  assign y15626 = ~1'b0 ;
  assign y15627 = ~1'b0 ;
  assign y15628 = n25688 ;
  assign y15629 = 1'b0 ;
  assign y15630 = ~1'b0 ;
  assign y15631 = n25690 ;
  assign y15632 = n25691 ;
  assign y15633 = 1'b0 ;
  assign y15634 = ~n25693 ;
  assign y15635 = ~1'b0 ;
  assign y15636 = n21297 ;
  assign y15637 = n19058 ;
  assign y15638 = n25695 ;
  assign y15639 = n25696 ;
  assign y15640 = ~1'b0 ;
  assign y15641 = n25703 ;
  assign y15642 = n11330 ;
  assign y15643 = ~n25705 ;
  assign y15644 = ~1'b0 ;
  assign y15645 = ~1'b0 ;
  assign y15646 = n25706 ;
  assign y15647 = n25712 ;
  assign y15648 = ~n25713 ;
  assign y15649 = n25714 ;
  assign y15650 = ~1'b0 ;
  assign y15651 = n25725 ;
  assign y15652 = n25727 ;
  assign y15653 = n25728 ;
  assign y15654 = ~1'b0 ;
  assign y15655 = ~1'b0 ;
  assign y15656 = ~1'b0 ;
  assign y15657 = ~n25732 ;
  assign y15658 = n25733 ;
  assign y15659 = ~x12 ;
  assign y15660 = ~1'b0 ;
  assign y15661 = ~n25735 ;
  assign y15662 = ~1'b0 ;
  assign y15663 = ~1'b0 ;
  assign y15664 = ~1'b0 ;
  assign y15665 = ~n25736 ;
  assign y15666 = n25741 ;
  assign y15667 = n25744 ;
  assign y15668 = ~1'b0 ;
  assign y15669 = ~n25745 ;
  assign y15670 = ~1'b0 ;
  assign y15671 = ~1'b0 ;
  assign y15672 = ~n25746 ;
  assign y15673 = n25747 ;
  assign y15674 = ~1'b0 ;
  assign y15675 = ~n25749 ;
  assign y15676 = n25750 ;
  assign y15677 = ~1'b0 ;
  assign y15678 = n25751 ;
  assign y15679 = ~1'b0 ;
  assign y15680 = ~1'b0 ;
  assign y15681 = ~n25753 ;
  assign y15682 = n25754 ;
  assign y15683 = n25755 ;
  assign y15684 = ~1'b0 ;
  assign y15685 = n20538 ;
  assign y15686 = ~n25758 ;
  assign y15687 = ~n8058 ;
  assign y15688 = ~1'b0 ;
  assign y15689 = ~n12018 ;
  assign y15690 = 1'b0 ;
  assign y15691 = ~n25761 ;
  assign y15692 = ~1'b0 ;
  assign y15693 = ~1'b0 ;
  assign y15694 = n25763 ;
  assign y15695 = n12694 ;
  assign y15696 = ~1'b0 ;
  assign y15697 = n25765 ;
  assign y15698 = n25769 ;
  assign y15699 = n25771 ;
  assign y15700 = n25495 ;
  assign y15701 = n6640 ;
  assign y15702 = ~n25779 ;
  assign y15703 = ~n25781 ;
  assign y15704 = ~n25787 ;
  assign y15705 = ~n25789 ;
  assign y15706 = n25791 ;
  assign y15707 = ~n25792 ;
  assign y15708 = n6517 ;
  assign y15709 = ~1'b0 ;
  assign y15710 = ~n25794 ;
  assign y15711 = ~n25795 ;
  assign y15712 = n2263 ;
  assign y15713 = ~n25796 ;
  assign y15714 = ~n25800 ;
  assign y15715 = ~1'b0 ;
  assign y15716 = ~n25804 ;
  assign y15717 = ~1'b0 ;
  assign y15718 = ~n25807 ;
  assign y15719 = ~1'b0 ;
  assign y15720 = n12576 ;
  assign y15721 = ~n25809 ;
  assign y15722 = ~1'b0 ;
  assign y15723 = ~n25810 ;
  assign y15724 = ~n25813 ;
  assign y15725 = ~1'b0 ;
  assign y15726 = ~n25815 ;
  assign y15727 = 1'b0 ;
  assign y15728 = ~n5422 ;
  assign y15729 = ~1'b0 ;
  assign y15730 = ~1'b0 ;
  assign y15731 = ~1'b0 ;
  assign y15732 = ~1'b0 ;
  assign y15733 = n25816 ;
  assign y15734 = ~1'b0 ;
  assign y15735 = ~1'b0 ;
  assign y15736 = n20310 ;
  assign y15737 = ~n25819 ;
  assign y15738 = n25823 ;
  assign y15739 = ~1'b0 ;
  assign y15740 = n25824 ;
  assign y15741 = ~n25825 ;
  assign y15742 = n25826 ;
  assign y15743 = ~1'b0 ;
  assign y15744 = ~n25827 ;
  assign y15745 = n25829 ;
  assign y15746 = ~1'b0 ;
  assign y15747 = n25831 ;
  assign y15748 = n14924 ;
  assign y15749 = n25832 ;
  assign y15750 = ~n25833 ;
  assign y15751 = ~n25837 ;
  assign y15752 = 1'b0 ;
  assign y15753 = n25838 ;
  assign y15754 = ~1'b0 ;
  assign y15755 = ~n25839 ;
  assign y15756 = ~1'b0 ;
  assign y15757 = ~n1337 ;
  assign y15758 = n25849 ;
  assign y15759 = n5419 ;
  assign y15760 = n25851 ;
  assign y15761 = ~1'b0 ;
  assign y15762 = ~1'b0 ;
  assign y15763 = 1'b0 ;
  assign y15764 = ~1'b0 ;
  assign y15765 = 1'b0 ;
  assign y15766 = ~1'b0 ;
  assign y15767 = ~1'b0 ;
  assign y15768 = n16285 ;
  assign y15769 = ~1'b0 ;
  assign y15770 = n25863 ;
  assign y15771 = ~1'b0 ;
  assign y15772 = ~1'b0 ;
  assign y15773 = ~n25865 ;
  assign y15774 = ~n25866 ;
  assign y15775 = ~1'b0 ;
  assign y15776 = n25867 ;
  assign y15777 = 1'b0 ;
  assign y15778 = n25873 ;
  assign y15779 = 1'b0 ;
  assign y15780 = ~n25875 ;
  assign y15781 = ~n25876 ;
  assign y15782 = n25877 ;
  assign y15783 = ~1'b0 ;
  assign y15784 = ~1'b0 ;
  assign y15785 = ~1'b0 ;
  assign y15786 = ~1'b0 ;
  assign y15787 = n25879 ;
  assign y15788 = ~n25881 ;
  assign y15789 = ~n20160 ;
  assign y15790 = ~n25883 ;
  assign y15791 = ~1'b0 ;
  assign y15792 = n25890 ;
  assign y15793 = ~n25891 ;
  assign y15794 = n25893 ;
  assign y15795 = ~1'b0 ;
  assign y15796 = 1'b0 ;
  assign y15797 = n25901 ;
  assign y15798 = n25902 ;
  assign y15799 = ~n25905 ;
  assign y15800 = ~1'b0 ;
  assign y15801 = ~1'b0 ;
  assign y15802 = ~n25909 ;
  assign y15803 = ~1'b0 ;
  assign y15804 = ~1'b0 ;
  assign y15805 = ~n14942 ;
  assign y15806 = ~1'b0 ;
  assign y15807 = n25910 ;
  assign y15808 = n25912 ;
  assign y15809 = ~1'b0 ;
  assign y15810 = ~1'b0 ;
  assign y15811 = ~n25914 ;
  assign y15812 = ~n24094 ;
  assign y15813 = ~n25916 ;
  assign y15814 = ~1'b0 ;
  assign y15815 = ~n2157 ;
  assign y15816 = ~n25918 ;
  assign y15817 = ~1'b0 ;
  assign y15818 = ~n1865 ;
  assign y15819 = ~1'b0 ;
  assign y15820 = n25921 ;
  assign y15821 = n25922 ;
  assign y15822 = ~1'b0 ;
  assign y15823 = n25925 ;
  assign y15824 = n25926 ;
  assign y15825 = n11884 ;
  assign y15826 = n19803 ;
  assign y15827 = n25929 ;
  assign y15828 = ~1'b0 ;
  assign y15829 = ~1'b0 ;
  assign y15830 = n25930 ;
  assign y15831 = ~1'b0 ;
  assign y15832 = ~1'b0 ;
  assign y15833 = ~1'b0 ;
  assign y15834 = ~n25935 ;
  assign y15835 = ~1'b0 ;
  assign y15836 = n25936 ;
  assign y15837 = ~1'b0 ;
  assign y15838 = n25938 ;
  assign y15839 = ~n25941 ;
  assign y15840 = ~1'b0 ;
  assign y15841 = ~1'b0 ;
  assign y15842 = 1'b0 ;
  assign y15843 = ~1'b0 ;
  assign y15844 = ~n25946 ;
  assign y15845 = ~n25949 ;
  assign y15846 = ~1'b0 ;
  assign y15847 = ~n25950 ;
  assign y15848 = ~1'b0 ;
  assign y15849 = ~n25951 ;
  assign y15850 = ~1'b0 ;
  assign y15851 = n25953 ;
  assign y15852 = ~n25954 ;
  assign y15853 = ~n25958 ;
  assign y15854 = ~1'b0 ;
  assign y15855 = ~n25962 ;
  assign y15856 = ~n25964 ;
  assign y15857 = ~x226 ;
  assign y15858 = n25965 ;
  assign y15859 = n25967 ;
  assign y15860 = ~1'b0 ;
  assign y15861 = ~1'b0 ;
  assign y15862 = ~1'b0 ;
  assign y15863 = n25968 ;
  assign y15864 = n25969 ;
  assign y15865 = ~1'b0 ;
  assign y15866 = ~1'b0 ;
  assign y15867 = ~1'b0 ;
  assign y15868 = 1'b0 ;
  assign y15869 = n25971 ;
  assign y15870 = ~n25974 ;
  assign y15871 = ~1'b0 ;
  assign y15872 = ~n25979 ;
  assign y15873 = n25982 ;
  assign y15874 = n25984 ;
  assign y15875 = ~n25986 ;
  assign y15876 = ~n25987 ;
  assign y15877 = n25990 ;
  assign y15878 = 1'b0 ;
  assign y15879 = n21117 ;
  assign y15880 = ~n25991 ;
  assign y15881 = ~n25993 ;
  assign y15882 = n25994 ;
  assign y15883 = ~1'b0 ;
  assign y15884 = 1'b0 ;
  assign y15885 = n25995 ;
  assign y15886 = n25997 ;
  assign y15887 = n26000 ;
  assign y15888 = ~n26005 ;
  assign y15889 = ~1'b0 ;
  assign y15890 = n26006 ;
  assign y15891 = n26008 ;
  assign y15892 = ~n26009 ;
  assign y15893 = ~1'b0 ;
  assign y15894 = ~1'b0 ;
  assign y15895 = ~n26013 ;
  assign y15896 = n26018 ;
  assign y15897 = ~n26019 ;
  assign y15898 = n7083 ;
  assign y15899 = ~1'b0 ;
  assign y15900 = ~1'b0 ;
  assign y15901 = n26023 ;
  assign y15902 = n26025 ;
  assign y15903 = ~1'b0 ;
  assign y15904 = ~1'b0 ;
  assign y15905 = n26027 ;
  assign y15906 = ~1'b0 ;
  assign y15907 = ~1'b0 ;
  assign y15908 = ~1'b0 ;
  assign y15909 = 1'b0 ;
  assign y15910 = ~n26028 ;
  assign y15911 = n26029 ;
  assign y15912 = ~n26032 ;
  assign y15913 = n2185 ;
  assign y15914 = ~1'b0 ;
  assign y15915 = ~n22876 ;
  assign y15916 = n3842 ;
  assign y15917 = n26034 ;
  assign y15918 = ~1'b0 ;
  assign y15919 = ~n26043 ;
  assign y15920 = ~n26044 ;
  assign y15921 = ~n26047 ;
  assign y15922 = ~1'b0 ;
  assign y15923 = ~n26054 ;
  assign y15924 = ~1'b0 ;
  assign y15925 = ~n26059 ;
  assign y15926 = n26062 ;
  assign y15927 = ~1'b0 ;
  assign y15928 = ~n26069 ;
  assign y15929 = ~n18717 ;
  assign y15930 = ~1'b0 ;
  assign y15931 = ~1'b0 ;
  assign y15932 = ~n26070 ;
  assign y15933 = ~1'b0 ;
  assign y15934 = ~n4678 ;
  assign y15935 = ~n26074 ;
  assign y15936 = ~1'b0 ;
  assign y15937 = ~n26075 ;
  assign y15938 = n26076 ;
  assign y15939 = ~n26077 ;
  assign y15940 = ~n26080 ;
  assign y15941 = n26088 ;
  assign y15942 = n26089 ;
  assign y15943 = ~n26094 ;
  assign y15944 = ~n26096 ;
  assign y15945 = ~x20 ;
  assign y15946 = ~1'b0 ;
  assign y15947 = n26097 ;
  assign y15948 = ~n26098 ;
  assign y15949 = ~1'b0 ;
  assign y15950 = n26105 ;
  assign y15951 = ~1'b0 ;
  assign y15952 = n26106 ;
  assign y15953 = ~n26107 ;
  assign y15954 = ~n26108 ;
  assign y15955 = ~1'b0 ;
  assign y15956 = ~1'b0 ;
  assign y15957 = n26113 ;
  assign y15958 = n26116 ;
  assign y15959 = ~n1772 ;
  assign y15960 = ~1'b0 ;
  assign y15961 = ~1'b0 ;
  assign y15962 = n26118 ;
  assign y15963 = ~1'b0 ;
  assign y15964 = n26119 ;
  assign y15965 = ~n26120 ;
  assign y15966 = ~n26122 ;
  assign y15967 = ~1'b0 ;
  assign y15968 = n26127 ;
  assign y15969 = ~1'b0 ;
  assign y15970 = ~n26128 ;
  assign y15971 = ~n26135 ;
  assign y15972 = ~1'b0 ;
  assign y15973 = n16018 ;
  assign y15974 = n26136 ;
  assign y15975 = ~n26137 ;
  assign y15976 = n26146 ;
  assign y15977 = n26150 ;
  assign y15978 = ~1'b0 ;
  assign y15979 = ~n26152 ;
  assign y15980 = n26154 ;
  assign y15981 = n26166 ;
  assign y15982 = ~1'b0 ;
  assign y15983 = ~n26170 ;
  assign y15984 = ~n26171 ;
  assign y15985 = 1'b0 ;
  assign y15986 = ~n26176 ;
  assign y15987 = n26177 ;
  assign y15988 = ~1'b0 ;
  assign y15989 = ~1'b0 ;
  assign y15990 = ~1'b0 ;
  assign y15991 = ~n26182 ;
  assign y15992 = ~n26184 ;
  assign y15993 = n26185 ;
  assign y15994 = ~n26189 ;
  assign y15995 = ~n26190 ;
  assign y15996 = n26194 ;
  assign y15997 = n26198 ;
  assign y15998 = 1'b0 ;
  assign y15999 = ~n26199 ;
  assign y16000 = ~n26202 ;
  assign y16001 = ~1'b0 ;
  assign y16002 = n26205 ;
  assign y16003 = n26215 ;
  assign y16004 = n26220 ;
  assign y16005 = ~n24147 ;
  assign y16006 = ~1'b0 ;
  assign y16007 = ~1'b0 ;
  assign y16008 = n26222 ;
  assign y16009 = ~n26223 ;
  assign y16010 = ~n26226 ;
  assign y16011 = ~n26232 ;
  assign y16012 = ~n26237 ;
  assign y16013 = n26240 ;
  assign y16014 = ~n26242 ;
  assign y16015 = n26246 ;
  assign y16016 = n26247 ;
  assign y16017 = ~n26250 ;
  assign y16018 = n26252 ;
  assign y16019 = n26255 ;
  assign y16020 = ~n26257 ;
  assign y16021 = n26260 ;
  assign y16022 = ~1'b0 ;
  assign y16023 = ~1'b0 ;
  assign y16024 = n26266 ;
  assign y16025 = 1'b0 ;
  assign y16026 = ~n26267 ;
  assign y16027 = n26270 ;
  assign y16028 = ~1'b0 ;
  assign y16029 = ~n26271 ;
  assign y16030 = n26272 ;
  assign y16031 = ~1'b0 ;
  assign y16032 = ~1'b0 ;
  assign y16033 = n1952 ;
  assign y16034 = ~n26273 ;
  assign y16035 = ~1'b0 ;
  assign y16036 = ~n26274 ;
  assign y16037 = ~n26275 ;
  assign y16038 = ~1'b0 ;
  assign y16039 = ~n26277 ;
  assign y16040 = ~n26278 ;
  assign y16041 = ~n26281 ;
  assign y16042 = ~n26283 ;
  assign y16043 = n26285 ;
  assign y16044 = n26287 ;
  assign y16045 = ~n26289 ;
  assign y16046 = n26290 ;
  assign y16047 = ~1'b0 ;
  assign y16048 = n26294 ;
  assign y16049 = n18077 ;
  assign y16050 = ~n26296 ;
  assign y16051 = ~n6328 ;
  assign y16052 = 1'b0 ;
  assign y16053 = ~1'b0 ;
  assign y16054 = ~1'b0 ;
  assign y16055 = ~1'b0 ;
  assign y16056 = n26298 ;
  assign y16057 = ~n26300 ;
  assign y16058 = ~n26302 ;
  assign y16059 = n26305 ;
  assign y16060 = ~1'b0 ;
  assign y16061 = ~n26307 ;
  assign y16062 = n26309 ;
  assign y16063 = n26310 ;
  assign y16064 = ~n26314 ;
  assign y16065 = ~n26315 ;
  assign y16066 = n26318 ;
  assign y16067 = n26320 ;
  assign y16068 = ~1'b0 ;
  assign y16069 = ~n26322 ;
  assign y16070 = ~1'b0 ;
  assign y16071 = ~n26323 ;
  assign y16072 = ~1'b0 ;
  assign y16073 = n26324 ;
  assign y16074 = ~1'b0 ;
  assign y16075 = n15654 ;
  assign y16076 = n26329 ;
  assign y16077 = ~1'b0 ;
  assign y16078 = n26330 ;
  assign y16079 = ~n26333 ;
  assign y16080 = ~1'b0 ;
  assign y16081 = ~1'b0 ;
  assign y16082 = ~1'b0 ;
  assign y16083 = ~1'b0 ;
  assign y16084 = ~1'b0 ;
  assign y16085 = n26334 ;
  assign y16086 = ~1'b0 ;
  assign y16087 = ~1'b0 ;
  assign y16088 = ~1'b0 ;
  assign y16089 = ~1'b0 ;
  assign y16090 = ~n26335 ;
  assign y16091 = ~n18341 ;
  assign y16092 = ~1'b0 ;
  assign y16093 = ~1'b0 ;
  assign y16094 = ~n26336 ;
  assign y16095 = n26338 ;
  assign y16096 = ~1'b0 ;
  assign y16097 = n26339 ;
  assign y16098 = 1'b0 ;
  assign y16099 = ~1'b0 ;
  assign y16100 = ~n26341 ;
  assign y16101 = n26342 ;
  assign y16102 = ~n26345 ;
  assign y16103 = n8824 ;
  assign y16104 = n26347 ;
  assign y16105 = n26348 ;
  assign y16106 = n26349 ;
  assign y16107 = ~1'b0 ;
  assign y16108 = ~1'b0 ;
  assign y16109 = ~n26356 ;
  assign y16110 = ~1'b0 ;
  assign y16111 = n26358 ;
  assign y16112 = n4341 ;
  assign y16113 = n26360 ;
  assign y16114 = ~1'b0 ;
  assign y16115 = ~n26361 ;
  assign y16116 = ~n1628 ;
  assign y16117 = n26372 ;
  assign y16118 = ~1'b0 ;
  assign y16119 = n6786 ;
  assign y16120 = n26374 ;
  assign y16121 = ~n26378 ;
  assign y16122 = n26379 ;
  assign y16123 = ~1'b0 ;
  assign y16124 = ~n26381 ;
  assign y16125 = n20959 ;
  assign y16126 = ~n26391 ;
  assign y16127 = n26392 ;
  assign y16128 = ~n26393 ;
  assign y16129 = ~n26399 ;
  assign y16130 = ~1'b0 ;
  assign y16131 = ~1'b0 ;
  assign y16132 = n26401 ;
  assign y16133 = ~n26403 ;
  assign y16134 = n26406 ;
  assign y16135 = n26407 ;
  assign y16136 = ~n26409 ;
  assign y16137 = 1'b0 ;
  assign y16138 = ~n26413 ;
  assign y16139 = n26416 ;
  assign y16140 = n26418 ;
  assign y16141 = ~1'b0 ;
  assign y16142 = 1'b0 ;
  assign y16143 = ~n26420 ;
  assign y16144 = n26421 ;
  assign y16145 = ~n26423 ;
  assign y16146 = n26428 ;
  assign y16147 = 1'b0 ;
  assign y16148 = ~n26434 ;
  assign y16149 = ~n26439 ;
  assign y16150 = ~1'b0 ;
  assign y16151 = ~n16284 ;
  assign y16152 = ~1'b0 ;
  assign y16153 = n26442 ;
  assign y16154 = ~1'b0 ;
  assign y16155 = ~1'b0 ;
  assign y16156 = ~n26445 ;
  assign y16157 = n14530 ;
  assign y16158 = ~n11125 ;
  assign y16159 = n5758 ;
  assign y16160 = ~1'b0 ;
  assign y16161 = n26448 ;
  assign y16162 = ~1'b0 ;
  assign y16163 = n26450 ;
  assign y16164 = ~n26454 ;
  assign y16165 = n26457 ;
  assign y16166 = n3895 ;
  assign y16167 = n26459 ;
  assign y16168 = ~n26460 ;
  assign y16169 = n26469 ;
  assign y16170 = ~n26473 ;
  assign y16171 = n26474 ;
  assign y16172 = n26476 ;
  assign y16173 = ~1'b0 ;
  assign y16174 = ~n26480 ;
  assign y16175 = n26481 ;
  assign y16176 = ~1'b0 ;
  assign y16177 = ~1'b0 ;
  assign y16178 = ~n26483 ;
  assign y16179 = ~n26485 ;
  assign y16180 = ~1'b0 ;
  assign y16181 = ~n26492 ;
  assign y16182 = ~1'b0 ;
  assign y16183 = ~n26493 ;
  assign y16184 = ~x219 ;
  assign y16185 = n26494 ;
  assign y16186 = n26495 ;
  assign y16187 = ~1'b0 ;
  assign y16188 = ~n26496 ;
  assign y16189 = ~1'b0 ;
  assign y16190 = ~n26500 ;
  assign y16191 = ~1'b0 ;
  assign y16192 = ~1'b0 ;
  assign y16193 = n5559 ;
  assign y16194 = 1'b0 ;
  assign y16195 = ~1'b0 ;
  assign y16196 = ~1'b0 ;
  assign y16197 = ~n26504 ;
  assign y16198 = ~1'b0 ;
  assign y16199 = ~n4047 ;
  assign y16200 = ~n26505 ;
  assign y16201 = n23386 ;
  assign y16202 = ~1'b0 ;
  assign y16203 = ~n26507 ;
  assign y16204 = ~1'b0 ;
  assign y16205 = ~n26510 ;
  assign y16206 = n26511 ;
  assign y16207 = ~n4726 ;
  assign y16208 = ~1'b0 ;
  assign y16209 = n26514 ;
  assign y16210 = ~n26515 ;
  assign y16211 = ~1'b0 ;
  assign y16212 = ~1'b0 ;
  assign y16213 = ~n26516 ;
  assign y16214 = ~n26517 ;
  assign y16215 = ~1'b0 ;
  assign y16216 = n10514 ;
  assign y16217 = ~1'b0 ;
  assign y16218 = 1'b0 ;
  assign y16219 = ~1'b0 ;
  assign y16220 = ~1'b0 ;
  assign y16221 = n12346 ;
  assign y16222 = ~1'b0 ;
  assign y16223 = ~n26521 ;
  assign y16224 = 1'b0 ;
  assign y16225 = ~n26523 ;
  assign y16226 = n26529 ;
  assign y16227 = ~1'b0 ;
  assign y16228 = ~n26533 ;
  assign y16229 = n26534 ;
  assign y16230 = ~n26537 ;
  assign y16231 = ~n26542 ;
  assign y16232 = n26544 ;
  assign y16233 = n26546 ;
  assign y16234 = ~1'b0 ;
  assign y16235 = n26549 ;
  assign y16236 = ~1'b0 ;
  assign y16237 = ~1'b0 ;
  assign y16238 = n26550 ;
  assign y16239 = n7701 ;
  assign y16240 = n26551 ;
  assign y16241 = n26554 ;
  assign y16242 = ~1'b0 ;
  assign y16243 = n26555 ;
  assign y16244 = ~1'b0 ;
  assign y16245 = ~n26557 ;
  assign y16246 = ~n26560 ;
  assign y16247 = n26565 ;
  assign y16248 = ~n26566 ;
  assign y16249 = n13095 ;
  assign y16250 = n13297 ;
  assign y16251 = ~1'b0 ;
  assign y16252 = ~1'b0 ;
  assign y16253 = ~n26570 ;
  assign y16254 = n26571 ;
  assign y16255 = ~1'b0 ;
  assign y16256 = ~1'b0 ;
  assign y16257 = ~n26577 ;
  assign y16258 = ~1'b0 ;
  assign y16259 = ~1'b0 ;
  assign y16260 = ~1'b0 ;
  assign y16261 = ~n26579 ;
  assign y16262 = n26581 ;
  assign y16263 = ~n2071 ;
  assign y16264 = 1'b0 ;
  assign y16265 = ~n26582 ;
  assign y16266 = ~n26588 ;
  assign y16267 = ~n26591 ;
  assign y16268 = ~n26593 ;
  assign y16269 = ~n26595 ;
  assign y16270 = ~1'b0 ;
  assign y16271 = ~n26596 ;
  assign y16272 = ~n26597 ;
  assign y16273 = ~1'b0 ;
  assign y16274 = n26598 ;
  assign y16275 = n21748 ;
  assign y16276 = ~n26600 ;
  assign y16277 = ~1'b0 ;
  assign y16278 = ~1'b0 ;
  assign y16279 = ~n26601 ;
  assign y16280 = n26605 ;
  assign y16281 = ~n26606 ;
  assign y16282 = ~1'b0 ;
  assign y16283 = ~1'b0 ;
  assign y16284 = ~1'b0 ;
  assign y16285 = ~1'b0 ;
  assign y16286 = ~1'b0 ;
  assign y16287 = ~1'b0 ;
  assign y16288 = ~1'b0 ;
  assign y16289 = n26609 ;
  assign y16290 = ~1'b0 ;
  assign y16291 = 1'b0 ;
  assign y16292 = 1'b0 ;
  assign y16293 = ~n26612 ;
  assign y16294 = ~1'b0 ;
  assign y16295 = n26615 ;
  assign y16296 = n26619 ;
  assign y16297 = n26624 ;
  assign y16298 = ~1'b0 ;
  assign y16299 = ~n26626 ;
  assign y16300 = ~n26628 ;
  assign y16301 = ~1'b0 ;
  assign y16302 = ~n26629 ;
  assign y16303 = n26634 ;
  assign y16304 = n26639 ;
  assign y16305 = ~1'b0 ;
  assign y16306 = n16681 ;
  assign y16307 = n26640 ;
  assign y16308 = n26643 ;
  assign y16309 = n26644 ;
  assign y16310 = n26645 ;
  assign y16311 = ~1'b0 ;
  assign y16312 = ~n26646 ;
  assign y16313 = ~1'b0 ;
  assign y16314 = n26647 ;
  assign y16315 = ~1'b0 ;
  assign y16316 = ~1'b0 ;
  assign y16317 = ~1'b0 ;
  assign y16318 = n26653 ;
  assign y16319 = n26654 ;
  assign y16320 = ~1'b0 ;
  assign y16321 = ~1'b0 ;
  assign y16322 = ~1'b0 ;
  assign y16323 = ~n26655 ;
  assign y16324 = n26659 ;
  assign y16325 = ~1'b0 ;
  assign y16326 = ~1'b0 ;
  assign y16327 = n26660 ;
  assign y16328 = ~1'b0 ;
  assign y16329 = ~1'b0 ;
  assign y16330 = ~n8056 ;
  assign y16331 = ~n26661 ;
  assign y16332 = ~1'b0 ;
  assign y16333 = ~1'b0 ;
  assign y16334 = ~n26666 ;
  assign y16335 = n26667 ;
  assign y16336 = ~1'b0 ;
  assign y16337 = ~n26668 ;
  assign y16338 = ~n26669 ;
  assign y16339 = ~1'b0 ;
  assign y16340 = n26670 ;
  assign y16341 = ~1'b0 ;
  assign y16342 = n26671 ;
  assign y16343 = ~1'b0 ;
  assign y16344 = ~1'b0 ;
  assign y16345 = ~1'b0 ;
  assign y16346 = ~n26673 ;
  assign y16347 = ~n26675 ;
  assign y16348 = ~1'b0 ;
  assign y16349 = n26676 ;
  assign y16350 = ~1'b0 ;
  assign y16351 = ~1'b0 ;
  assign y16352 = n26679 ;
  assign y16353 = ~n16135 ;
  assign y16354 = 1'b0 ;
  assign y16355 = ~1'b0 ;
  assign y16356 = ~n26684 ;
  assign y16357 = n26686 ;
  assign y16358 = ~n26688 ;
  assign y16359 = ~n20430 ;
  assign y16360 = ~n26689 ;
  assign y16361 = ~n26698 ;
  assign y16362 = 1'b0 ;
  assign y16363 = ~1'b0 ;
  assign y16364 = ~1'b0 ;
  assign y16365 = ~1'b0 ;
  assign y16366 = ~n26699 ;
  assign y16367 = n26701 ;
  assign y16368 = n26704 ;
  assign y16369 = n26708 ;
  assign y16370 = ~n26709 ;
  assign y16371 = n26713 ;
  assign y16372 = n26715 ;
  assign y16373 = ~n20619 ;
  assign y16374 = ~n26718 ;
  assign y16375 = n26723 ;
  assign y16376 = n4423 ;
  assign y16377 = ~n26724 ;
  assign y16378 = n26730 ;
  assign y16379 = n22161 ;
  assign y16380 = n26734 ;
  assign y16381 = ~1'b0 ;
  assign y16382 = 1'b0 ;
  assign y16383 = n26736 ;
  assign y16384 = ~n26737 ;
  assign y16385 = n26740 ;
  assign y16386 = n26743 ;
  assign y16387 = n26748 ;
  assign y16388 = n26750 ;
  assign y16389 = n26755 ;
  assign y16390 = ~n26756 ;
  assign y16391 = ~n26760 ;
  assign y16392 = ~n26762 ;
  assign y16393 = ~n26768 ;
  assign y16394 = ~n838 ;
  assign y16395 = ~1'b0 ;
  assign y16396 = ~n26770 ;
  assign y16397 = ~1'b0 ;
  assign y16398 = ~n26771 ;
  assign y16399 = ~n26777 ;
  assign y16400 = ~n26779 ;
  assign y16401 = ~n26781 ;
  assign y16402 = n26783 ;
  assign y16403 = ~1'b0 ;
  assign y16404 = ~1'b0 ;
  assign y16405 = ~n20430 ;
  assign y16406 = n26791 ;
  assign y16407 = n5189 ;
  assign y16408 = ~n26795 ;
  assign y16409 = ~1'b0 ;
  assign y16410 = ~n26798 ;
  assign y16411 = n26802 ;
  assign y16412 = ~1'b0 ;
  assign y16413 = ~1'b0 ;
  assign y16414 = n26803 ;
  assign y16415 = ~n26804 ;
  assign y16416 = ~1'b0 ;
  assign y16417 = n26806 ;
  assign y16418 = ~n26808 ;
  assign y16419 = ~1'b0 ;
  assign y16420 = ~n26809 ;
  assign y16421 = ~n16039 ;
  assign y16422 = n9326 ;
  assign y16423 = n25376 ;
  assign y16424 = ~1'b0 ;
  assign y16425 = ~1'b0 ;
  assign y16426 = ~1'b0 ;
  assign y16427 = ~n26812 ;
  assign y16428 = ~1'b0 ;
  assign y16429 = n26813 ;
  assign y16430 = ~1'b0 ;
  assign y16431 = ~1'b0 ;
  assign y16432 = n26695 ;
  assign y16433 = ~1'b0 ;
  assign y16434 = ~n26815 ;
  assign y16435 = n26819 ;
  assign y16436 = ~1'b0 ;
  assign y16437 = ~n26823 ;
  assign y16438 = n26830 ;
  assign y16439 = n26833 ;
  assign y16440 = ~n26834 ;
  assign y16441 = ~1'b0 ;
  assign y16442 = n26835 ;
  assign y16443 = ~1'b0 ;
  assign y16444 = n26836 ;
  assign y16445 = ~n26837 ;
  assign y16446 = n26841 ;
  assign y16447 = n26842 ;
  assign y16448 = n10531 ;
  assign y16449 = n26843 ;
  assign y16450 = ~n26844 ;
  assign y16451 = n26848 ;
  assign y16452 = n26850 ;
  assign y16453 = ~1'b0 ;
  assign y16454 = n26852 ;
  assign y16455 = ~n20220 ;
  assign y16456 = 1'b0 ;
  assign y16457 = ~1'b0 ;
  assign y16458 = ~1'b0 ;
  assign y16459 = 1'b0 ;
  assign y16460 = ~n26856 ;
  assign y16461 = ~n26858 ;
  assign y16462 = n26862 ;
  assign y16463 = n26864 ;
  assign y16464 = n26865 ;
  assign y16465 = n12225 ;
  assign y16466 = n26867 ;
  assign y16467 = ~n26871 ;
  assign y16468 = n26876 ;
  assign y16469 = ~1'b0 ;
  assign y16470 = ~n26879 ;
  assign y16471 = ~n26881 ;
  assign y16472 = n26882 ;
  assign y16473 = ~n12928 ;
  assign y16474 = n26884 ;
  assign y16475 = n26885 ;
  assign y16476 = n26888 ;
  assign y16477 = ~n26893 ;
  assign y16478 = n26894 ;
  assign y16479 = ~n26896 ;
  assign y16480 = ~n20626 ;
  assign y16481 = ~1'b0 ;
  assign y16482 = ~n26899 ;
  assign y16483 = n26901 ;
  assign y16484 = ~1'b0 ;
  assign y16485 = 1'b0 ;
  assign y16486 = n26903 ;
  assign y16487 = n13449 ;
  assign y16488 = ~1'b0 ;
  assign y16489 = ~n12721 ;
  assign y16490 = n26905 ;
  assign y16491 = ~n26907 ;
  assign y16492 = ~n26916 ;
  assign y16493 = ~1'b0 ;
  assign y16494 = ~n26919 ;
  assign y16495 = ~n26923 ;
  assign y16496 = ~1'b0 ;
  assign y16497 = ~n14995 ;
  assign y16498 = n26926 ;
  assign y16499 = ~n26927 ;
  assign y16500 = n26928 ;
  assign y16501 = ~n26929 ;
  assign y16502 = n26932 ;
  assign y16503 = ~1'b0 ;
  assign y16504 = ~1'b0 ;
  assign y16505 = n26934 ;
  assign y16506 = ~1'b0 ;
  assign y16507 = n26939 ;
  assign y16508 = ~n14279 ;
  assign y16509 = ~n26941 ;
  assign y16510 = ~1'b0 ;
  assign y16511 = ~1'b0 ;
  assign y16512 = n26946 ;
  assign y16513 = ~n26948 ;
  assign y16514 = ~n26949 ;
  assign y16515 = n26950 ;
  assign y16516 = ~n26952 ;
  assign y16517 = n26955 ;
  assign y16518 = ~n26957 ;
  assign y16519 = ~1'b0 ;
  assign y16520 = ~n26964 ;
  assign y16521 = ~1'b0 ;
  assign y16522 = ~n26966 ;
  assign y16523 = ~1'b0 ;
  assign y16524 = ~1'b0 ;
  assign y16525 = n571 ;
  assign y16526 = ~1'b0 ;
  assign y16527 = ~1'b0 ;
  assign y16528 = ~n26968 ;
  assign y16529 = n26970 ;
  assign y16530 = ~1'b0 ;
  assign y16531 = n26973 ;
  assign y16532 = ~n26975 ;
  assign y16533 = n26976 ;
  assign y16534 = ~1'b0 ;
  assign y16535 = n26978 ;
  assign y16536 = ~n26980 ;
  assign y16537 = ~n26982 ;
  assign y16538 = ~n26983 ;
  assign y16539 = n26986 ;
  assign y16540 = ~n26989 ;
  assign y16541 = n26990 ;
  assign y16542 = ~n26994 ;
  assign y16543 = ~1'b0 ;
  assign y16544 = ~n26995 ;
  assign y16545 = ~1'b0 ;
  assign y16546 = ~1'b0 ;
  assign y16547 = n10646 ;
  assign y16548 = n26996 ;
  assign y16549 = 1'b0 ;
  assign y16550 = ~1'b0 ;
  assign y16551 = n26997 ;
  assign y16552 = ~n27001 ;
  assign y16553 = n27003 ;
  assign y16554 = ~1'b0 ;
  assign y16555 = ~n27004 ;
  assign y16556 = n27012 ;
  assign y16557 = ~n27013 ;
  assign y16558 = ~n27019 ;
  assign y16559 = n27024 ;
  assign y16560 = ~1'b0 ;
  assign y16561 = n27031 ;
  assign y16562 = ~n27032 ;
  assign y16563 = n27035 ;
  assign y16564 = ~n27039 ;
  assign y16565 = ~n9385 ;
  assign y16566 = ~1'b0 ;
  assign y16567 = ~1'b0 ;
  assign y16568 = n27045 ;
  assign y16569 = ~n27048 ;
  assign y16570 = ~n27049 ;
  assign y16571 = n27050 ;
  assign y16572 = n27052 ;
  assign y16573 = 1'b0 ;
  assign y16574 = n27054 ;
  assign y16575 = n27056 ;
  assign y16576 = n27057 ;
  assign y16577 = n6076 ;
  assign y16578 = ~1'b0 ;
  assign y16579 = ~1'b0 ;
  assign y16580 = ~1'b0 ;
  assign y16581 = ~n27066 ;
  assign y16582 = n21062 ;
  assign y16583 = ~n27067 ;
  assign y16584 = n261 ;
  assign y16585 = ~n27071 ;
  assign y16586 = ~n27072 ;
  assign y16587 = n1867 ;
  assign y16588 = ~1'b0 ;
  assign y16589 = n27073 ;
  assign y16590 = n27074 ;
  assign y16591 = ~1'b0 ;
  assign y16592 = n27079 ;
  assign y16593 = ~1'b0 ;
  assign y16594 = ~n23051 ;
  assign y16595 = ~n27083 ;
  assign y16596 = ~1'b0 ;
  assign y16597 = ~1'b0 ;
  assign y16598 = ~n27084 ;
  assign y16599 = ~1'b0 ;
  assign y16600 = n14449 ;
  assign y16601 = 1'b0 ;
  assign y16602 = ~1'b0 ;
  assign y16603 = n5305 ;
  assign y16604 = n27085 ;
  assign y16605 = ~n27086 ;
  assign y16606 = ~n27088 ;
  assign y16607 = ~1'b0 ;
  assign y16608 = ~n27089 ;
  assign y16609 = ~1'b0 ;
  assign y16610 = n27090 ;
  assign y16611 = ~1'b0 ;
  assign y16612 = ~n27091 ;
  assign y16613 = ~n27092 ;
  assign y16614 = ~n27093 ;
  assign y16615 = ~1'b0 ;
  assign y16616 = ~1'b0 ;
  assign y16617 = ~n27099 ;
  assign y16618 = ~1'b0 ;
  assign y16619 = n27101 ;
  assign y16620 = ~1'b0 ;
  assign y16621 = 1'b0 ;
  assign y16622 = n22795 ;
  assign y16623 = n2436 ;
  assign y16624 = ~1'b0 ;
  assign y16625 = n27106 ;
  assign y16626 = n27107 ;
  assign y16627 = ~1'b0 ;
  assign y16628 = ~n27108 ;
  assign y16629 = ~1'b0 ;
  assign y16630 = ~1'b0 ;
  assign y16631 = ~n27109 ;
  assign y16632 = ~n27115 ;
  assign y16633 = ~1'b0 ;
  assign y16634 = ~n27117 ;
  assign y16635 = 1'b0 ;
  assign y16636 = n27120 ;
  assign y16637 = n27121 ;
  assign y16638 = n27122 ;
  assign y16639 = ~1'b0 ;
  assign y16640 = ~n27123 ;
  assign y16641 = n27127 ;
  assign y16642 = ~1'b0 ;
  assign y16643 = ~n27131 ;
  assign y16644 = ~1'b0 ;
  assign y16645 = n27132 ;
  assign y16646 = ~n27136 ;
  assign y16647 = ~n7613 ;
  assign y16648 = n27142 ;
  assign y16649 = ~n27145 ;
  assign y16650 = ~1'b0 ;
  assign y16651 = n27146 ;
  assign y16652 = ~1'b0 ;
  assign y16653 = n5631 ;
  assign y16654 = n27147 ;
  assign y16655 = ~n6357 ;
  assign y16656 = ~n27148 ;
  assign y16657 = n15248 ;
  assign y16658 = n27149 ;
  assign y16659 = ~n27151 ;
  assign y16660 = ~n6582 ;
  assign y16661 = n27153 ;
  assign y16662 = n27160 ;
  assign y16663 = ~1'b0 ;
  assign y16664 = ~n27161 ;
  assign y16665 = ~1'b0 ;
  assign y16666 = ~1'b0 ;
  assign y16667 = ~n27163 ;
  assign y16668 = ~n3581 ;
  assign y16669 = ~n27165 ;
  assign y16670 = ~n27174 ;
  assign y16671 = ~1'b0 ;
  assign y16672 = n27177 ;
  assign y16673 = ~1'b0 ;
  assign y16674 = ~1'b0 ;
  assign y16675 = ~1'b0 ;
  assign y16676 = n27181 ;
  assign y16677 = ~1'b0 ;
  assign y16678 = n27182 ;
  assign y16679 = ~n27184 ;
  assign y16680 = 1'b0 ;
  assign y16681 = n27185 ;
  assign y16682 = ~1'b0 ;
  assign y16683 = n12691 ;
  assign y16684 = ~1'b0 ;
  assign y16685 = ~1'b0 ;
  assign y16686 = n27190 ;
  assign y16687 = ~n27192 ;
  assign y16688 = n27195 ;
  assign y16689 = n16882 ;
  assign y16690 = 1'b0 ;
  assign y16691 = ~1'b0 ;
  assign y16692 = ~n27202 ;
  assign y16693 = n27204 ;
  assign y16694 = n27206 ;
  assign y16695 = n27210 ;
  assign y16696 = ~n27213 ;
  assign y16697 = n27216 ;
  assign y16698 = n27219 ;
  assign y16699 = ~n27221 ;
  assign y16700 = ~1'b0 ;
  assign y16701 = n27224 ;
  assign y16702 = ~n27226 ;
  assign y16703 = ~1'b0 ;
  assign y16704 = ~1'b0 ;
  assign y16705 = ~n27228 ;
  assign y16706 = ~1'b0 ;
  assign y16707 = ~1'b0 ;
  assign y16708 = ~1'b0 ;
  assign y16709 = n14131 ;
  assign y16710 = n27229 ;
  assign y16711 = 1'b0 ;
  assign y16712 = ~n683 ;
  assign y16713 = n27230 ;
  assign y16714 = ~1'b0 ;
  assign y16715 = ~1'b0 ;
  assign y16716 = n4848 ;
  assign y16717 = ~1'b0 ;
  assign y16718 = ~1'b0 ;
  assign y16719 = ~1'b0 ;
  assign y16720 = n27232 ;
  assign y16721 = n27233 ;
  assign y16722 = n27243 ;
  assign y16723 = ~n27245 ;
  assign y16724 = ~n27247 ;
  assign y16725 = ~1'b0 ;
  assign y16726 = ~1'b0 ;
  assign y16727 = n27251 ;
  assign y16728 = ~1'b0 ;
  assign y16729 = ~1'b0 ;
  assign y16730 = ~n27254 ;
  assign y16731 = ~n27259 ;
  assign y16732 = ~1'b0 ;
  assign y16733 = ~n27264 ;
  assign y16734 = ~1'b0 ;
  assign y16735 = ~n27266 ;
  assign y16736 = ~1'b0 ;
  assign y16737 = n27267 ;
  assign y16738 = ~n27268 ;
  assign y16739 = ~1'b0 ;
  assign y16740 = n27269 ;
  assign y16741 = ~1'b0 ;
  assign y16742 = n27273 ;
  assign y16743 = ~1'b0 ;
  assign y16744 = ~n12330 ;
  assign y16745 = ~n27274 ;
  assign y16746 = ~1'b0 ;
  assign y16747 = ~n425 ;
  assign y16748 = ~n307 ;
  assign y16749 = n27276 ;
  assign y16750 = 1'b0 ;
  assign y16751 = ~1'b0 ;
  assign y16752 = n27280 ;
  assign y16753 = ~1'b0 ;
  assign y16754 = n27285 ;
  assign y16755 = n27287 ;
  assign y16756 = ~n27290 ;
  assign y16757 = n27291 ;
  assign y16758 = ~n15927 ;
  assign y16759 = ~n7892 ;
  assign y16760 = n27298 ;
  assign y16761 = n27299 ;
  assign y16762 = n27302 ;
  assign y16763 = n27303 ;
  assign y16764 = ~n27304 ;
  assign y16765 = ~1'b0 ;
  assign y16766 = 1'b0 ;
  assign y16767 = ~n27307 ;
  assign y16768 = ~n27311 ;
  assign y16769 = n27318 ;
  assign y16770 = ~n27323 ;
  assign y16771 = ~n27327 ;
  assign y16772 = n27328 ;
  assign y16773 = ~n27330 ;
  assign y16774 = ~1'b0 ;
  assign y16775 = ~n27334 ;
  assign y16776 = n5050 ;
  assign y16777 = ~n27337 ;
  assign y16778 = ~1'b0 ;
  assign y16779 = ~n5282 ;
  assign y16780 = ~1'b0 ;
  assign y16781 = n27344 ;
  assign y16782 = ~1'b0 ;
  assign y16783 = ~1'b0 ;
  assign y16784 = ~n27346 ;
  assign y16785 = ~n27347 ;
  assign y16786 = n2357 ;
  assign y16787 = n27348 ;
  assign y16788 = n27353 ;
  assign y16789 = n27355 ;
  assign y16790 = n25138 ;
  assign y16791 = n27359 ;
  assign y16792 = ~1'b0 ;
  assign y16793 = n27360 ;
  assign y16794 = ~n27365 ;
  assign y16795 = ~1'b0 ;
  assign y16796 = n27368 ;
  assign y16797 = ~n27372 ;
  assign y16798 = ~n14523 ;
  assign y16799 = ~1'b0 ;
  assign y16800 = ~n27375 ;
  assign y16801 = n27377 ;
  assign y16802 = ~1'b0 ;
  assign y16803 = n27380 ;
  assign y16804 = n27386 ;
  assign y16805 = ~1'b0 ;
  assign y16806 = n27389 ;
  assign y16807 = n27390 ;
  assign y16808 = n27395 ;
  assign y16809 = n27397 ;
  assign y16810 = ~n27399 ;
  assign y16811 = ~1'b0 ;
  assign y16812 = n27400 ;
  assign y16813 = ~n27401 ;
  assign y16814 = 1'b0 ;
  assign y16815 = ~1'b0 ;
  assign y16816 = ~n27402 ;
  assign y16817 = ~n27404 ;
  assign y16818 = 1'b0 ;
  assign y16819 = ~n27405 ;
  assign y16820 = ~1'b0 ;
  assign y16821 = ~1'b0 ;
  assign y16822 = ~1'b0 ;
  assign y16823 = n27406 ;
  assign y16824 = ~1'b0 ;
  assign y16825 = n27409 ;
  assign y16826 = ~n27413 ;
  assign y16827 = ~n27416 ;
  assign y16828 = n27417 ;
  assign y16829 = ~1'b0 ;
  assign y16830 = ~n27421 ;
  assign y16831 = ~n27423 ;
  assign y16832 = ~1'b0 ;
  assign y16833 = 1'b0 ;
  assign y16834 = ~n27424 ;
  assign y16835 = n27428 ;
  assign y16836 = ~1'b0 ;
  assign y16837 = ~n27430 ;
  assign y16838 = ~n5489 ;
  assign y16839 = n27437 ;
  assign y16840 = ~n9779 ;
  assign y16841 = ~1'b0 ;
  assign y16842 = ~n27439 ;
  assign y16843 = ~n27442 ;
  assign y16844 = ~1'b0 ;
  assign y16845 = ~1'b0 ;
  assign y16846 = ~n27448 ;
  assign y16847 = ~1'b0 ;
  assign y16848 = n27451 ;
  assign y16849 = ~1'b0 ;
  assign y16850 = ~1'b0 ;
  assign y16851 = ~1'b0 ;
  assign y16852 = n27452 ;
  assign y16853 = ~1'b0 ;
  assign y16854 = ~1'b0 ;
  assign y16855 = n27453 ;
  assign y16856 = ~n3499 ;
  assign y16857 = n27455 ;
  assign y16858 = ~n27457 ;
  assign y16859 = ~n27459 ;
  assign y16860 = ~1'b0 ;
  assign y16861 = ~1'b0 ;
  assign y16862 = n27464 ;
  assign y16863 = ~n27465 ;
  assign y16864 = n27466 ;
  assign y16865 = ~n27467 ;
  assign y16866 = ~n27471 ;
  assign y16867 = ~n24480 ;
  assign y16868 = n27473 ;
  assign y16869 = n27474 ;
  assign y16870 = ~1'b0 ;
  assign y16871 = ~1'b0 ;
  assign y16872 = n27477 ;
  assign y16873 = ~1'b0 ;
  assign y16874 = n11001 ;
  assign y16875 = ~n27478 ;
  assign y16876 = n27479 ;
  assign y16877 = ~1'b0 ;
  assign y16878 = ~1'b0 ;
  assign y16879 = ~1'b0 ;
  assign y16880 = ~n27480 ;
  assign y16881 = ~1'b0 ;
  assign y16882 = n27482 ;
  assign y16883 = ~n27484 ;
  assign y16884 = n27485 ;
  assign y16885 = ~n27487 ;
  assign y16886 = ~1'b0 ;
  assign y16887 = ~n23280 ;
  assign y16888 = ~n27488 ;
  assign y16889 = n27491 ;
  assign y16890 = ~n27492 ;
  assign y16891 = n25105 ;
  assign y16892 = n9339 ;
  assign y16893 = n27493 ;
  assign y16894 = n5744 ;
  assign y16895 = ~1'b0 ;
  assign y16896 = ~1'b0 ;
  assign y16897 = ~n27494 ;
  assign y16898 = ~n1658 ;
  assign y16899 = ~n27496 ;
  assign y16900 = n27497 ;
  assign y16901 = ~1'b0 ;
  assign y16902 = ~n27498 ;
  assign y16903 = ~1'b0 ;
  assign y16904 = ~n27499 ;
  assign y16905 = ~1'b0 ;
  assign y16906 = ~1'b0 ;
  assign y16907 = n27500 ;
  assign y16908 = n27501 ;
  assign y16909 = ~n27504 ;
  assign y16910 = ~n27505 ;
  assign y16911 = ~n27506 ;
  assign y16912 = ~1'b0 ;
  assign y16913 = ~1'b0 ;
  assign y16914 = ~1'b0 ;
  assign y16915 = n6944 ;
  assign y16916 = ~n27508 ;
  assign y16917 = ~n27511 ;
  assign y16918 = ~1'b0 ;
  assign y16919 = ~n27512 ;
  assign y16920 = n27513 ;
  assign y16921 = ~n27514 ;
  assign y16922 = ~n13331 ;
  assign y16923 = n20931 ;
  assign y16924 = ~1'b0 ;
  assign y16925 = ~n27517 ;
  assign y16926 = ~1'b0 ;
  assign y16927 = ~n27519 ;
  assign y16928 = n24139 ;
  assign y16929 = ~n27523 ;
  assign y16930 = ~n27526 ;
  assign y16931 = ~1'b0 ;
  assign y16932 = n27527 ;
  assign y16933 = ~1'b0 ;
  assign y16934 = ~n27529 ;
  assign y16935 = ~1'b0 ;
  assign y16936 = ~n27531 ;
  assign y16937 = ~1'b0 ;
  assign y16938 = ~1'b0 ;
  assign y16939 = ~n27532 ;
  assign y16940 = n27533 ;
  assign y16941 = ~1'b0 ;
  assign y16942 = ~1'b0 ;
  assign y16943 = ~1'b0 ;
  assign y16944 = ~n27534 ;
  assign y16945 = ~1'b0 ;
  assign y16946 = ~n27536 ;
  assign y16947 = ~1'b0 ;
  assign y16948 = ~n27540 ;
  assign y16949 = ~1'b0 ;
  assign y16950 = ~1'b0 ;
  assign y16951 = n27544 ;
  assign y16952 = ~1'b0 ;
  assign y16953 = ~x76 ;
  assign y16954 = ~n27545 ;
  assign y16955 = ~n27546 ;
  assign y16956 = n27547 ;
  assign y16957 = n27551 ;
  assign y16958 = ~1'b0 ;
  assign y16959 = n27553 ;
  assign y16960 = n27555 ;
  assign y16961 = 1'b0 ;
  assign y16962 = ~1'b0 ;
  assign y16963 = n27556 ;
  assign y16964 = ~n27558 ;
  assign y16965 = n27559 ;
  assign y16966 = 1'b0 ;
  assign y16967 = ~1'b0 ;
  assign y16968 = n25101 ;
  assign y16969 = ~n27560 ;
  assign y16970 = ~n27562 ;
  assign y16971 = ~n27568 ;
  assign y16972 = ~n27569 ;
  assign y16973 = ~1'b0 ;
  assign y16974 = ~n27571 ;
  assign y16975 = 1'b0 ;
  assign y16976 = ~1'b0 ;
  assign y16977 = n27575 ;
  assign y16978 = ~1'b0 ;
  assign y16979 = n27577 ;
  assign y16980 = ~n27578 ;
  assign y16981 = n27580 ;
  assign y16982 = ~n27584 ;
  assign y16983 = n27586 ;
  assign y16984 = ~n27588 ;
  assign y16985 = n27590 ;
  assign y16986 = n27593 ;
  assign y16987 = ~n27594 ;
  assign y16988 = n27595 ;
  assign y16989 = ~n27598 ;
  assign y16990 = ~n27601 ;
  assign y16991 = ~n27602 ;
  assign y16992 = ~n27606 ;
  assign y16993 = ~n10174 ;
  assign y16994 = ~n27607 ;
  assign y16995 = ~1'b0 ;
  assign y16996 = n27608 ;
  assign y16997 = ~n27610 ;
  assign y16998 = ~1'b0 ;
  assign y16999 = ~n27611 ;
  assign y17000 = ~1'b0 ;
  assign y17001 = n7061 ;
  assign y17002 = ~n27612 ;
  assign y17003 = n27623 ;
  assign y17004 = ~1'b0 ;
  assign y17005 = ~n27626 ;
  assign y17006 = n27630 ;
  assign y17007 = ~1'b0 ;
  assign y17008 = n27633 ;
  assign y17009 = n27634 ;
  assign y17010 = ~n27637 ;
  assign y17011 = ~1'b0 ;
  assign y17012 = n27641 ;
  assign y17013 = ~1'b0 ;
  assign y17014 = ~1'b0 ;
  assign y17015 = n27642 ;
  assign y17016 = ~1'b0 ;
  assign y17017 = n27647 ;
  assign y17018 = ~1'b0 ;
  assign y17019 = ~1'b0 ;
  assign y17020 = n27649 ;
  assign y17021 = n27650 ;
  assign y17022 = ~1'b0 ;
  assign y17023 = ~n27653 ;
  assign y17024 = ~1'b0 ;
  assign y17025 = n27656 ;
  assign y17026 = n27657 ;
  assign y17027 = n27661 ;
  assign y17028 = n23236 ;
  assign y17029 = n27663 ;
  assign y17030 = ~1'b0 ;
  assign y17031 = ~1'b0 ;
  assign y17032 = ~n27664 ;
  assign y17033 = ~n27670 ;
  assign y17034 = ~n27672 ;
  assign y17035 = ~n27676 ;
  assign y17036 = n25252 ;
  assign y17037 = ~1'b0 ;
  assign y17038 = ~1'b0 ;
  assign y17039 = n27678 ;
  assign y17040 = ~n27679 ;
  assign y17041 = ~1'b0 ;
  assign y17042 = ~1'b0 ;
  assign y17043 = ~1'b0 ;
  assign y17044 = ~n27682 ;
  assign y17045 = n27685 ;
  assign y17046 = n27686 ;
  assign y17047 = n27688 ;
  assign y17048 = 1'b0 ;
  assign y17049 = ~n27689 ;
  assign y17050 = ~1'b0 ;
  assign y17051 = ~n27691 ;
  assign y17052 = ~n27693 ;
  assign y17053 = n27696 ;
  assign y17054 = ~n27699 ;
  assign y17055 = ~n27700 ;
  assign y17056 = ~1'b0 ;
  assign y17057 = ~n27702 ;
  assign y17058 = ~n27704 ;
  assign y17059 = ~n27707 ;
  assign y17060 = ~n27709 ;
  assign y17061 = ~1'b0 ;
  assign y17062 = ~1'b0 ;
  assign y17063 = ~n27711 ;
  assign y17064 = ~1'b0 ;
  assign y17065 = n27712 ;
  assign y17066 = ~1'b0 ;
  assign y17067 = ~n27716 ;
  assign y17068 = ~n27718 ;
  assign y17069 = n27720 ;
  assign y17070 = ~1'b0 ;
  assign y17071 = n27722 ;
  assign y17072 = n27723 ;
  assign y17073 = n27725 ;
  assign y17074 = ~1'b0 ;
  assign y17075 = ~1'b0 ;
  assign y17076 = ~n27726 ;
  assign y17077 = n27727 ;
  assign y17078 = ~n27730 ;
  assign y17079 = ~1'b0 ;
  assign y17080 = n27732 ;
  assign y17081 = ~n27733 ;
  assign y17082 = ~n27735 ;
  assign y17083 = n27736 ;
  assign y17084 = ~1'b0 ;
  assign y17085 = ~1'b0 ;
  assign y17086 = ~n27738 ;
  assign y17087 = n27741 ;
  assign y17088 = ~n27743 ;
  assign y17089 = ~1'b0 ;
  assign y17090 = n27746 ;
  assign y17091 = n27747 ;
  assign y17092 = n27748 ;
  assign y17093 = ~1'b0 ;
  assign y17094 = ~n27750 ;
  assign y17095 = n27753 ;
  assign y17096 = ~1'b0 ;
  assign y17097 = ~1'b0 ;
  assign y17098 = ~1'b0 ;
  assign y17099 = ~n27757 ;
  assign y17100 = ~1'b0 ;
  assign y17101 = ~1'b0 ;
  assign y17102 = 1'b0 ;
  assign y17103 = 1'b0 ;
  assign y17104 = ~1'b0 ;
  assign y17105 = ~n574 ;
  assign y17106 = ~1'b0 ;
  assign y17107 = n27758 ;
  assign y17108 = ~n27767 ;
  assign y17109 = n6991 ;
  assign y17110 = n27769 ;
  assign y17111 = n27771 ;
  assign y17112 = ~n27772 ;
  assign y17113 = ~1'b0 ;
  assign y17114 = ~1'b0 ;
  assign y17115 = ~1'b0 ;
  assign y17116 = ~n27775 ;
  assign y17117 = ~x162 ;
  assign y17118 = n11357 ;
  assign y17119 = ~n27778 ;
  assign y17120 = 1'b0 ;
  assign y17121 = n27779 ;
  assign y17122 = ~n27781 ;
  assign y17123 = n27782 ;
  assign y17124 = ~1'b0 ;
  assign y17125 = ~1'b0 ;
  assign y17126 = ~1'b0 ;
  assign y17127 = n27785 ;
  assign y17128 = ~n27787 ;
  assign y17129 = ~n27790 ;
  assign y17130 = ~1'b0 ;
  assign y17131 = ~n27794 ;
  assign y17132 = ~1'b0 ;
  assign y17133 = ~1'b0 ;
  assign y17134 = ~n27795 ;
  assign y17135 = ~1'b0 ;
  assign y17136 = ~n27800 ;
  assign y17137 = ~n27805 ;
  assign y17138 = ~n2466 ;
  assign y17139 = ~1'b0 ;
  assign y17140 = ~1'b0 ;
  assign y17141 = ~1'b0 ;
  assign y17142 = ~1'b0 ;
  assign y17143 = ~n27808 ;
  assign y17144 = n26500 ;
  assign y17145 = ~n27809 ;
  assign y17146 = ~1'b0 ;
  assign y17147 = ~n27810 ;
  assign y17148 = ~n27811 ;
  assign y17149 = ~1'b0 ;
  assign y17150 = ~1'b0 ;
  assign y17151 = ~n27812 ;
  assign y17152 = ~n27817 ;
  assign y17153 = n15085 ;
  assign y17154 = ~1'b0 ;
  assign y17155 = ~n27819 ;
  assign y17156 = n27820 ;
  assign y17157 = n27821 ;
  assign y17158 = n27823 ;
  assign y17159 = ~1'b0 ;
  assign y17160 = n8131 ;
  assign y17161 = ~n27826 ;
  assign y17162 = ~1'b0 ;
  assign y17163 = ~1'b0 ;
  assign y17164 = n27827 ;
  assign y17165 = n27828 ;
  assign y17166 = ~n27830 ;
  assign y17167 = ~n27831 ;
  assign y17168 = 1'b0 ;
  assign y17169 = ~1'b0 ;
  assign y17170 = ~n27836 ;
  assign y17171 = ~1'b0 ;
  assign y17172 = ~n27840 ;
  assign y17173 = ~1'b0 ;
  assign y17174 = ~1'b0 ;
  assign y17175 = n27841 ;
  assign y17176 = ~1'b0 ;
  assign y17177 = ~1'b0 ;
  assign y17178 = ~n27842 ;
  assign y17179 = ~1'b0 ;
  assign y17180 = ~n27844 ;
  assign y17181 = ~n27846 ;
  assign y17182 = n27848 ;
  assign y17183 = ~n27851 ;
  assign y17184 = ~1'b0 ;
  assign y17185 = ~n27852 ;
  assign y17186 = ~1'b0 ;
  assign y17187 = ~1'b0 ;
  assign y17188 = ~1'b0 ;
  assign y17189 = n27854 ;
  assign y17190 = ~1'b0 ;
  assign y17191 = n27855 ;
  assign y17192 = n27887 ;
  assign y17193 = ~n27891 ;
  assign y17194 = ~n27895 ;
  assign y17195 = n27897 ;
  assign y17196 = n27898 ;
  assign y17197 = n27899 ;
  assign y17198 = ~n27900 ;
  assign y17199 = ~1'b0 ;
  assign y17200 = ~1'b0 ;
  assign y17201 = ~1'b0 ;
  assign y17202 = ~n27907 ;
  assign y17203 = n27908 ;
  assign y17204 = n25249 ;
  assign y17205 = ~1'b0 ;
  assign y17206 = ~1'b0 ;
  assign y17207 = n27909 ;
  assign y17208 = ~n9380 ;
  assign y17209 = n27910 ;
  assign y17210 = ~1'b0 ;
  assign y17211 = n27913 ;
  assign y17212 = 1'b0 ;
  assign y17213 = ~1'b0 ;
  assign y17214 = n8470 ;
  assign y17215 = ~n27914 ;
  assign y17216 = ~1'b0 ;
  assign y17217 = ~n27916 ;
  assign y17218 = ~1'b0 ;
  assign y17219 = ~n27917 ;
  assign y17220 = ~n27919 ;
  assign y17221 = ~n27920 ;
  assign y17222 = ~1'b0 ;
  assign y17223 = ~1'b0 ;
  assign y17224 = ~1'b0 ;
  assign y17225 = ~1'b0 ;
  assign y17226 = ~n27922 ;
  assign y17227 = n27924 ;
  assign y17228 = ~1'b0 ;
  assign y17229 = n27926 ;
  assign y17230 = ~n27927 ;
  assign y17231 = ~1'b0 ;
  assign y17232 = n3302 ;
  assign y17233 = ~n8436 ;
  assign y17234 = n27928 ;
  assign y17235 = n27930 ;
  assign y17236 = 1'b0 ;
  assign y17237 = 1'b0 ;
  assign y17238 = ~1'b0 ;
  assign y17239 = ~1'b0 ;
  assign y17240 = 1'b0 ;
  assign y17241 = ~1'b0 ;
  assign y17242 = ~n27932 ;
  assign y17243 = ~1'b0 ;
  assign y17244 = n27934 ;
  assign y17245 = ~n13197 ;
  assign y17246 = ~1'b0 ;
  assign y17247 = ~1'b0 ;
  assign y17248 = ~1'b0 ;
  assign y17249 = ~n7246 ;
  assign y17250 = n19507 ;
  assign y17251 = n27938 ;
  assign y17252 = ~n27939 ;
  assign y17253 = ~1'b0 ;
  assign y17254 = n27943 ;
  assign y17255 = n27944 ;
  assign y17256 = ~n27948 ;
  assign y17257 = ~n27952 ;
  assign y17258 = ~1'b0 ;
  assign y17259 = n27954 ;
  assign y17260 = n27959 ;
  assign y17261 = ~1'b0 ;
  assign y17262 = ~n27965 ;
  assign y17263 = ~1'b0 ;
  assign y17264 = ~1'b0 ;
  assign y17265 = n27967 ;
  assign y17266 = ~n27971 ;
  assign y17267 = ~1'b0 ;
  assign y17268 = ~n27973 ;
  assign y17269 = ~1'b0 ;
  assign y17270 = ~1'b0 ;
  assign y17271 = ~1'b0 ;
  assign y17272 = ~n27977 ;
  assign y17273 = ~n27978 ;
  assign y17274 = ~n27980 ;
  assign y17275 = ~1'b0 ;
  assign y17276 = ~1'b0 ;
  assign y17277 = n20177 ;
  assign y17278 = ~1'b0 ;
  assign y17279 = ~1'b0 ;
  assign y17280 = ~n27982 ;
  assign y17281 = n27984 ;
  assign y17282 = n27985 ;
  assign y17283 = n27989 ;
  assign y17284 = ~n27990 ;
  assign y17285 = 1'b0 ;
  assign y17286 = n27991 ;
  assign y17287 = ~1'b0 ;
  assign y17288 = n10364 ;
  assign y17289 = ~n27992 ;
  assign y17290 = ~1'b0 ;
  assign y17291 = ~n27993 ;
  assign y17292 = ~n23210 ;
  assign y17293 = n27996 ;
  assign y17294 = ~1'b0 ;
  assign y17295 = n27998 ;
  assign y17296 = ~1'b0 ;
  assign y17297 = ~n28000 ;
  assign y17298 = n28001 ;
  assign y17299 = ~n28003 ;
  assign y17300 = n28006 ;
  assign y17301 = ~1'b0 ;
  assign y17302 = ~n28010 ;
  assign y17303 = ~n28012 ;
  assign y17304 = n28014 ;
  assign y17305 = n28015 ;
  assign y17306 = n28017 ;
  assign y17307 = n28018 ;
  assign y17308 = n27698 ;
  assign y17309 = n28021 ;
  assign y17310 = ~1'b0 ;
  assign y17311 = ~1'b0 ;
  assign y17312 = ~1'b0 ;
  assign y17313 = ~1'b0 ;
  assign y17314 = ~n28024 ;
  assign y17315 = n28027 ;
  assign y17316 = n28028 ;
  assign y17317 = n28032 ;
  assign y17318 = ~1'b0 ;
  assign y17319 = ~n28035 ;
  assign y17320 = ~n28038 ;
  assign y17321 = ~n28041 ;
  assign y17322 = n28044 ;
  assign y17323 = n28045 ;
  assign y17324 = ~1'b0 ;
  assign y17325 = n10334 ;
  assign y17326 = n28047 ;
  assign y17327 = n28049 ;
  assign y17328 = ~1'b0 ;
  assign y17329 = ~n28052 ;
  assign y17330 = ~1'b0 ;
  assign y17331 = ~n28054 ;
  assign y17332 = n28059 ;
  assign y17333 = n28060 ;
  assign y17334 = n28062 ;
  assign y17335 = ~1'b0 ;
  assign y17336 = ~n28065 ;
  assign y17337 = ~1'b0 ;
  assign y17338 = n28066 ;
  assign y17339 = n28067 ;
  assign y17340 = n28068 ;
  assign y17341 = 1'b0 ;
  assign y17342 = ~n28069 ;
  assign y17343 = ~n9168 ;
  assign y17344 = ~1'b0 ;
  assign y17345 = ~1'b0 ;
  assign y17346 = ~n28071 ;
  assign y17347 = ~n28074 ;
  assign y17348 = ~n28075 ;
  assign y17349 = n28077 ;
  assign y17350 = ~1'b0 ;
  assign y17351 = n2457 ;
  assign y17352 = n7083 ;
  assign y17353 = ~1'b0 ;
  assign y17354 = ~1'b0 ;
  assign y17355 = ~n28081 ;
  assign y17356 = n28085 ;
  assign y17357 = ~1'b0 ;
  assign y17358 = n28086 ;
  assign y17359 = ~1'b0 ;
  assign y17360 = ~n28091 ;
  assign y17361 = ~n28092 ;
  assign y17362 = n28108 ;
  assign y17363 = ~n28109 ;
  assign y17364 = n28111 ;
  assign y17365 = ~n28114 ;
  assign y17366 = ~n28115 ;
  assign y17367 = n28116 ;
  assign y17368 = n28124 ;
  assign y17369 = n28125 ;
  assign y17370 = ~n28128 ;
  assign y17371 = ~n14248 ;
  assign y17372 = ~1'b0 ;
  assign y17373 = n28132 ;
  assign y17374 = ~n28133 ;
  assign y17375 = ~n28136 ;
  assign y17376 = n28138 ;
  assign y17377 = ~n2766 ;
  assign y17378 = ~n28140 ;
  assign y17379 = ~n28150 ;
  assign y17380 = n28152 ;
  assign y17381 = ~1'b0 ;
  assign y17382 = ~n28154 ;
  assign y17383 = n28155 ;
  assign y17384 = n28159 ;
  assign y17385 = ~1'b0 ;
  assign y17386 = 1'b0 ;
  assign y17387 = n28160 ;
  assign y17388 = ~n28161 ;
  assign y17389 = ~1'b0 ;
  assign y17390 = ~1'b0 ;
  assign y17391 = ~1'b0 ;
  assign y17392 = ~n28163 ;
  assign y17393 = ~1'b0 ;
  assign y17394 = ~1'b0 ;
  assign y17395 = ~n28169 ;
  assign y17396 = ~1'b0 ;
  assign y17397 = ~1'b0 ;
  assign y17398 = ~1'b0 ;
  assign y17399 = ~n9135 ;
  assign y17400 = ~1'b0 ;
  assign y17401 = n28171 ;
  assign y17402 = ~1'b0 ;
  assign y17403 = n4993 ;
  assign y17404 = ~1'b0 ;
  assign y17405 = ~n28174 ;
  assign y17406 = ~1'b0 ;
  assign y17407 = ~1'b0 ;
  assign y17408 = 1'b0 ;
  assign y17409 = ~1'b0 ;
  assign y17410 = n12011 ;
  assign y17411 = n28177 ;
  assign y17412 = n28184 ;
  assign y17413 = n28187 ;
  assign y17414 = n538 ;
  assign y17415 = ~n28188 ;
  assign y17416 = ~n28195 ;
  assign y17417 = ~1'b0 ;
  assign y17418 = ~1'b0 ;
  assign y17419 = ~n28202 ;
  assign y17420 = ~1'b0 ;
  assign y17421 = n28203 ;
  assign y17422 = ~1'b0 ;
  assign y17423 = ~n28209 ;
  assign y17424 = ~1'b0 ;
  assign y17425 = ~1'b0 ;
  assign y17426 = ~1'b0 ;
  assign y17427 = n28211 ;
  assign y17428 = ~1'b0 ;
  assign y17429 = ~1'b0 ;
  assign y17430 = ~n28212 ;
  assign y17431 = n28216 ;
  assign y17432 = n28219 ;
  assign y17433 = n28225 ;
  assign y17434 = n28236 ;
  assign y17435 = ~n12359 ;
  assign y17436 = ~1'b0 ;
  assign y17437 = ~1'b0 ;
  assign y17438 = ~1'b0 ;
  assign y17439 = ~1'b0 ;
  assign y17440 = ~n28238 ;
  assign y17441 = ~n28242 ;
  assign y17442 = ~n28243 ;
  assign y17443 = n28245 ;
  assign y17444 = ~1'b0 ;
  assign y17445 = ~n28246 ;
  assign y17446 = n28248 ;
  assign y17447 = n28249 ;
  assign y17448 = ~n15267 ;
  assign y17449 = ~n28250 ;
  assign y17450 = n28254 ;
  assign y17451 = ~n9225 ;
  assign y17452 = n28256 ;
  assign y17453 = ~1'b0 ;
  assign y17454 = ~n28260 ;
  assign y17455 = ~1'b0 ;
  assign y17456 = ~1'b0 ;
  assign y17457 = ~n28262 ;
  assign y17458 = n28265 ;
  assign y17459 = ~1'b0 ;
  assign y17460 = ~n28266 ;
  assign y17461 = n10175 ;
  assign y17462 = n28267 ;
  assign y17463 = ~n28270 ;
  assign y17464 = n28271 ;
  assign y17465 = n5568 ;
  assign y17466 = ~n28276 ;
  assign y17467 = n28278 ;
  assign y17468 = ~n28279 ;
  assign y17469 = n28284 ;
  assign y17470 = ~n15867 ;
  assign y17471 = ~1'b0 ;
  assign y17472 = ~n28286 ;
  assign y17473 = n28291 ;
  assign y17474 = ~1'b0 ;
  assign y17475 = n28293 ;
  assign y17476 = n28296 ;
  assign y17477 = n28298 ;
  assign y17478 = n28301 ;
  assign y17479 = ~1'b0 ;
  assign y17480 = n28303 ;
  assign y17481 = ~n28305 ;
  assign y17482 = n28307 ;
  assign y17483 = n28308 ;
  assign y17484 = ~n20799 ;
  assign y17485 = ~1'b0 ;
  assign y17486 = ~n28309 ;
  assign y17487 = n28313 ;
  assign y17488 = ~1'b0 ;
  assign y17489 = n28316 ;
  assign y17490 = n28317 ;
  assign y17491 = ~n12427 ;
  assign y17492 = ~n28327 ;
  assign y17493 = ~n28330 ;
  assign y17494 = ~n9377 ;
  assign y17495 = ~n28335 ;
  assign y17496 = ~1'b0 ;
  assign y17497 = n28341 ;
  assign y17498 = ~n28344 ;
  assign y17499 = ~1'b0 ;
  assign y17500 = n28345 ;
  assign y17501 = ~1'b0 ;
  assign y17502 = ~n28349 ;
  assign y17503 = n28351 ;
  assign y17504 = ~n28353 ;
  assign y17505 = ~1'b0 ;
  assign y17506 = n28354 ;
  assign y17507 = ~n28357 ;
  assign y17508 = ~1'b0 ;
  assign y17509 = ~n28362 ;
  assign y17510 = n28363 ;
  assign y17511 = ~1'b0 ;
  assign y17512 = ~1'b0 ;
  assign y17513 = n28367 ;
  assign y17514 = n28374 ;
  assign y17515 = ~1'b0 ;
  assign y17516 = ~1'b0 ;
  assign y17517 = n28377 ;
  assign y17518 = n28381 ;
  assign y17519 = ~n28384 ;
  assign y17520 = n28385 ;
  assign y17521 = ~n28387 ;
  assign y17522 = n28392 ;
  assign y17523 = ~1'b0 ;
  assign y17524 = ~1'b0 ;
  assign y17525 = ~1'b0 ;
  assign y17526 = ~n28394 ;
  assign y17527 = ~1'b0 ;
  assign y17528 = ~n28398 ;
  assign y17529 = ~n28400 ;
  assign y17530 = n28405 ;
  assign y17531 = n28410 ;
  assign y17532 = ~n28412 ;
  assign y17533 = ~n28413 ;
  assign y17534 = n28414 ;
  assign y17535 = ~1'b0 ;
  assign y17536 = n28421 ;
  assign y17537 = ~1'b0 ;
  assign y17538 = ~n28422 ;
  assign y17539 = ~1'b0 ;
  assign y17540 = ~n28425 ;
  assign y17541 = ~n28429 ;
  assign y17542 = n28433 ;
  assign y17543 = ~n28434 ;
  assign y17544 = 1'b0 ;
  assign y17545 = ~n28436 ;
  assign y17546 = ~1'b0 ;
  assign y17547 = ~1'b0 ;
  assign y17548 = ~n28438 ;
  assign y17549 = ~1'b0 ;
  assign y17550 = ~n28439 ;
  assign y17551 = n20023 ;
  assign y17552 = x101 ;
  assign y17553 = ~1'b0 ;
  assign y17554 = ~1'b0 ;
  assign y17555 = n28440 ;
  assign y17556 = ~1'b0 ;
  assign y17557 = n28441 ;
  assign y17558 = ~1'b0 ;
  assign y17559 = ~n28445 ;
  assign y17560 = ~1'b0 ;
  assign y17561 = ~n28446 ;
  assign y17562 = n28447 ;
  assign y17563 = n28449 ;
  assign y17564 = ~n28453 ;
  assign y17565 = n28456 ;
  assign y17566 = n28462 ;
  assign y17567 = n28463 ;
  assign y17568 = ~1'b0 ;
  assign y17569 = ~1'b0 ;
  assign y17570 = ~n28476 ;
  assign y17571 = ~1'b0 ;
  assign y17572 = n28477 ;
  assign y17573 = ~n28480 ;
  assign y17574 = ~1'b0 ;
  assign y17575 = n20811 ;
  assign y17576 = ~1'b0 ;
  assign y17577 = ~1'b0 ;
  assign y17578 = ~1'b0 ;
  assign y17579 = ~n28483 ;
  assign y17580 = ~n28484 ;
  assign y17581 = n28485 ;
  assign y17582 = ~1'b0 ;
  assign y17583 = ~n28491 ;
  assign y17584 = n28498 ;
  assign y17585 = n28503 ;
  assign y17586 = ~1'b0 ;
  assign y17587 = ~1'b0 ;
  assign y17588 = ~n28506 ;
  assign y17589 = ~n14157 ;
  assign y17590 = n28513 ;
  assign y17591 = 1'b0 ;
  assign y17592 = ~n28514 ;
  assign y17593 = n28515 ;
  assign y17594 = n28517 ;
  assign y17595 = ~1'b0 ;
  assign y17596 = ~n28518 ;
  assign y17597 = ~1'b0 ;
  assign y17598 = 1'b0 ;
  assign y17599 = n28520 ;
  assign y17600 = ~1'b0 ;
  assign y17601 = ~n28523 ;
  assign y17602 = n28525 ;
  assign y17603 = n28527 ;
  assign y17604 = ~1'b0 ;
  assign y17605 = n28531 ;
  assign y17606 = n28532 ;
  assign y17607 = ~1'b0 ;
  assign y17608 = n28533 ;
  assign y17609 = ~1'b0 ;
  assign y17610 = ~n27283 ;
  assign y17611 = ~n28535 ;
  assign y17612 = ~1'b0 ;
  assign y17613 = ~1'b0 ;
  assign y17614 = n28537 ;
  assign y17615 = n25083 ;
  assign y17616 = ~n28541 ;
  assign y17617 = n28542 ;
  assign y17618 = ~1'b0 ;
  assign y17619 = n17038 ;
  assign y17620 = n28543 ;
  assign y17621 = ~1'b0 ;
  assign y17622 = ~1'b0 ;
  assign y17623 = n28546 ;
  assign y17624 = ~n28548 ;
  assign y17625 = ~1'b0 ;
  assign y17626 = n28554 ;
  assign y17627 = ~1'b0 ;
  assign y17628 = ~1'b0 ;
  assign y17629 = n28558 ;
  assign y17630 = ~n28564 ;
  assign y17631 = ~1'b0 ;
  assign y17632 = ~n28568 ;
  assign y17633 = ~n4617 ;
  assign y17634 = n20764 ;
  assign y17635 = ~n28569 ;
  assign y17636 = n28577 ;
  assign y17637 = ~1'b0 ;
  assign y17638 = ~n28581 ;
  assign y17639 = ~1'b0 ;
  assign y17640 = n28582 ;
  assign y17641 = ~n28583 ;
  assign y17642 = ~1'b0 ;
  assign y17643 = n28585 ;
  assign y17644 = n28586 ;
  assign y17645 = ~n28591 ;
  assign y17646 = ~1'b0 ;
  assign y17647 = ~n26089 ;
  assign y17648 = ~n28593 ;
  assign y17649 = n28597 ;
  assign y17650 = ~n28598 ;
  assign y17651 = ~1'b0 ;
  assign y17652 = ~1'b0 ;
  assign y17653 = ~1'b0 ;
  assign y17654 = ~n28599 ;
  assign y17655 = ~1'b0 ;
  assign y17656 = n28600 ;
  assign y17657 = n7679 ;
  assign y17658 = n28602 ;
  assign y17659 = n28603 ;
  assign y17660 = ~n28606 ;
  assign y17661 = ~n28609 ;
  assign y17662 = ~1'b0 ;
  assign y17663 = ~1'b0 ;
  assign y17664 = ~n28611 ;
  assign y17665 = ~n3091 ;
  assign y17666 = ~1'b0 ;
  assign y17667 = ~n28613 ;
  assign y17668 = n28614 ;
  assign y17669 = ~1'b0 ;
  assign y17670 = ~1'b0 ;
  assign y17671 = ~n28615 ;
  assign y17672 = ~n28617 ;
  assign y17673 = n28619 ;
  assign y17674 = ~n28620 ;
  assign y17675 = ~n28622 ;
  assign y17676 = n28623 ;
  assign y17677 = ~n19366 ;
  assign y17678 = n28625 ;
  assign y17679 = ~n855 ;
  assign y17680 = ~n28633 ;
  assign y17681 = n25872 ;
  assign y17682 = ~n28637 ;
  assign y17683 = ~n28640 ;
  assign y17684 = ~n28641 ;
  assign y17685 = ~1'b0 ;
  assign y17686 = ~n28643 ;
  assign y17687 = ~n1572 ;
  assign y17688 = ~1'b0 ;
  assign y17689 = n28645 ;
  assign y17690 = ~1'b0 ;
  assign y17691 = n28650 ;
  assign y17692 = ~n28651 ;
  assign y17693 = ~1'b0 ;
  assign y17694 = n28653 ;
  assign y17695 = ~n28657 ;
  assign y17696 = ~n28658 ;
  assign y17697 = ~1'b0 ;
  assign y17698 = n28660 ;
  assign y17699 = ~n28665 ;
  assign y17700 = ~1'b0 ;
  assign y17701 = ~1'b0 ;
  assign y17702 = ~1'b0 ;
  assign y17703 = ~n28667 ;
  assign y17704 = n1544 ;
  assign y17705 = n28668 ;
  assign y17706 = ~n28673 ;
  assign y17707 = ~1'b0 ;
  assign y17708 = ~n28674 ;
  assign y17709 = ~1'b0 ;
  assign y17710 = n28677 ;
  assign y17711 = ~1'b0 ;
  assign y17712 = ~1'b0 ;
  assign y17713 = n28678 ;
  assign y17714 = ~1'b0 ;
  assign y17715 = ~n28680 ;
  assign y17716 = ~1'b0 ;
  assign y17717 = ~1'b0 ;
  assign y17718 = ~n28681 ;
  assign y17719 = 1'b0 ;
  assign y17720 = ~n28682 ;
  assign y17721 = ~1'b0 ;
  assign y17722 = ~1'b0 ;
  assign y17723 = n28685 ;
  assign y17724 = ~n28686 ;
  assign y17725 = n28690 ;
  assign y17726 = ~n9233 ;
  assign y17727 = ~1'b0 ;
  assign y17728 = ~1'b0 ;
  assign y17729 = n28693 ;
  assign y17730 = 1'b0 ;
  assign y17731 = ~n28695 ;
  assign y17732 = ~1'b0 ;
  assign y17733 = ~n28697 ;
  assign y17734 = n28698 ;
  assign y17735 = ~n28700 ;
  assign y17736 = ~1'b0 ;
  assign y17737 = n28704 ;
  assign y17738 = ~1'b0 ;
  assign y17739 = 1'b0 ;
  assign y17740 = ~n28706 ;
  assign y17741 = ~1'b0 ;
  assign y17742 = n28707 ;
  assign y17743 = 1'b0 ;
  assign y17744 = n28708 ;
  assign y17745 = n28711 ;
  assign y17746 = ~1'b0 ;
  assign y17747 = ~1'b0 ;
  assign y17748 = ~1'b0 ;
  assign y17749 = ~n28712 ;
  assign y17750 = ~1'b0 ;
  assign y17751 = ~n28714 ;
  assign y17752 = ~1'b0 ;
  assign y17753 = ~1'b0 ;
  assign y17754 = 1'b0 ;
  assign y17755 = n3910 ;
  assign y17756 = ~n28715 ;
  assign y17757 = ~1'b0 ;
  assign y17758 = n28718 ;
  assign y17759 = ~n28720 ;
  assign y17760 = ~n28721 ;
  assign y17761 = ~n28723 ;
  assign y17762 = ~n28728 ;
  assign y17763 = ~n28730 ;
  assign y17764 = ~1'b0 ;
  assign y17765 = ~n28735 ;
  assign y17766 = ~1'b0 ;
  assign y17767 = ~n28736 ;
  assign y17768 = n28739 ;
  assign y17769 = n28742 ;
  assign y17770 = n28743 ;
  assign y17771 = 1'b0 ;
  assign y17772 = ~1'b0 ;
  assign y17773 = n28745 ;
  assign y17774 = n28746 ;
  assign y17775 = n21475 ;
  assign y17776 = ~n4791 ;
  assign y17777 = ~1'b0 ;
  assign y17778 = n28747 ;
  assign y17779 = ~n7675 ;
  assign y17780 = n28748 ;
  assign y17781 = n28749 ;
  assign y17782 = ~n28751 ;
  assign y17783 = ~1'b0 ;
  assign y17784 = ~n28752 ;
  assign y17785 = ~1'b0 ;
  assign y17786 = n28753 ;
  assign y17787 = n28757 ;
  assign y17788 = ~n28759 ;
  assign y17789 = ~n28761 ;
  assign y17790 = n28763 ;
  assign y17791 = ~1'b0 ;
  assign y17792 = n28767 ;
  assign y17793 = n28768 ;
  assign y17794 = n28772 ;
  assign y17795 = n28773 ;
  assign y17796 = ~1'b0 ;
  assign y17797 = ~n28774 ;
  assign y17798 = ~1'b0 ;
  assign y17799 = n3186 ;
  assign y17800 = ~n10669 ;
  assign y17801 = ~1'b0 ;
  assign y17802 = n28775 ;
  assign y17803 = ~n28779 ;
  assign y17804 = ~n28781 ;
  assign y17805 = ~n5959 ;
  assign y17806 = ~n259 ;
  assign y17807 = ~1'b0 ;
  assign y17808 = ~1'b0 ;
  assign y17809 = ~n28782 ;
  assign y17810 = n28783 ;
  assign y17811 = n28784 ;
  assign y17812 = ~n5852 ;
  assign y17813 = 1'b0 ;
  assign y17814 = ~1'b0 ;
  assign y17815 = ~n28785 ;
  assign y17816 = ~1'b0 ;
  assign y17817 = 1'b0 ;
  assign y17818 = n836 ;
  assign y17819 = n28786 ;
  assign y17820 = ~n28788 ;
  assign y17821 = ~1'b0 ;
  assign y17822 = ~1'b0 ;
  assign y17823 = ~1'b0 ;
  assign y17824 = ~1'b0 ;
  assign y17825 = ~1'b0 ;
  assign y17826 = 1'b0 ;
  assign y17827 = ~1'b0 ;
  assign y17828 = n28792 ;
  assign y17829 = n28798 ;
  assign y17830 = 1'b0 ;
  assign y17831 = n3825 ;
  assign y17832 = ~1'b0 ;
  assign y17833 = ~n28801 ;
  assign y17834 = n28803 ;
  assign y17835 = ~n28807 ;
  assign y17836 = ~1'b0 ;
  assign y17837 = n13029 ;
  assign y17838 = ~n28810 ;
  assign y17839 = ~n28815 ;
  assign y17840 = ~1'b0 ;
  assign y17841 = n28816 ;
  assign y17842 = ~1'b0 ;
  assign y17843 = n28817 ;
  assign y17844 = n4853 ;
  assign y17845 = ~n28819 ;
  assign y17846 = ~n28824 ;
  assign y17847 = ~n28825 ;
  assign y17848 = ~1'b0 ;
  assign y17849 = n28826 ;
  assign y17850 = ~1'b0 ;
  assign y17851 = ~1'b0 ;
  assign y17852 = ~1'b0 ;
  assign y17853 = ~n28828 ;
  assign y17854 = ~1'b0 ;
  assign y17855 = ~1'b0 ;
  assign y17856 = ~n28831 ;
  assign y17857 = n28832 ;
  assign y17858 = ~n14907 ;
  assign y17859 = ~1'b0 ;
  assign y17860 = ~1'b0 ;
  assign y17861 = ~1'b0 ;
  assign y17862 = n28834 ;
  assign y17863 = n28836 ;
  assign y17864 = ~n25249 ;
  assign y17865 = ~1'b0 ;
  assign y17866 = ~1'b0 ;
  assign y17867 = ~1'b0 ;
  assign y17868 = n28839 ;
  assign y17869 = n28840 ;
  assign y17870 = ~n28841 ;
  assign y17871 = n28842 ;
  assign y17872 = 1'b0 ;
  assign y17873 = ~1'b0 ;
  assign y17874 = ~n28843 ;
  assign y17875 = ~1'b0 ;
  assign y17876 = ~n28844 ;
  assign y17877 = n28849 ;
  assign y17878 = n28850 ;
  assign y17879 = ~1'b0 ;
  assign y17880 = ~1'b0 ;
  assign y17881 = n28853 ;
  assign y17882 = ~n28855 ;
  assign y17883 = n28856 ;
  assign y17884 = ~n415 ;
  assign y17885 = n28857 ;
  assign y17886 = n28859 ;
  assign y17887 = ~n28860 ;
  assign y17888 = ~n28861 ;
  assign y17889 = n18299 ;
  assign y17890 = ~1'b0 ;
  assign y17891 = ~n28862 ;
  assign y17892 = ~n28863 ;
  assign y17893 = ~1'b0 ;
  assign y17894 = ~n28864 ;
  assign y17895 = n28866 ;
  assign y17896 = ~1'b0 ;
  assign y17897 = n8536 ;
  assign y17898 = n28868 ;
  assign y17899 = ~n28875 ;
  assign y17900 = n28876 ;
  assign y17901 = ~n28877 ;
  assign y17902 = ~1'b0 ;
  assign y17903 = ~1'b0 ;
  assign y17904 = ~n28878 ;
  assign y17905 = ~1'b0 ;
  assign y17906 = ~n28882 ;
  assign y17907 = n13896 ;
  assign y17908 = ~n28884 ;
  assign y17909 = n28885 ;
  assign y17910 = ~1'b0 ;
  assign y17911 = 1'b0 ;
  assign y17912 = ~1'b0 ;
  assign y17913 = n28891 ;
  assign y17914 = ~n28896 ;
  assign y17915 = ~1'b0 ;
  assign y17916 = ~1'b0 ;
  assign y17917 = n28897 ;
  assign y17918 = ~1'b0 ;
  assign y17919 = n28899 ;
  assign y17920 = ~1'b0 ;
  assign y17921 = ~n28900 ;
  assign y17922 = ~n28904 ;
  assign y17923 = n28907 ;
  assign y17924 = n28909 ;
  assign y17925 = ~1'b0 ;
  assign y17926 = 1'b0 ;
  assign y17927 = n28911 ;
  assign y17928 = ~1'b0 ;
  assign y17929 = ~n28912 ;
  assign y17930 = ~n13139 ;
  assign y17931 = n28913 ;
  assign y17932 = ~n28914 ;
  assign y17933 = ~n28916 ;
  assign y17934 = ~1'b0 ;
  assign y17935 = n4899 ;
  assign y17936 = n28917 ;
  assign y17937 = n28918 ;
  assign y17938 = ~n19595 ;
  assign y17939 = ~1'b0 ;
  assign y17940 = n28919 ;
  assign y17941 = n15417 ;
  assign y17942 = ~n28923 ;
  assign y17943 = n28927 ;
  assign y17944 = ~n28930 ;
  assign y17945 = ~1'b0 ;
  assign y17946 = n28932 ;
  assign y17947 = n28933 ;
  assign y17948 = n28935 ;
  assign y17949 = n28938 ;
  assign y17950 = ~n28940 ;
  assign y17951 = ~n28942 ;
  assign y17952 = n28943 ;
  assign y17953 = ~n4701 ;
  assign y17954 = n28944 ;
  assign y17955 = 1'b0 ;
  assign y17956 = ~1'b0 ;
  assign y17957 = ~n7524 ;
  assign y17958 = ~n28947 ;
  assign y17959 = n28951 ;
  assign y17960 = n28952 ;
  assign y17961 = 1'b0 ;
  assign y17962 = ~n20676 ;
  assign y17963 = ~n28955 ;
  assign y17964 = ~n28958 ;
  assign y17965 = 1'b0 ;
  assign y17966 = n11308 ;
  assign y17967 = n28961 ;
  assign y17968 = n28965 ;
  assign y17969 = ~n28967 ;
  assign y17970 = n28968 ;
  assign y17971 = n28984 ;
  assign y17972 = ~1'b0 ;
  assign y17973 = ~n28987 ;
  assign y17974 = ~1'b0 ;
  assign y17975 = ~n28989 ;
  assign y17976 = ~n28992 ;
  assign y17977 = n28998 ;
  assign y17978 = n29001 ;
  assign y17979 = ~n29005 ;
  assign y17980 = ~n29007 ;
  assign y17981 = ~n12839 ;
  assign y17982 = n29008 ;
  assign y17983 = ~1'b0 ;
  assign y17984 = ~1'b0 ;
  assign y17985 = ~n29009 ;
  assign y17986 = ~n29011 ;
  assign y17987 = n29015 ;
  assign y17988 = ~n29018 ;
  assign y17989 = ~1'b0 ;
  assign y17990 = n29019 ;
  assign y17991 = ~n29021 ;
  assign y17992 = ~n29024 ;
  assign y17993 = n29026 ;
  assign y17994 = ~n29030 ;
  assign y17995 = ~n29035 ;
  assign y17996 = n29036 ;
  assign y17997 = ~n29040 ;
  assign y17998 = ~1'b0 ;
  assign y17999 = ~1'b0 ;
  assign y18000 = ~n29041 ;
  assign y18001 = ~1'b0 ;
  assign y18002 = ~n29046 ;
  assign y18003 = ~n29048 ;
  assign y18004 = ~1'b0 ;
  assign y18005 = ~n29049 ;
  assign y18006 = ~1'b0 ;
  assign y18007 = ~1'b0 ;
  assign y18008 = ~1'b0 ;
  assign y18009 = n29050 ;
  assign y18010 = ~1'b0 ;
  assign y18011 = ~1'b0 ;
  assign y18012 = n29052 ;
  assign y18013 = ~n27370 ;
  assign y18014 = n29053 ;
  assign y18015 = ~n29055 ;
  assign y18016 = ~n29057 ;
  assign y18017 = ~n26252 ;
  assign y18018 = n29058 ;
  assign y18019 = ~1'b0 ;
  assign y18020 = ~n29059 ;
  assign y18021 = ~n29060 ;
  assign y18022 = ~n29068 ;
  assign y18023 = ~n7829 ;
  assign y18024 = 1'b0 ;
  assign y18025 = ~n29069 ;
  assign y18026 = ~1'b0 ;
  assign y18027 = ~n2807 ;
  assign y18028 = n29071 ;
  assign y18029 = ~1'b0 ;
  assign y18030 = ~1'b0 ;
  assign y18031 = n26737 ;
  assign y18032 = n29072 ;
  assign y18033 = ~n29073 ;
  assign y18034 = n18047 ;
  assign y18035 = n6184 ;
  assign y18036 = ~1'b0 ;
  assign y18037 = ~1'b0 ;
  assign y18038 = n29074 ;
  assign y18039 = ~1'b0 ;
  assign y18040 = ~1'b0 ;
  assign y18041 = ~n27638 ;
  assign y18042 = ~n29080 ;
  assign y18043 = ~1'b0 ;
  assign y18044 = n29082 ;
  assign y18045 = n29083 ;
  assign y18046 = ~n12467 ;
  assign y18047 = ~1'b0 ;
  assign y18048 = ~1'b0 ;
  assign y18049 = n29089 ;
  assign y18050 = ~n29091 ;
  assign y18051 = n29092 ;
  assign y18052 = ~1'b0 ;
  assign y18053 = ~n29094 ;
  assign y18054 = n29097 ;
  assign y18055 = n29101 ;
  assign y18056 = n29104 ;
  assign y18057 = n29105 ;
  assign y18058 = ~n29106 ;
  assign y18059 = 1'b0 ;
  assign y18060 = n29109 ;
  assign y18061 = ~n29113 ;
  assign y18062 = ~1'b0 ;
  assign y18063 = n29115 ;
  assign y18064 = ~1'b0 ;
  assign y18065 = ~n29118 ;
  assign y18066 = ~n29119 ;
  assign y18067 = n29122 ;
  assign y18068 = ~1'b0 ;
  assign y18069 = ~n29128 ;
  assign y18070 = ~1'b0 ;
  assign y18071 = ~n29129 ;
  assign y18072 = ~n29131 ;
  assign y18073 = n29134 ;
  assign y18074 = ~1'b0 ;
  assign y18075 = ~n29137 ;
  assign y18076 = ~1'b0 ;
  assign y18077 = ~n29138 ;
  assign y18078 = ~1'b0 ;
  assign y18079 = 1'b0 ;
  assign y18080 = n833 ;
  assign y18081 = ~1'b0 ;
  assign y18082 = ~1'b0 ;
  assign y18083 = ~1'b0 ;
  assign y18084 = ~1'b0 ;
  assign y18085 = ~1'b0 ;
  assign y18086 = ~1'b0 ;
  assign y18087 = n29139 ;
  assign y18088 = n7100 ;
  assign y18089 = n29140 ;
  assign y18090 = ~n22449 ;
  assign y18091 = ~n29142 ;
  assign y18092 = ~n29146 ;
  assign y18093 = n29148 ;
  assign y18094 = n29152 ;
  assign y18095 = ~1'b0 ;
  assign y18096 = n6608 ;
  assign y18097 = ~n29160 ;
  assign y18098 = ~1'b0 ;
  assign y18099 = 1'b0 ;
  assign y18100 = n2296 ;
  assign y18101 = ~1'b0 ;
  assign y18102 = n29165 ;
  assign y18103 = ~1'b0 ;
  assign y18104 = ~n29175 ;
  assign y18105 = ~1'b0 ;
  assign y18106 = ~1'b0 ;
  assign y18107 = ~1'b0 ;
  assign y18108 = n3329 ;
  assign y18109 = ~n29181 ;
  assign y18110 = ~1'b0 ;
  assign y18111 = n29183 ;
  assign y18112 = n29185 ;
  assign y18113 = ~1'b0 ;
  assign y18114 = n29188 ;
  assign y18115 = ~1'b0 ;
  assign y18116 = ~1'b0 ;
  assign y18117 = n23308 ;
  assign y18118 = n29190 ;
  assign y18119 = ~1'b0 ;
  assign y18120 = n29194 ;
  assign y18121 = n29195 ;
  assign y18122 = 1'b0 ;
  assign y18123 = ~1'b0 ;
  assign y18124 = ~1'b0 ;
  assign y18125 = ~n29200 ;
  assign y18126 = ~n29201 ;
  assign y18127 = n7940 ;
  assign y18128 = ~1'b0 ;
  assign y18129 = ~1'b0 ;
  assign y18130 = ~1'b0 ;
  assign y18131 = ~1'b0 ;
  assign y18132 = ~1'b0 ;
  assign y18133 = ~1'b0 ;
  assign y18134 = ~n29202 ;
  assign y18135 = ~1'b0 ;
  assign y18136 = ~1'b0 ;
  assign y18137 = n6253 ;
  assign y18138 = ~1'b0 ;
  assign y18139 = ~1'b0 ;
  assign y18140 = n10364 ;
  assign y18141 = n29206 ;
  assign y18142 = ~1'b0 ;
  assign y18143 = ~1'b0 ;
  assign y18144 = ~n29211 ;
  assign y18145 = n29216 ;
  assign y18146 = ~n7367 ;
  assign y18147 = ~1'b0 ;
  assign y18148 = n29218 ;
  assign y18149 = ~1'b0 ;
  assign y18150 = ~1'b0 ;
  assign y18151 = ~1'b0 ;
  assign y18152 = ~n27585 ;
  assign y18153 = ~n29220 ;
  assign y18154 = n29221 ;
  assign y18155 = ~1'b0 ;
  assign y18156 = ~n29225 ;
  assign y18157 = ~n29227 ;
  assign y18158 = ~1'b0 ;
  assign y18159 = ~1'b0 ;
  assign y18160 = n29230 ;
  assign y18161 = ~n29231 ;
  assign y18162 = n29234 ;
  assign y18163 = n29236 ;
  assign y18164 = n29239 ;
  assign y18165 = ~n29241 ;
  assign y18166 = n29245 ;
  assign y18167 = n29249 ;
  assign y18168 = n28057 ;
  assign y18169 = ~n29254 ;
  assign y18170 = n5190 ;
  assign y18171 = ~1'b0 ;
  assign y18172 = ~1'b0 ;
  assign y18173 = n14641 ;
  assign y18174 = ~n29256 ;
  assign y18175 = ~1'b0 ;
  assign y18176 = ~n29258 ;
  assign y18177 = ~1'b0 ;
  assign y18178 = n29260 ;
  assign y18179 = ~n29261 ;
  assign y18180 = n29265 ;
  assign y18181 = ~1'b0 ;
  assign y18182 = ~1'b0 ;
  assign y18183 = ~n29267 ;
  assign y18184 = ~1'b0 ;
  assign y18185 = ~1'b0 ;
  assign y18186 = ~1'b0 ;
  assign y18187 = n28790 ;
  assign y18188 = ~n29269 ;
  assign y18189 = ~1'b0 ;
  assign y18190 = n29271 ;
  assign y18191 = ~n29275 ;
  assign y18192 = ~n29277 ;
  assign y18193 = ~n29279 ;
  assign y18194 = ~n29282 ;
  assign y18195 = ~n29283 ;
  assign y18196 = ~1'b0 ;
  assign y18197 = n29284 ;
  assign y18198 = ~n29286 ;
  assign y18199 = ~1'b0 ;
  assign y18200 = ~1'b0 ;
  assign y18201 = n29291 ;
  assign y18202 = n29294 ;
  assign y18203 = n29297 ;
  assign y18204 = ~n26072 ;
  assign y18205 = ~n18028 ;
  assign y18206 = ~n29299 ;
  assign y18207 = ~1'b0 ;
  assign y18208 = ~n29301 ;
  assign y18209 = ~n29303 ;
  assign y18210 = ~n29304 ;
  assign y18211 = ~1'b0 ;
  assign y18212 = n29307 ;
  assign y18213 = ~n29308 ;
  assign y18214 = n29312 ;
  assign y18215 = n29314 ;
  assign y18216 = n29315 ;
  assign y18217 = n29316 ;
  assign y18218 = ~1'b0 ;
  assign y18219 = n29319 ;
  assign y18220 = n29320 ;
  assign y18221 = ~n29322 ;
  assign y18222 = n29323 ;
  assign y18223 = n29327 ;
  assign y18224 = 1'b0 ;
  assign y18225 = ~n29328 ;
  assign y18226 = n29329 ;
  assign y18227 = ~n7895 ;
  assign y18228 = ~n29333 ;
  assign y18229 = ~1'b0 ;
  assign y18230 = ~n29334 ;
  assign y18231 = n1634 ;
  assign y18232 = n29335 ;
  assign y18233 = ~n29337 ;
  assign y18234 = ~n1680 ;
  assign y18235 = ~1'b0 ;
  assign y18236 = ~n29338 ;
  assign y18237 = ~n6779 ;
  assign y18238 = ~1'b0 ;
  assign y18239 = n29340 ;
  assign y18240 = ~n29341 ;
  assign y18241 = ~n29347 ;
  assign y18242 = ~n24337 ;
  assign y18243 = ~n29348 ;
  assign y18244 = n29349 ;
  assign y18245 = n29350 ;
  assign y18246 = ~1'b0 ;
  assign y18247 = n29353 ;
  assign y18248 = n29354 ;
  assign y18249 = 1'b0 ;
  assign y18250 = ~n29355 ;
  assign y18251 = ~n29359 ;
  assign y18252 = ~n29361 ;
  assign y18253 = ~n29363 ;
  assign y18254 = ~n10488 ;
  assign y18255 = ~1'b0 ;
  assign y18256 = ~n9287 ;
  assign y18257 = n29365 ;
  assign y18258 = ~n29368 ;
  assign y18259 = n29370 ;
  assign y18260 = ~1'b0 ;
  assign y18261 = ~1'b0 ;
  assign y18262 = n29371 ;
  assign y18263 = ~1'b0 ;
  assign y18264 = n29372 ;
  assign y18265 = ~1'b0 ;
  assign y18266 = ~1'b0 ;
  assign y18267 = ~1'b0 ;
  assign y18268 = ~n29373 ;
  assign y18269 = ~1'b0 ;
  assign y18270 = n5918 ;
  assign y18271 = n29375 ;
  assign y18272 = ~n29377 ;
  assign y18273 = ~n29379 ;
  assign y18274 = n29380 ;
  assign y18275 = ~n3462 ;
  assign y18276 = n6576 ;
  assign y18277 = ~n29381 ;
  assign y18278 = n29382 ;
  assign y18279 = ~1'b0 ;
  assign y18280 = ~1'b0 ;
  assign y18281 = ~1'b0 ;
  assign y18282 = ~1'b0 ;
  assign y18283 = n29385 ;
  assign y18284 = ~n29388 ;
  assign y18285 = ~n29389 ;
  assign y18286 = ~n29393 ;
  assign y18287 = ~1'b0 ;
  assign y18288 = ~n29395 ;
  assign y18289 = ~n29402 ;
  assign y18290 = ~n29407 ;
  assign y18291 = ~n29410 ;
  assign y18292 = ~n29413 ;
  assign y18293 = ~n29416 ;
  assign y18294 = ~n29419 ;
  assign y18295 = n29420 ;
  assign y18296 = ~1'b0 ;
  assign y18297 = ~n29424 ;
  assign y18298 = ~n29426 ;
  assign y18299 = n29429 ;
  assign y18300 = n29432 ;
  assign y18301 = n29434 ;
  assign y18302 = ~1'b0 ;
  assign y18303 = n29436 ;
  assign y18304 = ~1'b0 ;
  assign y18305 = ~n29439 ;
  assign y18306 = n29440 ;
  assign y18307 = ~n29441 ;
  assign y18308 = ~n29443 ;
  assign y18309 = n29444 ;
  assign y18310 = ~n29445 ;
  assign y18311 = n29447 ;
  assign y18312 = n29448 ;
  assign y18313 = ~1'b0 ;
  assign y18314 = n29450 ;
  assign y18315 = n29452 ;
  assign y18316 = n29453 ;
  assign y18317 = n15334 ;
  assign y18318 = n29456 ;
  assign y18319 = n29457 ;
  assign y18320 = ~n14452 ;
  assign y18321 = ~1'b0 ;
  assign y18322 = ~n29460 ;
  assign y18323 = ~1'b0 ;
  assign y18324 = ~1'b0 ;
  assign y18325 = ~n29461 ;
  assign y18326 = ~1'b0 ;
  assign y18327 = ~1'b0 ;
  assign y18328 = n29463 ;
  assign y18329 = n29464 ;
  assign y18330 = n29465 ;
  assign y18331 = ~1'b0 ;
  assign y18332 = ~n29468 ;
  assign y18333 = ~1'b0 ;
  assign y18334 = ~1'b0 ;
  assign y18335 = 1'b0 ;
  assign y18336 = n29469 ;
  assign y18337 = ~1'b0 ;
  assign y18338 = ~1'b0 ;
  assign y18339 = ~n6801 ;
  assign y18340 = 1'b0 ;
  assign y18341 = ~1'b0 ;
  assign y18342 = ~1'b0 ;
  assign y18343 = ~n7571 ;
  assign y18344 = ~n29471 ;
  assign y18345 = n29474 ;
  assign y18346 = ~n29475 ;
  assign y18347 = n29476 ;
  assign y18348 = ~1'b0 ;
  assign y18349 = n29479 ;
  assign y18350 = n29480 ;
  assign y18351 = n20438 ;
  assign y18352 = ~1'b0 ;
  assign y18353 = ~n29483 ;
  assign y18354 = ~1'b0 ;
  assign y18355 = n29485 ;
  assign y18356 = ~n29486 ;
  assign y18357 = n29487 ;
  assign y18358 = n29488 ;
  assign y18359 = n29489 ;
  assign y18360 = 1'b0 ;
  assign y18361 = ~n29490 ;
  assign y18362 = ~n29491 ;
  assign y18363 = ~1'b0 ;
  assign y18364 = n3533 ;
  assign y18365 = ~1'b0 ;
  assign y18366 = ~1'b0 ;
  assign y18367 = ~n29493 ;
  assign y18368 = ~n29494 ;
  assign y18369 = n11720 ;
  assign y18370 = ~1'b0 ;
  assign y18371 = n9654 ;
  assign y18372 = n29495 ;
  assign y18373 = ~1'b0 ;
  assign y18374 = ~1'b0 ;
  assign y18375 = ~n29497 ;
  assign y18376 = ~n13261 ;
  assign y18377 = ~n29503 ;
  assign y18378 = n29505 ;
  assign y18379 = n29508 ;
  assign y18380 = n29510 ;
  assign y18381 = ~1'b0 ;
  assign y18382 = n29512 ;
  assign y18383 = ~n532 ;
  assign y18384 = n29520 ;
  assign y18385 = n29522 ;
  assign y18386 = ~n29524 ;
  assign y18387 = n6025 ;
  assign y18388 = ~1'b0 ;
  assign y18389 = ~1'b0 ;
  assign y18390 = ~n29527 ;
  assign y18391 = n29529 ;
  assign y18392 = ~1'b0 ;
  assign y18393 = ~1'b0 ;
  assign y18394 = ~n29530 ;
  assign y18395 = ~1'b0 ;
  assign y18396 = n29531 ;
  assign y18397 = ~n29533 ;
  assign y18398 = n29536 ;
  assign y18399 = ~1'b0 ;
  assign y18400 = ~n29537 ;
  assign y18401 = ~1'b0 ;
  assign y18402 = ~n29538 ;
  assign y18403 = 1'b0 ;
  assign y18404 = ~1'b0 ;
  assign y18405 = n29539 ;
  assign y18406 = ~1'b0 ;
  assign y18407 = 1'b0 ;
  assign y18408 = n29540 ;
  assign y18409 = ~n29541 ;
  assign y18410 = ~n29546 ;
  assign y18411 = ~1'b0 ;
  assign y18412 = ~n29547 ;
  assign y18413 = ~1'b0 ;
  assign y18414 = ~1'b0 ;
  assign y18415 = ~1'b0 ;
  assign y18416 = ~1'b0 ;
  assign y18417 = n29551 ;
  assign y18418 = ~n29552 ;
  assign y18419 = ~1'b0 ;
  assign y18420 = ~1'b0 ;
  assign y18421 = n29553 ;
  assign y18422 = ~n29554 ;
  assign y18423 = ~n29558 ;
  assign y18424 = n29559 ;
  assign y18425 = ~1'b0 ;
  assign y18426 = n29564 ;
  assign y18427 = ~n29565 ;
  assign y18428 = ~n29567 ;
  assign y18429 = ~n29568 ;
  assign y18430 = ~1'b0 ;
  assign y18431 = ~n29570 ;
  assign y18432 = ~n29574 ;
  assign y18433 = ~n29576 ;
  assign y18434 = ~n29578 ;
  assign y18435 = ~n29581 ;
  assign y18436 = n29586 ;
  assign y18437 = ~1'b0 ;
  assign y18438 = n29587 ;
  assign y18439 = ~n29589 ;
  assign y18440 = ~n29595 ;
  assign y18441 = n25118 ;
  assign y18442 = ~n29597 ;
  assign y18443 = n29599 ;
  assign y18444 = ~n29600 ;
  assign y18445 = ~1'b0 ;
  assign y18446 = ~n29602 ;
  assign y18447 = ~1'b0 ;
  assign y18448 = ~1'b0 ;
  assign y18449 = ~n29604 ;
  assign y18450 = ~n29606 ;
  assign y18451 = n29607 ;
  assign y18452 = ~1'b0 ;
  assign y18453 = ~1'b0 ;
  assign y18454 = n29612 ;
  assign y18455 = ~n29621 ;
  assign y18456 = 1'b0 ;
  assign y18457 = ~1'b0 ;
  assign y18458 = ~n29624 ;
  assign y18459 = n29627 ;
  assign y18460 = ~1'b0 ;
  assign y18461 = ~n29630 ;
  assign y18462 = ~n29632 ;
  assign y18463 = ~n29636 ;
  assign y18464 = n29637 ;
  assign y18465 = ~n14442 ;
  assign y18466 = ~n29460 ;
  assign y18467 = ~1'b0 ;
  assign y18468 = ~1'b0 ;
  assign y18469 = n29640 ;
  assign y18470 = ~n29647 ;
  assign y18471 = n29651 ;
  assign y18472 = n12018 ;
  assign y18473 = ~1'b0 ;
  assign y18474 = n29655 ;
  assign y18475 = ~n29657 ;
  assign y18476 = ~1'b0 ;
  assign y18477 = ~1'b0 ;
  assign y18478 = ~n17009 ;
  assign y18479 = ~n29658 ;
  assign y18480 = n29661 ;
  assign y18481 = ~n29665 ;
  assign y18482 = ~1'b0 ;
  assign y18483 = ~n29670 ;
  assign y18484 = ~n29671 ;
  assign y18485 = n29675 ;
  assign y18486 = ~n29682 ;
  assign y18487 = ~n29684 ;
  assign y18488 = ~n29687 ;
  assign y18489 = n29688 ;
  assign y18490 = ~1'b0 ;
  assign y18491 = ~1'b0 ;
  assign y18492 = ~1'b0 ;
  assign y18493 = 1'b0 ;
  assign y18494 = ~1'b0 ;
  assign y18495 = ~1'b0 ;
  assign y18496 = ~n29689 ;
  assign y18497 = n29690 ;
  assign y18498 = n29692 ;
  assign y18499 = ~1'b0 ;
  assign y18500 = n29697 ;
  assign y18501 = n29701 ;
  assign y18502 = n29702 ;
  assign y18503 = n29707 ;
  assign y18504 = ~1'b0 ;
  assign y18505 = n29712 ;
  assign y18506 = ~n29713 ;
  assign y18507 = n13438 ;
  assign y18508 = ~n29715 ;
  assign y18509 = ~1'b0 ;
  assign y18510 = ~n29716 ;
  assign y18511 = ~1'b0 ;
  assign y18512 = n29719 ;
  assign y18513 = n29721 ;
  assign y18514 = ~1'b0 ;
  assign y18515 = 1'b0 ;
  assign y18516 = ~n29732 ;
  assign y18517 = n29740 ;
  assign y18518 = n6193 ;
  assign y18519 = ~n29741 ;
  assign y18520 = n29743 ;
  assign y18521 = ~n29744 ;
  assign y18522 = ~1'b0 ;
  assign y18523 = n29745 ;
  assign y18524 = ~1'b0 ;
  assign y18525 = ~1'b0 ;
  assign y18526 = ~n4592 ;
  assign y18527 = n3858 ;
  assign y18528 = ~n29747 ;
  assign y18529 = ~1'b0 ;
  assign y18530 = ~1'b0 ;
  assign y18531 = n27943 ;
  assign y18532 = n29750 ;
  assign y18533 = ~1'b0 ;
  assign y18534 = ~n29751 ;
  assign y18535 = n29754 ;
  assign y18536 = n29755 ;
  assign y18537 = ~1'b0 ;
  assign y18538 = ~n29756 ;
  assign y18539 = ~1'b0 ;
  assign y18540 = n29757 ;
  assign y18541 = n29759 ;
  assign y18542 = n29762 ;
  assign y18543 = ~n29763 ;
  assign y18544 = ~1'b0 ;
  assign y18545 = ~1'b0 ;
  assign y18546 = n29768 ;
  assign y18547 = 1'b0 ;
  assign y18548 = n29770 ;
  assign y18549 = n29773 ;
  assign y18550 = ~n29774 ;
  assign y18551 = ~1'b0 ;
  assign y18552 = ~n29778 ;
  assign y18553 = n10195 ;
  assign y18554 = 1'b0 ;
  assign y18555 = ~1'b0 ;
  assign y18556 = ~n8837 ;
  assign y18557 = 1'b0 ;
  assign y18558 = ~n29780 ;
  assign y18559 = ~1'b0 ;
  assign y18560 = n29784 ;
  assign y18561 = ~n29786 ;
  assign y18562 = ~n28402 ;
  assign y18563 = ~n29787 ;
  assign y18564 = ~n29788 ;
  assign y18565 = ~n29790 ;
  assign y18566 = ~1'b0 ;
  assign y18567 = n29794 ;
  assign y18568 = n29796 ;
  assign y18569 = ~1'b0 ;
  assign y18570 = n29799 ;
  assign y18571 = ~n6934 ;
  assign y18572 = ~n29806 ;
  assign y18573 = ~n29807 ;
  assign y18574 = ~1'b0 ;
  assign y18575 = ~n29808 ;
  assign y18576 = ~1'b0 ;
  assign y18577 = ~1'b0 ;
  assign y18578 = ~n29811 ;
  assign y18579 = ~1'b0 ;
  assign y18580 = ~1'b0 ;
  assign y18581 = ~n29812 ;
  assign y18582 = ~n29814 ;
  assign y18583 = ~n3566 ;
  assign y18584 = ~1'b0 ;
  assign y18585 = ~1'b0 ;
  assign y18586 = n29817 ;
  assign y18587 = 1'b0 ;
  assign y18588 = ~n29818 ;
  assign y18589 = ~n29820 ;
  assign y18590 = n29824 ;
  assign y18591 = ~1'b0 ;
  assign y18592 = ~n29825 ;
  assign y18593 = ~1'b0 ;
  assign y18594 = ~1'b0 ;
  assign y18595 = ~1'b0 ;
  assign y18596 = ~1'b0 ;
  assign y18597 = n29829 ;
  assign y18598 = ~n29833 ;
  assign y18599 = ~n29835 ;
  assign y18600 = ~1'b0 ;
  assign y18601 = ~n29838 ;
  assign y18602 = n29839 ;
  assign y18603 = ~1'b0 ;
  assign y18604 = ~n4727 ;
  assign y18605 = n29840 ;
  assign y18606 = n3499 ;
  assign y18607 = ~1'b0 ;
  assign y18608 = ~1'b0 ;
  assign y18609 = n21852 ;
  assign y18610 = ~n29841 ;
  assign y18611 = ~1'b0 ;
  assign y18612 = n29842 ;
  assign y18613 = ~1'b0 ;
  assign y18614 = n29843 ;
  assign y18615 = n29845 ;
  assign y18616 = n29847 ;
  assign y18617 = ~1'b0 ;
  assign y18618 = ~1'b0 ;
  assign y18619 = n29848 ;
  assign y18620 = 1'b0 ;
  assign y18621 = ~n29849 ;
  assign y18622 = ~1'b0 ;
  assign y18623 = ~1'b0 ;
  assign y18624 = n29852 ;
  assign y18625 = ~1'b0 ;
  assign y18626 = n29854 ;
  assign y18627 = n2750 ;
  assign y18628 = n29857 ;
  assign y18629 = ~n29859 ;
  assign y18630 = n19800 ;
  assign y18631 = ~n29874 ;
  assign y18632 = ~1'b0 ;
  assign y18633 = ~n4505 ;
  assign y18634 = ~1'b0 ;
  assign y18635 = n29875 ;
  assign y18636 = ~n29877 ;
  assign y18637 = ~n29879 ;
  assign y18638 = ~n17969 ;
  assign y18639 = ~n29881 ;
  assign y18640 = ~1'b0 ;
  assign y18641 = ~n29883 ;
  assign y18642 = n29884 ;
  assign y18643 = ~n10329 ;
  assign y18644 = ~n29886 ;
  assign y18645 = ~n12227 ;
  assign y18646 = n29887 ;
  assign y18647 = ~1'b0 ;
  assign y18648 = ~1'b0 ;
  assign y18649 = ~1'b0 ;
  assign y18650 = n29888 ;
  assign y18651 = n1278 ;
  assign y18652 = ~1'b0 ;
  assign y18653 = ~1'b0 ;
  assign y18654 = n17505 ;
  assign y18655 = n29889 ;
  assign y18656 = ~1'b0 ;
  assign y18657 = ~1'b0 ;
  assign y18658 = ~1'b0 ;
  assign y18659 = ~n29890 ;
  assign y18660 = ~n29893 ;
  assign y18661 = ~1'b0 ;
  assign y18662 = ~n29895 ;
  assign y18663 = ~1'b0 ;
  assign y18664 = ~1'b0 ;
  assign y18665 = n29897 ;
  assign y18666 = n29900 ;
  assign y18667 = ~1'b0 ;
  assign y18668 = ~n29901 ;
  assign y18669 = ~1'b0 ;
  assign y18670 = ~1'b0 ;
  assign y18671 = ~1'b0 ;
  assign y18672 = ~n29903 ;
  assign y18673 = ~n29908 ;
  assign y18674 = ~1'b0 ;
  assign y18675 = ~n29910 ;
  assign y18676 = ~n29913 ;
  assign y18677 = 1'b0 ;
  assign y18678 = 1'b0 ;
  assign y18679 = n29916 ;
  assign y18680 = ~n29918 ;
  assign y18681 = ~n29919 ;
  assign y18682 = ~n29920 ;
  assign y18683 = n29921 ;
  assign y18684 = ~1'b0 ;
  assign y18685 = ~n29923 ;
  assign y18686 = n29924 ;
  assign y18687 = ~1'b0 ;
  assign y18688 = n29925 ;
  assign y18689 = ~n29928 ;
  assign y18690 = ~n18581 ;
  assign y18691 = ~1'b0 ;
  assign y18692 = ~1'b0 ;
  assign y18693 = n11456 ;
  assign y18694 = ~1'b0 ;
  assign y18695 = n29929 ;
  assign y18696 = ~n29932 ;
  assign y18697 = n29934 ;
  assign y18698 = ~1'b0 ;
  assign y18699 = n29940 ;
  assign y18700 = n29941 ;
  assign y18701 = ~1'b0 ;
  assign y18702 = ~n29942 ;
  assign y18703 = ~1'b0 ;
  assign y18704 = 1'b0 ;
  assign y18705 = ~1'b0 ;
  assign y18706 = ~1'b0 ;
  assign y18707 = ~n29946 ;
  assign y18708 = ~1'b0 ;
  assign y18709 = ~n29948 ;
  assign y18710 = 1'b0 ;
  assign y18711 = 1'b0 ;
  assign y18712 = ~n29949 ;
  assign y18713 = ~n29950 ;
  assign y18714 = ~n29953 ;
  assign y18715 = ~n10575 ;
  assign y18716 = ~1'b0 ;
  assign y18717 = n29955 ;
  assign y18718 = ~n29956 ;
  assign y18719 = 1'b0 ;
  assign y18720 = ~1'b0 ;
  assign y18721 = ~n29966 ;
  assign y18722 = n1487 ;
  assign y18723 = ~n29968 ;
  assign y18724 = ~1'b0 ;
  assign y18725 = ~n15380 ;
  assign y18726 = ~n29972 ;
  assign y18727 = ~n29978 ;
  assign y18728 = ~1'b0 ;
  assign y18729 = n29981 ;
  assign y18730 = ~1'b0 ;
  assign y18731 = n29982 ;
  assign y18732 = ~n29987 ;
  assign y18733 = ~1'b0 ;
  assign y18734 = ~n29988 ;
  assign y18735 = ~n27341 ;
  assign y18736 = ~n29992 ;
  assign y18737 = n29993 ;
  assign y18738 = n700 ;
  assign y18739 = ~1'b0 ;
  assign y18740 = ~1'b0 ;
  assign y18741 = ~n29994 ;
  assign y18742 = ~n29995 ;
  assign y18743 = ~1'b0 ;
  assign y18744 = ~n29998 ;
  assign y18745 = ~n30000 ;
  assign y18746 = ~1'b0 ;
  assign y18747 = ~n30002 ;
  assign y18748 = ~1'b0 ;
  assign y18749 = ~n30003 ;
  assign y18750 = ~n30005 ;
  assign y18751 = ~1'b0 ;
  assign y18752 = ~1'b0 ;
  assign y18753 = ~1'b0 ;
  assign y18754 = ~1'b0 ;
  assign y18755 = ~1'b0 ;
  assign y18756 = n30006 ;
  assign y18757 = ~1'b0 ;
  assign y18758 = n30009 ;
  assign y18759 = ~n30017 ;
  assign y18760 = ~1'b0 ;
  assign y18761 = ~n30018 ;
  assign y18762 = ~n30022 ;
  assign y18763 = ~n30024 ;
  assign y18764 = ~1'b0 ;
  assign y18765 = n30026 ;
  assign y18766 = ~n30028 ;
  assign y18767 = n30029 ;
  assign y18768 = n30030 ;
  assign y18769 = ~1'b0 ;
  assign y18770 = ~1'b0 ;
  assign y18771 = n30031 ;
  assign y18772 = ~n3549 ;
  assign y18773 = ~n30033 ;
  assign y18774 = ~1'b0 ;
  assign y18775 = n23519 ;
  assign y18776 = n6034 ;
  assign y18777 = ~n30035 ;
  assign y18778 = n28584 ;
  assign y18779 = 1'b0 ;
  assign y18780 = ~1'b0 ;
  assign y18781 = ~1'b0 ;
  assign y18782 = n361 ;
  assign y18783 = ~1'b0 ;
  assign y18784 = n16628 ;
  assign y18785 = 1'b0 ;
  assign y18786 = n30038 ;
  assign y18787 = ~1'b0 ;
  assign y18788 = ~n30040 ;
  assign y18789 = n30043 ;
  assign y18790 = ~n30046 ;
  assign y18791 = ~n30048 ;
  assign y18792 = ~1'b0 ;
  assign y18793 = ~n30050 ;
  assign y18794 = n30052 ;
  assign y18795 = 1'b0 ;
  assign y18796 = ~1'b0 ;
  assign y18797 = ~1'b0 ;
  assign y18798 = n30053 ;
  assign y18799 = ~1'b0 ;
  assign y18800 = ~n30055 ;
  assign y18801 = ~1'b0 ;
  assign y18802 = ~n30056 ;
  assign y18803 = n30060 ;
  assign y18804 = ~n30061 ;
  assign y18805 = n30062 ;
  assign y18806 = ~n30064 ;
  assign y18807 = n30066 ;
  assign y18808 = 1'b0 ;
  assign y18809 = ~1'b0 ;
  assign y18810 = ~1'b0 ;
  assign y18811 = n11226 ;
  assign y18812 = 1'b0 ;
  assign y18813 = ~1'b0 ;
  assign y18814 = ~1'b0 ;
  assign y18815 = ~1'b0 ;
  assign y18816 = n2099 ;
  assign y18817 = ~1'b0 ;
  assign y18818 = n30068 ;
  assign y18819 = ~n30069 ;
  assign y18820 = ~1'b0 ;
  assign y18821 = ~n20435 ;
  assign y18822 = ~n10018 ;
  assign y18823 = n30070 ;
  assign y18824 = ~1'b0 ;
  assign y18825 = ~n30073 ;
  assign y18826 = ~1'b0 ;
  assign y18827 = ~1'b0 ;
  assign y18828 = ~1'b0 ;
  assign y18829 = ~1'b0 ;
  assign y18830 = ~1'b0 ;
  assign y18831 = ~1'b0 ;
  assign y18832 = ~n30074 ;
  assign y18833 = ~1'b0 ;
  assign y18834 = ~1'b0 ;
  assign y18835 = n30075 ;
  assign y18836 = ~n30080 ;
  assign y18837 = n30081 ;
  assign y18838 = n30082 ;
  assign y18839 = n30085 ;
  assign y18840 = ~1'b0 ;
  assign y18841 = ~n30087 ;
  assign y18842 = n30088 ;
  assign y18843 = ~1'b0 ;
  assign y18844 = n30089 ;
  assign y18845 = 1'b0 ;
  assign y18846 = ~n25107 ;
  assign y18847 = n30092 ;
  assign y18848 = ~1'b0 ;
  assign y18849 = n30093 ;
  assign y18850 = ~1'b0 ;
  assign y18851 = n30099 ;
  assign y18852 = n4326 ;
  assign y18853 = n5067 ;
  assign y18854 = ~1'b0 ;
  assign y18855 = ~1'b0 ;
  assign y18856 = ~n30103 ;
  assign y18857 = ~1'b0 ;
  assign y18858 = ~n30105 ;
  assign y18859 = n30107 ;
  assign y18860 = ~n30110 ;
  assign y18861 = ~n30112 ;
  assign y18862 = ~1'b0 ;
  assign y18863 = ~1'b0 ;
  assign y18864 = n30115 ;
  assign y18865 = n30116 ;
  assign y18866 = ~1'b0 ;
  assign y18867 = n30118 ;
  assign y18868 = ~1'b0 ;
  assign y18869 = ~1'b0 ;
  assign y18870 = n30119 ;
  assign y18871 = ~n30127 ;
  assign y18872 = n30128 ;
  assign y18873 = ~1'b0 ;
  assign y18874 = ~n30129 ;
  assign y18875 = ~1'b0 ;
  assign y18876 = n7305 ;
  assign y18877 = ~1'b0 ;
  assign y18878 = ~n30130 ;
  assign y18879 = ~1'b0 ;
  assign y18880 = ~n11164 ;
  assign y18881 = ~n30135 ;
  assign y18882 = ~1'b0 ;
  assign y18883 = ~n30136 ;
  assign y18884 = n30138 ;
  assign y18885 = ~n30156 ;
  assign y18886 = ~n30162 ;
  assign y18887 = ~n30164 ;
  assign y18888 = ~n30166 ;
  assign y18889 = ~n19924 ;
  assign y18890 = n30167 ;
  assign y18891 = ~1'b0 ;
  assign y18892 = n30169 ;
  assign y18893 = ~1'b0 ;
  assign y18894 = ~1'b0 ;
  assign y18895 = n30174 ;
  assign y18896 = ~n30175 ;
  assign y18897 = n30177 ;
  assign y18898 = ~1'b0 ;
  assign y18899 = ~n30179 ;
  assign y18900 = n30180 ;
  assign y18901 = ~1'b0 ;
  assign y18902 = n30181 ;
  assign y18903 = ~1'b0 ;
  assign y18904 = ~n30184 ;
  assign y18905 = ~1'b0 ;
  assign y18906 = n30187 ;
  assign y18907 = n30188 ;
  assign y18908 = ~1'b0 ;
  assign y18909 = ~n30191 ;
  assign y18910 = 1'b0 ;
  assign y18911 = n30192 ;
  assign y18912 = ~n30193 ;
  assign y18913 = ~n30194 ;
  assign y18914 = n30198 ;
  assign y18915 = n27869 ;
  assign y18916 = ~n30201 ;
  assign y18917 = ~1'b0 ;
  assign y18918 = n30204 ;
  assign y18919 = n30205 ;
  assign y18920 = n30207 ;
  assign y18921 = ~1'b0 ;
  assign y18922 = n30208 ;
  assign y18923 = ~1'b0 ;
  assign y18924 = ~1'b0 ;
  assign y18925 = ~1'b0 ;
  assign y18926 = ~n30209 ;
  assign y18927 = ~1'b0 ;
  assign y18928 = n30210 ;
  assign y18929 = ~n30212 ;
  assign y18930 = ~1'b0 ;
  assign y18931 = ~1'b0 ;
  assign y18932 = ~n30215 ;
  assign y18933 = ~n30219 ;
  assign y18934 = 1'b0 ;
  assign y18935 = ~n30224 ;
  assign y18936 = n30225 ;
  assign y18937 = ~n30229 ;
  assign y18938 = ~1'b0 ;
  assign y18939 = n7037 ;
  assign y18940 = ~n30230 ;
  assign y18941 = 1'b0 ;
  assign y18942 = ~n30232 ;
  assign y18943 = n30236 ;
  assign y18944 = ~1'b0 ;
  assign y18945 = ~n30237 ;
  assign y18946 = n30240 ;
  assign y18947 = ~n23135 ;
  assign y18948 = n30241 ;
  assign y18949 = ~1'b0 ;
  assign y18950 = n30242 ;
  assign y18951 = n30244 ;
  assign y18952 = ~n7996 ;
  assign y18953 = ~1'b0 ;
  assign y18954 = ~n30248 ;
  assign y18955 = ~1'b0 ;
  assign y18956 = ~n30259 ;
  assign y18957 = n30260 ;
  assign y18958 = n30261 ;
  assign y18959 = n8396 ;
  assign y18960 = ~1'b0 ;
  assign y18961 = n30263 ;
  assign y18962 = ~1'b0 ;
  assign y18963 = ~n30265 ;
  assign y18964 = ~n30267 ;
  assign y18965 = ~1'b0 ;
  assign y18966 = ~1'b0 ;
  assign y18967 = ~n30270 ;
  assign y18968 = n30272 ;
  assign y18969 = ~n30273 ;
  assign y18970 = ~1'b0 ;
  assign y18971 = ~1'b0 ;
  assign y18972 = ~1'b0 ;
  assign y18973 = n30274 ;
  assign y18974 = ~n30275 ;
  assign y18975 = ~1'b0 ;
  assign y18976 = n30278 ;
  assign y18977 = n13636 ;
  assign y18978 = ~1'b0 ;
  assign y18979 = n30280 ;
  assign y18980 = ~n30281 ;
  assign y18981 = n30285 ;
  assign y18982 = ~n4325 ;
  assign y18983 = n30287 ;
  assign y18984 = ~1'b0 ;
  assign y18985 = ~n30288 ;
  assign y18986 = ~n30291 ;
  assign y18987 = ~n30295 ;
  assign y18988 = ~1'b0 ;
  assign y18989 = n30298 ;
  assign y18990 = ~n30306 ;
  assign y18991 = ~1'b0 ;
  assign y18992 = ~n30307 ;
  assign y18993 = n30309 ;
  assign y18994 = ~n30313 ;
  assign y18995 = n30318 ;
  assign y18996 = n30319 ;
  assign y18997 = ~1'b0 ;
  assign y18998 = n30321 ;
  assign y18999 = ~1'b0 ;
  assign y19000 = ~n30323 ;
  assign y19001 = ~n30324 ;
  assign y19002 = ~1'b0 ;
  assign y19003 = n30329 ;
  assign y19004 = ~1'b0 ;
  assign y19005 = ~n30333 ;
  assign y19006 = 1'b0 ;
  assign y19007 = ~1'b0 ;
  assign y19008 = ~n30341 ;
  assign y19009 = n30344 ;
  assign y19010 = ~n14694 ;
  assign y19011 = ~n30346 ;
  assign y19012 = ~1'b0 ;
  assign y19013 = n8713 ;
  assign y19014 = ~n30347 ;
  assign y19015 = ~n30348 ;
  assign y19016 = 1'b0 ;
  assign y19017 = n30350 ;
  assign y19018 = ~n30352 ;
  assign y19019 = ~1'b0 ;
  assign y19020 = ~n13895 ;
  assign y19021 = n30353 ;
  assign y19022 = ~n30355 ;
  assign y19023 = n30356 ;
  assign y19024 = n30357 ;
  assign y19025 = ~1'b0 ;
  assign y19026 = ~1'b0 ;
  assign y19027 = ~1'b0 ;
  assign y19028 = n30358 ;
  assign y19029 = ~n30363 ;
  assign y19030 = n5054 ;
  assign y19031 = n6195 ;
  assign y19032 = ~n30375 ;
  assign y19033 = ~1'b0 ;
  assign y19034 = n30376 ;
  assign y19035 = ~1'b0 ;
  assign y19036 = n30378 ;
  assign y19037 = ~1'b0 ;
  assign y19038 = ~1'b0 ;
  assign y19039 = ~n30385 ;
  assign y19040 = ~n30387 ;
  assign y19041 = ~1'b0 ;
  assign y19042 = ~1'b0 ;
  assign y19043 = ~1'b0 ;
  assign y19044 = ~n30392 ;
  assign y19045 = 1'b0 ;
  assign y19046 = ~n30393 ;
  assign y19047 = ~n30396 ;
  assign y19048 = ~1'b0 ;
  assign y19049 = ~n30398 ;
  assign y19050 = n30399 ;
  assign y19051 = 1'b0 ;
  assign y19052 = ~n30400 ;
  assign y19053 = ~n30402 ;
  assign y19054 = ~n30403 ;
  assign y19055 = ~n30405 ;
  assign y19056 = ~1'b0 ;
  assign y19057 = ~1'b0 ;
  assign y19058 = ~1'b0 ;
  assign y19059 = ~n30406 ;
  assign y19060 = ~n30408 ;
  assign y19061 = ~n30409 ;
  assign y19062 = ~1'b0 ;
  assign y19063 = ~1'b0 ;
  assign y19064 = ~n30412 ;
  assign y19065 = ~n30413 ;
  assign y19066 = n30414 ;
  assign y19067 = ~n30416 ;
  assign y19068 = ~1'b0 ;
  assign y19069 = 1'b0 ;
  assign y19070 = n30417 ;
  assign y19071 = ~1'b0 ;
  assign y19072 = ~n30424 ;
  assign y19073 = ~1'b0 ;
  assign y19074 = ~1'b0 ;
  assign y19075 = ~1'b0 ;
  assign y19076 = n30425 ;
  assign y19077 = ~n30426 ;
  assign y19078 = ~1'b0 ;
  assign y19079 = ~1'b0 ;
  assign y19080 = ~1'b0 ;
  assign y19081 = n30429 ;
  assign y19082 = n30433 ;
  assign y19083 = ~1'b0 ;
  assign y19084 = ~n30436 ;
  assign y19085 = ~1'b0 ;
  assign y19086 = n30448 ;
  assign y19087 = n24789 ;
  assign y19088 = n30450 ;
  assign y19089 = ~n30456 ;
  assign y19090 = ~1'b0 ;
  assign y19091 = ~n30458 ;
  assign y19092 = ~n30459 ;
  assign y19093 = ~1'b0 ;
  assign y19094 = ~n30461 ;
  assign y19095 = n30462 ;
  assign y19096 = ~1'b0 ;
  assign y19097 = n30463 ;
  assign y19098 = n17182 ;
  assign y19099 = n30465 ;
  assign y19100 = n30466 ;
  assign y19101 = n30467 ;
  assign y19102 = ~1'b0 ;
  assign y19103 = ~n30470 ;
  assign y19104 = ~n30472 ;
  assign y19105 = ~n30474 ;
  assign y19106 = ~1'b0 ;
  assign y19107 = 1'b0 ;
  assign y19108 = ~1'b0 ;
  assign y19109 = n7822 ;
  assign y19110 = n30475 ;
  assign y19111 = n8633 ;
  assign y19112 = ~1'b0 ;
  assign y19113 = ~n30477 ;
  assign y19114 = ~1'b0 ;
  assign y19115 = ~n30480 ;
  assign y19116 = ~n30483 ;
  assign y19117 = n30487 ;
  assign y19118 = ~1'b0 ;
  assign y19119 = n30488 ;
  assign y19120 = ~n30490 ;
  assign y19121 = n30491 ;
  assign y19122 = n30493 ;
  assign y19123 = ~n30495 ;
  assign y19124 = ~1'b0 ;
  assign y19125 = ~1'b0 ;
  assign y19126 = ~1'b0 ;
  assign y19127 = n8646 ;
  assign y19128 = n30496 ;
  assign y19129 = ~1'b0 ;
  assign y19130 = ~n30504 ;
  assign y19131 = ~n30505 ;
  assign y19132 = ~n30506 ;
  assign y19133 = n30507 ;
  assign y19134 = ~n30508 ;
  assign y19135 = ~1'b0 ;
  assign y19136 = ~n30509 ;
  assign y19137 = ~n30512 ;
  assign y19138 = n30513 ;
  assign y19139 = n30514 ;
  assign y19140 = ~n30517 ;
  assign y19141 = ~n30522 ;
  assign y19142 = n26866 ;
  assign y19143 = ~n30526 ;
  assign y19144 = n30528 ;
  assign y19145 = ~1'b0 ;
  assign y19146 = n30531 ;
  assign y19147 = ~n30533 ;
  assign y19148 = ~n30534 ;
  assign y19149 = ~n30535 ;
  assign y19150 = n30537 ;
  assign y19151 = n30538 ;
  assign y19152 = ~1'b0 ;
  assign y19153 = ~1'b0 ;
  assign y19154 = ~n30539 ;
  assign y19155 = ~1'b0 ;
  assign y19156 = ~n30542 ;
  assign y19157 = ~n30545 ;
  assign y19158 = ~n257 ;
  assign y19159 = n30549 ;
  assign y19160 = n30552 ;
  assign y19161 = ~n271 ;
  assign y19162 = n29709 ;
  assign y19163 = ~n30558 ;
  assign y19164 = n30560 ;
  assign y19165 = ~n30562 ;
  assign y19166 = ~n30565 ;
  assign y19167 = ~1'b0 ;
  assign y19168 = ~1'b0 ;
  assign y19169 = ~n30566 ;
  assign y19170 = n30568 ;
  assign y19171 = ~1'b0 ;
  assign y19172 = n30569 ;
  assign y19173 = ~1'b0 ;
  assign y19174 = ~n30574 ;
  assign y19175 = ~1'b0 ;
  assign y19176 = ~n10396 ;
  assign y19177 = n30577 ;
  assign y19178 = ~1'b0 ;
  assign y19179 = ~n17550 ;
  assign y19180 = n30579 ;
  assign y19181 = ~n30583 ;
  assign y19182 = n30584 ;
  assign y19183 = ~n11341 ;
  assign y19184 = ~n30587 ;
  assign y19185 = ~1'b0 ;
  assign y19186 = n30588 ;
  assign y19187 = n30593 ;
  assign y19188 = n30594 ;
  assign y19189 = ~1'b0 ;
  assign y19190 = ~1'b0 ;
  assign y19191 = ~n30595 ;
  assign y19192 = ~1'b0 ;
  assign y19193 = ~1'b0 ;
  assign y19194 = ~1'b0 ;
  assign y19195 = ~n30596 ;
  assign y19196 = ~n30600 ;
  assign y19197 = n30602 ;
  assign y19198 = ~n30604 ;
  assign y19199 = ~1'b0 ;
  assign y19200 = n30605 ;
  assign y19201 = ~1'b0 ;
  assign y19202 = ~n30608 ;
  assign y19203 = n30609 ;
  assign y19204 = ~n30610 ;
  assign y19205 = ~n30612 ;
  assign y19206 = ~n30620 ;
  assign y19207 = ~1'b0 ;
  assign y19208 = n30621 ;
  assign y19209 = ~n30623 ;
  assign y19210 = ~n30624 ;
  assign y19211 = ~n30625 ;
  assign y19212 = ~n30627 ;
  assign y19213 = ~n30628 ;
  assign y19214 = ~1'b0 ;
  assign y19215 = 1'b0 ;
  assign y19216 = ~n13313 ;
  assign y19217 = n30631 ;
  assign y19218 = 1'b0 ;
  assign y19219 = ~1'b0 ;
  assign y19220 = ~n30636 ;
  assign y19221 = ~1'b0 ;
  assign y19222 = ~n30638 ;
  assign y19223 = ~1'b0 ;
  assign y19224 = ~1'b0 ;
  assign y19225 = ~n30639 ;
  assign y19226 = ~n30640 ;
  assign y19227 = n21658 ;
  assign y19228 = ~n30641 ;
  assign y19229 = n30642 ;
  assign y19230 = ~n20715 ;
  assign y19231 = ~1'b0 ;
  assign y19232 = ~1'b0 ;
  assign y19233 = n30644 ;
  assign y19234 = ~n30645 ;
  assign y19235 = ~1'b0 ;
  assign y19236 = ~1'b0 ;
  assign y19237 = ~1'b0 ;
  assign y19238 = ~1'b0 ;
  assign y19239 = n30647 ;
  assign y19240 = 1'b0 ;
  assign y19241 = ~1'b0 ;
  assign y19242 = 1'b0 ;
  assign y19243 = n30649 ;
  assign y19244 = ~n10724 ;
  assign y19245 = n30650 ;
  assign y19246 = ~1'b0 ;
  assign y19247 = n30652 ;
  assign y19248 = ~1'b0 ;
  assign y19249 = n6625 ;
  assign y19250 = ~n30653 ;
  assign y19251 = n30655 ;
  assign y19252 = ~n30658 ;
  assign y19253 = n30660 ;
  assign y19254 = n1688 ;
  assign y19255 = n30662 ;
  assign y19256 = 1'b0 ;
  assign y19257 = ~1'b0 ;
  assign y19258 = ~n30663 ;
  assign y19259 = ~n29762 ;
  assign y19260 = ~n30665 ;
  assign y19261 = n23737 ;
  assign y19262 = n30667 ;
  assign y19263 = ~n30669 ;
  assign y19264 = ~n30670 ;
  assign y19265 = n30672 ;
  assign y19266 = n30675 ;
  assign y19267 = ~1'b0 ;
  assign y19268 = n30677 ;
  assign y19269 = ~n1791 ;
  assign y19270 = n30679 ;
  assign y19271 = ~n30680 ;
  assign y19272 = ~n27098 ;
  assign y19273 = ~1'b0 ;
  assign y19274 = ~1'b0 ;
  assign y19275 = n30681 ;
  assign y19276 = ~1'b0 ;
  assign y19277 = ~1'b0 ;
  assign y19278 = ~1'b0 ;
  assign y19279 = ~n30687 ;
  assign y19280 = n30688 ;
  assign y19281 = ~1'b0 ;
  assign y19282 = ~n30689 ;
  assign y19283 = 1'b0 ;
  assign y19284 = n30691 ;
  assign y19285 = ~1'b0 ;
  assign y19286 = n30692 ;
  assign y19287 = n30694 ;
  assign y19288 = ~1'b0 ;
  assign y19289 = 1'b0 ;
  assign y19290 = n30697 ;
  assign y19291 = ~1'b0 ;
  assign y19292 = ~1'b0 ;
  assign y19293 = ~1'b0 ;
  assign y19294 = n30698 ;
  assign y19295 = ~1'b0 ;
  assign y19296 = n30699 ;
  assign y19297 = n30700 ;
  assign y19298 = 1'b0 ;
  assign y19299 = ~1'b0 ;
  assign y19300 = ~1'b0 ;
  assign y19301 = n30701 ;
  assign y19302 = ~n30702 ;
  assign y19303 = ~n23739 ;
  assign y19304 = n30704 ;
  assign y19305 = ~1'b0 ;
  assign y19306 = n30707 ;
  assign y19307 = n30709 ;
  assign y19308 = ~n30710 ;
  assign y19309 = n30711 ;
  assign y19310 = n30717 ;
  assign y19311 = ~1'b0 ;
  assign y19312 = ~1'b0 ;
  assign y19313 = n1404 ;
  assign y19314 = n30205 ;
  assign y19315 = n30719 ;
  assign y19316 = ~1'b0 ;
  assign y19317 = ~1'b0 ;
  assign y19318 = ~1'b0 ;
  assign y19319 = ~1'b0 ;
  assign y19320 = n30723 ;
  assign y19321 = ~1'b0 ;
  assign y19322 = n30725 ;
  assign y19323 = n30728 ;
  assign y19324 = ~n30731 ;
  assign y19325 = ~1'b0 ;
  assign y19326 = ~1'b0 ;
  assign y19327 = 1'b0 ;
  assign y19328 = n30732 ;
  assign y19329 = ~n30734 ;
  assign y19330 = ~1'b0 ;
  assign y19331 = ~1'b0 ;
  assign y19332 = n30735 ;
  assign y19333 = ~n8816 ;
  assign y19334 = n4727 ;
  assign y19335 = n15123 ;
  assign y19336 = ~n30737 ;
  assign y19337 = ~n30739 ;
  assign y19338 = ~n30740 ;
  assign y19339 = ~n30743 ;
  assign y19340 = ~n30744 ;
  assign y19341 = n30745 ;
  assign y19342 = n17322 ;
  assign y19343 = ~n30746 ;
  assign y19344 = n27766 ;
  assign y19345 = ~1'b0 ;
  assign y19346 = ~1'b0 ;
  assign y19347 = ~1'b0 ;
  assign y19348 = ~1'b0 ;
  assign y19349 = ~n30747 ;
  assign y19350 = n30748 ;
  assign y19351 = ~1'b0 ;
  assign y19352 = ~1'b0 ;
  assign y19353 = ~n7984 ;
  assign y19354 = ~n30751 ;
  assign y19355 = n30752 ;
  assign y19356 = ~n11465 ;
  assign y19357 = n26207 ;
  assign y19358 = ~1'b0 ;
  assign y19359 = n30753 ;
  assign y19360 = 1'b0 ;
  assign y19361 = ~n30754 ;
  assign y19362 = ~1'b0 ;
  assign y19363 = ~1'b0 ;
  assign y19364 = ~n30755 ;
  assign y19365 = n30757 ;
  assign y19366 = ~1'b0 ;
  assign y19367 = ~1'b0 ;
  assign y19368 = ~n30759 ;
  assign y19369 = ~n6068 ;
  assign y19370 = ~1'b0 ;
  assign y19371 = ~1'b0 ;
  assign y19372 = ~1'b0 ;
  assign y19373 = 1'b0 ;
  assign y19374 = ~n30760 ;
  assign y19375 = ~1'b0 ;
  assign y19376 = ~1'b0 ;
  assign y19377 = ~n17714 ;
  assign y19378 = ~1'b0 ;
  assign y19379 = ~n30766 ;
  assign y19380 = ~n30768 ;
  assign y19381 = n30769 ;
  assign y19382 = n16489 ;
  assign y19383 = ~n30770 ;
  assign y19384 = n30771 ;
  assign y19385 = ~1'b0 ;
  assign y19386 = n30775 ;
  assign y19387 = ~n22533 ;
  assign y19388 = n30779 ;
  assign y19389 = ~n30782 ;
  assign y19390 = ~n17322 ;
  assign y19391 = ~1'b0 ;
  assign y19392 = 1'b0 ;
  assign y19393 = ~1'b0 ;
  assign y19394 = ~1'b0 ;
  assign y19395 = n30785 ;
  assign y19396 = ~n30788 ;
  assign y19397 = ~n30791 ;
  assign y19398 = n25708 ;
  assign y19399 = n30795 ;
  assign y19400 = ~n30798 ;
  assign y19401 = ~1'b0 ;
  assign y19402 = ~1'b0 ;
  assign y19403 = ~1'b0 ;
  assign y19404 = n30801 ;
  assign y19405 = ~n30802 ;
  assign y19406 = 1'b0 ;
  assign y19407 = ~1'b0 ;
  assign y19408 = ~n30805 ;
  assign y19409 = ~1'b0 ;
  assign y19410 = ~1'b0 ;
  assign y19411 = ~1'b0 ;
  assign y19412 = ~1'b0 ;
  assign y19413 = n30807 ;
  assign y19414 = ~1'b0 ;
  assign y19415 = ~n26040 ;
  assign y19416 = ~1'b0 ;
  assign y19417 = n30809 ;
  assign y19418 = ~1'b0 ;
  assign y19419 = 1'b0 ;
  assign y19420 = ~n30811 ;
  assign y19421 = ~n30812 ;
  assign y19422 = n30814 ;
  assign y19423 = ~n30816 ;
  assign y19424 = ~1'b0 ;
  assign y19425 = n21989 ;
  assign y19426 = ~n30820 ;
  assign y19427 = n24140 ;
  assign y19428 = n30821 ;
  assign y19429 = n30824 ;
  assign y19430 = ~n30827 ;
  assign y19431 = ~n30828 ;
  assign y19432 = 1'b0 ;
  assign y19433 = ~n30829 ;
  assign y19434 = ~n4578 ;
  assign y19435 = ~n30830 ;
  assign y19436 = ~1'b0 ;
  assign y19437 = ~n18137 ;
  assign y19438 = ~n30832 ;
  assign y19439 = ~1'b0 ;
  assign y19440 = ~1'b0 ;
  assign y19441 = n30835 ;
  assign y19442 = ~1'b0 ;
  assign y19443 = ~n24622 ;
  assign y19444 = ~1'b0 ;
  assign y19445 = n30836 ;
  assign y19446 = ~1'b0 ;
  assign y19447 = ~n26269 ;
  assign y19448 = ~1'b0 ;
  assign y19449 = ~1'b0 ;
  assign y19450 = n30839 ;
  assign y19451 = ~1'b0 ;
  assign y19452 = n30841 ;
  assign y19453 = n30842 ;
  assign y19454 = n30844 ;
  assign y19455 = ~1'b0 ;
  assign y19456 = n30846 ;
  assign y19457 = ~n30848 ;
  assign y19458 = ~n1511 ;
  assign y19459 = ~1'b0 ;
  assign y19460 = ~n30849 ;
  assign y19461 = ~1'b0 ;
  assign y19462 = ~1'b0 ;
  assign y19463 = ~n30851 ;
  assign y19464 = ~n12136 ;
  assign y19465 = n30852 ;
  assign y19466 = ~n30855 ;
  assign y19467 = ~1'b0 ;
  assign y19468 = n30857 ;
  assign y19469 = n30862 ;
  assign y19470 = n30864 ;
  assign y19471 = ~n30866 ;
  assign y19472 = ~n30870 ;
  assign y19473 = ~1'b0 ;
  assign y19474 = ~1'b0 ;
  assign y19475 = ~1'b0 ;
  assign y19476 = ~1'b0 ;
  assign y19477 = ~1'b0 ;
  assign y19478 = ~1'b0 ;
  assign y19479 = ~n30872 ;
  assign y19480 = n2517 ;
  assign y19481 = ~1'b0 ;
  assign y19482 = ~n30873 ;
  assign y19483 = 1'b0 ;
  assign y19484 = ~1'b0 ;
  assign y19485 = ~n30875 ;
  assign y19486 = n30877 ;
  assign y19487 = ~n30880 ;
  assign y19488 = ~1'b0 ;
  assign y19489 = ~1'b0 ;
  assign y19490 = ~n13649 ;
  assign y19491 = n30883 ;
  assign y19492 = n30885 ;
  assign y19493 = ~n30887 ;
  assign y19494 = ~1'b0 ;
  assign y19495 = ~1'b0 ;
  assign y19496 = ~1'b0 ;
  assign y19497 = n30889 ;
  assign y19498 = n30891 ;
  assign y19499 = n30892 ;
  assign y19500 = ~1'b0 ;
  assign y19501 = n30894 ;
  assign y19502 = ~1'b0 ;
  assign y19503 = ~n30899 ;
  assign y19504 = n30900 ;
  assign y19505 = n30901 ;
  assign y19506 = ~n30905 ;
  assign y19507 = ~n30906 ;
  assign y19508 = ~1'b0 ;
  assign y19509 = ~1'b0 ;
  assign y19510 = ~n30908 ;
  assign y19511 = ~n30915 ;
  assign y19512 = n30916 ;
  assign y19513 = ~n27029 ;
  assign y19514 = n1922 ;
  assign y19515 = ~1'b0 ;
  assign y19516 = ~1'b0 ;
  assign y19517 = ~1'b0 ;
  assign y19518 = ~1'b0 ;
  assign y19519 = ~1'b0 ;
  assign y19520 = n30920 ;
  assign y19521 = n30921 ;
  assign y19522 = ~n30923 ;
  assign y19523 = ~n30925 ;
  assign y19524 = ~n30926 ;
  assign y19525 = ~n30929 ;
  assign y19526 = n30932 ;
  assign y19527 = ~n30934 ;
  assign y19528 = ~1'b0 ;
  assign y19529 = n30935 ;
  assign y19530 = n30939 ;
  assign y19531 = ~n30940 ;
  assign y19532 = n30942 ;
  assign y19533 = ~1'b0 ;
  assign y19534 = ~1'b0 ;
  assign y19535 = ~n30944 ;
  assign y19536 = ~1'b0 ;
  assign y19537 = ~1'b0 ;
  assign y19538 = ~n30946 ;
  assign y19539 = ~1'b0 ;
  assign y19540 = ~1'b0 ;
  assign y19541 = ~n30949 ;
  assign y19542 = ~1'b0 ;
  assign y19543 = ~1'b0 ;
  assign y19544 = ~1'b0 ;
  assign y19545 = ~1'b0 ;
  assign y19546 = n30950 ;
  assign y19547 = ~n27905 ;
  assign y19548 = ~n30952 ;
  assign y19549 = n30958 ;
  assign y19550 = ~1'b0 ;
  assign y19551 = ~n30960 ;
  assign y19552 = ~n30963 ;
  assign y19553 = n30964 ;
  assign y19554 = ~n30967 ;
  assign y19555 = ~1'b0 ;
  assign y19556 = n30968 ;
  assign y19557 = n30969 ;
  assign y19558 = ~n30970 ;
  assign y19559 = ~1'b0 ;
  assign y19560 = n30972 ;
  assign y19561 = ~n30974 ;
  assign y19562 = ~n30976 ;
  assign y19563 = ~n30977 ;
  assign y19564 = 1'b0 ;
  assign y19565 = n30979 ;
  assign y19566 = n7744 ;
  assign y19567 = n30981 ;
  assign y19568 = ~1'b0 ;
  assign y19569 = n30986 ;
  assign y19570 = n30987 ;
  assign y19571 = n30988 ;
  assign y19572 = ~n30989 ;
  assign y19573 = n30990 ;
  assign y19574 = ~1'b0 ;
  assign y19575 = ~1'b0 ;
  assign y19576 = n30993 ;
  assign y19577 = ~n30994 ;
  assign y19578 = ~1'b0 ;
  assign y19579 = 1'b0 ;
  assign y19580 = ~n30995 ;
  assign y19581 = ~1'b0 ;
  assign y19582 = ~n30997 ;
  assign y19583 = ~1'b0 ;
  assign y19584 = ~1'b0 ;
  assign y19585 = ~n31000 ;
  assign y19586 = ~1'b0 ;
  assign y19587 = ~n31002 ;
  assign y19588 = n31003 ;
  assign y19589 = ~n2318 ;
  assign y19590 = n21762 ;
  assign y19591 = n31005 ;
  assign y19592 = ~1'b0 ;
  assign y19593 = ~1'b0 ;
  assign y19594 = n31006 ;
  assign y19595 = n31008 ;
  assign y19596 = ~n31009 ;
  assign y19597 = ~n31011 ;
  assign y19598 = ~1'b0 ;
  assign y19599 = ~1'b0 ;
  assign y19600 = ~1'b0 ;
  assign y19601 = n31012 ;
  assign y19602 = ~n7766 ;
  assign y19603 = ~n31014 ;
  assign y19604 = ~1'b0 ;
  assign y19605 = ~n31018 ;
  assign y19606 = n31019 ;
  assign y19607 = n31024 ;
  assign y19608 = ~n31025 ;
  assign y19609 = n10298 ;
  assign y19610 = ~1'b0 ;
  assign y19611 = ~n31027 ;
  assign y19612 = n31028 ;
  assign y19613 = ~n31029 ;
  assign y19614 = ~1'b0 ;
  assign y19615 = n31031 ;
  assign y19616 = ~1'b0 ;
  assign y19617 = n4087 ;
  assign y19618 = n31032 ;
  assign y19619 = ~1'b0 ;
  assign y19620 = ~1'b0 ;
  assign y19621 = ~n31033 ;
  assign y19622 = n31035 ;
  assign y19623 = n31039 ;
  assign y19624 = ~1'b0 ;
  assign y19625 = 1'b0 ;
  assign y19626 = ~n31042 ;
  assign y19627 = ~n31044 ;
  assign y19628 = ~1'b0 ;
  assign y19629 = 1'b0 ;
  assign y19630 = ~n31046 ;
  assign y19631 = n31047 ;
  assign y19632 = ~1'b0 ;
  assign y19633 = ~n31056 ;
  assign y19634 = ~1'b0 ;
  assign y19635 = ~n31063 ;
  assign y19636 = ~1'b0 ;
  assign y19637 = ~1'b0 ;
  assign y19638 = ~n31066 ;
  assign y19639 = ~n12207 ;
  assign y19640 = 1'b0 ;
  assign y19641 = ~1'b0 ;
  assign y19642 = ~n21712 ;
  assign y19643 = 1'b0 ;
  assign y19644 = ~1'b0 ;
  assign y19645 = ~1'b0 ;
  assign y19646 = n31067 ;
  assign y19647 = ~n31071 ;
  assign y19648 = ~n23185 ;
  assign y19649 = n1952 ;
  assign y19650 = ~1'b0 ;
  assign y19651 = ~1'b0 ;
  assign y19652 = ~n31072 ;
  assign y19653 = ~n31073 ;
  assign y19654 = ~n31074 ;
  assign y19655 = n31076 ;
  assign y19656 = n31077 ;
  assign y19657 = ~1'b0 ;
  assign y19658 = ~1'b0 ;
  assign y19659 = ~1'b0 ;
  assign y19660 = 1'b0 ;
  assign y19661 = ~n31079 ;
  assign y19662 = ~1'b0 ;
  assign y19663 = ~n31082 ;
  assign y19664 = ~n31084 ;
  assign y19665 = ~1'b0 ;
  assign y19666 = n2269 ;
  assign y19667 = ~1'b0 ;
  assign y19668 = n31088 ;
  assign y19669 = n31090 ;
  assign y19670 = ~n31096 ;
  assign y19671 = ~1'b0 ;
  assign y19672 = ~n31098 ;
  assign y19673 = n503 ;
  assign y19674 = ~1'b0 ;
  assign y19675 = n2097 ;
  assign y19676 = n31100 ;
  assign y19677 = ~1'b0 ;
  assign y19678 = n31101 ;
  assign y19679 = n31102 ;
  assign y19680 = ~n31103 ;
  assign y19681 = n31108 ;
  assign y19682 = ~n31109 ;
  assign y19683 = ~1'b0 ;
  assign y19684 = ~1'b0 ;
  assign y19685 = n31110 ;
  assign y19686 = ~1'b0 ;
  assign y19687 = ~1'b0 ;
  assign y19688 = ~1'b0 ;
  assign y19689 = ~1'b0 ;
  assign y19690 = ~n31112 ;
  assign y19691 = ~1'b0 ;
  assign y19692 = n31113 ;
  assign y19693 = ~1'b0 ;
  assign y19694 = ~n31114 ;
  assign y19695 = ~n31116 ;
  assign y19696 = ~1'b0 ;
  assign y19697 = 1'b0 ;
  assign y19698 = ~1'b0 ;
  assign y19699 = n1031 ;
  assign y19700 = ~n31117 ;
  assign y19701 = ~n31119 ;
  assign y19702 = ~1'b0 ;
  assign y19703 = ~1'b0 ;
  assign y19704 = n31121 ;
  assign y19705 = n31122 ;
  assign y19706 = ~n31127 ;
  assign y19707 = ~1'b0 ;
  assign y19708 = ~1'b0 ;
  assign y19709 = ~n31133 ;
  assign y19710 = n9700 ;
  assign y19711 = ~n31136 ;
  assign y19712 = ~n31137 ;
  assign y19713 = ~n31139 ;
  assign y19714 = ~n31141 ;
  assign y19715 = ~n31143 ;
  assign y19716 = ~n31145 ;
  assign y19717 = ~n31147 ;
  assign y19718 = ~n31148 ;
  assign y19719 = ~1'b0 ;
  assign y19720 = n31150 ;
  assign y19721 = ~n31151 ;
  assign y19722 = n31153 ;
  assign y19723 = ~1'b0 ;
  assign y19724 = 1'b0 ;
  assign y19725 = ~n31155 ;
  assign y19726 = ~1'b0 ;
  assign y19727 = ~1'b0 ;
  assign y19728 = n31158 ;
  assign y19729 = n2879 ;
  assign y19730 = ~1'b0 ;
  assign y19731 = n31161 ;
  assign y19732 = ~n31162 ;
  assign y19733 = ~n31165 ;
  assign y19734 = n31167 ;
  assign y19735 = n31168 ;
  assign y19736 = ~1'b0 ;
  assign y19737 = n31173 ;
  assign y19738 = ~1'b0 ;
  assign y19739 = n6644 ;
  assign y19740 = ~1'b0 ;
  assign y19741 = n28374 ;
  assign y19742 = ~n23065 ;
  assign y19743 = ~1'b0 ;
  assign y19744 = ~1'b0 ;
  assign y19745 = ~1'b0 ;
  assign y19746 = ~1'b0 ;
  assign y19747 = ~n31175 ;
  assign y19748 = n31178 ;
  assign y19749 = ~n31181 ;
  assign y19750 = ~1'b0 ;
  assign y19751 = 1'b0 ;
  assign y19752 = n31182 ;
  assign y19753 = n20310 ;
  assign y19754 = n31183 ;
  assign y19755 = ~1'b0 ;
  assign y19756 = ~n31186 ;
  assign y19757 = ~n31187 ;
  assign y19758 = ~1'b0 ;
  assign y19759 = ~1'b0 ;
  assign y19760 = ~1'b0 ;
  assign y19761 = ~n31190 ;
  assign y19762 = ~n31192 ;
  assign y19763 = n19682 ;
  assign y19764 = n31194 ;
  assign y19765 = ~n31196 ;
  assign y19766 = ~n31198 ;
  assign y19767 = ~n31199 ;
  assign y19768 = ~n23273 ;
  assign y19769 = n31200 ;
  assign y19770 = ~n31201 ;
  assign y19771 = n31202 ;
  assign y19772 = ~n31203 ;
  assign y19773 = ~n31207 ;
  assign y19774 = 1'b0 ;
  assign y19775 = ~n31208 ;
  assign y19776 = ~n31210 ;
  assign y19777 = ~n31211 ;
  assign y19778 = ~1'b0 ;
  assign y19779 = ~n31213 ;
  assign y19780 = n31214 ;
  assign y19781 = n31219 ;
  assign y19782 = ~1'b0 ;
  assign y19783 = ~n31223 ;
  assign y19784 = ~n31225 ;
  assign y19785 = ~1'b0 ;
  assign y19786 = ~1'b0 ;
  assign y19787 = ~1'b0 ;
  assign y19788 = n31226 ;
  assign y19789 = ~n31227 ;
  assign y19790 = ~1'b0 ;
  assign y19791 = ~n31229 ;
  assign y19792 = n31232 ;
  assign y19793 = ~1'b0 ;
  assign y19794 = n31233 ;
  assign y19795 = n31234 ;
  assign y19796 = n31247 ;
  assign y19797 = ~1'b0 ;
  assign y19798 = ~n31249 ;
  assign y19799 = n31251 ;
  assign y19800 = ~1'b0 ;
  assign y19801 = ~n31257 ;
  assign y19802 = ~1'b0 ;
  assign y19803 = n18952 ;
  assign y19804 = n31260 ;
  assign y19805 = n31262 ;
  assign y19806 = ~n31268 ;
  assign y19807 = ~1'b0 ;
  assign y19808 = ~n31275 ;
  assign y19809 = n31277 ;
  assign y19810 = ~n31280 ;
  assign y19811 = n31281 ;
  assign y19812 = ~n3678 ;
  assign y19813 = n31290 ;
  assign y19814 = ~n31294 ;
  assign y19815 = n31295 ;
  assign y19816 = ~n31296 ;
  assign y19817 = n31297 ;
  assign y19818 = ~n31301 ;
  assign y19819 = ~1'b0 ;
  assign y19820 = ~1'b0 ;
  assign y19821 = ~n31303 ;
  assign y19822 = ~n31305 ;
  assign y19823 = ~n31307 ;
  assign y19824 = n31308 ;
  assign y19825 = ~n2450 ;
  assign y19826 = ~1'b0 ;
  assign y19827 = n31311 ;
  assign y19828 = n31315 ;
  assign y19829 = 1'b0 ;
  assign y19830 = n31316 ;
  assign y19831 = ~n31318 ;
  assign y19832 = n31320 ;
  assign y19833 = ~n31324 ;
  assign y19834 = n31326 ;
  assign y19835 = n31328 ;
  assign y19836 = ~n31330 ;
  assign y19837 = ~n31331 ;
  assign y19838 = n2175 ;
  assign y19839 = ~1'b0 ;
  assign y19840 = ~1'b0 ;
  assign y19841 = ~n31333 ;
  assign y19842 = n31334 ;
  assign y19843 = ~n31336 ;
  assign y19844 = n31337 ;
  assign y19845 = n31338 ;
  assign y19846 = ~n31347 ;
  assign y19847 = ~1'b0 ;
  assign y19848 = ~n31348 ;
  assign y19849 = ~1'b0 ;
  assign y19850 = ~1'b0 ;
  assign y19851 = ~1'b0 ;
  assign y19852 = ~1'b0 ;
  assign y19853 = n31350 ;
  assign y19854 = ~1'b0 ;
  assign y19855 = n31351 ;
  assign y19856 = ~n31352 ;
  assign y19857 = ~n31355 ;
  assign y19858 = ~1'b0 ;
  assign y19859 = 1'b0 ;
  assign y19860 = ~1'b0 ;
  assign y19861 = n31356 ;
  assign y19862 = ~n31358 ;
  assign y19863 = ~1'b0 ;
  assign y19864 = ~1'b0 ;
  assign y19865 = n31359 ;
  assign y19866 = ~1'b0 ;
  assign y19867 = ~1'b0 ;
  assign y19868 = ~1'b0 ;
  assign y19869 = ~1'b0 ;
  assign y19870 = ~1'b0 ;
  assign y19871 = ~1'b0 ;
  assign y19872 = n31362 ;
  assign y19873 = 1'b0 ;
  assign y19874 = ~1'b0 ;
  assign y19875 = ~n12621 ;
  assign y19876 = ~n31365 ;
  assign y19877 = n31366 ;
  assign y19878 = 1'b0 ;
  assign y19879 = ~1'b0 ;
  assign y19880 = ~n31372 ;
  assign y19881 = n360 ;
  assign y19882 = ~1'b0 ;
  assign y19883 = ~1'b0 ;
  assign y19884 = ~n31373 ;
  assign y19885 = ~1'b0 ;
  assign y19886 = n31381 ;
  assign y19887 = n31382 ;
  assign y19888 = ~n31383 ;
  assign y19889 = n31388 ;
  assign y19890 = ~n1810 ;
  assign y19891 = ~n31389 ;
  assign y19892 = 1'b0 ;
  assign y19893 = n31390 ;
  assign y19894 = ~1'b0 ;
  assign y19895 = ~n31393 ;
  assign y19896 = ~n31394 ;
  assign y19897 = ~1'b0 ;
  assign y19898 = ~1'b0 ;
  assign y19899 = ~1'b0 ;
  assign y19900 = n31395 ;
  assign y19901 = ~n31396 ;
  assign y19902 = ~n31398 ;
  assign y19903 = ~n10334 ;
  assign y19904 = n31402 ;
  assign y19905 = ~n31404 ;
  assign y19906 = ~1'b0 ;
  assign y19907 = ~n31408 ;
  assign y19908 = ~n31410 ;
  assign y19909 = ~n31414 ;
  assign y19910 = ~1'b0 ;
  assign y19911 = ~n31415 ;
  assign y19912 = ~n31417 ;
  assign y19913 = n31418 ;
  assign y19914 = ~1'b0 ;
  assign y19915 = n31419 ;
  assign y19916 = n31421 ;
  assign y19917 = ~n14604 ;
  assign y19918 = ~n31424 ;
  assign y19919 = ~1'b0 ;
  assign y19920 = ~n31426 ;
  assign y19921 = ~1'b0 ;
  assign y19922 = n31428 ;
  assign y19923 = ~n31430 ;
  assign y19924 = n10663 ;
  assign y19925 = ~1'b0 ;
  assign y19926 = ~n31432 ;
  assign y19927 = ~n31433 ;
  assign y19928 = ~n31434 ;
  assign y19929 = n31435 ;
  assign y19930 = ~1'b0 ;
  assign y19931 = ~1'b0 ;
  assign y19932 = ~1'b0 ;
  assign y19933 = ~1'b0 ;
  assign y19934 = ~1'b0 ;
  assign y19935 = n31436 ;
  assign y19936 = ~1'b0 ;
  assign y19937 = n31439 ;
  assign y19938 = n31441 ;
  assign y19939 = n31442 ;
  assign y19940 = ~1'b0 ;
  assign y19941 = 1'b0 ;
  assign y19942 = n31445 ;
  assign y19943 = 1'b0 ;
  assign y19944 = n20120 ;
  assign y19945 = ~n31447 ;
  assign y19946 = n31448 ;
  assign y19947 = ~n31449 ;
  assign y19948 = ~1'b0 ;
  assign y19949 = n31452 ;
  assign y19950 = ~n31453 ;
  assign y19951 = 1'b0 ;
  assign y19952 = ~n31454 ;
  assign y19953 = ~1'b0 ;
  assign y19954 = ~n31457 ;
  assign y19955 = ~n19095 ;
  assign y19956 = ~n31458 ;
  assign y19957 = n31459 ;
  assign y19958 = ~1'b0 ;
  assign y19959 = ~1'b0 ;
  assign y19960 = ~n9875 ;
  assign y19961 = ~n31460 ;
  assign y19962 = ~n31461 ;
  assign y19963 = ~n31464 ;
  assign y19964 = ~1'b0 ;
  assign y19965 = n31468 ;
  assign y19966 = n31469 ;
  assign y19967 = ~1'b0 ;
  assign y19968 = n31472 ;
  assign y19969 = ~1'b0 ;
  assign y19970 = ~n31473 ;
  assign y19971 = ~1'b0 ;
  assign y19972 = n31476 ;
  assign y19973 = 1'b0 ;
  assign y19974 = ~1'b0 ;
  assign y19975 = ~1'b0 ;
  assign y19976 = ~n31480 ;
  assign y19977 = n31483 ;
  assign y19978 = ~n12973 ;
  assign y19979 = n31484 ;
  assign y19980 = ~n29412 ;
  assign y19981 = ~1'b0 ;
  assign y19982 = ~1'b0 ;
  assign y19983 = n23451 ;
  assign y19984 = ~n29924 ;
  assign y19985 = ~1'b0 ;
  assign y19986 = ~n31486 ;
  assign y19987 = n31487 ;
  assign y19988 = ~n31488 ;
  assign y19989 = ~1'b0 ;
  assign y19990 = n31489 ;
  assign y19991 = n31490 ;
  assign y19992 = ~n31491 ;
  assign y19993 = ~n31493 ;
  assign y19994 = ~n31496 ;
  assign y19995 = ~n31499 ;
  assign y19996 = n9446 ;
  assign y19997 = n31503 ;
  assign y19998 = n31504 ;
  assign y19999 = ~1'b0 ;
  assign y20000 = ~1'b0 ;
  assign y20001 = ~n31505 ;
  assign y20002 = n31506 ;
  assign y20003 = ~n12874 ;
  assign y20004 = n31511 ;
  assign y20005 = ~n31513 ;
  assign y20006 = ~1'b0 ;
  assign y20007 = n31516 ;
  assign y20008 = n31518 ;
  assign y20009 = n31519 ;
  assign y20010 = n31520 ;
  assign y20011 = n31526 ;
  assign y20012 = ~1'b0 ;
  assign y20013 = ~n31529 ;
  assign y20014 = ~n31532 ;
  assign y20015 = ~1'b0 ;
  assign y20016 = n31534 ;
  assign y20017 = ~n31536 ;
  assign y20018 = ~n15773 ;
  assign y20019 = ~1'b0 ;
  assign y20020 = ~n31537 ;
  assign y20021 = n31539 ;
  assign y20022 = ~n31546 ;
  assign y20023 = ~n31548 ;
  assign y20024 = ~n31549 ;
  assign y20025 = ~n15183 ;
  assign y20026 = ~1'b0 ;
  assign y20027 = n31551 ;
  assign y20028 = ~n31553 ;
  assign y20029 = n31556 ;
  assign y20030 = ~1'b0 ;
  assign y20031 = n31557 ;
  assign y20032 = ~1'b0 ;
  assign y20033 = ~n21588 ;
  assign y20034 = ~1'b0 ;
  assign y20035 = ~1'b0 ;
  assign y20036 = n31558 ;
  assign y20037 = ~1'b0 ;
  assign y20038 = n31559 ;
  assign y20039 = n31565 ;
  assign y20040 = ~n31566 ;
  assign y20041 = n30139 ;
  assign y20042 = n9066 ;
  assign y20043 = n31567 ;
  assign y20044 = n31568 ;
  assign y20045 = n31574 ;
  assign y20046 = ~1'b0 ;
  assign y20047 = ~1'b0 ;
  assign y20048 = n31576 ;
  assign y20049 = ~n31578 ;
  assign y20050 = n31579 ;
  assign y20051 = ~1'b0 ;
  assign y20052 = n17143 ;
  assign y20053 = n31581 ;
  assign y20054 = n1689 ;
  assign y20055 = ~1'b0 ;
  assign y20056 = 1'b0 ;
  assign y20057 = n31582 ;
  assign y20058 = n31583 ;
  assign y20059 = n31586 ;
  assign y20060 = ~1'b0 ;
  assign y20061 = ~1'b0 ;
  assign y20062 = ~1'b0 ;
  assign y20063 = ~n31610 ;
  assign y20064 = 1'b0 ;
  assign y20065 = ~1'b0 ;
  assign y20066 = n31612 ;
  assign y20067 = ~n7888 ;
  assign y20068 = 1'b0 ;
  assign y20069 = ~1'b0 ;
  assign y20070 = ~1'b0 ;
  assign y20071 = ~1'b0 ;
  assign y20072 = n31615 ;
  assign y20073 = n31617 ;
  assign y20074 = ~n31618 ;
  assign y20075 = ~1'b0 ;
  assign y20076 = ~1'b0 ;
  assign y20077 = ~n31619 ;
  assign y20078 = n31620 ;
  assign y20079 = ~n31622 ;
  assign y20080 = ~n31626 ;
  assign y20081 = ~n14872 ;
  assign y20082 = ~1'b0 ;
  assign y20083 = n31628 ;
  assign y20084 = ~n31630 ;
  assign y20085 = ~1'b0 ;
  assign y20086 = ~1'b0 ;
  assign y20087 = n31631 ;
  assign y20088 = n31634 ;
  assign y20089 = ~n31635 ;
  assign y20090 = ~1'b0 ;
  assign y20091 = ~n2998 ;
  assign y20092 = ~n31640 ;
  assign y20093 = ~n3931 ;
  assign y20094 = n31642 ;
  assign y20095 = 1'b0 ;
  assign y20096 = ~1'b0 ;
  assign y20097 = n31643 ;
  assign y20098 = ~n31649 ;
  assign y20099 = ~1'b0 ;
  assign y20100 = ~n31653 ;
  assign y20101 = ~1'b0 ;
  assign y20102 = ~1'b0 ;
  assign y20103 = n31655 ;
  assign y20104 = ~n31657 ;
  assign y20105 = n31658 ;
  assign y20106 = ~1'b0 ;
  assign y20107 = ~1'b0 ;
  assign y20108 = ~1'b0 ;
  assign y20109 = n31659 ;
  assign y20110 = n31662 ;
  assign y20111 = n31663 ;
  assign y20112 = n31668 ;
  assign y20113 = ~1'b0 ;
  assign y20114 = ~n30202 ;
  assign y20115 = n31669 ;
  assign y20116 = n31670 ;
  assign y20117 = ~n31345 ;
  assign y20118 = n31672 ;
  assign y20119 = ~1'b0 ;
  assign y20120 = ~n31673 ;
  assign y20121 = ~1'b0 ;
  assign y20122 = ~n31676 ;
  assign y20123 = n31677 ;
  assign y20124 = ~n31680 ;
  assign y20125 = ~1'b0 ;
  assign y20126 = ~n31681 ;
  assign y20127 = ~1'b0 ;
  assign y20128 = n31683 ;
  assign y20129 = n31684 ;
  assign y20130 = ~n31687 ;
  assign y20131 = x155 ;
  assign y20132 = ~n31689 ;
  assign y20133 = n31691 ;
  assign y20134 = ~n31694 ;
  assign y20135 = ~1'b0 ;
  assign y20136 = ~n31696 ;
  assign y20137 = ~n31700 ;
  assign y20138 = ~n31702 ;
  assign y20139 = ~n3703 ;
  assign y20140 = ~n11448 ;
  assign y20141 = ~1'b0 ;
  assign y20142 = n31703 ;
  assign y20143 = ~n31708 ;
  assign y20144 = ~n31709 ;
  assign y20145 = ~n31710 ;
  assign y20146 = ~n27665 ;
  assign y20147 = ~n31713 ;
  assign y20148 = ~1'b0 ;
  assign y20149 = n31714 ;
  assign y20150 = ~1'b0 ;
  assign y20151 = n31717 ;
  assign y20152 = n31718 ;
  assign y20153 = n10806 ;
  assign y20154 = ~1'b0 ;
  assign y20155 = n31719 ;
  assign y20156 = ~1'b0 ;
  assign y20157 = n31720 ;
  assign y20158 = ~1'b0 ;
  assign y20159 = ~1'b0 ;
  assign y20160 = ~1'b0 ;
  assign y20161 = ~1'b0 ;
  assign y20162 = ~1'b0 ;
  assign y20163 = 1'b0 ;
  assign y20164 = ~n31721 ;
  assign y20165 = n31722 ;
  assign y20166 = ~n31723 ;
  assign y20167 = ~1'b0 ;
  assign y20168 = ~n31726 ;
  assign y20169 = ~1'b0 ;
  assign y20170 = n31727 ;
  assign y20171 = ~n31729 ;
  assign y20172 = ~n31730 ;
  assign y20173 = n31731 ;
  assign y20174 = ~n31732 ;
  assign y20175 = ~n31734 ;
  assign y20176 = ~1'b0 ;
  assign y20177 = ~1'b0 ;
  assign y20178 = ~1'b0 ;
  assign y20179 = n10292 ;
  assign y20180 = n31735 ;
  assign y20181 = ~n31736 ;
  assign y20182 = ~1'b0 ;
  assign y20183 = n31738 ;
  assign y20184 = ~1'b0 ;
  assign y20185 = n31745 ;
  assign y20186 = n31746 ;
  assign y20187 = ~n31750 ;
  assign y20188 = ~1'b0 ;
  assign y20189 = 1'b0 ;
  assign y20190 = n31754 ;
  assign y20191 = ~n31756 ;
  assign y20192 = ~n31759 ;
  assign y20193 = ~n2977 ;
  assign y20194 = n31760 ;
  assign y20195 = n31762 ;
  assign y20196 = n31766 ;
  assign y20197 = ~n31767 ;
  assign y20198 = ~1'b0 ;
  assign y20199 = n31772 ;
  assign y20200 = n31777 ;
  assign y20201 = n31782 ;
  assign y20202 = ~n31783 ;
  assign y20203 = n31789 ;
  assign y20204 = ~1'b0 ;
  assign y20205 = ~n31791 ;
  assign y20206 = ~n31792 ;
  assign y20207 = ~1'b0 ;
  assign y20208 = ~n31794 ;
  assign y20209 = ~n31804 ;
  assign y20210 = n31805 ;
  assign y20211 = ~1'b0 ;
  assign y20212 = ~n31808 ;
  assign y20213 = ~1'b0 ;
  assign y20214 = n31810 ;
  assign y20215 = n31817 ;
  assign y20216 = ~1'b0 ;
  assign y20217 = n31820 ;
  assign y20218 = ~1'b0 ;
  assign y20219 = n31821 ;
  assign y20220 = ~n31823 ;
  assign y20221 = ~1'b0 ;
  assign y20222 = n31144 ;
  assign y20223 = ~n31825 ;
  assign y20224 = n31827 ;
  assign y20225 = ~1'b0 ;
  assign y20226 = ~n31832 ;
  assign y20227 = n31835 ;
  assign y20228 = n31838 ;
  assign y20229 = ~n31841 ;
  assign y20230 = ~n31844 ;
  assign y20231 = ~1'b0 ;
  assign y20232 = ~n31847 ;
  assign y20233 = ~n23959 ;
  assign y20234 = ~1'b0 ;
  assign y20235 = ~n31851 ;
  assign y20236 = ~n10834 ;
  assign y20237 = ~1'b0 ;
  assign y20238 = n31853 ;
  assign y20239 = ~1'b0 ;
  assign y20240 = ~1'b0 ;
  assign y20241 = ~n31854 ;
  assign y20242 = ~n31855 ;
  assign y20243 = ~n31856 ;
  assign y20244 = ~1'b0 ;
  assign y20245 = ~n31858 ;
  assign y20246 = ~1'b0 ;
  assign y20247 = ~n20676 ;
  assign y20248 = n31862 ;
  assign y20249 = ~1'b0 ;
  assign y20250 = n1014 ;
  assign y20251 = n31865 ;
  assign y20252 = ~n31869 ;
  assign y20253 = ~n20396 ;
  assign y20254 = ~n31870 ;
  assign y20255 = ~1'b0 ;
  assign y20256 = n31872 ;
  assign y20257 = ~n31873 ;
  assign y20258 = ~n31875 ;
  assign y20259 = ~1'b0 ;
  assign y20260 = ~1'b0 ;
  assign y20261 = ~1'b0 ;
  assign y20262 = ~1'b0 ;
  assign y20263 = n18552 ;
  assign y20264 = ~1'b0 ;
  assign y20265 = n31876 ;
  assign y20266 = ~n31877 ;
  assign y20267 = ~n1139 ;
  assign y20268 = ~1'b0 ;
  assign y20269 = ~1'b0 ;
  assign y20270 = ~n31880 ;
  assign y20271 = ~n4319 ;
  assign y20272 = ~n31882 ;
  assign y20273 = ~n31886 ;
  assign y20274 = ~n31887 ;
  assign y20275 = ~n31890 ;
  assign y20276 = ~1'b0 ;
  assign y20277 = n31892 ;
  assign y20278 = ~n31893 ;
  assign y20279 = ~n31895 ;
  assign y20280 = ~n31896 ;
  assign y20281 = ~n31898 ;
  assign y20282 = ~n4375 ;
  assign y20283 = ~1'b0 ;
  assign y20284 = ~1'b0 ;
  assign y20285 = ~1'b0 ;
  assign y20286 = ~n31899 ;
  assign y20287 = n31900 ;
  assign y20288 = ~1'b0 ;
  assign y20289 = ~n31902 ;
  assign y20290 = ~n31904 ;
  assign y20291 = ~n31909 ;
  assign y20292 = n31911 ;
  assign y20293 = n31913 ;
  assign y20294 = ~1'b0 ;
  assign y20295 = ~n31914 ;
  assign y20296 = ~n31916 ;
  assign y20297 = n31919 ;
  assign y20298 = n31920 ;
  assign y20299 = ~n4295 ;
  assign y20300 = n31924 ;
  assign y20301 = ~1'b0 ;
  assign y20302 = ~1'b0 ;
  assign y20303 = ~1'b0 ;
  assign y20304 = ~1'b0 ;
  assign y20305 = ~n31925 ;
  assign y20306 = ~1'b0 ;
  assign y20307 = n31926 ;
  assign y20308 = ~1'b0 ;
  assign y20309 = ~n31927 ;
  assign y20310 = ~1'b0 ;
  assign y20311 = n31932 ;
  assign y20312 = ~n31937 ;
  assign y20313 = ~n31941 ;
  assign y20314 = ~1'b0 ;
  assign y20315 = ~1'b0 ;
  assign y20316 = ~1'b0 ;
  assign y20317 = ~n15292 ;
  assign y20318 = n31942 ;
  assign y20319 = n31943 ;
  assign y20320 = ~n31945 ;
  assign y20321 = n31946 ;
  assign y20322 = n31947 ;
  assign y20323 = ~1'b0 ;
  assign y20324 = 1'b0 ;
  assign y20325 = n31949 ;
  assign y20326 = ~1'b0 ;
  assign y20327 = n31950 ;
  assign y20328 = ~n31952 ;
  assign y20329 = ~1'b0 ;
  assign y20330 = n31956 ;
  assign y20331 = n31958 ;
  assign y20332 = n14069 ;
  assign y20333 = ~1'b0 ;
  assign y20334 = ~n24139 ;
  assign y20335 = n31960 ;
  assign y20336 = n31962 ;
  assign y20337 = ~1'b0 ;
  assign y20338 = ~n31964 ;
  assign y20339 = ~n31968 ;
  assign y20340 = n31969 ;
  assign y20341 = n31971 ;
  assign y20342 = n7851 ;
  assign y20343 = ~1'b0 ;
  assign y20344 = n27784 ;
  assign y20345 = ~1'b0 ;
  assign y20346 = ~1'b0 ;
  assign y20347 = ~1'b0 ;
  assign y20348 = ~1'b0 ;
  assign y20349 = ~n31972 ;
  assign y20350 = n13479 ;
  assign y20351 = ~1'b0 ;
  assign y20352 = n31973 ;
  assign y20353 = n31974 ;
  assign y20354 = n31976 ;
  assign y20355 = ~1'b0 ;
  assign y20356 = ~n27010 ;
  assign y20357 = n31983 ;
  assign y20358 = ~1'b0 ;
  assign y20359 = ~1'b0 ;
  assign y20360 = ~1'b0 ;
  assign y20361 = n31984 ;
  assign y20362 = n31989 ;
  assign y20363 = 1'b0 ;
  assign y20364 = ~n31992 ;
  assign y20365 = ~1'b0 ;
  assign y20366 = ~n28702 ;
  assign y20367 = ~1'b0 ;
  assign y20368 = ~n15423 ;
  assign y20369 = 1'b0 ;
  assign y20370 = ~1'b0 ;
  assign y20371 = ~n22993 ;
  assign y20372 = ~1'b0 ;
  assign y20373 = ~n31994 ;
  assign y20374 = ~n31995 ;
  assign y20375 = n32000 ;
  assign y20376 = ~1'b0 ;
  assign y20377 = n32003 ;
  assign y20378 = ~1'b0 ;
  assign y20379 = n32004 ;
  assign y20380 = n21055 ;
  assign y20381 = ~n32006 ;
  assign y20382 = n32007 ;
  assign y20383 = n32008 ;
  assign y20384 = ~1'b0 ;
  assign y20385 = ~1'b0 ;
  assign y20386 = ~1'b0 ;
  assign y20387 = ~1'b0 ;
  assign y20388 = ~n17591 ;
  assign y20389 = n32010 ;
  assign y20390 = n32013 ;
  assign y20391 = n32014 ;
  assign y20392 = ~1'b0 ;
  assign y20393 = ~n32015 ;
  assign y20394 = ~n32016 ;
  assign y20395 = ~n32017 ;
  assign y20396 = ~1'b0 ;
  assign y20397 = ~1'b0 ;
  assign y20398 = ~1'b0 ;
  assign y20399 = n32018 ;
  assign y20400 = ~n32021 ;
  assign y20401 = n32022 ;
  assign y20402 = ~1'b0 ;
  assign y20403 = ~1'b0 ;
  assign y20404 = n32026 ;
  assign y20405 = n14871 ;
  assign y20406 = ~1'b0 ;
  assign y20407 = ~1'b0 ;
  assign y20408 = n19841 ;
  assign y20409 = n32027 ;
  assign y20410 = ~n32028 ;
  assign y20411 = ~1'b0 ;
  assign y20412 = ~n32031 ;
  assign y20413 = ~n32038 ;
  assign y20414 = ~1'b0 ;
  assign y20415 = 1'b0 ;
  assign y20416 = n32040 ;
  assign y20417 = n15411 ;
  assign y20418 = ~1'b0 ;
  assign y20419 = ~1'b0 ;
  assign y20420 = ~1'b0 ;
  assign y20421 = ~1'b0 ;
  assign y20422 = ~n32041 ;
  assign y20423 = ~n32042 ;
  assign y20424 = 1'b0 ;
  assign y20425 = ~n17109 ;
  assign y20426 = ~n32043 ;
  assign y20427 = ~n32047 ;
  assign y20428 = 1'b0 ;
  assign y20429 = ~1'b0 ;
  assign y20430 = ~1'b0 ;
  assign y20431 = n32049 ;
  assign y20432 = ~1'b0 ;
  assign y20433 = ~n32051 ;
  assign y20434 = ~n29285 ;
  assign y20435 = ~1'b0 ;
  assign y20436 = ~1'b0 ;
  assign y20437 = ~n32057 ;
  assign y20438 = ~n10116 ;
  assign y20439 = ~1'b0 ;
  assign y20440 = n32058 ;
  assign y20441 = ~n32059 ;
  assign y20442 = ~1'b0 ;
  assign y20443 = n17789 ;
  assign y20444 = n16797 ;
  assign y20445 = n32062 ;
  assign y20446 = ~n32066 ;
  assign y20447 = n32067 ;
  assign y20448 = n32068 ;
  assign y20449 = ~n32069 ;
  assign y20450 = ~1'b0 ;
  assign y20451 = n3181 ;
  assign y20452 = ~1'b0 ;
  assign y20453 = ~1'b0 ;
  assign y20454 = ~n32072 ;
  assign y20455 = n32073 ;
  assign y20456 = ~1'b0 ;
  assign y20457 = ~1'b0 ;
  assign y20458 = ~1'b0 ;
  assign y20459 = n32076 ;
  assign y20460 = 1'b0 ;
  assign y20461 = n32078 ;
  assign y20462 = n32080 ;
  assign y20463 = ~1'b0 ;
  assign y20464 = ~n32082 ;
  assign y20465 = n32083 ;
  assign y20466 = n305 ;
  assign y20467 = ~n32084 ;
  assign y20468 = n32087 ;
  assign y20469 = ~n32089 ;
  assign y20470 = n32090 ;
  assign y20471 = ~n32091 ;
  assign y20472 = ~n32092 ;
  assign y20473 = n32093 ;
  assign y20474 = ~n32094 ;
  assign y20475 = n32095 ;
  assign y20476 = 1'b0 ;
  assign y20477 = 1'b0 ;
  assign y20478 = ~1'b0 ;
  assign y20479 = ~1'b0 ;
  assign y20480 = ~n32099 ;
  assign y20481 = ~n32103 ;
  assign y20482 = n32105 ;
  assign y20483 = 1'b0 ;
  assign y20484 = n32107 ;
  assign y20485 = ~n7234 ;
  assign y20486 = ~n32109 ;
  assign y20487 = n32111 ;
  assign y20488 = n20256 ;
  assign y20489 = n32114 ;
  assign y20490 = ~1'b0 ;
  assign y20491 = n32116 ;
  assign y20492 = ~1'b0 ;
  assign y20493 = n32117 ;
  assign y20494 = n32118 ;
  assign y20495 = ~1'b0 ;
  assign y20496 = ~1'b0 ;
  assign y20497 = n32119 ;
  assign y20498 = ~1'b0 ;
  assign y20499 = n32120 ;
  assign y20500 = n4582 ;
  assign y20501 = n32121 ;
  assign y20502 = n32123 ;
  assign y20503 = n32130 ;
  assign y20504 = ~n32132 ;
  assign y20505 = ~n7508 ;
  assign y20506 = ~n32133 ;
  assign y20507 = n32136 ;
  assign y20508 = ~n32138 ;
  assign y20509 = ~n32143 ;
  assign y20510 = ~n32148 ;
  assign y20511 = ~n32149 ;
  assign y20512 = n29368 ;
  assign y20513 = ~1'b0 ;
  assign y20514 = ~1'b0 ;
  assign y20515 = ~1'b0 ;
  assign y20516 = ~n32150 ;
  assign y20517 = ~n32152 ;
  assign y20518 = n32154 ;
  assign y20519 = ~n32158 ;
  assign y20520 = ~n32163 ;
  assign y20521 = ~n32169 ;
  assign y20522 = ~n32171 ;
  assign y20523 = ~n32173 ;
  assign y20524 = n32174 ;
  assign y20525 = n32175 ;
  assign y20526 = ~1'b0 ;
  assign y20527 = ~1'b0 ;
  assign y20528 = n6473 ;
  assign y20529 = ~1'b0 ;
  assign y20530 = ~1'b0 ;
  assign y20531 = n20393 ;
  assign y20532 = ~1'b0 ;
  assign y20533 = ~n32176 ;
  assign y20534 = ~n32177 ;
  assign y20535 = n32178 ;
  assign y20536 = n32179 ;
  assign y20537 = n32182 ;
  assign y20538 = ~n7951 ;
  assign y20539 = ~n3473 ;
  assign y20540 = n32183 ;
  assign y20541 = ~n32184 ;
  assign y20542 = ~1'b0 ;
  assign y20543 = ~n32188 ;
  assign y20544 = ~n32192 ;
  assign y20545 = n32195 ;
  assign y20546 = ~n32196 ;
  assign y20547 = n32201 ;
  assign y20548 = n32203 ;
  assign y20549 = ~n32205 ;
  assign y20550 = ~n32206 ;
  assign y20551 = ~1'b0 ;
  assign y20552 = ~1'b0 ;
  assign y20553 = n32210 ;
  assign y20554 = ~1'b0 ;
  assign y20555 = n32213 ;
  assign y20556 = n32215 ;
  assign y20557 = ~n32217 ;
  assign y20558 = ~1'b0 ;
  assign y20559 = ~n32218 ;
  assign y20560 = 1'b0 ;
  assign y20561 = ~n32219 ;
  assign y20562 = ~1'b0 ;
  assign y20563 = ~n32220 ;
  assign y20564 = n26049 ;
  assign y20565 = ~1'b0 ;
  assign y20566 = n32225 ;
  assign y20567 = ~1'b0 ;
  assign y20568 = n32226 ;
  assign y20569 = n32234 ;
  assign y20570 = ~1'b0 ;
  assign y20571 = 1'b0 ;
  assign y20572 = n32236 ;
  assign y20573 = ~n13589 ;
  assign y20574 = ~1'b0 ;
  assign y20575 = ~n32238 ;
  assign y20576 = ~n32251 ;
  assign y20577 = n32253 ;
  assign y20578 = ~1'b0 ;
  assign y20579 = ~n32255 ;
  assign y20580 = ~n32259 ;
  assign y20581 = ~n32261 ;
  assign y20582 = ~1'b0 ;
  assign y20583 = ~1'b0 ;
  assign y20584 = ~n32265 ;
  assign y20585 = ~n14485 ;
  assign y20586 = ~1'b0 ;
  assign y20587 = n32267 ;
  assign y20588 = n32268 ;
  assign y20589 = ~1'b0 ;
  assign y20590 = ~n32270 ;
  assign y20591 = ~1'b0 ;
  assign y20592 = ~n32272 ;
  assign y20593 = ~n32275 ;
  assign y20594 = ~n32276 ;
  assign y20595 = n32277 ;
  assign y20596 = ~n13066 ;
  assign y20597 = n32279 ;
  assign y20598 = ~n32280 ;
  assign y20599 = n32281 ;
  assign y20600 = ~n32283 ;
  assign y20601 = ~1'b0 ;
  assign y20602 = n32284 ;
  assign y20603 = ~n32287 ;
  assign y20604 = ~1'b0 ;
  assign y20605 = ~1'b0 ;
  assign y20606 = ~1'b0 ;
  assign y20607 = n32290 ;
  assign y20608 = ~1'b0 ;
  assign y20609 = n32291 ;
  assign y20610 = ~n8448 ;
  assign y20611 = n32297 ;
  assign y20612 = ~n32301 ;
  assign y20613 = ~n32305 ;
  assign y20614 = ~n27249 ;
  assign y20615 = ~n32307 ;
  assign y20616 = ~n32311 ;
  assign y20617 = n32313 ;
  assign y20618 = ~n32315 ;
  assign y20619 = ~1'b0 ;
  assign y20620 = ~1'b0 ;
  assign y20621 = n32317 ;
  assign y20622 = n32320 ;
  assign y20623 = n32323 ;
  assign y20624 = ~1'b0 ;
  assign y20625 = ~n32335 ;
  assign y20626 = n32336 ;
  assign y20627 = ~n32339 ;
  assign y20628 = 1'b0 ;
  assign y20629 = n32340 ;
  assign y20630 = ~1'b0 ;
  assign y20631 = ~n32341 ;
  assign y20632 = ~n32349 ;
  assign y20633 = n32353 ;
  assign y20634 = 1'b0 ;
  assign y20635 = n32356 ;
  assign y20636 = ~n32358 ;
  assign y20637 = ~1'b0 ;
  assign y20638 = ~1'b0 ;
  assign y20639 = ~n32360 ;
  assign y20640 = ~n32364 ;
  assign y20641 = ~n32366 ;
  assign y20642 = ~n32367 ;
  assign y20643 = n32369 ;
  assign y20644 = ~n32370 ;
  assign y20645 = ~1'b0 ;
  assign y20646 = ~n32372 ;
  assign y20647 = ~n32374 ;
  assign y20648 = ~1'b0 ;
  assign y20649 = ~1'b0 ;
  assign y20650 = ~n32376 ;
  assign y20651 = ~n32378 ;
  assign y20652 = ~n32380 ;
  assign y20653 = ~n32382 ;
  assign y20654 = ~1'b0 ;
  assign y20655 = ~n32386 ;
  assign y20656 = ~1'b0 ;
  assign y20657 = ~1'b0 ;
  assign y20658 = n32387 ;
  assign y20659 = 1'b0 ;
  assign y20660 = ~1'b0 ;
  assign y20661 = n32388 ;
  assign y20662 = n32390 ;
  assign y20663 = ~1'b0 ;
  assign y20664 = n32391 ;
  assign y20665 = ~n32392 ;
  assign y20666 = n32393 ;
  assign y20667 = ~n13134 ;
  assign y20668 = n32395 ;
  assign y20669 = ~n32396 ;
  assign y20670 = ~n32398 ;
  assign y20671 = ~n32407 ;
  assign y20672 = ~n32409 ;
  assign y20673 = ~1'b0 ;
  assign y20674 = ~1'b0 ;
  assign y20675 = ~n32416 ;
  assign y20676 = n32418 ;
  assign y20677 = ~n27062 ;
  assign y20678 = ~1'b0 ;
  assign y20679 = ~n32419 ;
  assign y20680 = n32421 ;
  assign y20681 = ~n32422 ;
  assign y20682 = ~n13871 ;
  assign y20683 = ~n12769 ;
  assign y20684 = ~n32424 ;
  assign y20685 = n32426 ;
  assign y20686 = ~1'b0 ;
  assign y20687 = n32428 ;
  assign y20688 = ~n32430 ;
  assign y20689 = n32431 ;
  assign y20690 = ~n32436 ;
  assign y20691 = n13761 ;
  assign y20692 = ~1'b0 ;
  assign y20693 = ~n32438 ;
  assign y20694 = ~1'b0 ;
  assign y20695 = 1'b0 ;
  assign y20696 = n32439 ;
  assign y20697 = n32440 ;
  assign y20698 = ~1'b0 ;
  assign y20699 = 1'b0 ;
  assign y20700 = ~n32443 ;
  assign y20701 = ~1'b0 ;
  assign y20702 = n32452 ;
  assign y20703 = ~1'b0 ;
  assign y20704 = n32456 ;
  assign y20705 = ~n32457 ;
  assign y20706 = n32458 ;
  assign y20707 = ~1'b0 ;
  assign y20708 = ~1'b0 ;
  assign y20709 = ~n32463 ;
  assign y20710 = n32466 ;
  assign y20711 = ~1'b0 ;
  assign y20712 = ~n32469 ;
  assign y20713 = ~n32471 ;
  assign y20714 = n32473 ;
  assign y20715 = ~1'b0 ;
  assign y20716 = ~1'b0 ;
  assign y20717 = ~1'b0 ;
  assign y20718 = n32477 ;
  assign y20719 = n32481 ;
  assign y20720 = n32482 ;
  assign y20721 = ~1'b0 ;
  assign y20722 = 1'b0 ;
  assign y20723 = ~1'b0 ;
  assign y20724 = n32484 ;
  assign y20725 = ~1'b0 ;
  assign y20726 = ~1'b0 ;
  assign y20727 = ~n32487 ;
  assign y20728 = ~1'b0 ;
  assign y20729 = ~1'b0 ;
  assign y20730 = ~n32488 ;
  assign y20731 = ~n5783 ;
  assign y20732 = n1761 ;
  assign y20733 = ~1'b0 ;
  assign y20734 = ~n32492 ;
  assign y20735 = n32493 ;
  assign y20736 = ~1'b0 ;
  assign y20737 = ~1'b0 ;
  assign y20738 = n9321 ;
  assign y20739 = ~n32495 ;
  assign y20740 = ~n32499 ;
  assign y20741 = n32501 ;
  assign y20742 = n32502 ;
  assign y20743 = n32504 ;
  assign y20744 = ~n32507 ;
  assign y20745 = ~n32513 ;
  assign y20746 = n32516 ;
  assign y20747 = ~1'b0 ;
  assign y20748 = ~n32518 ;
  assign y20749 = n32520 ;
  assign y20750 = n32521 ;
  assign y20751 = ~n32525 ;
  assign y20752 = ~1'b0 ;
  assign y20753 = ~n32528 ;
  assign y20754 = ~1'b0 ;
  assign y20755 = n32529 ;
  assign y20756 = 1'b0 ;
  assign y20757 = n32534 ;
  assign y20758 = n32535 ;
  assign y20759 = ~1'b0 ;
  assign y20760 = n32537 ;
  assign y20761 = ~n32540 ;
  assign y20762 = ~1'b0 ;
  assign y20763 = ~n32541 ;
  assign y20764 = ~n32545 ;
  assign y20765 = ~n32552 ;
  assign y20766 = n32553 ;
  assign y20767 = ~n14424 ;
  assign y20768 = n32554 ;
  assign y20769 = ~1'b0 ;
  assign y20770 = ~1'b0 ;
  assign y20771 = ~1'b0 ;
  assign y20772 = n32555 ;
  assign y20773 = n32556 ;
  assign y20774 = ~1'b0 ;
  assign y20775 = ~n32557 ;
  assign y20776 = ~1'b0 ;
  assign y20777 = ~n32558 ;
  assign y20778 = ~n5918 ;
  assign y20779 = n6158 ;
  assign y20780 = ~n32559 ;
  assign y20781 = n32560 ;
  assign y20782 = ~1'b0 ;
  assign y20783 = ~1'b0 ;
  assign y20784 = ~n32561 ;
  assign y20785 = n32565 ;
  assign y20786 = ~n32567 ;
  assign y20787 = n32569 ;
  assign y20788 = n32572 ;
  assign y20789 = ~n2921 ;
  assign y20790 = ~1'b0 ;
  assign y20791 = ~n32575 ;
  assign y20792 = ~n32576 ;
  assign y20793 = ~n32577 ;
  assign y20794 = ~1'b0 ;
  assign y20795 = n32578 ;
  assign y20796 = ~1'b0 ;
  assign y20797 = 1'b0 ;
  assign y20798 = ~1'b0 ;
  assign y20799 = ~n30470 ;
  assign y20800 = n32579 ;
  assign y20801 = ~n9179 ;
  assign y20802 = ~1'b0 ;
  assign y20803 = n32580 ;
  assign y20804 = n32582 ;
  assign y20805 = n32585 ;
  assign y20806 = ~n4204 ;
  assign y20807 = ~n12238 ;
  assign y20808 = ~n32586 ;
  assign y20809 = n24404 ;
  assign y20810 = ~n32587 ;
  assign y20811 = ~1'b0 ;
  assign y20812 = ~n32590 ;
  assign y20813 = n32591 ;
  assign y20814 = n32595 ;
  assign y20815 = n32598 ;
  assign y20816 = ~1'b0 ;
  assign y20817 = n13708 ;
  assign y20818 = ~1'b0 ;
  assign y20819 = n32599 ;
  assign y20820 = ~1'b0 ;
  assign y20821 = ~n32607 ;
  assign y20822 = ~n32608 ;
  assign y20823 = 1'b0 ;
  assign y20824 = n32609 ;
  assign y20825 = n32611 ;
  assign y20826 = ~n6300 ;
  assign y20827 = n32613 ;
  assign y20828 = ~1'b0 ;
  assign y20829 = ~n32615 ;
  assign y20830 = ~1'b0 ;
  assign y20831 = n3625 ;
  assign y20832 = ~n32617 ;
  assign y20833 = n28684 ;
  assign y20834 = ~1'b0 ;
  assign y20835 = ~1'b0 ;
  assign y20836 = ~n32623 ;
  assign y20837 = ~n32624 ;
  assign y20838 = n32626 ;
  assign y20839 = ~n32627 ;
  assign y20840 = n31838 ;
  assign y20841 = n2042 ;
  assign y20842 = n23010 ;
  assign y20843 = ~1'b0 ;
  assign y20844 = ~n32630 ;
  assign y20845 = ~n32639 ;
  assign y20846 = n32642 ;
  assign y20847 = ~n32645 ;
  assign y20848 = n32647 ;
  assign y20849 = ~n32649 ;
  assign y20850 = ~n32650 ;
  assign y20851 = n32651 ;
  assign y20852 = ~1'b0 ;
  assign y20853 = n32652 ;
  assign y20854 = ~1'b0 ;
  assign y20855 = ~1'b0 ;
  assign y20856 = ~n32653 ;
  assign y20857 = ~n32654 ;
  assign y20858 = ~n32657 ;
  assign y20859 = ~1'b0 ;
  assign y20860 = ~n32660 ;
  assign y20861 = ~n32661 ;
  assign y20862 = ~n32662 ;
  assign y20863 = n32664 ;
  assign y20864 = ~1'b0 ;
  assign y20865 = n32667 ;
  assign y20866 = n32670 ;
  assign y20867 = n32674 ;
  assign y20868 = ~1'b0 ;
  assign y20869 = ~1'b0 ;
  assign y20870 = n32675 ;
  assign y20871 = n32678 ;
  assign y20872 = ~n32679 ;
  assign y20873 = ~n19165 ;
  assign y20874 = ~n32682 ;
  assign y20875 = ~1'b0 ;
  assign y20876 = n12496 ;
  assign y20877 = ~n32684 ;
  assign y20878 = ~n32685 ;
  assign y20879 = ~1'b0 ;
  assign y20880 = ~1'b0 ;
  assign y20881 = ~n32686 ;
  assign y20882 = ~n32691 ;
  assign y20883 = ~n32693 ;
  assign y20884 = n32694 ;
  assign y20885 = ~1'b0 ;
  assign y20886 = ~n21675 ;
  assign y20887 = 1'b0 ;
  assign y20888 = n32695 ;
  assign y20889 = ~n32710 ;
  assign y20890 = 1'b0 ;
  assign y20891 = ~1'b0 ;
  assign y20892 = n14089 ;
  assign y20893 = ~1'b0 ;
  assign y20894 = ~1'b0 ;
  assign y20895 = ~n32713 ;
  assign y20896 = ~1'b0 ;
  assign y20897 = ~1'b0 ;
  assign y20898 = ~n32715 ;
  assign y20899 = n32716 ;
  assign y20900 = n13995 ;
  assign y20901 = ~n14487 ;
  assign y20902 = 1'b0 ;
  assign y20903 = n32719 ;
  assign y20904 = ~1'b0 ;
  assign y20905 = ~n32720 ;
  assign y20906 = ~n32721 ;
  assign y20907 = ~1'b0 ;
  assign y20908 = ~n32724 ;
  assign y20909 = ~n32728 ;
  assign y20910 = ~n32731 ;
  assign y20911 = ~n32732 ;
  assign y20912 = ~n32733 ;
  assign y20913 = ~1'b0 ;
  assign y20914 = ~n32734 ;
  assign y20915 = 1'b0 ;
  assign y20916 = ~n32739 ;
  assign y20917 = ~n32741 ;
  assign y20918 = n32744 ;
  assign y20919 = n32746 ;
  assign y20920 = n32748 ;
  assign y20921 = ~1'b0 ;
  assign y20922 = ~1'b0 ;
  assign y20923 = ~n32750 ;
  assign y20924 = ~n32752 ;
  assign y20925 = ~1'b0 ;
  assign y20926 = ~n32756 ;
  assign y20927 = ~n32758 ;
  assign y20928 = n32759 ;
  assign y20929 = n32761 ;
  assign y20930 = ~1'b0 ;
  assign y20931 = ~1'b0 ;
  assign y20932 = n32762 ;
  assign y20933 = n10075 ;
  assign y20934 = ~n10086 ;
  assign y20935 = n32764 ;
  assign y20936 = n32767 ;
  assign y20937 = 1'b0 ;
  assign y20938 = ~n32769 ;
  assign y20939 = ~n32780 ;
  assign y20940 = ~1'b0 ;
  assign y20941 = ~n32781 ;
  assign y20942 = ~1'b0 ;
  assign y20943 = ~n32786 ;
  assign y20944 = ~n2678 ;
  assign y20945 = ~n32787 ;
  assign y20946 = ~1'b0 ;
  assign y20947 = ~n32791 ;
  assign y20948 = ~1'b0 ;
  assign y20949 = ~n1389 ;
  assign y20950 = n32794 ;
  assign y20951 = ~1'b0 ;
  assign y20952 = n26374 ;
  assign y20953 = ~n32796 ;
  assign y20954 = n32797 ;
  assign y20955 = n3832 ;
  assign y20956 = ~n32798 ;
  assign y20957 = n28175 ;
  assign y20958 = ~1'b0 ;
  assign y20959 = ~n32800 ;
  assign y20960 = n32802 ;
  assign y20961 = ~n32807 ;
  assign y20962 = n32810 ;
  assign y20963 = ~n32817 ;
  assign y20964 = ~n32818 ;
  assign y20965 = n27253 ;
  assign y20966 = 1'b0 ;
  assign y20967 = n32820 ;
  assign y20968 = n32822 ;
  assign y20969 = ~n32823 ;
  assign y20970 = n20820 ;
  assign y20971 = ~1'b0 ;
  assign y20972 = n32826 ;
  assign y20973 = ~n32828 ;
  assign y20974 = ~n32829 ;
  assign y20975 = ~1'b0 ;
  assign y20976 = ~1'b0 ;
  assign y20977 = ~n32830 ;
  assign y20978 = ~n29386 ;
  assign y20979 = ~1'b0 ;
  assign y20980 = ~n32834 ;
  assign y20981 = ~n32835 ;
  assign y20982 = ~n32837 ;
  assign y20983 = n21666 ;
  assign y20984 = ~1'b0 ;
  assign y20985 = ~1'b0 ;
  assign y20986 = ~1'b0 ;
  assign y20987 = n32838 ;
  assign y20988 = ~n32840 ;
  assign y20989 = n32842 ;
  assign y20990 = ~n32843 ;
  assign y20991 = ~n5506 ;
  assign y20992 = n32844 ;
  assign y20993 = ~n25872 ;
  assign y20994 = ~n32846 ;
  assign y20995 = ~n32849 ;
  assign y20996 = n32850 ;
  assign y20997 = ~1'b0 ;
  assign y20998 = ~n32852 ;
  assign y20999 = n32855 ;
  assign y21000 = ~n32858 ;
  assign y21001 = 1'b0 ;
  assign y21002 = ~1'b0 ;
  assign y21003 = n32860 ;
  assign y21004 = ~n32861 ;
  assign y21005 = ~n32865 ;
  assign y21006 = ~1'b0 ;
  assign y21007 = n32868 ;
  assign y21008 = ~n18095 ;
  assign y21009 = n32869 ;
  assign y21010 = ~1'b0 ;
  assign y21011 = ~1'b0 ;
  assign y21012 = ~1'b0 ;
  assign y21013 = ~n32871 ;
  assign y21014 = ~1'b0 ;
  assign y21015 = ~1'b0 ;
  assign y21016 = ~1'b0 ;
  assign y21017 = ~1'b0 ;
  assign y21018 = ~1'b0 ;
  assign y21019 = ~1'b0 ;
  assign y21020 = ~1'b0 ;
  assign y21021 = ~n32874 ;
  assign y21022 = ~1'b0 ;
  assign y21023 = n32877 ;
  assign y21024 = ~1'b0 ;
  assign y21025 = ~1'b0 ;
  assign y21026 = n32879 ;
  assign y21027 = ~n32881 ;
  assign y21028 = ~n32883 ;
  assign y21029 = ~n32884 ;
  assign y21030 = n32885 ;
  assign y21031 = ~n32892 ;
  assign y21032 = ~n32895 ;
  assign y21033 = ~1'b0 ;
  assign y21034 = ~n32896 ;
  assign y21035 = 1'b0 ;
  assign y21036 = ~1'b0 ;
  assign y21037 = ~n32898 ;
  assign y21038 = ~1'b0 ;
  assign y21039 = ~1'b0 ;
  assign y21040 = ~n32900 ;
  assign y21041 = n32904 ;
  assign y21042 = ~n32905 ;
  assign y21043 = ~n32907 ;
  assign y21044 = n32908 ;
  assign y21045 = n580 ;
  assign y21046 = ~1'b0 ;
  assign y21047 = ~1'b0 ;
  assign y21048 = n32910 ;
  assign y21049 = n32912 ;
  assign y21050 = ~n32913 ;
  assign y21051 = n32915 ;
  assign y21052 = n32916 ;
  assign y21053 = n32305 ;
  assign y21054 = ~1'b0 ;
  assign y21055 = ~1'b0 ;
  assign y21056 = ~1'b0 ;
  assign y21057 = n32928 ;
  assign y21058 = ~n32929 ;
  assign y21059 = ~1'b0 ;
  assign y21060 = ~n32931 ;
  assign y21061 = ~n32932 ;
  assign y21062 = ~n32935 ;
  assign y21063 = n32941 ;
  assign y21064 = ~n32944 ;
  assign y21065 = n32946 ;
  assign y21066 = ~1'b0 ;
  assign y21067 = n16768 ;
  assign y21068 = ~n32947 ;
  assign y21069 = ~n32950 ;
  assign y21070 = ~1'b0 ;
  assign y21071 = ~n32951 ;
  assign y21072 = ~n4111 ;
  assign y21073 = n32956 ;
  assign y21074 = ~n4851 ;
  assign y21075 = ~n9764 ;
  assign y21076 = n32957 ;
  assign y21077 = ~1'b0 ;
  assign y21078 = n15600 ;
  assign y21079 = ~n32958 ;
  assign y21080 = n32964 ;
  assign y21081 = ~n32965 ;
  assign y21082 = ~n32969 ;
  assign y21083 = ~1'b0 ;
  assign y21084 = ~1'b0 ;
  assign y21085 = n32973 ;
  assign y21086 = ~1'b0 ;
  assign y21087 = ~1'b0 ;
  assign y21088 = ~1'b0 ;
  assign y21089 = 1'b0 ;
  assign y21090 = ~n32974 ;
  assign y21091 = ~1'b0 ;
  assign y21092 = n2334 ;
  assign y21093 = ~n32975 ;
  assign y21094 = ~1'b0 ;
  assign y21095 = ~1'b0 ;
  assign y21096 = ~1'b0 ;
  assign y21097 = ~n32976 ;
  assign y21098 = ~n32979 ;
  assign y21099 = ~n32988 ;
  assign y21100 = 1'b0 ;
  assign y21101 = n32991 ;
  assign y21102 = n32995 ;
  assign y21103 = ~n33000 ;
  assign y21104 = n33001 ;
  assign y21105 = ~n33003 ;
  assign y21106 = ~1'b0 ;
  assign y21107 = ~1'b0 ;
  assign y21108 = ~1'b0 ;
  assign y21109 = n33006 ;
  assign y21110 = ~1'b0 ;
  assign y21111 = ~n33007 ;
  assign y21112 = ~1'b0 ;
  assign y21113 = ~1'b0 ;
  assign y21114 = ~n33009 ;
  assign y21115 = ~1'b0 ;
  assign y21116 = ~n33011 ;
  assign y21117 = ~n33014 ;
  assign y21118 = n33019 ;
  assign y21119 = n33020 ;
  assign y21120 = n14376 ;
  assign y21121 = ~1'b0 ;
  assign y21122 = ~1'b0 ;
  assign y21123 = ~n33027 ;
  assign y21124 = 1'b0 ;
  assign y21125 = 1'b0 ;
  assign y21126 = ~n12386 ;
  assign y21127 = ~n33028 ;
  assign y21128 = ~1'b0 ;
  assign y21129 = ~1'b0 ;
  assign y21130 = ~n7463 ;
  assign y21131 = n33030 ;
  assign y21132 = ~n33032 ;
  assign y21133 = n33033 ;
  assign y21134 = ~1'b0 ;
  assign y21135 = n25410 ;
  assign y21136 = ~n17004 ;
  assign y21137 = ~n33035 ;
  assign y21138 = ~n33037 ;
  assign y21139 = ~1'b0 ;
  assign y21140 = 1'b0 ;
  assign y21141 = ~1'b0 ;
  assign y21142 = n33038 ;
  assign y21143 = n33039 ;
  assign y21144 = n33042 ;
  assign y21145 = ~n33046 ;
  assign y21146 = ~n33050 ;
  assign y21147 = ~n12616 ;
  assign y21148 = ~1'b0 ;
  assign y21149 = ~n33053 ;
  assign y21150 = ~n33055 ;
  assign y21151 = ~1'b0 ;
  assign y21152 = n17372 ;
  assign y21153 = ~n33059 ;
  assign y21154 = ~n27571 ;
  assign y21155 = ~1'b0 ;
  assign y21156 = n17312 ;
  assign y21157 = n33060 ;
  assign y21158 = n33062 ;
  assign y21159 = ~n10087 ;
  assign y21160 = ~n8702 ;
  assign y21161 = ~1'b0 ;
  assign y21162 = n33063 ;
  assign y21163 = n33065 ;
  assign y21164 = ~1'b0 ;
  assign y21165 = ~n33066 ;
  assign y21166 = ~1'b0 ;
  assign y21167 = ~1'b0 ;
  assign y21168 = ~1'b0 ;
  assign y21169 = n33067 ;
  assign y21170 = ~n33068 ;
  assign y21171 = n3694 ;
  assign y21172 = n33069 ;
  assign y21173 = ~1'b0 ;
  assign y21174 = ~1'b0 ;
  assign y21175 = ~1'b0 ;
  assign y21176 = ~n33072 ;
  assign y21177 = n33073 ;
  assign y21178 = n28595 ;
  assign y21179 = ~1'b0 ;
  assign y21180 = n33074 ;
  assign y21181 = ~n3611 ;
  assign y21182 = ~1'b0 ;
  assign y21183 = ~n33075 ;
  assign y21184 = ~n33076 ;
  assign y21185 = ~1'b0 ;
  assign y21186 = n33078 ;
  assign y21187 = n33079 ;
  assign y21188 = ~n33081 ;
  assign y21189 = n3703 ;
  assign y21190 = ~1'b0 ;
  assign y21191 = ~n33082 ;
  assign y21192 = ~n33085 ;
  assign y21193 = ~1'b0 ;
  assign y21194 = n33086 ;
  assign y21195 = n33087 ;
  assign y21196 = ~1'b0 ;
  assign y21197 = ~1'b0 ;
  assign y21198 = ~n10684 ;
  assign y21199 = ~1'b0 ;
  assign y21200 = ~n33088 ;
  assign y21201 = ~n33090 ;
  assign y21202 = ~n33092 ;
  assign y21203 = ~1'b0 ;
  assign y21204 = ~n33095 ;
  assign y21205 = ~n33099 ;
  assign y21206 = n33100 ;
  assign y21207 = ~1'b0 ;
  assign y21208 = n33103 ;
  assign y21209 = ~n33104 ;
  assign y21210 = ~n33106 ;
  assign y21211 = 1'b0 ;
  assign y21212 = ~n33113 ;
  assign y21213 = n33117 ;
  assign y21214 = n33121 ;
  assign y21215 = n33125 ;
  assign y21216 = n33128 ;
  assign y21217 = n33129 ;
  assign y21218 = ~n33133 ;
  assign y21219 = ~n33134 ;
  assign y21220 = ~n33135 ;
  assign y21221 = ~1'b0 ;
  assign y21222 = ~n33137 ;
  assign y21223 = n12455 ;
  assign y21224 = ~1'b0 ;
  assign y21225 = ~1'b0 ;
  assign y21226 = ~n2806 ;
  assign y21227 = n33141 ;
  assign y21228 = ~1'b0 ;
  assign y21229 = n33142 ;
  assign y21230 = ~1'b0 ;
  assign y21231 = ~n33143 ;
  assign y21232 = ~1'b0 ;
  assign y21233 = ~1'b0 ;
  assign y21234 = ~1'b0 ;
  assign y21235 = n33145 ;
  assign y21236 = 1'b0 ;
  assign y21237 = ~1'b0 ;
  assign y21238 = n33147 ;
  assign y21239 = ~n33149 ;
  assign y21240 = ~n3850 ;
  assign y21241 = ~1'b0 ;
  assign y21242 = ~1'b0 ;
  assign y21243 = ~n33152 ;
  assign y21244 = ~1'b0 ;
  assign y21245 = ~1'b0 ;
  assign y21246 = ~n33153 ;
  assign y21247 = ~n33158 ;
  assign y21248 = n33159 ;
  assign y21249 = 1'b0 ;
  assign y21250 = ~n33165 ;
  assign y21251 = ~1'b0 ;
  assign y21252 = n7653 ;
  assign y21253 = n33169 ;
  assign y21254 = ~n3694 ;
  assign y21255 = n33171 ;
  assign y21256 = ~1'b0 ;
  assign y21257 = n33173 ;
  assign y21258 = n33177 ;
  assign y21259 = ~1'b0 ;
  assign y21260 = ~1'b0 ;
  assign y21261 = ~n22310 ;
  assign y21262 = ~1'b0 ;
  assign y21263 = n33181 ;
  assign y21264 = ~n33183 ;
  assign y21265 = ~1'b0 ;
  assign y21266 = n21209 ;
  assign y21267 = ~n33186 ;
  assign y21268 = n33191 ;
  assign y21269 = ~1'b0 ;
  assign y21270 = ~n33195 ;
  assign y21271 = n33198 ;
  assign y21272 = ~n33202 ;
  assign y21273 = ~1'b0 ;
  assign y21274 = ~n9854 ;
  assign y21275 = n33204 ;
  assign y21276 = n33207 ;
  assign y21277 = ~n33209 ;
  assign y21278 = ~n33210 ;
  assign y21279 = ~1'b0 ;
  assign y21280 = ~1'b0 ;
  assign y21281 = n33211 ;
  assign y21282 = ~n33215 ;
  assign y21283 = ~n33217 ;
  assign y21284 = ~1'b0 ;
  assign y21285 = ~1'b0 ;
  assign y21286 = ~1'b0 ;
  assign y21287 = n33219 ;
  assign y21288 = ~n33220 ;
  assign y21289 = n17936 ;
  assign y21290 = ~n33221 ;
  assign y21291 = ~1'b0 ;
  assign y21292 = ~1'b0 ;
  assign y21293 = n33223 ;
  assign y21294 = n33227 ;
  assign y21295 = n33232 ;
  assign y21296 = n33233 ;
  assign y21297 = ~1'b0 ;
  assign y21298 = n33235 ;
  assign y21299 = ~1'b0 ;
  assign y21300 = n33236 ;
  assign y21301 = n33241 ;
  assign y21302 = 1'b0 ;
  assign y21303 = ~n33243 ;
  assign y21304 = n33244 ;
  assign y21305 = ~1'b0 ;
  assign y21306 = n33245 ;
  assign y21307 = ~1'b0 ;
  assign y21308 = ~1'b0 ;
  assign y21309 = n33246 ;
  assign y21310 = n33250 ;
  assign y21311 = ~n33251 ;
  assign y21312 = ~n33252 ;
  assign y21313 = ~n33253 ;
  assign y21314 = n33256 ;
  assign y21315 = ~n33257 ;
  assign y21316 = n33262 ;
  assign y21317 = n33265 ;
  assign y21318 = ~n33269 ;
  assign y21319 = ~1'b0 ;
  assign y21320 = ~n33270 ;
  assign y21321 = ~n15328 ;
  assign y21322 = ~1'b0 ;
  assign y21323 = n33271 ;
  assign y21324 = n23162 ;
  assign y21325 = ~n33272 ;
  assign y21326 = n25535 ;
  assign y21327 = ~1'b0 ;
  assign y21328 = 1'b0 ;
  assign y21329 = ~n33274 ;
  assign y21330 = n33279 ;
  assign y21331 = ~1'b0 ;
  assign y21332 = ~1'b0 ;
  assign y21333 = n33280 ;
  assign y21334 = n33283 ;
  assign y21335 = ~1'b0 ;
  assign y21336 = ~n33285 ;
  assign y21337 = ~n33289 ;
  assign y21338 = n33290 ;
  assign y21339 = ~n33292 ;
  assign y21340 = ~1'b0 ;
  assign y21341 = n33293 ;
  assign y21342 = 1'b0 ;
  assign y21343 = ~1'b0 ;
  assign y21344 = ~n33294 ;
  assign y21345 = ~1'b0 ;
  assign y21346 = n5675 ;
  assign y21347 = n33295 ;
  assign y21348 = ~1'b0 ;
  assign y21349 = ~1'b0 ;
  assign y21350 = 1'b0 ;
  assign y21351 = n11241 ;
  assign y21352 = 1'b0 ;
  assign y21353 = 1'b0 ;
  assign y21354 = n33299 ;
  assign y21355 = n33302 ;
  assign y21356 = ~1'b0 ;
  assign y21357 = ~1'b0 ;
  assign y21358 = n33304 ;
  assign y21359 = ~1'b0 ;
  assign y21360 = n33306 ;
  assign y21361 = n33310 ;
  assign y21362 = n33313 ;
  assign y21363 = ~1'b0 ;
  assign y21364 = n33315 ;
  assign y21365 = ~1'b0 ;
  assign y21366 = n3521 ;
  assign y21367 = ~1'b0 ;
  assign y21368 = ~1'b0 ;
  assign y21369 = ~1'b0 ;
  assign y21370 = n33317 ;
  assign y21371 = ~1'b0 ;
  assign y21372 = n25793 ;
  assign y21373 = ~1'b0 ;
  assign y21374 = n19439 ;
  assign y21375 = ~1'b0 ;
  assign y21376 = ~1'b0 ;
  assign y21377 = ~n33319 ;
  assign y21378 = ~n33321 ;
  assign y21379 = ~1'b0 ;
  assign y21380 = ~1'b0 ;
  assign y21381 = ~1'b0 ;
  assign y21382 = ~n33322 ;
  assign y21383 = ~n33323 ;
  assign y21384 = ~1'b0 ;
  assign y21385 = ~1'b0 ;
  assign y21386 = ~1'b0 ;
  assign y21387 = n33327 ;
  assign y21388 = ~1'b0 ;
  assign y21389 = n33328 ;
  assign y21390 = ~n33330 ;
  assign y21391 = n33331 ;
  assign y21392 = ~1'b0 ;
  assign y21393 = ~1'b0 ;
  assign y21394 = ~n33332 ;
  assign y21395 = n7544 ;
  assign y21396 = ~1'b0 ;
  assign y21397 = ~1'b0 ;
  assign y21398 = n33336 ;
  assign y21399 = ~1'b0 ;
  assign y21400 = n33338 ;
  assign y21401 = n9947 ;
  assign y21402 = ~1'b0 ;
  assign y21403 = ~n33339 ;
  assign y21404 = ~n33340 ;
  assign y21405 = ~n21427 ;
  assign y21406 = ~1'b0 ;
  assign y21407 = n33341 ;
  assign y21408 = ~1'b0 ;
  assign y21409 = ~1'b0 ;
  assign y21410 = ~1'b0 ;
  assign y21411 = ~n33343 ;
  assign y21412 = n33346 ;
  assign y21413 = n3397 ;
  assign y21414 = ~n33347 ;
  assign y21415 = ~n33351 ;
  assign y21416 = ~n33354 ;
  assign y21417 = ~1'b0 ;
  assign y21418 = ~1'b0 ;
  assign y21419 = ~n33357 ;
  assign y21420 = ~n33359 ;
  assign y21421 = ~1'b0 ;
  assign y21422 = n33362 ;
  assign y21423 = 1'b0 ;
  assign y21424 = ~n33363 ;
  assign y21425 = ~n33364 ;
  assign y21426 = ~n33366 ;
  assign y21427 = ~n20616 ;
  assign y21428 = ~n33367 ;
  assign y21429 = ~1'b0 ;
  assign y21430 = n33371 ;
  assign y21431 = ~1'b0 ;
  assign y21432 = ~1'b0 ;
  assign y21433 = ~1'b0 ;
  assign y21434 = ~n33372 ;
  assign y21435 = ~1'b0 ;
  assign y21436 = n33375 ;
  assign y21437 = ~n33377 ;
  assign y21438 = ~n33378 ;
  assign y21439 = ~1'b0 ;
  assign y21440 = ~n33381 ;
  assign y21441 = ~n33382 ;
  assign y21442 = ~1'b0 ;
  assign y21443 = ~n31194 ;
  assign y21444 = ~n33387 ;
  assign y21445 = ~1'b0 ;
  assign y21446 = ~1'b0 ;
  assign y21447 = n33389 ;
  assign y21448 = ~1'b0 ;
  assign y21449 = ~1'b0 ;
  assign y21450 = n33390 ;
  assign y21451 = ~1'b0 ;
  assign y21452 = n33391 ;
  assign y21453 = ~n33392 ;
  assign y21454 = n33394 ;
  assign y21455 = n33396 ;
  assign y21456 = n33398 ;
  assign y21457 = ~n33399 ;
  assign y21458 = ~n11211 ;
  assign y21459 = ~n33406 ;
  assign y21460 = ~1'b0 ;
  assign y21461 = ~1'b0 ;
  assign y21462 = ~1'b0 ;
  assign y21463 = n33408 ;
  assign y21464 = n33409 ;
  assign y21465 = ~n33410 ;
  assign y21466 = ~1'b0 ;
  assign y21467 = ~1'b0 ;
  assign y21468 = n33412 ;
  assign y21469 = n33413 ;
  assign y21470 = ~1'b0 ;
  assign y21471 = ~n4460 ;
  assign y21472 = n33414 ;
  assign y21473 = n33416 ;
  assign y21474 = n33417 ;
  assign y21475 = ~n33424 ;
  assign y21476 = ~n33425 ;
  assign y21477 = ~n33430 ;
  assign y21478 = n33432 ;
  assign y21479 = ~1'b0 ;
  assign y21480 = ~n33437 ;
  assign y21481 = ~1'b0 ;
  assign y21482 = ~1'b0 ;
  assign y21483 = ~1'b0 ;
  assign y21484 = ~n33438 ;
  assign y21485 = n33440 ;
  assign y21486 = ~1'b0 ;
  assign y21487 = ~1'b0 ;
  assign y21488 = ~n33442 ;
  assign y21489 = n33445 ;
  assign y21490 = 1'b0 ;
  assign y21491 = ~n33446 ;
  assign y21492 = n33449 ;
  assign y21493 = ~n33452 ;
  assign y21494 = ~n33454 ;
  assign y21495 = ~1'b0 ;
  assign y21496 = ~n33457 ;
  assign y21497 = ~n33458 ;
  assign y21498 = ~1'b0 ;
  assign y21499 = n33459 ;
  assign y21500 = ~n33460 ;
  assign y21501 = n33461 ;
  assign y21502 = ~n33464 ;
  assign y21503 = n33465 ;
  assign y21504 = ~n33467 ;
  assign y21505 = ~n33468 ;
  assign y21506 = n4957 ;
  assign y21507 = ~n33473 ;
  assign y21508 = ~1'b0 ;
  assign y21509 = n33474 ;
  assign y21510 = ~n24647 ;
  assign y21511 = n33476 ;
  assign y21512 = ~1'b0 ;
  assign y21513 = 1'b0 ;
  assign y21514 = n33481 ;
  assign y21515 = n33484 ;
  assign y21516 = ~n33485 ;
  assign y21517 = ~n33487 ;
  assign y21518 = n33488 ;
  assign y21519 = n25615 ;
  assign y21520 = ~1'b0 ;
  assign y21521 = n33490 ;
  assign y21522 = ~n33494 ;
  assign y21523 = ~1'b0 ;
  assign y21524 = ~1'b0 ;
  assign y21525 = ~1'b0 ;
  assign y21526 = ~1'b0 ;
  assign y21527 = n33496 ;
  assign y21528 = ~n18541 ;
  assign y21529 = ~1'b0 ;
  assign y21530 = ~1'b0 ;
  assign y21531 = ~1'b0 ;
  assign y21532 = ~n14591 ;
  assign y21533 = n33498 ;
  assign y21534 = ~n33499 ;
  assign y21535 = ~n33501 ;
  assign y21536 = n33506 ;
  assign y21537 = ~1'b0 ;
  assign y21538 = n33507 ;
  assign y21539 = ~n33508 ;
  assign y21540 = 1'b0 ;
  assign y21541 = ~n33509 ;
  assign y21542 = ~1'b0 ;
  assign y21543 = ~n33510 ;
  assign y21544 = ~1'b0 ;
  assign y21545 = ~1'b0 ;
  assign y21546 = ~n33515 ;
  assign y21547 = n33517 ;
  assign y21548 = ~1'b0 ;
  assign y21549 = ~1'b0 ;
  assign y21550 = ~1'b0 ;
  assign y21551 = n8157 ;
  assign y21552 = n33519 ;
  assign y21553 = ~1'b0 ;
  assign y21554 = n11093 ;
  assign y21555 = ~n33521 ;
  assign y21556 = ~1'b0 ;
  assign y21557 = ~1'b0 ;
  assign y21558 = n33531 ;
  assign y21559 = 1'b0 ;
  assign y21560 = ~1'b0 ;
  assign y21561 = ~1'b0 ;
  assign y21562 = ~1'b0 ;
  assign y21563 = ~n33534 ;
  assign y21564 = n33536 ;
  assign y21565 = n33538 ;
  assign y21566 = n33541 ;
  assign y21567 = n33542 ;
  assign y21568 = ~1'b0 ;
  assign y21569 = n33546 ;
  assign y21570 = ~n5334 ;
  assign y21571 = 1'b0 ;
  assign y21572 = ~1'b0 ;
  assign y21573 = n33547 ;
  assign y21574 = n28543 ;
  assign y21575 = n33550 ;
  assign y21576 = ~n33552 ;
  assign y21577 = ~n33553 ;
  assign y21578 = ~n6351 ;
  assign y21579 = n33554 ;
  assign y21580 = ~1'b0 ;
  assign y21581 = ~n33555 ;
  assign y21582 = ~1'b0 ;
  assign y21583 = n20272 ;
  assign y21584 = ~1'b0 ;
  assign y21585 = ~n33556 ;
  assign y21586 = ~n33557 ;
  assign y21587 = ~n24351 ;
  assign y21588 = n33558 ;
  assign y21589 = ~n33559 ;
  assign y21590 = n33562 ;
  assign y21591 = ~n33563 ;
  assign y21592 = ~1'b0 ;
  assign y21593 = ~1'b0 ;
  assign y21594 = ~1'b0 ;
  assign y21595 = ~n33569 ;
  assign y21596 = n33571 ;
  assign y21597 = n33572 ;
  assign y21598 = ~n33574 ;
  assign y21599 = n33575 ;
  assign y21600 = ~1'b0 ;
  assign y21601 = n33578 ;
  assign y21602 = ~1'b0 ;
  assign y21603 = ~n33579 ;
  assign y21604 = n33584 ;
  assign y21605 = 1'b0 ;
  assign y21606 = ~1'b0 ;
  assign y21607 = ~n33590 ;
  assign y21608 = n12245 ;
  assign y21609 = ~1'b0 ;
  assign y21610 = ~1'b0 ;
  assign y21611 = ~1'b0 ;
  assign y21612 = ~n33592 ;
  assign y21613 = ~1'b0 ;
  assign y21614 = ~1'b0 ;
  assign y21615 = ~n33593 ;
  assign y21616 = ~n33595 ;
  assign y21617 = ~1'b0 ;
  assign y21618 = ~n33597 ;
  assign y21619 = ~1'b0 ;
  assign y21620 = ~n33604 ;
  assign y21621 = ~1'b0 ;
  assign y21622 = n33606 ;
  assign y21623 = ~n33608 ;
  assign y21624 = ~n33609 ;
  assign y21625 = ~n33610 ;
  assign y21626 = ~n33614 ;
  assign y21627 = ~n33616 ;
  assign y21628 = ~1'b0 ;
  assign y21629 = ~n10078 ;
  assign y21630 = ~1'b0 ;
  assign y21631 = n33620 ;
  assign y21632 = n33623 ;
  assign y21633 = ~n33625 ;
  assign y21634 = n33626 ;
  assign y21635 = ~1'b0 ;
  assign y21636 = n33627 ;
  assign y21637 = n33628 ;
  assign y21638 = ~n33629 ;
  assign y21639 = ~n9618 ;
  assign y21640 = ~n33630 ;
  assign y21641 = ~n33631 ;
  assign y21642 = ~n33636 ;
  assign y21643 = n33639 ;
  assign y21644 = ~1'b0 ;
  assign y21645 = ~n33640 ;
  assign y21646 = ~n33642 ;
  assign y21647 = ~n33643 ;
  assign y21648 = 1'b0 ;
  assign y21649 = 1'b0 ;
  assign y21650 = n33644 ;
  assign y21651 = n33649 ;
  assign y21652 = n33651 ;
  assign y21653 = n33652 ;
  assign y21654 = n33656 ;
  assign y21655 = n33657 ;
  assign y21656 = ~n10522 ;
  assign y21657 = n33665 ;
  assign y21658 = ~n33667 ;
  assign y21659 = n20756 ;
  assign y21660 = ~1'b0 ;
  assign y21661 = ~n33669 ;
  assign y21662 = ~n33671 ;
  assign y21663 = ~n4094 ;
  assign y21664 = ~n33673 ;
  assign y21665 = ~1'b0 ;
  assign y21666 = n33679 ;
  assign y21667 = ~n33683 ;
  assign y21668 = ~n33685 ;
  assign y21669 = 1'b0 ;
  assign y21670 = n33686 ;
  assign y21671 = n33689 ;
  assign y21672 = n33690 ;
  assign y21673 = ~1'b0 ;
  assign y21674 = ~n33697 ;
  assign y21675 = ~1'b0 ;
  assign y21676 = ~n33699 ;
  assign y21677 = ~n33700 ;
  assign y21678 = n33701 ;
  assign y21679 = ~n32648 ;
  assign y21680 = ~n32796 ;
  assign y21681 = ~1'b0 ;
  assign y21682 = ~1'b0 ;
  assign y21683 = ~1'b0 ;
  assign y21684 = ~n33702 ;
  assign y21685 = ~1'b0 ;
  assign y21686 = ~1'b0 ;
  assign y21687 = 1'b0 ;
  assign y21688 = ~n33703 ;
  assign y21689 = ~1'b0 ;
  assign y21690 = ~1'b0 ;
  assign y21691 = ~n33704 ;
  assign y21692 = ~n33708 ;
  assign y21693 = ~1'b0 ;
  assign y21694 = ~1'b0 ;
  assign y21695 = ~1'b0 ;
  assign y21696 = ~1'b0 ;
  assign y21697 = ~n33709 ;
  assign y21698 = n33710 ;
  assign y21699 = n25000 ;
  assign y21700 = ~1'b0 ;
  assign y21701 = ~n33711 ;
  assign y21702 = ~n33712 ;
  assign y21703 = n33713 ;
  assign y21704 = n33715 ;
  assign y21705 = ~1'b0 ;
  assign y21706 = n33717 ;
  assign y21707 = 1'b0 ;
  assign y21708 = ~1'b0 ;
  assign y21709 = n33721 ;
  assign y21710 = ~1'b0 ;
  assign y21711 = ~n33724 ;
  assign y21712 = ~1'b0 ;
  assign y21713 = n33726 ;
  assign y21714 = ~n22756 ;
  assign y21715 = n33727 ;
  assign y21716 = n33729 ;
  assign y21717 = ~1'b0 ;
  assign y21718 = n33730 ;
  assign y21719 = ~1'b0 ;
  assign y21720 = ~1'b0 ;
  assign y21721 = ~n33731 ;
  assign y21722 = ~1'b0 ;
  assign y21723 = n33734 ;
  assign y21724 = ~1'b0 ;
  assign y21725 = ~n33736 ;
  assign y21726 = 1'b0 ;
  assign y21727 = n33737 ;
  assign y21728 = ~1'b0 ;
  assign y21729 = n33739 ;
  assign y21730 = ~1'b0 ;
  assign y21731 = ~1'b0 ;
  assign y21732 = ~n33741 ;
  assign y21733 = 1'b0 ;
  assign y21734 = 1'b0 ;
  assign y21735 = ~1'b0 ;
  assign y21736 = ~1'b0 ;
  assign y21737 = ~1'b0 ;
  assign y21738 = ~1'b0 ;
  assign y21739 = ~n33742 ;
  assign y21740 = n33747 ;
  assign y21741 = n33748 ;
  assign y21742 = ~n33752 ;
  assign y21743 = n33753 ;
  assign y21744 = n33755 ;
  assign y21745 = ~1'b0 ;
  assign y21746 = n33759 ;
  assign y21747 = ~n33763 ;
  assign y21748 = ~1'b0 ;
  assign y21749 = ~1'b0 ;
  assign y21750 = n33766 ;
  assign y21751 = ~1'b0 ;
  assign y21752 = n33768 ;
  assign y21753 = n33769 ;
  assign y21754 = n26997 ;
  assign y21755 = n33771 ;
  assign y21756 = n33772 ;
  assign y21757 = n33773 ;
  assign y21758 = ~n7236 ;
  assign y21759 = ~1'b0 ;
  assign y21760 = ~n33777 ;
  assign y21761 = ~1'b0 ;
  assign y21762 = ~n33778 ;
  assign y21763 = ~n33780 ;
  assign y21764 = n33782 ;
  assign y21765 = n3466 ;
  assign y21766 = ~n33784 ;
  assign y21767 = ~1'b0 ;
  assign y21768 = ~n15716 ;
  assign y21769 = ~n33786 ;
  assign y21770 = ~1'b0 ;
  assign y21771 = 1'b0 ;
  assign y21772 = ~n33789 ;
  assign y21773 = ~n33791 ;
  assign y21774 = ~n33792 ;
  assign y21775 = n33793 ;
  assign y21776 = 1'b0 ;
  assign y21777 = ~1'b0 ;
  assign y21778 = ~1'b0 ;
  assign y21779 = ~n33794 ;
  assign y21780 = n33795 ;
  assign y21781 = ~n21630 ;
  assign y21782 = ~1'b0 ;
  assign y21783 = ~n33797 ;
  assign y21784 = ~n33802 ;
  assign y21785 = ~n33806 ;
  assign y21786 = ~1'b0 ;
  assign y21787 = ~n33808 ;
  assign y21788 = ~n33809 ;
  assign y21789 = ~n1443 ;
  assign y21790 = n6211 ;
  assign y21791 = n33817 ;
  assign y21792 = n26598 ;
  assign y21793 = n33821 ;
  assign y21794 = ~1'b0 ;
  assign y21795 = ~n33822 ;
  assign y21796 = ~1'b0 ;
  assign y21797 = ~n6344 ;
  assign y21798 = ~1'b0 ;
  assign y21799 = ~1'b0 ;
  assign y21800 = ~1'b0 ;
  assign y21801 = ~n33824 ;
  assign y21802 = ~1'b0 ;
  assign y21803 = ~n21944 ;
  assign y21804 = n1327 ;
  assign y21805 = n33828 ;
  assign y21806 = n33829 ;
  assign y21807 = n33830 ;
  assign y21808 = ~n33831 ;
  assign y21809 = ~1'b0 ;
  assign y21810 = n33834 ;
  assign y21811 = ~n33837 ;
  assign y21812 = n33840 ;
  assign y21813 = ~1'b0 ;
  assign y21814 = ~1'b0 ;
  assign y21815 = n33841 ;
  assign y21816 = ~1'b0 ;
  assign y21817 = ~1'b0 ;
  assign y21818 = n33843 ;
  assign y21819 = ~n33845 ;
  assign y21820 = ~n33846 ;
  assign y21821 = ~n33848 ;
  assign y21822 = n33849 ;
  assign y21823 = ~n4428 ;
  assign y21824 = ~1'b0 ;
  assign y21825 = ~n33851 ;
  assign y21826 = n33853 ;
  assign y21827 = n33855 ;
  assign y21828 = n33857 ;
  assign y21829 = n33858 ;
  assign y21830 = n2071 ;
  assign y21831 = ~1'b0 ;
  assign y21832 = ~n9380 ;
  assign y21833 = n33859 ;
  assign y21834 = ~1'b0 ;
  assign y21835 = ~1'b0 ;
  assign y21836 = ~n33862 ;
  assign y21837 = n4569 ;
  assign y21838 = n8286 ;
  assign y21839 = ~n33863 ;
  assign y21840 = n33865 ;
  assign y21841 = n33866 ;
  assign y21842 = ~1'b0 ;
  assign y21843 = ~1'b0 ;
  assign y21844 = ~1'b0 ;
  assign y21845 = ~1'b0 ;
  assign y21846 = n884 ;
  assign y21847 = n33869 ;
  assign y21848 = n4982 ;
  assign y21849 = ~1'b0 ;
  assign y21850 = n33872 ;
  assign y21851 = ~1'b0 ;
  assign y21852 = ~n33873 ;
  assign y21853 = ~1'b0 ;
  assign y21854 = ~n33876 ;
  assign y21855 = n33885 ;
  assign y21856 = ~1'b0 ;
  assign y21857 = ~1'b0 ;
  assign y21858 = 1'b0 ;
  assign y21859 = n4582 ;
  assign y21860 = ~1'b0 ;
  assign y21861 = ~n33888 ;
  assign y21862 = ~n33890 ;
  assign y21863 = ~n33895 ;
  assign y21864 = ~1'b0 ;
  assign y21865 = ~n33896 ;
  assign y21866 = ~n33898 ;
  assign y21867 = n33900 ;
  assign y21868 = ~n33906 ;
  assign y21869 = n33907 ;
  assign y21870 = ~n33911 ;
  assign y21871 = n33913 ;
  assign y21872 = ~1'b0 ;
  assign y21873 = n33916 ;
  assign y21874 = n33917 ;
  assign y21875 = ~1'b0 ;
  assign y21876 = ~1'b0 ;
  assign y21877 = ~1'b0 ;
  assign y21878 = 1'b0 ;
  assign y21879 = ~n20608 ;
  assign y21880 = ~n33925 ;
  assign y21881 = ~n33927 ;
  assign y21882 = ~n33929 ;
  assign y21883 = n33933 ;
  assign y21884 = ~1'b0 ;
  assign y21885 = ~1'b0 ;
  assign y21886 = n33937 ;
  assign y21887 = ~n33946 ;
  assign y21888 = ~1'b0 ;
  assign y21889 = ~1'b0 ;
  assign y21890 = ~n33950 ;
  assign y21891 = n33952 ;
  assign y21892 = n33953 ;
  assign y21893 = ~1'b0 ;
  assign y21894 = ~1'b0 ;
  assign y21895 = ~1'b0 ;
  assign y21896 = ~1'b0 ;
  assign y21897 = n33954 ;
  assign y21898 = ~n33956 ;
  assign y21899 = ~1'b0 ;
  assign y21900 = ~1'b0 ;
  assign y21901 = ~1'b0 ;
  assign y21902 = ~1'b0 ;
  assign y21903 = ~n33959 ;
  assign y21904 = ~1'b0 ;
  assign y21905 = n33961 ;
  assign y21906 = n33963 ;
  assign y21907 = ~1'b0 ;
  assign y21908 = ~n33965 ;
  assign y21909 = ~n33971 ;
  assign y21910 = ~n33973 ;
  assign y21911 = ~n33976 ;
  assign y21912 = ~n33979 ;
  assign y21913 = ~1'b0 ;
  assign y21914 = n33980 ;
  assign y21915 = ~1'b0 ;
  assign y21916 = n33982 ;
  assign y21917 = ~1'b0 ;
  assign y21918 = ~1'b0 ;
  assign y21919 = ~1'b0 ;
  assign y21920 = ~1'b0 ;
  assign y21921 = ~1'b0 ;
  assign y21922 = ~n33983 ;
  assign y21923 = ~1'b0 ;
  assign y21924 = ~1'b0 ;
  assign y21925 = ~1'b0 ;
  assign y21926 = ~x29 ;
  assign y21927 = ~1'b0 ;
  assign y21928 = ~n33987 ;
  assign y21929 = ~1'b0 ;
  assign y21930 = n26252 ;
  assign y21931 = n33989 ;
  assign y21932 = n806 ;
  assign y21933 = n33991 ;
  assign y21934 = ~1'b0 ;
  assign y21935 = n33993 ;
  assign y21936 = ~1'b0 ;
  assign y21937 = ~n33995 ;
  assign y21938 = ~1'b0 ;
  assign y21939 = ~n33997 ;
  assign y21940 = ~n18126 ;
  assign y21941 = ~1'b0 ;
  assign y21942 = n1757 ;
  assign y21943 = ~1'b0 ;
  assign y21944 = n34000 ;
  assign y21945 = ~1'b0 ;
  assign y21946 = ~n34003 ;
  assign y21947 = n16821 ;
  assign y21948 = ~n34004 ;
  assign y21949 = ~1'b0 ;
  assign y21950 = ~n34006 ;
  assign y21951 = ~1'b0 ;
  assign y21952 = n34007 ;
  assign y21953 = n34008 ;
  assign y21954 = ~1'b0 ;
  assign y21955 = ~n11148 ;
  assign y21956 = ~1'b0 ;
  assign y21957 = ~1'b0 ;
  assign y21958 = ~1'b0 ;
  assign y21959 = ~1'b0 ;
  assign y21960 = ~n34011 ;
  assign y21961 = ~1'b0 ;
  assign y21962 = ~n34013 ;
  assign y21963 = ~n34015 ;
  assign y21964 = ~1'b0 ;
  assign y21965 = n34017 ;
  assign y21966 = n33696 ;
  assign y21967 = ~1'b0 ;
  assign y21968 = 1'b0 ;
  assign y21969 = n34018 ;
  assign y21970 = ~n12721 ;
  assign y21971 = ~n34020 ;
  assign y21972 = ~1'b0 ;
  assign y21973 = n34021 ;
  assign y21974 = ~n34025 ;
  assign y21975 = n34026 ;
  assign y21976 = n34028 ;
  assign y21977 = n34029 ;
  assign y21978 = ~1'b0 ;
  assign y21979 = ~1'b0 ;
  assign y21980 = ~1'b0 ;
  assign y21981 = ~1'b0 ;
  assign y21982 = ~n1663 ;
  assign y21983 = ~1'b0 ;
  assign y21984 = n34030 ;
  assign y21985 = n15328 ;
  assign y21986 = ~n2029 ;
  assign y21987 = n34032 ;
  assign y21988 = ~n34033 ;
  assign y21989 = ~1'b0 ;
  assign y21990 = n34034 ;
  assign y21991 = n34035 ;
  assign y21992 = ~n34036 ;
  assign y21993 = ~1'b0 ;
  assign y21994 = ~1'b0 ;
  assign y21995 = n34038 ;
  assign y21996 = n34039 ;
  assign y21997 = n23245 ;
  assign y21998 = n34044 ;
  assign y21999 = ~1'b0 ;
  assign y22000 = ~1'b0 ;
  assign y22001 = ~n34046 ;
  assign y22002 = ~1'b0 ;
  assign y22003 = ~n34049 ;
  assign y22004 = n34053 ;
  assign y22005 = 1'b0 ;
  assign y22006 = ~n34056 ;
  assign y22007 = 1'b0 ;
  assign y22008 = ~n21854 ;
  assign y22009 = n34058 ;
  assign y22010 = ~1'b0 ;
  assign y22011 = ~n34061 ;
  assign y22012 = ~n34068 ;
  assign y22013 = 1'b0 ;
  assign y22014 = ~n34070 ;
  assign y22015 = 1'b0 ;
  assign y22016 = ~n34072 ;
  assign y22017 = n34073 ;
  assign y22018 = ~1'b0 ;
  assign y22019 = ~n12324 ;
  assign y22020 = ~n34078 ;
  assign y22021 = ~n34082 ;
  assign y22022 = ~1'b0 ;
  assign y22023 = ~n26116 ;
  assign y22024 = n34086 ;
  assign y22025 = n23825 ;
  assign y22026 = ~1'b0 ;
  assign y22027 = ~1'b0 ;
  assign y22028 = x17 ;
  assign y22029 = n34087 ;
  assign y22030 = n34088 ;
  assign y22031 = n34094 ;
  assign y22032 = ~1'b0 ;
  assign y22033 = ~n34096 ;
  assign y22034 = ~1'b0 ;
  assign y22035 = ~n34097 ;
  assign y22036 = n34100 ;
  assign y22037 = ~n34101 ;
  assign y22038 = ~1'b0 ;
  assign y22039 = ~n34102 ;
  assign y22040 = ~1'b0 ;
  assign y22041 = ~n34103 ;
  assign y22042 = n34104 ;
  assign y22043 = n4810 ;
  assign y22044 = n1223 ;
  assign y22045 = ~1'b0 ;
  assign y22046 = 1'b0 ;
  assign y22047 = ~1'b0 ;
  assign y22048 = 1'b0 ;
  assign y22049 = ~1'b0 ;
  assign y22050 = ~n34105 ;
  assign y22051 = ~1'b0 ;
  assign y22052 = n34106 ;
  assign y22053 = ~n34108 ;
  assign y22054 = n34109 ;
  assign y22055 = ~1'b0 ;
  assign y22056 = ~n34111 ;
  assign y22057 = ~1'b0 ;
  assign y22058 = n34113 ;
  assign y22059 = ~1'b0 ;
  assign y22060 = ~n34115 ;
  assign y22061 = ~n34119 ;
  assign y22062 = ~1'b0 ;
  assign y22063 = n34125 ;
  assign y22064 = n34128 ;
  assign y22065 = ~n34131 ;
  assign y22066 = ~1'b0 ;
  assign y22067 = ~1'b0 ;
  assign y22068 = ~1'b0 ;
  assign y22069 = ~1'b0 ;
  assign y22070 = ~n34132 ;
  assign y22071 = ~1'b0 ;
  assign y22072 = n34133 ;
  assign y22073 = ~1'b0 ;
  assign y22074 = n12474 ;
  assign y22075 = ~n34135 ;
  assign y22076 = ~n21960 ;
  assign y22077 = ~n34137 ;
  assign y22078 = ~n34141 ;
  assign y22079 = ~1'b0 ;
  assign y22080 = ~1'b0 ;
  assign y22081 = n34142 ;
  assign y22082 = n34143 ;
  assign y22083 = ~n34145 ;
  assign y22084 = 1'b0 ;
  assign y22085 = ~n34146 ;
  assign y22086 = n34147 ;
  assign y22087 = ~n34149 ;
  assign y22088 = n34150 ;
  assign y22089 = n20459 ;
  assign y22090 = n34151 ;
  assign y22091 = ~1'b0 ;
  assign y22092 = ~1'b0 ;
  assign y22093 = ~1'b0 ;
  assign y22094 = n34153 ;
  assign y22095 = n34155 ;
  assign y22096 = ~1'b0 ;
  assign y22097 = ~1'b0 ;
  assign y22098 = ~1'b0 ;
  assign y22099 = n15423 ;
  assign y22100 = ~n34158 ;
  assign y22101 = ~1'b0 ;
  assign y22102 = ~1'b0 ;
  assign y22103 = n34159 ;
  assign y22104 = n34164 ;
  assign y22105 = ~n9339 ;
  assign y22106 = ~n34174 ;
  assign y22107 = ~n34176 ;
  assign y22108 = ~1'b0 ;
  assign y22109 = n34177 ;
  assign y22110 = n34179 ;
  assign y22111 = ~1'b0 ;
  assign y22112 = ~1'b0 ;
  assign y22113 = ~n34181 ;
  assign y22114 = ~n34183 ;
  assign y22115 = ~1'b0 ;
  assign y22116 = n34184 ;
  assign y22117 = n16744 ;
  assign y22118 = ~1'b0 ;
  assign y22119 = n34185 ;
  assign y22120 = ~1'b0 ;
  assign y22121 = n34188 ;
  assign y22122 = ~1'b0 ;
  assign y22123 = n34189 ;
  assign y22124 = n34190 ;
  assign y22125 = ~n34193 ;
  assign y22126 = ~1'b0 ;
  assign y22127 = ~n34197 ;
  assign y22128 = n34198 ;
  assign y22129 = ~1'b0 ;
  assign y22130 = ~n28689 ;
  assign y22131 = n34202 ;
  assign y22132 = n34205 ;
  assign y22133 = ~1'b0 ;
  assign y22134 = n34206 ;
  assign y22135 = ~n29404 ;
  assign y22136 = n15456 ;
  assign y22137 = ~1'b0 ;
  assign y22138 = ~n34207 ;
  assign y22139 = n34210 ;
  assign y22140 = ~n34213 ;
  assign y22141 = ~1'b0 ;
  assign y22142 = ~1'b0 ;
  assign y22143 = ~1'b0 ;
  assign y22144 = ~n5778 ;
  assign y22145 = ~n34214 ;
  assign y22146 = ~n16942 ;
  assign y22147 = ~1'b0 ;
  assign y22148 = n34215 ;
  assign y22149 = n34217 ;
  assign y22150 = 1'b0 ;
  assign y22151 = ~1'b0 ;
  assign y22152 = ~n34220 ;
  assign y22153 = ~1'b0 ;
  assign y22154 = ~1'b0 ;
  assign y22155 = ~n34221 ;
  assign y22156 = n34222 ;
  assign y22157 = ~1'b0 ;
  assign y22158 = ~n34223 ;
  assign y22159 = n34227 ;
  assign y22160 = n34235 ;
  assign y22161 = ~1'b0 ;
  assign y22162 = n34236 ;
  assign y22163 = n34242 ;
  assign y22164 = ~1'b0 ;
  assign y22165 = ~1'b0 ;
  assign y22166 = ~n34244 ;
  assign y22167 = ~n34247 ;
  assign y22168 = ~1'b0 ;
  assign y22169 = ~n34249 ;
  assign y22170 = ~n34250 ;
  assign y22171 = ~1'b0 ;
  assign y22172 = n34253 ;
  assign y22173 = ~n34258 ;
  assign y22174 = n1443 ;
  assign y22175 = ~1'b0 ;
  assign y22176 = n5077 ;
  assign y22177 = n34259 ;
  assign y22178 = ~n34261 ;
  assign y22179 = n34263 ;
  assign y22180 = ~1'b0 ;
  assign y22181 = n34267 ;
  assign y22182 = n34271 ;
  assign y22183 = ~n16129 ;
  assign y22184 = n34273 ;
  assign y22185 = ~n34279 ;
  assign y22186 = ~1'b0 ;
  assign y22187 = ~1'b0 ;
  assign y22188 = n34281 ;
  assign y22189 = ~1'b0 ;
  assign y22190 = n34284 ;
  assign y22191 = ~1'b0 ;
  assign y22192 = ~n34288 ;
  assign y22193 = ~1'b0 ;
  assign y22194 = ~n14438 ;
  assign y22195 = n34292 ;
  assign y22196 = ~n34298 ;
  assign y22197 = ~1'b0 ;
  assign y22198 = ~n34299 ;
  assign y22199 = ~n34300 ;
  assign y22200 = n34302 ;
  assign y22201 = ~1'b0 ;
  assign y22202 = n34311 ;
  assign y22203 = ~1'b0 ;
  assign y22204 = ~1'b0 ;
  assign y22205 = ~1'b0 ;
  assign y22206 = ~n34312 ;
  assign y22207 = n34313 ;
  assign y22208 = ~1'b0 ;
  assign y22209 = n34314 ;
  assign y22210 = ~1'b0 ;
  assign y22211 = ~1'b0 ;
  assign y22212 = n34318 ;
  assign y22213 = n34319 ;
  assign y22214 = ~n34322 ;
  assign y22215 = ~n34329 ;
  assign y22216 = ~n34331 ;
  assign y22217 = n34332 ;
  assign y22218 = ~1'b0 ;
  assign y22219 = ~n34334 ;
  assign y22220 = n34335 ;
  assign y22221 = ~1'b0 ;
  assign y22222 = ~1'b0 ;
  assign y22223 = ~n34336 ;
  assign y22224 = ~1'b0 ;
  assign y22225 = n34337 ;
  assign y22226 = n34338 ;
  assign y22227 = n34340 ;
  assign y22228 = n34345 ;
  assign y22229 = ~n34347 ;
  assign y22230 = ~n16552 ;
  assign y22231 = ~1'b0 ;
  assign y22232 = ~n2223 ;
  assign y22233 = ~n34349 ;
  assign y22234 = n34352 ;
  assign y22235 = ~1'b0 ;
  assign y22236 = ~1'b0 ;
  assign y22237 = ~n34353 ;
  assign y22238 = n34355 ;
  assign y22239 = ~1'b0 ;
  assign y22240 = ~n34356 ;
  assign y22241 = n34358 ;
  assign y22242 = ~n34360 ;
  assign y22243 = ~n27575 ;
  assign y22244 = ~1'b0 ;
  assign y22245 = ~1'b0 ;
  assign y22246 = n34361 ;
  assign y22247 = n34368 ;
  assign y22248 = ~1'b0 ;
  assign y22249 = n20529 ;
  assign y22250 = ~1'b0 ;
  assign y22251 = ~n34371 ;
  assign y22252 = ~n34375 ;
  assign y22253 = x250 ;
  assign y22254 = n34377 ;
  assign y22255 = n34380 ;
  assign y22256 = ~1'b0 ;
  assign y22257 = n34383 ;
  assign y22258 = n34384 ;
  assign y22259 = n34386 ;
  assign y22260 = ~n20859 ;
  assign y22261 = ~1'b0 ;
  assign y22262 = n34388 ;
  assign y22263 = ~n34390 ;
  assign y22264 = ~n34392 ;
  assign y22265 = ~n34395 ;
  assign y22266 = n34400 ;
  assign y22267 = ~n2809 ;
  assign y22268 = n34404 ;
  assign y22269 = ~n34406 ;
  assign y22270 = ~n34408 ;
  assign y22271 = n34410 ;
  assign y22272 = ~n34422 ;
  assign y22273 = ~1'b0 ;
  assign y22274 = ~1'b0 ;
  assign y22275 = n25154 ;
  assign y22276 = n34425 ;
  assign y22277 = n34428 ;
  assign y22278 = ~n34434 ;
  assign y22279 = ~1'b0 ;
  assign y22280 = n34436 ;
  assign y22281 = ~n34437 ;
  assign y22282 = ~n34439 ;
  assign y22283 = ~n34441 ;
  assign y22284 = ~n34448 ;
  assign y22285 = n34449 ;
  assign y22286 = n34451 ;
  assign y22287 = ~1'b0 ;
  assign y22288 = 1'b0 ;
  assign y22289 = n34452 ;
  assign y22290 = n34453 ;
  assign y22291 = 1'b0 ;
  assign y22292 = n34455 ;
  assign y22293 = ~1'b0 ;
  assign y22294 = ~1'b0 ;
  assign y22295 = n34456 ;
  assign y22296 = n34457 ;
  assign y22297 = ~n34459 ;
  assign y22298 = ~n34460 ;
  assign y22299 = n34463 ;
  assign y22300 = ~n34467 ;
  assign y22301 = n34473 ;
  assign y22302 = ~1'b0 ;
  assign y22303 = ~n34475 ;
  assign y22304 = ~1'b0 ;
  assign y22305 = n34476 ;
  assign y22306 = ~n34480 ;
  assign y22307 = ~1'b0 ;
  assign y22308 = ~1'b0 ;
  assign y22309 = ~n34481 ;
  assign y22310 = n34482 ;
  assign y22311 = ~n34484 ;
  assign y22312 = ~1'b0 ;
  assign y22313 = n34486 ;
  assign y22314 = ~1'b0 ;
  assign y22315 = ~1'b0 ;
  assign y22316 = ~n34488 ;
  assign y22317 = n34489 ;
  assign y22318 = ~n34491 ;
  assign y22319 = ~n34493 ;
  assign y22320 = ~n34494 ;
  assign y22321 = ~n34496 ;
  assign y22322 = ~1'b0 ;
  assign y22323 = ~n34501 ;
  assign y22324 = ~n34504 ;
  assign y22325 = n34506 ;
  assign y22326 = n34510 ;
  assign y22327 = n34512 ;
  assign y22328 = ~n34514 ;
  assign y22329 = 1'b0 ;
  assign y22330 = n24530 ;
  assign y22331 = n34517 ;
  assign y22332 = ~n34519 ;
  assign y22333 = 1'b0 ;
  assign y22334 = n26971 ;
  assign y22335 = ~n34520 ;
  assign y22336 = ~1'b0 ;
  assign y22337 = n34525 ;
  assign y22338 = n28826 ;
  assign y22339 = ~n34526 ;
  assign y22340 = 1'b0 ;
  assign y22341 = n34530 ;
  assign y22342 = n11454 ;
  assign y22343 = ~1'b0 ;
  assign y22344 = ~1'b0 ;
  assign y22345 = 1'b0 ;
  assign y22346 = 1'b0 ;
  assign y22347 = n34534 ;
  assign y22348 = ~1'b0 ;
  assign y22349 = ~n34535 ;
  assign y22350 = ~n34539 ;
  assign y22351 = ~1'b0 ;
  assign y22352 = n34540 ;
  assign y22353 = ~1'b0 ;
  assign y22354 = n34541 ;
  assign y22355 = n34544 ;
  assign y22356 = n15768 ;
  assign y22357 = n34547 ;
  assign y22358 = 1'b0 ;
  assign y22359 = n34548 ;
  assign y22360 = n34549 ;
  assign y22361 = n3333 ;
  assign y22362 = ~1'b0 ;
  assign y22363 = n34551 ;
  assign y22364 = ~1'b0 ;
  assign y22365 = n34552 ;
  assign y22366 = n34554 ;
  assign y22367 = n32584 ;
  assign y22368 = ~1'b0 ;
  assign y22369 = n34555 ;
  assign y22370 = n34556 ;
  assign y22371 = ~n34559 ;
  assign y22372 = 1'b0 ;
  assign y22373 = ~1'b0 ;
  assign y22374 = n34560 ;
  assign y22375 = ~n34563 ;
  assign y22376 = ~1'b0 ;
  assign y22377 = ~n34564 ;
  assign y22378 = n34566 ;
  assign y22379 = ~1'b0 ;
  assign y22380 = ~1'b0 ;
  assign y22381 = n34571 ;
  assign y22382 = n1324 ;
  assign y22383 = ~n34573 ;
  assign y22384 = ~1'b0 ;
  assign y22385 = n34574 ;
  assign y22386 = ~n34575 ;
  assign y22387 = ~1'b0 ;
  assign y22388 = ~1'b0 ;
  assign y22389 = ~n34580 ;
  assign y22390 = n34582 ;
  assign y22391 = n34583 ;
  assign y22392 = n34584 ;
  assign y22393 = n34586 ;
  assign y22394 = ~n34588 ;
  assign y22395 = 1'b0 ;
  assign y22396 = n34589 ;
  assign y22397 = ~n34591 ;
  assign y22398 = ~1'b0 ;
  assign y22399 = n34593 ;
  assign y22400 = ~n8959 ;
  assign y22401 = n6119 ;
  assign y22402 = ~n34595 ;
  assign y22403 = ~1'b0 ;
  assign y22404 = ~n34598 ;
  assign y22405 = ~n34599 ;
  assign y22406 = 1'b0 ;
  assign y22407 = n34602 ;
  assign y22408 = n15477 ;
  assign y22409 = ~1'b0 ;
  assign y22410 = ~1'b0 ;
  assign y22411 = ~1'b0 ;
  assign y22412 = ~1'b0 ;
  assign y22413 = ~1'b0 ;
  assign y22414 = ~1'b0 ;
  assign y22415 = n4261 ;
  assign y22416 = ~n34604 ;
  assign y22417 = n34609 ;
  assign y22418 = ~n34610 ;
  assign y22419 = ~n34611 ;
  assign y22420 = n34612 ;
  assign y22421 = ~n34614 ;
  assign y22422 = ~1'b0 ;
  assign y22423 = ~1'b0 ;
  assign y22424 = ~1'b0 ;
  assign y22425 = n34617 ;
  assign y22426 = ~n34621 ;
  assign y22427 = n34622 ;
  assign y22428 = 1'b0 ;
  assign y22429 = ~n34623 ;
  assign y22430 = n15161 ;
  assign y22431 = ~1'b0 ;
  assign y22432 = n34624 ;
  assign y22433 = ~n34628 ;
  assign y22434 = ~1'b0 ;
  assign y22435 = n34629 ;
  assign y22436 = ~n34630 ;
  assign y22437 = ~n34631 ;
  assign y22438 = n8959 ;
  assign y22439 = ~1'b0 ;
  assign y22440 = ~1'b0 ;
  assign y22441 = ~n34635 ;
  assign y22442 = 1'b0 ;
  assign y22443 = ~1'b0 ;
  assign y22444 = ~n34638 ;
  assign y22445 = ~n34640 ;
  assign y22446 = ~n34641 ;
  assign y22447 = n34642 ;
  assign y22448 = ~n34643 ;
  assign y22449 = n34644 ;
  assign y22450 = ~1'b0 ;
  assign y22451 = ~1'b0 ;
  assign y22452 = 1'b0 ;
  assign y22453 = ~n34645 ;
  assign y22454 = n34647 ;
  assign y22455 = n34648 ;
  assign y22456 = ~1'b0 ;
  assign y22457 = ~n34649 ;
  assign y22458 = n34653 ;
  assign y22459 = 1'b0 ;
  assign y22460 = n14407 ;
  assign y22461 = n34657 ;
  assign y22462 = ~1'b0 ;
  assign y22463 = ~n34665 ;
  assign y22464 = ~1'b0 ;
  assign y22465 = ~n34666 ;
  assign y22466 = ~1'b0 ;
  assign y22467 = n24321 ;
  assign y22468 = ~1'b0 ;
  assign y22469 = n34667 ;
  assign y22470 = n34669 ;
  assign y22471 = ~1'b0 ;
  assign y22472 = ~1'b0 ;
  assign y22473 = ~1'b0 ;
  assign y22474 = n34671 ;
  assign y22475 = ~n15531 ;
  assign y22476 = ~1'b0 ;
  assign y22477 = ~1'b0 ;
  assign y22478 = n34675 ;
  assign y22479 = n34683 ;
  assign y22480 = n34688 ;
  assign y22481 = n34689 ;
  assign y22482 = ~1'b0 ;
  assign y22483 = ~1'b0 ;
  assign y22484 = n26937 ;
  assign y22485 = ~n34690 ;
  assign y22486 = n34692 ;
  assign y22487 = n34695 ;
  assign y22488 = n34696 ;
  assign y22489 = n34697 ;
  assign y22490 = ~n34701 ;
  assign y22491 = ~1'b0 ;
  assign y22492 = n34702 ;
  assign y22493 = ~1'b0 ;
  assign y22494 = n8873 ;
  assign y22495 = ~1'b0 ;
  assign y22496 = ~n11711 ;
  assign y22497 = n34706 ;
  assign y22498 = 1'b0 ;
  assign y22499 = 1'b0 ;
  assign y22500 = n34707 ;
  assign y22501 = ~1'b0 ;
  assign y22502 = ~n34709 ;
  assign y22503 = ~n34710 ;
  assign y22504 = n34711 ;
  assign y22505 = ~n34714 ;
  assign y22506 = n34717 ;
  assign y22507 = ~1'b0 ;
  assign y22508 = n34718 ;
  assign y22509 = ~1'b0 ;
  assign y22510 = n34721 ;
  assign y22511 = ~n34723 ;
  assign y22512 = ~1'b0 ;
  assign y22513 = ~n4755 ;
  assign y22514 = n34725 ;
  assign y22515 = n34728 ;
  assign y22516 = ~1'b0 ;
  assign y22517 = ~1'b0 ;
  assign y22518 = 1'b0 ;
  assign y22519 = ~n34729 ;
  assign y22520 = ~n34734 ;
  assign y22521 = ~n34735 ;
  assign y22522 = ~n25640 ;
  assign y22523 = ~1'b0 ;
  assign y22524 = ~1'b0 ;
  assign y22525 = ~n31179 ;
  assign y22526 = ~n31161 ;
  assign y22527 = ~n34737 ;
  assign y22528 = ~1'b0 ;
  assign y22529 = ~1'b0 ;
  assign y22530 = ~n14073 ;
  assign y22531 = n34743 ;
  assign y22532 = ~n34744 ;
  assign y22533 = ~n34745 ;
  assign y22534 = n34747 ;
  assign y22535 = ~n34751 ;
  assign y22536 = ~1'b0 ;
  assign y22537 = n34752 ;
  assign y22538 = ~n13491 ;
  assign y22539 = n34754 ;
  assign y22540 = 1'b0 ;
  assign y22541 = ~1'b0 ;
  assign y22542 = ~1'b0 ;
  assign y22543 = ~n34761 ;
  assign y22544 = 1'b0 ;
  assign y22545 = n34765 ;
  assign y22546 = ~1'b0 ;
  assign y22547 = ~1'b0 ;
  assign y22548 = ~n33803 ;
  assign y22549 = ~n34767 ;
  assign y22550 = n34768 ;
  assign y22551 = ~n34769 ;
  assign y22552 = n34771 ;
  assign y22553 = ~1'b0 ;
  assign y22554 = ~1'b0 ;
  assign y22555 = ~1'b0 ;
  assign y22556 = ~1'b0 ;
  assign y22557 = ~n34773 ;
  assign y22558 = ~n34776 ;
  assign y22559 = n34778 ;
  assign y22560 = ~1'b0 ;
  assign y22561 = ~1'b0 ;
  assign y22562 = n34779 ;
  assign y22563 = ~1'b0 ;
  assign y22564 = ~n34781 ;
  assign y22565 = ~1'b0 ;
  assign y22566 = n34783 ;
  assign y22567 = ~1'b0 ;
  assign y22568 = ~n34785 ;
  assign y22569 = ~n34787 ;
  assign y22570 = ~n22897 ;
  assign y22571 = ~1'b0 ;
  assign y22572 = ~n34788 ;
  assign y22573 = ~1'b0 ;
  assign y22574 = ~1'b0 ;
  assign y22575 = ~1'b0 ;
  assign y22576 = ~1'b0 ;
  assign y22577 = ~1'b0 ;
  assign y22578 = n30430 ;
  assign y22579 = ~n34792 ;
  assign y22580 = ~n34796 ;
  assign y22581 = ~1'b0 ;
  assign y22582 = n34797 ;
  assign y22583 = ~1'b0 ;
  assign y22584 = ~1'b0 ;
  assign y22585 = 1'b0 ;
  assign y22586 = n34798 ;
  assign y22587 = ~1'b0 ;
  assign y22588 = n34799 ;
  assign y22589 = n34801 ;
  assign y22590 = n34802 ;
  assign y22591 = n34803 ;
  assign y22592 = ~1'b0 ;
  assign y22593 = n34806 ;
  assign y22594 = ~1'b0 ;
  assign y22595 = n24429 ;
  assign y22596 = ~n34810 ;
  assign y22597 = ~1'b0 ;
  assign y22598 = n34811 ;
  assign y22599 = n34812 ;
  assign y22600 = n34814 ;
  assign y22601 = n20804 ;
  assign y22602 = ~1'b0 ;
  assign y22603 = ~1'b0 ;
  assign y22604 = ~n28241 ;
  assign y22605 = ~1'b0 ;
  assign y22606 = n34815 ;
  assign y22607 = n34818 ;
  assign y22608 = n34822 ;
  assign y22609 = ~1'b0 ;
  assign y22610 = n34824 ;
  assign y22611 = n34826 ;
  assign y22612 = ~n34828 ;
  assign y22613 = ~1'b0 ;
  assign y22614 = ~1'b0 ;
  assign y22615 = n34834 ;
  assign y22616 = n34838 ;
  assign y22617 = ~1'b0 ;
  assign y22618 = n34840 ;
  assign y22619 = n34842 ;
  assign y22620 = ~n34844 ;
  assign y22621 = n34848 ;
  assign y22622 = ~1'b0 ;
  assign y22623 = ~n34851 ;
  assign y22624 = n732 ;
  assign y22625 = ~n34852 ;
  assign y22626 = ~n18028 ;
  assign y22627 = n34853 ;
  assign y22628 = n34856 ;
  assign y22629 = ~n34858 ;
  assign y22630 = ~n19966 ;
  assign y22631 = ~1'b0 ;
  assign y22632 = n34860 ;
  assign y22633 = ~n34862 ;
  assign y22634 = ~n34865 ;
  assign y22635 = ~n34866 ;
  assign y22636 = n34872 ;
  assign y22637 = ~n34878 ;
  assign y22638 = ~n34881 ;
  assign y22639 = ~n34882 ;
  assign y22640 = ~n34885 ;
  assign y22641 = n34886 ;
  assign y22642 = ~n34887 ;
  assign y22643 = ~n34888 ;
  assign y22644 = ~1'b0 ;
  assign y22645 = n34890 ;
  assign y22646 = ~n34893 ;
  assign y22647 = ~n34894 ;
  assign y22648 = n13355 ;
  assign y22649 = ~n13833 ;
  assign y22650 = n34895 ;
  assign y22651 = ~1'b0 ;
  assign y22652 = n34899 ;
  assign y22653 = ~n25467 ;
  assign y22654 = ~1'b0 ;
  assign y22655 = ~1'b0 ;
  assign y22656 = n34901 ;
  assign y22657 = 1'b0 ;
  assign y22658 = ~1'b0 ;
  assign y22659 = ~1'b0 ;
  assign y22660 = ~1'b0 ;
  assign y22661 = ~n34906 ;
  assign y22662 = ~n34908 ;
  assign y22663 = ~n34909 ;
  assign y22664 = ~n34910 ;
  assign y22665 = ~1'b0 ;
  assign y22666 = ~n34916 ;
  assign y22667 = ~1'b0 ;
  assign y22668 = ~n34921 ;
  assign y22669 = ~1'b0 ;
  assign y22670 = n34924 ;
  assign y22671 = ~n34926 ;
  assign y22672 = n34927 ;
  assign y22673 = ~n34929 ;
  assign y22674 = n4236 ;
  assign y22675 = ~n34932 ;
  assign y22676 = ~n34937 ;
  assign y22677 = ~n34938 ;
  assign y22678 = ~n17507 ;
  assign y22679 = 1'b0 ;
  assign y22680 = ~n34940 ;
  assign y22681 = ~n34943 ;
  assign y22682 = ~1'b0 ;
  assign y22683 = n34947 ;
  assign y22684 = ~n34948 ;
  assign y22685 = ~1'b0 ;
  assign y22686 = ~n34952 ;
  assign y22687 = n34955 ;
  assign y22688 = n34958 ;
  assign y22689 = 1'b0 ;
  assign y22690 = ~n34959 ;
  assign y22691 = ~n34964 ;
  assign y22692 = ~n34966 ;
  assign y22693 = n34967 ;
  assign y22694 = ~n6258 ;
  assign y22695 = ~1'b0 ;
  assign y22696 = ~1'b0 ;
  assign y22697 = n34968 ;
  assign y22698 = ~1'b0 ;
  assign y22699 = ~1'b0 ;
  assign y22700 = ~n34970 ;
  assign y22701 = ~1'b0 ;
  assign y22702 = n10168 ;
  assign y22703 = ~1'b0 ;
  assign y22704 = n34973 ;
  assign y22705 = n10997 ;
  assign y22706 = ~n34976 ;
  assign y22707 = n13807 ;
  assign y22708 = n34977 ;
  assign y22709 = ~n34979 ;
  assign y22710 = ~1'b0 ;
  assign y22711 = ~n34980 ;
  assign y22712 = ~n34982 ;
  assign y22713 = n34983 ;
  assign y22714 = ~1'b0 ;
  assign y22715 = n34984 ;
  assign y22716 = ~1'b0 ;
  assign y22717 = ~n34986 ;
  assign y22718 = ~1'b0 ;
  assign y22719 = n34992 ;
  assign y22720 = ~n34998 ;
  assign y22721 = ~1'b0 ;
  assign y22722 = ~n35001 ;
  assign y22723 = n35003 ;
  assign y22724 = ~n35005 ;
  assign y22725 = ~n35006 ;
  assign y22726 = ~1'b0 ;
  assign y22727 = ~n35008 ;
  assign y22728 = ~1'b0 ;
  assign y22729 = n35010 ;
  assign y22730 = n35012 ;
  assign y22731 = ~n35015 ;
  assign y22732 = n35016 ;
  assign y22733 = ~1'b0 ;
  assign y22734 = n35020 ;
  assign y22735 = ~n35022 ;
  assign y22736 = n2741 ;
  assign y22737 = ~1'b0 ;
  assign y22738 = ~1'b0 ;
  assign y22739 = ~n35023 ;
  assign y22740 = ~1'b0 ;
  assign y22741 = ~n4039 ;
  assign y22742 = n30554 ;
  assign y22743 = ~n35025 ;
  assign y22744 = ~1'b0 ;
  assign y22745 = ~1'b0 ;
  assign y22746 = n35028 ;
  assign y22747 = ~1'b0 ;
  assign y22748 = ~n35032 ;
  assign y22749 = ~n35033 ;
  assign y22750 = ~1'b0 ;
  assign y22751 = ~n35037 ;
  assign y22752 = ~n35038 ;
  assign y22753 = ~1'b0 ;
  assign y22754 = ~n35041 ;
  assign y22755 = n14759 ;
  assign y22756 = ~n35043 ;
  assign y22757 = n35044 ;
  assign y22758 = ~n35046 ;
  assign y22759 = ~n35048 ;
  assign y22760 = ~n35049 ;
  assign y22761 = ~n35050 ;
  assign y22762 = n35052 ;
  assign y22763 = n35056 ;
  assign y22764 = n35059 ;
  assign y22765 = ~1'b0 ;
  assign y22766 = ~1'b0 ;
  assign y22767 = ~n35061 ;
  assign y22768 = n35065 ;
  assign y22769 = ~n35069 ;
  assign y22770 = ~n2685 ;
  assign y22771 = ~1'b0 ;
  assign y22772 = ~n35076 ;
  assign y22773 = ~1'b0 ;
  assign y22774 = ~n35078 ;
  assign y22775 = n33633 ;
  assign y22776 = ~1'b0 ;
  assign y22777 = ~n35082 ;
  assign y22778 = ~n35083 ;
  assign y22779 = ~1'b0 ;
  assign y22780 = ~n35085 ;
  assign y22781 = ~n35088 ;
  assign y22782 = n27806 ;
  assign y22783 = n35091 ;
  assign y22784 = ~n27172 ;
  assign y22785 = ~1'b0 ;
  assign y22786 = ~n35092 ;
  assign y22787 = ~1'b0 ;
  assign y22788 = ~1'b0 ;
  assign y22789 = n35094 ;
  assign y22790 = n35096 ;
  assign y22791 = 1'b0 ;
  assign y22792 = ~1'b0 ;
  assign y22793 = ~1'b0 ;
  assign y22794 = n35097 ;
  assign y22795 = n35099 ;
  assign y22796 = n35100 ;
  assign y22797 = n35101 ;
  assign y22798 = ~n35104 ;
  assign y22799 = ~1'b0 ;
  assign y22800 = ~n35105 ;
  assign y22801 = ~n35110 ;
  assign y22802 = ~n35112 ;
  assign y22803 = n35117 ;
  assign y22804 = ~1'b0 ;
  assign y22805 = ~n35121 ;
  assign y22806 = 1'b0 ;
  assign y22807 = ~1'b0 ;
  assign y22808 = n35127 ;
  assign y22809 = ~n35128 ;
  assign y22810 = ~n35129 ;
  assign y22811 = n35137 ;
  assign y22812 = n35139 ;
  assign y22813 = ~n35144 ;
  assign y22814 = ~n35145 ;
  assign y22815 = ~1'b0 ;
  assign y22816 = n35146 ;
  assign y22817 = ~n35148 ;
  assign y22818 = n4955 ;
  assign y22819 = ~n35149 ;
  assign y22820 = ~n35152 ;
  assign y22821 = n35154 ;
  assign y22822 = n35155 ;
  assign y22823 = ~n35158 ;
  assign y22824 = ~1'b0 ;
  assign y22825 = n35163 ;
  assign y22826 = ~1'b0 ;
  assign y22827 = ~1'b0 ;
  assign y22828 = n35166 ;
  assign y22829 = ~n22722 ;
  assign y22830 = ~1'b0 ;
  assign y22831 = ~n35167 ;
  assign y22832 = ~n35168 ;
  assign y22833 = ~1'b0 ;
  assign y22834 = ~1'b0 ;
  assign y22835 = n35170 ;
  assign y22836 = ~1'b0 ;
  assign y22837 = n35175 ;
  assign y22838 = ~1'b0 ;
  assign y22839 = ~1'b0 ;
  assign y22840 = ~n35176 ;
  assign y22841 = ~n35177 ;
  assign y22842 = ~1'b0 ;
  assign y22843 = ~n35180 ;
  assign y22844 = ~1'b0 ;
  assign y22845 = ~n35183 ;
  assign y22846 = n35185 ;
  assign y22847 = ~n35186 ;
  assign y22848 = ~1'b0 ;
  assign y22849 = ~1'b0 ;
  assign y22850 = n34955 ;
  assign y22851 = 1'b0 ;
  assign y22852 = n35187 ;
  assign y22853 = ~n35190 ;
  assign y22854 = ~1'b0 ;
  assign y22855 = ~n35193 ;
  assign y22856 = ~n35194 ;
  assign y22857 = ~n35198 ;
  assign y22858 = ~n35200 ;
  assign y22859 = n35203 ;
  assign y22860 = 1'b0 ;
  assign y22861 = ~n35204 ;
  assign y22862 = ~1'b0 ;
  assign y22863 = ~n31449 ;
  assign y22864 = ~n35207 ;
  assign y22865 = n35209 ;
  assign y22866 = ~1'b0 ;
  assign y22867 = ~1'b0 ;
  assign y22868 = n35215 ;
  assign y22869 = n35220 ;
  assign y22870 = n3781 ;
  assign y22871 = n17048 ;
  assign y22872 = n35221 ;
  assign y22873 = ~n35223 ;
  assign y22874 = ~1'b0 ;
  assign y22875 = ~1'b0 ;
  assign y22876 = ~n35225 ;
  assign y22877 = n35227 ;
  assign y22878 = ~1'b0 ;
  assign y22879 = n35228 ;
  assign y22880 = n35229 ;
  assign y22881 = ~1'b0 ;
  assign y22882 = 1'b0 ;
  assign y22883 = n35231 ;
  assign y22884 = n35232 ;
  assign y22885 = ~n35233 ;
  assign y22886 = ~n35235 ;
  assign y22887 = ~n35238 ;
  assign y22888 = ~n35240 ;
  assign y22889 = ~1'b0 ;
  assign y22890 = ~n35245 ;
  assign y22891 = ~1'b0 ;
  assign y22892 = ~n35246 ;
  assign y22893 = ~1'b0 ;
  assign y22894 = ~n35247 ;
  assign y22895 = n35248 ;
  assign y22896 = ~1'b0 ;
  assign y22897 = n35250 ;
  assign y22898 = ~n8937 ;
  assign y22899 = n35251 ;
  assign y22900 = ~1'b0 ;
  assign y22901 = ~1'b0 ;
  assign y22902 = 1'b0 ;
  assign y22903 = ~n35253 ;
  assign y22904 = ~1'b0 ;
  assign y22905 = ~1'b0 ;
  assign y22906 = ~1'b0 ;
  assign y22907 = ~1'b0 ;
  assign y22908 = n35255 ;
  assign y22909 = n35261 ;
  assign y22910 = ~1'b0 ;
  assign y22911 = ~n35267 ;
  assign y22912 = ~1'b0 ;
  assign y22913 = ~n35270 ;
  assign y22914 = n35273 ;
  assign y22915 = ~n35275 ;
  assign y22916 = ~1'b0 ;
  assign y22917 = ~1'b0 ;
  assign y22918 = n3635 ;
  assign y22919 = n35279 ;
  assign y22920 = ~1'b0 ;
  assign y22921 = ~n35281 ;
  assign y22922 = ~n14921 ;
  assign y22923 = ~n35282 ;
  assign y22924 = n35285 ;
  assign y22925 = ~n35290 ;
  assign y22926 = ~n35291 ;
  assign y22927 = ~1'b0 ;
  assign y22928 = ~1'b0 ;
  assign y22929 = ~n35294 ;
  assign y22930 = ~n35297 ;
  assign y22931 = n35300 ;
  assign y22932 = ~1'b0 ;
  assign y22933 = ~1'b0 ;
  assign y22934 = ~1'b0 ;
  assign y22935 = ~n35304 ;
  assign y22936 = ~n35305 ;
  assign y22937 = ~n6068 ;
  assign y22938 = n35306 ;
  assign y22939 = n35313 ;
  assign y22940 = ~1'b0 ;
  assign y22941 = ~n35314 ;
  assign y22942 = ~n35316 ;
  assign y22943 = ~1'b0 ;
  assign y22944 = ~n7679 ;
  assign y22945 = ~n35318 ;
  assign y22946 = ~n35320 ;
  assign y22947 = n35323 ;
  assign y22948 = ~n35324 ;
  assign y22949 = n35334 ;
  assign y22950 = ~1'b0 ;
  assign y22951 = ~1'b0 ;
  assign y22952 = n35335 ;
  assign y22953 = n35337 ;
  assign y22954 = ~n35338 ;
  assign y22955 = ~n35341 ;
  assign y22956 = ~n35343 ;
  assign y22957 = ~n35344 ;
  assign y22958 = ~n35345 ;
  assign y22959 = ~n35346 ;
  assign y22960 = ~1'b0 ;
  assign y22961 = ~1'b0 ;
  assign y22962 = ~n35348 ;
  assign y22963 = ~n35350 ;
  assign y22964 = ~1'b0 ;
  assign y22965 = ~n35352 ;
  assign y22966 = n35353 ;
  assign y22967 = ~n35354 ;
  assign y22968 = ~1'b0 ;
  assign y22969 = n35356 ;
  assign y22970 = ~n35357 ;
  assign y22971 = ~1'b0 ;
  assign y22972 = ~n35361 ;
  assign y22973 = ~1'b0 ;
  assign y22974 = ~n35364 ;
  assign y22975 = n35365 ;
  assign y22976 = ~n35367 ;
  assign y22977 = ~1'b0 ;
  assign y22978 = n753 ;
  assign y22979 = n35370 ;
  assign y22980 = n35373 ;
  assign y22981 = ~1'b0 ;
  assign y22982 = ~n35376 ;
  assign y22983 = ~n35380 ;
  assign y22984 = 1'b0 ;
  assign y22985 = n20511 ;
  assign y22986 = n14311 ;
  assign y22987 = ~1'b0 ;
  assign y22988 = n35381 ;
  assign y22989 = ~n35383 ;
  assign y22990 = ~1'b0 ;
  assign y22991 = ~n35386 ;
  assign y22992 = ~1'b0 ;
  assign y22993 = ~1'b0 ;
  assign y22994 = n35387 ;
  assign y22995 = n35390 ;
  assign y22996 = n35396 ;
  assign y22997 = n35398 ;
  assign y22998 = n35399 ;
  assign y22999 = n35400 ;
  assign y23000 = ~1'b0 ;
  assign y23001 = ~n35401 ;
  assign y23002 = ~n35403 ;
  assign y23003 = n35404 ;
  assign y23004 = n35406 ;
  assign y23005 = ~1'b0 ;
  assign y23006 = ~n35407 ;
  assign y23007 = n35408 ;
  assign y23008 = ~n31101 ;
  assign y23009 = ~n35410 ;
  assign y23010 = ~n21333 ;
  assign y23011 = ~n35411 ;
  assign y23012 = ~n35413 ;
  assign y23013 = n35418 ;
  assign y23014 = ~n26520 ;
  assign y23015 = n35421 ;
  assign y23016 = ~1'b0 ;
  assign y23017 = ~n9765 ;
  assign y23018 = ~1'b0 ;
  assign y23019 = ~n35422 ;
  assign y23020 = ~1'b0 ;
  assign y23021 = n35423 ;
  assign y23022 = ~1'b0 ;
  assign y23023 = n35425 ;
  assign y23024 = ~1'b0 ;
  assign y23025 = ~1'b0 ;
  assign y23026 = n35427 ;
  assign y23027 = ~1'b0 ;
  assign y23028 = n35432 ;
  assign y23029 = ~1'b0 ;
  assign y23030 = n35433 ;
  assign y23031 = n17361 ;
  assign y23032 = ~1'b0 ;
  assign y23033 = ~1'b0 ;
  assign y23034 = ~n35436 ;
  assign y23035 = ~1'b0 ;
  assign y23036 = ~n35438 ;
  assign y23037 = ~1'b0 ;
  assign y23038 = n35439 ;
  assign y23039 = ~n35442 ;
  assign y23040 = n35443 ;
  assign y23041 = n35445 ;
  assign y23042 = ~n35446 ;
  assign y23043 = ~1'b0 ;
  assign y23044 = n35448 ;
  assign y23045 = n35456 ;
  assign y23046 = n35457 ;
  assign y23047 = ~1'b0 ;
  assign y23048 = ~n35458 ;
  assign y23049 = ~1'b0 ;
  assign y23050 = n35460 ;
  assign y23051 = ~n35465 ;
  assign y23052 = ~1'b0 ;
  assign y23053 = ~n28539 ;
  assign y23054 = ~n35466 ;
  assign y23055 = ~1'b0 ;
  assign y23056 = ~n6064 ;
  assign y23057 = ~1'b0 ;
  assign y23058 = ~n35467 ;
  assign y23059 = ~n21736 ;
  assign y23060 = ~n35469 ;
  assign y23061 = n35473 ;
  assign y23062 = n35474 ;
  assign y23063 = n35476 ;
  assign y23064 = n35477 ;
  assign y23065 = n35479 ;
  assign y23066 = ~n27780 ;
  assign y23067 = ~1'b0 ;
  assign y23068 = n35480 ;
  assign y23069 = ~n10887 ;
  assign y23070 = ~n35481 ;
  assign y23071 = ~n35484 ;
  assign y23072 = ~1'b0 ;
  assign y23073 = ~n35485 ;
  assign y23074 = n35487 ;
  assign y23075 = ~n35488 ;
  assign y23076 = ~n35490 ;
  assign y23077 = ~1'b0 ;
  assign y23078 = n35491 ;
  assign y23079 = ~n35492 ;
  assign y23080 = ~1'b0 ;
  assign y23081 = ~1'b0 ;
  assign y23082 = n35493 ;
  assign y23083 = n35494 ;
  assign y23084 = n35497 ;
  assign y23085 = ~1'b0 ;
  assign y23086 = ~1'b0 ;
  assign y23087 = ~n35499 ;
  assign y23088 = 1'b0 ;
  assign y23089 = n35503 ;
  assign y23090 = ~n35505 ;
  assign y23091 = ~1'b0 ;
  assign y23092 = ~n35506 ;
  assign y23093 = n35507 ;
  assign y23094 = ~1'b0 ;
  assign y23095 = ~1'b0 ;
  assign y23096 = ~1'b0 ;
  assign y23097 = n35509 ;
  assign y23098 = n35511 ;
  assign y23099 = ~n35512 ;
  assign y23100 = ~n35514 ;
  assign y23101 = n35515 ;
  assign y23102 = ~n35516 ;
  assign y23103 = n35517 ;
  assign y23104 = ~1'b0 ;
  assign y23105 = n35518 ;
  assign y23106 = n35520 ;
  assign y23107 = ~n35527 ;
  assign y23108 = n35529 ;
  assign y23109 = n35533 ;
  assign y23110 = ~n25588 ;
  assign y23111 = ~n35534 ;
  assign y23112 = n35536 ;
  assign y23113 = ~n15028 ;
  assign y23114 = ~1'b0 ;
  assign y23115 = ~n30269 ;
  assign y23116 = n31868 ;
  assign y23117 = n35540 ;
  assign y23118 = 1'b0 ;
  assign y23119 = ~1'b0 ;
  assign y23120 = 1'b0 ;
  assign y23121 = ~1'b0 ;
  assign y23122 = ~n35544 ;
  assign y23123 = 1'b0 ;
  assign y23124 = ~n35545 ;
  assign y23125 = 1'b0 ;
  assign y23126 = ~n35547 ;
  assign y23127 = ~1'b0 ;
  assign y23128 = 1'b0 ;
  assign y23129 = n35548 ;
  assign y23130 = 1'b0 ;
  assign y23131 = ~n35553 ;
  assign y23132 = ~n13025 ;
  assign y23133 = ~1'b0 ;
  assign y23134 = n35554 ;
  assign y23135 = n6791 ;
  assign y23136 = ~n561 ;
  assign y23137 = ~n35555 ;
  assign y23138 = ~1'b0 ;
  assign y23139 = ~n35557 ;
  assign y23140 = ~1'b0 ;
  assign y23141 = ~1'b0 ;
  assign y23142 = ~n35562 ;
  assign y23143 = ~n25023 ;
  assign y23144 = ~n19957 ;
  assign y23145 = n4888 ;
  assign y23146 = n35564 ;
  assign y23147 = ~1'b0 ;
  assign y23148 = ~1'b0 ;
  assign y23149 = ~1'b0 ;
  assign y23150 = x202 ;
  assign y23151 = ~n35565 ;
  assign y23152 = ~1'b0 ;
  assign y23153 = ~1'b0 ;
  assign y23154 = ~n3891 ;
  assign y23155 = ~n35566 ;
  assign y23156 = n35567 ;
  assign y23157 = n35568 ;
  assign y23158 = ~n35570 ;
  assign y23159 = ~1'b0 ;
  assign y23160 = n35574 ;
  assign y23161 = ~1'b0 ;
  assign y23162 = ~1'b0 ;
  assign y23163 = ~n35576 ;
  assign y23164 = n35577 ;
  assign y23165 = ~n35578 ;
  assign y23166 = ~1'b0 ;
  assign y23167 = ~1'b0 ;
  assign y23168 = ~1'b0 ;
  assign y23169 = ~n35580 ;
  assign y23170 = ~n1508 ;
  assign y23171 = ~n35581 ;
  assign y23172 = n35582 ;
  assign y23173 = n35584 ;
  assign y23174 = n35588 ;
  assign y23175 = ~n35589 ;
  assign y23176 = ~n35590 ;
  assign y23177 = n35592 ;
  assign y23178 = ~n35597 ;
  assign y23179 = ~1'b0 ;
  assign y23180 = ~n24663 ;
  assign y23181 = ~n35601 ;
  assign y23182 = n35604 ;
  assign y23183 = n35605 ;
  assign y23184 = n35607 ;
  assign y23185 = n35611 ;
  assign y23186 = ~n35612 ;
  assign y23187 = ~1'b0 ;
  assign y23188 = ~1'b0 ;
  assign y23189 = ~1'b0 ;
  assign y23190 = ~n7953 ;
  assign y23191 = 1'b0 ;
  assign y23192 = ~1'b0 ;
  assign y23193 = n35620 ;
  assign y23194 = ~n35621 ;
  assign y23195 = ~n35628 ;
  assign y23196 = ~n35631 ;
  assign y23197 = ~1'b0 ;
  assign y23198 = ~1'b0 ;
  assign y23199 = ~1'b0 ;
  assign y23200 = ~1'b0 ;
  assign y23201 = ~n15829 ;
  assign y23202 = ~n35633 ;
  assign y23203 = ~1'b0 ;
  assign y23204 = ~1'b0 ;
  assign y23205 = ~1'b0 ;
  assign y23206 = n35635 ;
  assign y23207 = ~n35637 ;
  assign y23208 = ~n35638 ;
  assign y23209 = ~n35642 ;
  assign y23210 = ~n35644 ;
  assign y23211 = ~1'b0 ;
  assign y23212 = ~1'b0 ;
  assign y23213 = n35648 ;
  assign y23214 = ~1'b0 ;
  assign y23215 = 1'b0 ;
  assign y23216 = ~n35650 ;
  assign y23217 = ~n35652 ;
  assign y23218 = ~n35653 ;
  assign y23219 = ~1'b0 ;
  assign y23220 = ~1'b0 ;
  assign y23221 = ~n35654 ;
  assign y23222 = ~1'b0 ;
  assign y23223 = ~1'b0 ;
  assign y23224 = n15720 ;
  assign y23225 = n35655 ;
  assign y23226 = ~n6689 ;
  assign y23227 = ~1'b0 ;
  assign y23228 = ~1'b0 ;
  assign y23229 = ~n35657 ;
  assign y23230 = 1'b0 ;
  assign y23231 = ~1'b0 ;
  assign y23232 = ~1'b0 ;
  assign y23233 = ~n35661 ;
  assign y23234 = ~n35662 ;
  assign y23235 = ~n29920 ;
  assign y23236 = ~n35666 ;
  assign y23237 = ~n35671 ;
  assign y23238 = 1'b0 ;
  assign y23239 = ~1'b0 ;
  assign y23240 = ~1'b0 ;
  assign y23241 = ~1'b0 ;
  assign y23242 = ~n35675 ;
  assign y23243 = ~1'b0 ;
  assign y23244 = ~n9771 ;
  assign y23245 = ~1'b0 ;
  assign y23246 = ~n35677 ;
  assign y23247 = ~n35678 ;
  assign y23248 = n956 ;
  assign y23249 = ~n35682 ;
  assign y23250 = ~1'b0 ;
  assign y23251 = n35685 ;
  assign y23252 = ~1'b0 ;
  assign y23253 = ~n35686 ;
  assign y23254 = n11914 ;
  assign y23255 = n35688 ;
  assign y23256 = ~n35690 ;
  assign y23257 = ~n35693 ;
  assign y23258 = ~1'b0 ;
  assign y23259 = ~1'b0 ;
  assign y23260 = ~1'b0 ;
  assign y23261 = ~1'b0 ;
  assign y23262 = ~n35694 ;
  assign y23263 = ~n35695 ;
  assign y23264 = ~1'b0 ;
  assign y23265 = n35696 ;
  assign y23266 = ~n35697 ;
  assign y23267 = ~n35702 ;
  assign y23268 = ~n14769 ;
  assign y23269 = n10346 ;
  assign y23270 = ~1'b0 ;
  assign y23271 = ~1'b0 ;
  assign y23272 = ~1'b0 ;
  assign y23273 = ~n35703 ;
  assign y23274 = ~1'b0 ;
  assign y23275 = ~1'b0 ;
  assign y23276 = ~n35704 ;
  assign y23277 = n35706 ;
  assign y23278 = ~1'b0 ;
  assign y23279 = n35707 ;
  assign y23280 = ~1'b0 ;
  assign y23281 = ~n35711 ;
  assign y23282 = ~1'b0 ;
  assign y23283 = ~1'b0 ;
  assign y23284 = ~n35712 ;
  assign y23285 = ~1'b0 ;
  assign y23286 = ~n35713 ;
  assign y23287 = n35714 ;
  assign y23288 = ~1'b0 ;
  assign y23289 = n5776 ;
  assign y23290 = n35718 ;
  assign y23291 = ~1'b0 ;
  assign y23292 = n35720 ;
  assign y23293 = ~1'b0 ;
  assign y23294 = ~1'b0 ;
  assign y23295 = ~1'b0 ;
  assign y23296 = ~n35722 ;
  assign y23297 = ~n35725 ;
  assign y23298 = n35727 ;
  assign y23299 = ~n30114 ;
  assign y23300 = ~1'b0 ;
  assign y23301 = ~1'b0 ;
  assign y23302 = ~n35729 ;
  assign y23303 = ~n35731 ;
  assign y23304 = n35736 ;
  assign y23305 = n35742 ;
  assign y23306 = n35746 ;
  assign y23307 = ~1'b0 ;
  assign y23308 = ~n35748 ;
  assign y23309 = ~1'b0 ;
  assign y23310 = ~1'b0 ;
  assign y23311 = ~1'b0 ;
  assign y23312 = ~1'b0 ;
  assign y23313 = ~1'b0 ;
  assign y23314 = 1'b0 ;
  assign y23315 = ~n35751 ;
  assign y23316 = n35752 ;
  assign y23317 = ~1'b0 ;
  assign y23318 = ~1'b0 ;
  assign y23319 = ~1'b0 ;
  assign y23320 = ~1'b0 ;
  assign y23321 = ~n35758 ;
  assign y23322 = ~1'b0 ;
  assign y23323 = n35761 ;
  assign y23324 = ~n35765 ;
  assign y23325 = ~1'b0 ;
  assign y23326 = 1'b0 ;
  assign y23327 = n35772 ;
  assign y23328 = n35774 ;
  assign y23329 = n35775 ;
  assign y23330 = 1'b0 ;
  assign y23331 = ~1'b0 ;
  assign y23332 = ~1'b0 ;
  assign y23333 = ~1'b0 ;
  assign y23334 = ~n35779 ;
  assign y23335 = ~1'b0 ;
  assign y23336 = ~n35782 ;
  assign y23337 = ~n35784 ;
  assign y23338 = n35785 ;
  assign y23339 = n35786 ;
  assign y23340 = ~n35787 ;
  assign y23341 = ~1'b0 ;
  assign y23342 = ~n35788 ;
  assign y23343 = ~n35790 ;
  assign y23344 = ~n35791 ;
  assign y23345 = ~n35793 ;
  assign y23346 = ~n35798 ;
  assign y23347 = ~1'b0 ;
  assign y23348 = n35799 ;
  assign y23349 = n12548 ;
  assign y23350 = ~n35800 ;
  assign y23351 = ~1'b0 ;
  assign y23352 = n35804 ;
  assign y23353 = n35805 ;
  assign y23354 = ~1'b0 ;
  assign y23355 = n35807 ;
  assign y23356 = ~n35808 ;
  assign y23357 = n35810 ;
  assign y23358 = n20162 ;
  assign y23359 = n15667 ;
  assign y23360 = ~1'b0 ;
  assign y23361 = ~1'b0 ;
  assign y23362 = ~1'b0 ;
  assign y23363 = ~n19138 ;
  assign y23364 = ~1'b0 ;
  assign y23365 = 1'b0 ;
  assign y23366 = n35811 ;
  assign y23367 = ~1'b0 ;
  assign y23368 = ~1'b0 ;
  assign y23369 = ~1'b0 ;
  assign y23370 = ~1'b0 ;
  assign y23371 = ~1'b0 ;
  assign y23372 = ~1'b0 ;
  assign y23373 = n35813 ;
  assign y23374 = n4501 ;
  assign y23375 = n35820 ;
  assign y23376 = n35824 ;
  assign y23377 = n35826 ;
  assign y23378 = n35827 ;
  assign y23379 = ~1'b0 ;
  assign y23380 = ~n35828 ;
  assign y23381 = ~1'b0 ;
  assign y23382 = ~1'b0 ;
  assign y23383 = ~n35829 ;
  assign y23384 = 1'b0 ;
  assign y23385 = 1'b0 ;
  assign y23386 = ~1'b0 ;
  assign y23387 = ~n35832 ;
  assign y23388 = ~n10164 ;
  assign y23389 = n35833 ;
  assign y23390 = ~n35834 ;
  assign y23391 = ~n35835 ;
  assign y23392 = n3364 ;
  assign y23393 = n35837 ;
  assign y23394 = ~1'b0 ;
  assign y23395 = ~n35839 ;
  assign y23396 = ~1'b0 ;
  assign y23397 = ~n35841 ;
  assign y23398 = ~n35843 ;
  assign y23399 = ~1'b0 ;
  assign y23400 = ~n35852 ;
  assign y23401 = 1'b0 ;
  assign y23402 = ~n35853 ;
  assign y23403 = n35855 ;
  assign y23404 = ~n35858 ;
  assign y23405 = n35861 ;
  assign y23406 = n35863 ;
  assign y23407 = n35865 ;
  assign y23408 = ~n26716 ;
  assign y23409 = ~1'b0 ;
  assign y23410 = ~n35867 ;
  assign y23411 = ~n35868 ;
  assign y23412 = ~n35873 ;
  assign y23413 = ~1'b0 ;
  assign y23414 = ~1'b0 ;
  assign y23415 = ~n35874 ;
  assign y23416 = ~n35876 ;
  assign y23417 = n35877 ;
  assign y23418 = ~n35878 ;
  assign y23419 = ~n9329 ;
  assign y23420 = ~n19697 ;
  assign y23421 = ~1'b0 ;
  assign y23422 = ~1'b0 ;
  assign y23423 = ~n35880 ;
  assign y23424 = ~n35881 ;
  assign y23425 = n35883 ;
  assign y23426 = ~1'b0 ;
  assign y23427 = ~1'b0 ;
  assign y23428 = n7882 ;
  assign y23429 = ~n35886 ;
  assign y23430 = 1'b0 ;
  assign y23431 = ~n35887 ;
  assign y23432 = ~1'b0 ;
  assign y23433 = ~1'b0 ;
  assign y23434 = ~1'b0 ;
  assign y23435 = ~1'b0 ;
  assign y23436 = n34745 ;
  assign y23437 = n35888 ;
  assign y23438 = ~1'b0 ;
  assign y23439 = ~n35889 ;
  assign y23440 = n35890 ;
  assign y23441 = n35891 ;
  assign y23442 = ~1'b0 ;
  assign y23443 = ~1'b0 ;
  assign y23444 = ~n35893 ;
  assign y23445 = ~n10702 ;
  assign y23446 = ~1'b0 ;
  assign y23447 = ~n35898 ;
  assign y23448 = ~n35901 ;
  assign y23449 = ~1'b0 ;
  assign y23450 = ~n35902 ;
  assign y23451 = n35904 ;
  assign y23452 = ~n35905 ;
  assign y23453 = ~n35906 ;
  assign y23454 = ~n35907 ;
  assign y23455 = ~n1345 ;
  assign y23456 = n35909 ;
  assign y23457 = n35910 ;
  assign y23458 = ~n35915 ;
  assign y23459 = n35919 ;
  assign y23460 = 1'b0 ;
  assign y23461 = n35920 ;
  assign y23462 = ~1'b0 ;
  assign y23463 = 1'b0 ;
  assign y23464 = ~1'b0 ;
  assign y23465 = ~1'b0 ;
  assign y23466 = n35925 ;
  assign y23467 = ~n35927 ;
  assign y23468 = ~1'b0 ;
  assign y23469 = ~1'b0 ;
  assign y23470 = ~n35932 ;
  assign y23471 = ~n35934 ;
  assign y23472 = n35937 ;
  assign y23473 = ~1'b0 ;
  assign y23474 = n35938 ;
  assign y23475 = ~1'b0 ;
  assign y23476 = n35939 ;
  assign y23477 = ~1'b0 ;
  assign y23478 = ~1'b0 ;
  assign y23479 = ~n35940 ;
  assign y23480 = ~n2342 ;
  assign y23481 = ~n35942 ;
  assign y23482 = n35948 ;
  assign y23483 = ~n35954 ;
  assign y23484 = ~n35955 ;
  assign y23485 = n35957 ;
  assign y23486 = ~1'b0 ;
  assign y23487 = ~1'b0 ;
  assign y23488 = 1'b0 ;
  assign y23489 = n35958 ;
  assign y23490 = n3756 ;
  assign y23491 = ~1'b0 ;
  assign y23492 = ~n5396 ;
  assign y23493 = ~1'b0 ;
  assign y23494 = ~n35959 ;
  assign y23495 = ~1'b0 ;
  assign y23496 = ~1'b0 ;
  assign y23497 = ~1'b0 ;
  assign y23498 = ~n35961 ;
  assign y23499 = n35962 ;
  assign y23500 = ~n35964 ;
  assign y23501 = n35965 ;
  assign y23502 = n35968 ;
  assign y23503 = ~n35969 ;
  assign y23504 = n35970 ;
  assign y23505 = ~n35972 ;
  assign y23506 = n35977 ;
  assign y23507 = ~n1402 ;
  assign y23508 = ~1'b0 ;
  assign y23509 = ~n35980 ;
  assign y23510 = n35982 ;
  assign y23511 = n35985 ;
  assign y23512 = ~1'b0 ;
  assign y23513 = n8334 ;
  assign y23514 = 1'b0 ;
  assign y23515 = n9508 ;
  assign y23516 = ~1'b0 ;
  assign y23517 = 1'b0 ;
  assign y23518 = ~n35986 ;
  assign y23519 = n35988 ;
  assign y23520 = n35989 ;
  assign y23521 = n35990 ;
  assign y23522 = n35993 ;
  assign y23523 = ~n35994 ;
  assign y23524 = n35995 ;
  assign y23525 = ~1'b0 ;
  assign y23526 = n6428 ;
  assign y23527 = n21397 ;
  assign y23528 = ~1'b0 ;
  assign y23529 = ~1'b0 ;
  assign y23530 = ~n35996 ;
  assign y23531 = n35998 ;
  assign y23532 = n35999 ;
  assign y23533 = n36001 ;
  assign y23534 = ~1'b0 ;
  assign y23535 = n36002 ;
  assign y23536 = ~1'b0 ;
  assign y23537 = ~1'b0 ;
  assign y23538 = n36003 ;
  assign y23539 = ~n6371 ;
  assign y23540 = n4257 ;
  assign y23541 = n36004 ;
  assign y23542 = ~1'b0 ;
  assign y23543 = n36006 ;
  assign y23544 = ~n13297 ;
  assign y23545 = ~n36008 ;
  assign y23546 = ~n15033 ;
  assign y23547 = ~1'b0 ;
  assign y23548 = ~1'b0 ;
  assign y23549 = ~n36009 ;
  assign y23550 = n36011 ;
  assign y23551 = ~n36012 ;
  assign y23552 = ~n36014 ;
  assign y23553 = n36016 ;
  assign y23554 = n36020 ;
  assign y23555 = ~n36023 ;
  assign y23556 = ~1'b0 ;
  assign y23557 = n36027 ;
  assign y23558 = ~1'b0 ;
  assign y23559 = ~n36028 ;
  assign y23560 = ~1'b0 ;
  assign y23561 = n36030 ;
  assign y23562 = n36031 ;
  assign y23563 = ~1'b0 ;
  assign y23564 = ~n36033 ;
  assign y23565 = n36036 ;
  assign y23566 = ~n36037 ;
  assign y23567 = ~n36038 ;
  assign y23568 = n36039 ;
  assign y23569 = n36040 ;
  assign y23570 = ~1'b0 ;
  assign y23571 = ~n36042 ;
  assign y23572 = ~n36043 ;
  assign y23573 = ~n36045 ;
  assign y23574 = ~1'b0 ;
  assign y23575 = ~1'b0 ;
  assign y23576 = n36047 ;
  assign y23577 = ~n36050 ;
  assign y23578 = ~1'b0 ;
  assign y23579 = n36051 ;
  assign y23580 = ~n36053 ;
  assign y23581 = n36054 ;
  assign y23582 = 1'b0 ;
  assign y23583 = ~n36058 ;
  assign y23584 = n36060 ;
  assign y23585 = ~1'b0 ;
  assign y23586 = ~1'b0 ;
  assign y23587 = ~n36061 ;
  assign y23588 = 1'b0 ;
  assign y23589 = n36063 ;
  assign y23590 = ~n36065 ;
  assign y23591 = n24484 ;
  assign y23592 = ~1'b0 ;
  assign y23593 = ~n36067 ;
  assign y23594 = ~1'b0 ;
  assign y23595 = ~1'b0 ;
  assign y23596 = n36069 ;
  assign y23597 = ~n19831 ;
  assign y23598 = n36070 ;
  assign y23599 = ~1'b0 ;
  assign y23600 = ~1'b0 ;
  assign y23601 = ~1'b0 ;
  assign y23602 = ~n36073 ;
  assign y23603 = n36075 ;
  assign y23604 = n36078 ;
  assign y23605 = ~n36082 ;
  assign y23606 = ~n36085 ;
  assign y23607 = ~n36088 ;
  assign y23608 = ~n36091 ;
  assign y23609 = n36092 ;
  assign y23610 = n36094 ;
  assign y23611 = ~1'b0 ;
  assign y23612 = ~n36096 ;
  assign y23613 = n36097 ;
  assign y23614 = n36099 ;
  assign y23615 = ~1'b0 ;
  assign y23616 = ~1'b0 ;
  assign y23617 = ~1'b0 ;
  assign y23618 = n36103 ;
  assign y23619 = ~1'b0 ;
  assign y23620 = n36104 ;
  assign y23621 = ~n36106 ;
  assign y23622 = ~1'b0 ;
  assign y23623 = ~1'b0 ;
  assign y23624 = n36107 ;
  assign y23625 = ~n36110 ;
  assign y23626 = n36117 ;
  assign y23627 = n36119 ;
  assign y23628 = n36121 ;
  assign y23629 = ~n36122 ;
  assign y23630 = ~n36123 ;
  assign y23631 = ~n36125 ;
  assign y23632 = ~1'b0 ;
  assign y23633 = ~n36126 ;
  assign y23634 = ~n36130 ;
  assign y23635 = ~1'b0 ;
  assign y23636 = ~n36133 ;
  assign y23637 = n36137 ;
  assign y23638 = n36138 ;
  assign y23639 = n25990 ;
  assign y23640 = ~n36139 ;
  assign y23641 = ~1'b0 ;
  assign y23642 = ~1'b0 ;
  assign y23643 = ~1'b0 ;
  assign y23644 = ~1'b0 ;
  assign y23645 = n36143 ;
  assign y23646 = n19794 ;
  assign y23647 = ~1'b0 ;
  assign y23648 = ~1'b0 ;
  assign y23649 = n36147 ;
  assign y23650 = ~n8718 ;
  assign y23651 = n34854 ;
  assign y23652 = ~1'b0 ;
  assign y23653 = ~n36148 ;
  assign y23654 = ~n36149 ;
  assign y23655 = ~1'b0 ;
  assign y23656 = ~1'b0 ;
  assign y23657 = ~n36150 ;
  assign y23658 = ~1'b0 ;
  assign y23659 = n36160 ;
  assign y23660 = ~1'b0 ;
  assign y23661 = ~n28057 ;
  assign y23662 = ~1'b0 ;
  assign y23663 = ~n36161 ;
  assign y23664 = ~n36162 ;
  assign y23665 = ~1'b0 ;
  assign y23666 = ~n36166 ;
  assign y23667 = ~1'b0 ;
  assign y23668 = ~1'b0 ;
  assign y23669 = ~1'b0 ;
  assign y23670 = n15050 ;
  assign y23671 = n36167 ;
  assign y23672 = ~1'b0 ;
  assign y23673 = n36169 ;
  assign y23674 = ~n36170 ;
  assign y23675 = ~1'b0 ;
  assign y23676 = n36173 ;
  assign y23677 = ~n36175 ;
  assign y23678 = ~n36176 ;
  assign y23679 = ~1'b0 ;
  assign y23680 = ~n36177 ;
  assign y23681 = ~n36186 ;
  assign y23682 = ~1'b0 ;
  assign y23683 = n36187 ;
  assign y23684 = n36189 ;
  assign y23685 = ~1'b0 ;
  assign y23686 = ~1'b0 ;
  assign y23687 = n36190 ;
  assign y23688 = ~n36191 ;
  assign y23689 = ~n36196 ;
  assign y23690 = 1'b0 ;
  assign y23691 = ~1'b0 ;
  assign y23692 = 1'b0 ;
  assign y23693 = n36197 ;
  assign y23694 = n8580 ;
  assign y23695 = n36199 ;
  assign y23696 = ~n36205 ;
  assign y23697 = ~1'b0 ;
  assign y23698 = n36206 ;
  assign y23699 = ~n36210 ;
  assign y23700 = ~n36212 ;
  assign y23701 = ~n14224 ;
  assign y23702 = ~1'b0 ;
  assign y23703 = ~n36215 ;
  assign y23704 = n36216 ;
  assign y23705 = ~1'b0 ;
  assign y23706 = ~n36217 ;
  assign y23707 = n36218 ;
  assign y23708 = n36219 ;
  assign y23709 = ~n36221 ;
  assign y23710 = n20312 ;
  assign y23711 = ~n36222 ;
  assign y23712 = ~n36224 ;
  assign y23713 = ~1'b0 ;
  assign y23714 = n36225 ;
  assign y23715 = ~n36226 ;
  assign y23716 = ~1'b0 ;
  assign y23717 = n36227 ;
  assign y23718 = ~n15312 ;
  assign y23719 = ~n36228 ;
  assign y23720 = ~n644 ;
  assign y23721 = ~n36230 ;
  assign y23722 = ~n36231 ;
  assign y23723 = ~n1192 ;
  assign y23724 = ~n36236 ;
  assign y23725 = ~n5943 ;
  assign y23726 = ~n20959 ;
  assign y23727 = n36238 ;
  assign y23728 = 1'b0 ;
  assign y23729 = ~n36239 ;
  assign y23730 = ~n36241 ;
  assign y23731 = ~n36242 ;
  assign y23732 = ~1'b0 ;
  assign y23733 = ~1'b0 ;
  assign y23734 = n36244 ;
  assign y23735 = n36246 ;
  assign y23736 = ~1'b0 ;
  assign y23737 = n36251 ;
  assign y23738 = n36253 ;
  assign y23739 = ~1'b0 ;
  assign y23740 = ~n36255 ;
  assign y23741 = n15896 ;
  assign y23742 = n36259 ;
  assign y23743 = ~1'b0 ;
  assign y23744 = n36260 ;
  assign y23745 = ~n34346 ;
  assign y23746 = 1'b0 ;
  assign y23747 = ~1'b0 ;
  assign y23748 = ~n36263 ;
  assign y23749 = n36265 ;
  assign y23750 = ~1'b0 ;
  assign y23751 = ~n36267 ;
  assign y23752 = n36270 ;
  assign y23753 = n36272 ;
  assign y23754 = n36273 ;
  assign y23755 = ~1'b0 ;
  assign y23756 = ~1'b0 ;
  assign y23757 = ~1'b0 ;
  assign y23758 = ~1'b0 ;
  assign y23759 = ~1'b0 ;
  assign y23760 = n36275 ;
  assign y23761 = ~1'b0 ;
  assign y23762 = ~n36276 ;
  assign y23763 = ~n36277 ;
  assign y23764 = ~n36278 ;
  assign y23765 = ~1'b0 ;
  assign y23766 = n9221 ;
  assign y23767 = n36281 ;
  assign y23768 = n36284 ;
  assign y23769 = ~n36285 ;
  assign y23770 = n36286 ;
  assign y23771 = n36288 ;
  assign y23772 = ~1'b0 ;
  assign y23773 = ~n25257 ;
  assign y23774 = ~1'b0 ;
  assign y23775 = ~n36292 ;
  assign y23776 = n36293 ;
  assign y23777 = ~n36294 ;
  assign y23778 = n36296 ;
  assign y23779 = n36297 ;
  assign y23780 = n36299 ;
  assign y23781 = ~n36303 ;
  assign y23782 = ~1'b0 ;
  assign y23783 = n2095 ;
  assign y23784 = ~n36304 ;
  assign y23785 = ~n36307 ;
  assign y23786 = ~1'b0 ;
  assign y23787 = ~n36308 ;
  assign y23788 = ~n36312 ;
  assign y23789 = ~n36314 ;
  assign y23790 = ~1'b0 ;
  assign y23791 = ~1'b0 ;
  assign y23792 = ~1'b0 ;
  assign y23793 = ~1'b0 ;
  assign y23794 = ~1'b0 ;
  assign y23795 = n36316 ;
  assign y23796 = ~n36318 ;
  assign y23797 = ~1'b0 ;
  assign y23798 = ~n36319 ;
  assign y23799 = ~n21105 ;
  assign y23800 = ~1'b0 ;
  assign y23801 = ~1'b0 ;
  assign y23802 = 1'b0 ;
  assign y23803 = ~1'b0 ;
  assign y23804 = n36320 ;
  assign y23805 = ~n36325 ;
  assign y23806 = ~n36329 ;
  assign y23807 = ~1'b0 ;
  assign y23808 = n36331 ;
  assign y23809 = ~n36332 ;
  assign y23810 = n36336 ;
  assign y23811 = ~n36337 ;
  assign y23812 = ~1'b0 ;
  assign y23813 = ~n36342 ;
  assign y23814 = n36347 ;
  assign y23815 = ~1'b0 ;
  assign y23816 = ~1'b0 ;
  assign y23817 = ~1'b0 ;
  assign y23818 = ~n36351 ;
  assign y23819 = ~1'b0 ;
  assign y23820 = n36352 ;
  assign y23821 = ~1'b0 ;
  assign y23822 = ~n36354 ;
  assign y23823 = ~n36357 ;
  assign y23824 = n36358 ;
  assign y23825 = n36362 ;
  assign y23826 = ~n36364 ;
  assign y23827 = n36368 ;
  assign y23828 = ~n5972 ;
  assign y23829 = ~n36371 ;
  assign y23830 = ~n36373 ;
  assign y23831 = ~1'b0 ;
  assign y23832 = ~n415 ;
  assign y23833 = ~n18140 ;
  assign y23834 = ~n36375 ;
  assign y23835 = n36378 ;
  assign y23836 = ~n36379 ;
  assign y23837 = ~1'b0 ;
  assign y23838 = ~n36381 ;
  assign y23839 = 1'b0 ;
  assign y23840 = ~n36385 ;
  assign y23841 = ~n36387 ;
  assign y23842 = ~n10672 ;
  assign y23843 = ~1'b0 ;
  assign y23844 = ~n36389 ;
  assign y23845 = ~n36391 ;
  assign y23846 = ~1'b0 ;
  assign y23847 = 1'b0 ;
  assign y23848 = ~1'b0 ;
  assign y23849 = ~n36392 ;
  assign y23850 = n36393 ;
  assign y23851 = n16600 ;
  assign y23852 = n36395 ;
  assign y23853 = n3376 ;
  assign y23854 = ~1'b0 ;
  assign y23855 = ~1'b0 ;
  assign y23856 = 1'b0 ;
  assign y23857 = n36396 ;
  assign y23858 = n36399 ;
  assign y23859 = n36402 ;
  assign y23860 = ~n36406 ;
  assign y23861 = n36408 ;
  assign y23862 = n27980 ;
  assign y23863 = n36409 ;
  assign y23864 = n36412 ;
  assign y23865 = 1'b0 ;
  assign y23866 = n36413 ;
  assign y23867 = ~1'b0 ;
  assign y23868 = ~n36418 ;
  assign y23869 = n19342 ;
  assign y23870 = ~n33568 ;
  assign y23871 = n36420 ;
  assign y23872 = ~1'b0 ;
  assign y23873 = ~n36422 ;
  assign y23874 = ~n11543 ;
  assign y23875 = n36423 ;
  assign y23876 = ~n36426 ;
  assign y23877 = ~1'b0 ;
  assign y23878 = ~1'b0 ;
  assign y23879 = ~n36429 ;
  assign y23880 = n36430 ;
  assign y23881 = n36431 ;
  assign y23882 = ~n36432 ;
  assign y23883 = ~n16684 ;
  assign y23884 = n36434 ;
  assign y23885 = ~1'b0 ;
  assign y23886 = n28784 ;
  assign y23887 = 1'b0 ;
  assign y23888 = ~n36437 ;
  assign y23889 = ~1'b0 ;
  assign y23890 = n19186 ;
  assign y23891 = ~n36438 ;
  assign y23892 = ~n36439 ;
  assign y23893 = ~n36440 ;
  assign y23894 = ~n36442 ;
  assign y23895 = ~1'b0 ;
  assign y23896 = 1'b0 ;
  assign y23897 = ~1'b0 ;
  assign y23898 = ~1'b0 ;
  assign y23899 = n36444 ;
  assign y23900 = ~1'b0 ;
  assign y23901 = ~n26871 ;
  assign y23902 = ~1'b0 ;
  assign y23903 = n1564 ;
  assign y23904 = n36445 ;
  assign y23905 = ~n36447 ;
  assign y23906 = 1'b0 ;
  assign y23907 = ~n36448 ;
  assign y23908 = n36449 ;
  assign y23909 = ~n36452 ;
  assign y23910 = ~1'b0 ;
  assign y23911 = ~1'b0 ;
  assign y23912 = n36453 ;
  assign y23913 = ~n3950 ;
  assign y23914 = n36455 ;
  assign y23915 = ~n36456 ;
  assign y23916 = ~1'b0 ;
  assign y23917 = n36457 ;
  assign y23918 = ~1'b0 ;
  assign y23919 = n36459 ;
  assign y23920 = ~1'b0 ;
  assign y23921 = n36461 ;
  assign y23922 = ~1'b0 ;
  assign y23923 = ~n6146 ;
  assign y23924 = n36463 ;
  assign y23925 = ~n36465 ;
  assign y23926 = ~n36467 ;
  assign y23927 = ~n36470 ;
  assign y23928 = 1'b0 ;
  assign y23929 = ~1'b0 ;
  assign y23930 = ~1'b0 ;
  assign y23931 = n36472 ;
  assign y23932 = n36476 ;
  assign y23933 = ~n36478 ;
  assign y23934 = ~n36481 ;
  assign y23935 = ~n36482 ;
  assign y23936 = ~n36487 ;
  assign y23937 = ~n36488 ;
  assign y23938 = ~1'b0 ;
  assign y23939 = n36490 ;
  assign y23940 = ~n36491 ;
  assign y23941 = ~1'b0 ;
  assign y23942 = ~n36494 ;
  assign y23943 = ~1'b0 ;
  assign y23944 = ~n36497 ;
  assign y23945 = ~1'b0 ;
  assign y23946 = n36500 ;
  assign y23947 = n1080 ;
  assign y23948 = ~n36510 ;
  assign y23949 = ~n36511 ;
  assign y23950 = ~n36532 ;
  assign y23951 = ~n36533 ;
  assign y23952 = 1'b0 ;
  assign y23953 = ~1'b0 ;
  assign y23954 = n36534 ;
  assign y23955 = ~1'b0 ;
  assign y23956 = n36537 ;
  assign y23957 = ~n36538 ;
  assign y23958 = ~n36539 ;
  assign y23959 = n36542 ;
  assign y23960 = n36543 ;
  assign y23961 = ~1'b0 ;
  assign y23962 = ~1'b0 ;
  assign y23963 = ~1'b0 ;
  assign y23964 = n36546 ;
  assign y23965 = n36551 ;
  assign y23966 = ~1'b0 ;
  assign y23967 = ~1'b0 ;
  assign y23968 = ~1'b0 ;
  assign y23969 = n36553 ;
  assign y23970 = ~1'b0 ;
  assign y23971 = ~n18786 ;
  assign y23972 = 1'b0 ;
  assign y23973 = ~n36562 ;
  assign y23974 = n36565 ;
  assign y23975 = n36567 ;
  assign y23976 = n36568 ;
  assign y23977 = ~1'b0 ;
  assign y23978 = ~1'b0 ;
  assign y23979 = ~n19910 ;
  assign y23980 = ~1'b0 ;
  assign y23981 = ~n36570 ;
  assign y23982 = ~n1657 ;
  assign y23983 = n5462 ;
  assign y23984 = ~1'b0 ;
  assign y23985 = ~n36572 ;
  assign y23986 = ~1'b0 ;
  assign y23987 = ~1'b0 ;
  assign y23988 = n36573 ;
  assign y23989 = 1'b0 ;
  assign y23990 = n36576 ;
  assign y23991 = ~n36578 ;
  assign y23992 = ~n36583 ;
  assign y23993 = ~1'b0 ;
  assign y23994 = 1'b0 ;
  assign y23995 = n36585 ;
  assign y23996 = n36587 ;
  assign y23997 = ~n36591 ;
  assign y23998 = ~1'b0 ;
  assign y23999 = ~n36597 ;
  assign y24000 = n36599 ;
  assign y24001 = ~n36600 ;
  assign y24002 = ~n36601 ;
  assign y24003 = ~1'b0 ;
  assign y24004 = ~n36603 ;
  assign y24005 = ~1'b0 ;
  assign y24006 = ~n36608 ;
  assign y24007 = ~n36612 ;
  assign y24008 = ~1'b0 ;
  assign y24009 = ~1'b0 ;
  assign y24010 = n36613 ;
  assign y24011 = ~1'b0 ;
  assign y24012 = ~n36616 ;
  assign y24013 = n3227 ;
  assign y24014 = ~n36620 ;
  assign y24015 = n36622 ;
  assign y24016 = ~1'b0 ;
  assign y24017 = ~1'b0 ;
  assign y24018 = n36623 ;
  assign y24019 = ~n36625 ;
  assign y24020 = n36627 ;
  assign y24021 = ~n36632 ;
  assign y24022 = ~n36638 ;
  assign y24023 = n36639 ;
  assign y24024 = ~n36643 ;
  assign y24025 = ~1'b0 ;
  assign y24026 = ~1'b0 ;
  assign y24027 = n36644 ;
  assign y24028 = ~1'b0 ;
  assign y24029 = ~1'b0 ;
  assign y24030 = 1'b0 ;
  assign y24031 = ~n36646 ;
  assign y24032 = ~1'b0 ;
  assign y24033 = n36650 ;
  assign y24034 = n36654 ;
  assign y24035 = ~n36656 ;
  assign y24036 = ~n7045 ;
  assign y24037 = ~1'b0 ;
  assign y24038 = ~n36658 ;
  assign y24039 = ~1'b0 ;
  assign y24040 = ~1'b0 ;
  assign y24041 = ~1'b0 ;
  assign y24042 = ~n18253 ;
  assign y24043 = ~1'b0 ;
  assign y24044 = 1'b0 ;
  assign y24045 = ~n22476 ;
  assign y24046 = ~n36660 ;
  assign y24047 = ~1'b0 ;
  assign y24048 = ~n36661 ;
  assign y24049 = n36662 ;
  assign y24050 = ~n36663 ;
  assign y24051 = ~n36666 ;
  assign y24052 = ~n7337 ;
  assign y24053 = n36668 ;
  assign y24054 = ~n36673 ;
  assign y24055 = ~1'b0 ;
  assign y24056 = ~n36674 ;
  assign y24057 = n36675 ;
  assign y24058 = n36679 ;
  assign y24059 = n36684 ;
  assign y24060 = ~n36685 ;
  assign y24061 = ~1'b0 ;
  assign y24062 = ~1'b0 ;
  assign y24063 = n36687 ;
  assign y24064 = ~1'b0 ;
  assign y24065 = n21965 ;
  assign y24066 = ~n36689 ;
  assign y24067 = ~n36693 ;
  assign y24068 = n36696 ;
  assign y24069 = n11895 ;
  assign y24070 = ~n36697 ;
  assign y24071 = ~n11616 ;
  assign y24072 = ~1'b0 ;
  assign y24073 = ~1'b0 ;
  assign y24074 = 1'b0 ;
  assign y24075 = n36701 ;
  assign y24076 = ~1'b0 ;
  assign y24077 = ~1'b0 ;
  assign y24078 = ~1'b0 ;
  assign y24079 = ~1'b0 ;
  assign y24080 = ~n36703 ;
  assign y24081 = ~n13643 ;
  assign y24082 = n36704 ;
  assign y24083 = ~n36707 ;
  assign y24084 = n36708 ;
  assign y24085 = n36709 ;
  assign y24086 = ~n36715 ;
  assign y24087 = ~n36720 ;
  assign y24088 = n36725 ;
  assign y24089 = ~1'b0 ;
  assign y24090 = ~1'b0 ;
  assign y24091 = ~1'b0 ;
  assign y24092 = ~n36728 ;
  assign y24093 = ~n36731 ;
  assign y24094 = n36732 ;
  assign y24095 = ~n1967 ;
  assign y24096 = ~n36735 ;
  assign y24097 = ~n8479 ;
  assign y24098 = ~n36738 ;
  assign y24099 = ~n36740 ;
  assign y24100 = n36744 ;
  assign y24101 = n36752 ;
  assign y24102 = n36754 ;
  assign y24103 = n36755 ;
  assign y24104 = ~1'b0 ;
  assign y24105 = 1'b0 ;
  assign y24106 = n36758 ;
  assign y24107 = 1'b0 ;
  assign y24108 = ~1'b0 ;
  assign y24109 = ~n36761 ;
  assign y24110 = n36763 ;
  assign y24111 = ~n36767 ;
  assign y24112 = ~n36769 ;
  assign y24113 = n36772 ;
  assign y24114 = n36773 ;
  assign y24115 = ~n36774 ;
  assign y24116 = ~n36775 ;
  assign y24117 = ~1'b0 ;
  assign y24118 = ~n36779 ;
  assign y24119 = n36781 ;
  assign y24120 = n6487 ;
  assign y24121 = ~1'b0 ;
  assign y24122 = ~1'b0 ;
  assign y24123 = ~1'b0 ;
  assign y24124 = ~1'b0 ;
  assign y24125 = n7051 ;
  assign y24126 = ~1'b0 ;
  assign y24127 = ~1'b0 ;
  assign y24128 = ~1'b0 ;
  assign y24129 = ~n1696 ;
  assign y24130 = ~n36782 ;
  assign y24131 = n36783 ;
  assign y24132 = ~n36788 ;
  assign y24133 = n10241 ;
  assign y24134 = ~1'b0 ;
  assign y24135 = ~1'b0 ;
  assign y24136 = n36791 ;
  assign y24137 = n36792 ;
  assign y24138 = ~1'b0 ;
  assign y24139 = ~n36795 ;
  assign y24140 = ~n36796 ;
  assign y24141 = ~1'b0 ;
  assign y24142 = ~n36797 ;
  assign y24143 = ~n4278 ;
  assign y24144 = 1'b0 ;
  assign y24145 = ~1'b0 ;
  assign y24146 = ~n36798 ;
  assign y24147 = ~1'b0 ;
  assign y24148 = ~1'b0 ;
  assign y24149 = ~1'b0 ;
  assign y24150 = ~n36799 ;
  assign y24151 = n36800 ;
  assign y24152 = ~n36803 ;
  assign y24153 = ~n36807 ;
  assign y24154 = n36809 ;
  assign y24155 = ~1'b0 ;
  assign y24156 = ~n36811 ;
  assign y24157 = ~n36813 ;
  assign y24158 = n36816 ;
  assign y24159 = n36817 ;
  assign y24160 = ~n633 ;
  assign y24161 = n36818 ;
  assign y24162 = ~n36820 ;
  assign y24163 = n36823 ;
  assign y24164 = ~1'b0 ;
  assign y24165 = ~1'b0 ;
  assign y24166 = ~n36824 ;
  assign y24167 = ~n36825 ;
  assign y24168 = ~1'b0 ;
  assign y24169 = ~n36826 ;
  assign y24170 = ~n36828 ;
  assign y24171 = ~1'b0 ;
  assign y24172 = n36831 ;
  assign y24173 = ~n36832 ;
  assign y24174 = 1'b0 ;
  assign y24175 = ~1'b0 ;
  assign y24176 = n36835 ;
  assign y24177 = n22450 ;
  assign y24178 = ~n36836 ;
  assign y24179 = ~n36838 ;
  assign y24180 = ~n36840 ;
  assign y24181 = ~1'b0 ;
  assign y24182 = 1'b0 ;
  assign y24183 = ~1'b0 ;
  assign y24184 = ~1'b0 ;
  assign y24185 = ~n36841 ;
  assign y24186 = n36846 ;
  assign y24187 = ~1'b0 ;
  assign y24188 = n36847 ;
  assign y24189 = ~n36849 ;
  assign y24190 = n36851 ;
  assign y24191 = ~n36853 ;
  assign y24192 = n36854 ;
  assign y24193 = ~1'b0 ;
  assign y24194 = ~n36855 ;
  assign y24195 = ~1'b0 ;
  assign y24196 = ~1'b0 ;
  assign y24197 = ~n36856 ;
  assign y24198 = ~1'b0 ;
  assign y24199 = n36864 ;
  assign y24200 = ~1'b0 ;
  assign y24201 = n36866 ;
  assign y24202 = ~1'b0 ;
  assign y24203 = ~1'b0 ;
  assign y24204 = ~n21386 ;
  assign y24205 = ~1'b0 ;
  assign y24206 = ~1'b0 ;
  assign y24207 = ~n36868 ;
  assign y24208 = n36871 ;
  assign y24209 = ~n36872 ;
  assign y24210 = ~n36876 ;
  assign y24211 = n36879 ;
  assign y24212 = ~1'b0 ;
  assign y24213 = ~1'b0 ;
  assign y24214 = 1'b0 ;
  assign y24215 = n36883 ;
  assign y24216 = ~n36886 ;
  assign y24217 = ~n4957 ;
  assign y24218 = ~n36889 ;
  assign y24219 = ~n6238 ;
  assign y24220 = n36891 ;
  assign y24221 = ~n36892 ;
  assign y24222 = ~1'b0 ;
  assign y24223 = ~n36895 ;
  assign y24224 = ~n36897 ;
  assign y24225 = ~n36899 ;
  assign y24226 = ~1'b0 ;
  assign y24227 = n36900 ;
  assign y24228 = ~1'b0 ;
  assign y24229 = n36901 ;
  assign y24230 = ~n36908 ;
  assign y24231 = ~1'b0 ;
  assign y24232 = ~n29024 ;
  assign y24233 = ~1'b0 ;
  assign y24234 = n36910 ;
  assign y24235 = ~1'b0 ;
  assign y24236 = ~n36912 ;
  assign y24237 = n36913 ;
  assign y24238 = n36914 ;
  assign y24239 = n36916 ;
  assign y24240 = ~n36921 ;
  assign y24241 = n36927 ;
  assign y24242 = 1'b0 ;
  assign y24243 = ~n36930 ;
  assign y24244 = ~n36931 ;
  assign y24245 = n36933 ;
  assign y24246 = ~1'b0 ;
  assign y24247 = ~1'b0 ;
  assign y24248 = ~n1769 ;
  assign y24249 = ~n36935 ;
  assign y24250 = ~n36936 ;
  assign y24251 = ~n36938 ;
  assign y24252 = ~n36939 ;
  assign y24253 = ~n36944 ;
  assign y24254 = ~1'b0 ;
  assign y24255 = ~n36948 ;
  assign y24256 = n2307 ;
  assign y24257 = ~1'b0 ;
  assign y24258 = n36949 ;
  assign y24259 = ~n36950 ;
  assign y24260 = ~1'b0 ;
  assign y24261 = ~n36951 ;
  assign y24262 = n36953 ;
  assign y24263 = n4315 ;
  assign y24264 = n36955 ;
  assign y24265 = ~1'b0 ;
  assign y24266 = ~n36957 ;
  assign y24267 = ~1'b0 ;
  assign y24268 = ~n20918 ;
  assign y24269 = ~n36962 ;
  assign y24270 = ~n36965 ;
  assign y24271 = n36966 ;
  assign y24272 = ~n36970 ;
  assign y24273 = ~1'b0 ;
  assign y24274 = ~1'b0 ;
  assign y24275 = 1'b0 ;
  assign y24276 = ~n36974 ;
  assign y24277 = ~n36978 ;
  assign y24278 = ~1'b0 ;
  assign y24279 = ~1'b0 ;
  assign y24280 = n36981 ;
  assign y24281 = ~n36984 ;
  assign y24282 = ~1'b0 ;
  assign y24283 = ~n36987 ;
  assign y24284 = ~1'b0 ;
  assign y24285 = ~1'b0 ;
  assign y24286 = ~n36990 ;
  assign y24287 = ~n36992 ;
  assign y24288 = ~n36997 ;
  assign y24289 = ~n37001 ;
  assign y24290 = ~n37002 ;
  assign y24291 = ~1'b0 ;
  assign y24292 = ~1'b0 ;
  assign y24293 = ~1'b0 ;
  assign y24294 = n37003 ;
  assign y24295 = ~n37004 ;
  assign y24296 = n37005 ;
  assign y24297 = ~1'b0 ;
  assign y24298 = ~n37010 ;
  assign y24299 = ~1'b0 ;
  assign y24300 = ~n836 ;
  assign y24301 = ~n37012 ;
  assign y24302 = n15651 ;
  assign y24303 = ~1'b0 ;
  assign y24304 = ~n37014 ;
  assign y24305 = ~n37017 ;
  assign y24306 = ~n37019 ;
  assign y24307 = ~n2325 ;
  assign y24308 = n37020 ;
  assign y24309 = 1'b0 ;
  assign y24310 = n37021 ;
  assign y24311 = ~n37022 ;
  assign y24312 = n37023 ;
  assign y24313 = ~n37025 ;
  assign y24314 = 1'b0 ;
  assign y24315 = 1'b0 ;
  assign y24316 = ~n37027 ;
  assign y24317 = ~1'b0 ;
  assign y24318 = ~1'b0 ;
  assign y24319 = n37028 ;
  assign y24320 = ~n5913 ;
  assign y24321 = n9652 ;
  assign y24322 = ~n37030 ;
  assign y24323 = ~n22174 ;
  assign y24324 = ~n37033 ;
  assign y24325 = 1'b0 ;
  assign y24326 = ~1'b0 ;
  assign y24327 = ~n37034 ;
  assign y24328 = ~1'b0 ;
  assign y24329 = n37035 ;
  assign y24330 = n27144 ;
  assign y24331 = ~n37036 ;
  assign y24332 = ~n37042 ;
  assign y24333 = ~n37044 ;
  assign y24334 = ~n37046 ;
  assign y24335 = ~n37048 ;
  assign y24336 = ~1'b0 ;
  assign y24337 = n37050 ;
  assign y24338 = ~n37052 ;
  assign y24339 = ~1'b0 ;
  assign y24340 = ~n37054 ;
  assign y24341 = ~1'b0 ;
  assign y24342 = n37055 ;
  assign y24343 = n37062 ;
  assign y24344 = 1'b0 ;
  assign y24345 = ~1'b0 ;
  assign y24346 = ~1'b0 ;
  assign y24347 = ~1'b0 ;
  assign y24348 = ~1'b0 ;
  assign y24349 = n5256 ;
  assign y24350 = ~1'b0 ;
  assign y24351 = ~1'b0 ;
  assign y24352 = ~n37063 ;
  assign y24353 = ~n37064 ;
  assign y24354 = ~n37066 ;
  assign y24355 = n37067 ;
  assign y24356 = ~n37070 ;
  assign y24357 = ~n37072 ;
  assign y24358 = ~n8173 ;
  assign y24359 = ~n37074 ;
  assign y24360 = n37075 ;
  assign y24361 = n6271 ;
  assign y24362 = ~1'b0 ;
  assign y24363 = ~1'b0 ;
  assign y24364 = ~n37079 ;
  assign y24365 = n37081 ;
  assign y24366 = ~n37082 ;
  assign y24367 = ~1'b0 ;
  assign y24368 = ~1'b0 ;
  assign y24369 = ~1'b0 ;
  assign y24370 = n37083 ;
  assign y24371 = n37088 ;
  assign y24372 = ~1'b0 ;
  assign y24373 = ~n37091 ;
  assign y24374 = ~1'b0 ;
  assign y24375 = ~n37092 ;
  assign y24376 = ~n37094 ;
  assign y24377 = n37096 ;
  assign y24378 = n11815 ;
  assign y24379 = ~n37098 ;
  assign y24380 = n37100 ;
  assign y24381 = n37101 ;
  assign y24382 = ~n37105 ;
  assign y24383 = ~1'b0 ;
  assign y24384 = ~n37106 ;
  assign y24385 = ~1'b0 ;
  assign y24386 = ~n37107 ;
  assign y24387 = n37108 ;
  assign y24388 = ~1'b0 ;
  assign y24389 = n27089 ;
  assign y24390 = n37109 ;
  assign y24391 = ~n5748 ;
  assign y24392 = n37110 ;
  assign y24393 = 1'b0 ;
  assign y24394 = n37112 ;
  assign y24395 = ~1'b0 ;
  assign y24396 = ~1'b0 ;
  assign y24397 = n37113 ;
  assign y24398 = ~1'b0 ;
  assign y24399 = ~n37114 ;
  assign y24400 = ~1'b0 ;
  assign y24401 = ~n1485 ;
  assign y24402 = ~1'b0 ;
  assign y24403 = n37115 ;
  assign y24404 = ~n8960 ;
  assign y24405 = n22771 ;
  assign y24406 = n37117 ;
  assign y24407 = ~1'b0 ;
  assign y24408 = n37120 ;
  assign y24409 = ~1'b0 ;
  assign y24410 = ~n17182 ;
  assign y24411 = ~1'b0 ;
  assign y24412 = ~1'b0 ;
  assign y24413 = n37122 ;
  assign y24414 = 1'b0 ;
  assign y24415 = ~n37126 ;
  assign y24416 = n37127 ;
  assign y24417 = ~n37137 ;
  assign y24418 = ~n37139 ;
  assign y24419 = n37140 ;
  assign y24420 = ~n37142 ;
  assign y24421 = ~n361 ;
  assign y24422 = ~1'b0 ;
  assign y24423 = ~n37145 ;
  assign y24424 = ~1'b0 ;
  assign y24425 = ~n28297 ;
  assign y24426 = n37146 ;
  assign y24427 = n21358 ;
  assign y24428 = ~1'b0 ;
  assign y24429 = ~n37147 ;
  assign y24430 = n37148 ;
  assign y24431 = ~1'b0 ;
  assign y24432 = ~1'b0 ;
  assign y24433 = ~n2991 ;
  assign y24434 = ~1'b0 ;
  assign y24435 = ~1'b0 ;
  assign y24436 = ~n37149 ;
  assign y24437 = ~n37150 ;
  assign y24438 = n37151 ;
  assign y24439 = ~n37154 ;
  assign y24440 = n37155 ;
  assign y24441 = ~1'b0 ;
  assign y24442 = ~n37156 ;
  assign y24443 = ~1'b0 ;
  assign y24444 = ~1'b0 ;
  assign y24445 = ~n24626 ;
  assign y24446 = ~1'b0 ;
  assign y24447 = ~n37157 ;
  assign y24448 = ~n1857 ;
  assign y24449 = ~1'b0 ;
  assign y24450 = ~1'b0 ;
  assign y24451 = n37159 ;
  assign y24452 = ~n37160 ;
  assign y24453 = ~1'b0 ;
  assign y24454 = ~1'b0 ;
  assign y24455 = ~1'b0 ;
  assign y24456 = n37162 ;
  assign y24457 = ~1'b0 ;
  assign y24458 = ~n37164 ;
  assign y24459 = n37165 ;
  assign y24460 = ~1'b0 ;
  assign y24461 = ~1'b0 ;
  assign y24462 = ~n20626 ;
  assign y24463 = ~1'b0 ;
  assign y24464 = ~n37166 ;
  assign y24465 = ~n37170 ;
  assign y24466 = ~n37172 ;
  assign y24467 = 1'b0 ;
  assign y24468 = ~n37173 ;
  assign y24469 = 1'b0 ;
  assign y24470 = n37175 ;
  assign y24471 = ~1'b0 ;
  assign y24472 = ~1'b0 ;
  assign y24473 = ~n37176 ;
  assign y24474 = ~1'b0 ;
  assign y24475 = n37178 ;
  assign y24476 = ~1'b0 ;
  assign y24477 = n37180 ;
  assign y24478 = ~1'b0 ;
  assign y24479 = ~1'b0 ;
  assign y24480 = n37181 ;
  assign y24481 = ~n37182 ;
  assign y24482 = n37184 ;
  assign y24483 = ~1'b0 ;
  assign y24484 = n37185 ;
  assign y24485 = n37186 ;
  assign y24486 = n37187 ;
  assign y24487 = ~1'b0 ;
  assign y24488 = n37188 ;
  assign y24489 = ~1'b0 ;
  assign y24490 = n37190 ;
  assign y24491 = ~1'b0 ;
  assign y24492 = ~n37192 ;
  assign y24493 = ~1'b0 ;
  assign y24494 = n5717 ;
  assign y24495 = n37194 ;
  assign y24496 = ~n37195 ;
  assign y24497 = 1'b0 ;
  assign y24498 = ~n37197 ;
  assign y24499 = n37200 ;
  assign y24500 = ~1'b0 ;
  assign y24501 = ~1'b0 ;
  assign y24502 = ~n37202 ;
  assign y24503 = ~n37205 ;
  assign y24504 = ~1'b0 ;
  assign y24505 = ~1'b0 ;
  assign y24506 = n6647 ;
  assign y24507 = ~n37207 ;
  assign y24508 = n37210 ;
  assign y24509 = ~n37213 ;
  assign y24510 = ~1'b0 ;
  assign y24511 = ~n37214 ;
  assign y24512 = ~n5675 ;
  assign y24513 = n37216 ;
  assign y24514 = ~1'b0 ;
  assign y24515 = n37218 ;
  assign y24516 = n37219 ;
  assign y24517 = n37221 ;
  assign y24518 = ~n37223 ;
  assign y24519 = ~n37225 ;
  assign y24520 = ~1'b0 ;
  assign y24521 = ~1'b0 ;
  assign y24522 = n8663 ;
  assign y24523 = ~1'b0 ;
  assign y24524 = ~1'b0 ;
  assign y24525 = ~n37226 ;
  assign y24526 = ~1'b0 ;
  assign y24527 = ~1'b0 ;
  assign y24528 = n37227 ;
  assign y24529 = n37228 ;
  assign y24530 = n37230 ;
  assign y24531 = ~n37231 ;
  assign y24532 = ~n37233 ;
  assign y24533 = ~1'b0 ;
  assign y24534 = ~1'b0 ;
  assign y24535 = ~n37234 ;
  assign y24536 = n37235 ;
  assign y24537 = n37239 ;
  assign y24538 = ~1'b0 ;
  assign y24539 = n37241 ;
  assign y24540 = n37242 ;
  assign y24541 = ~1'b0 ;
  assign y24542 = ~1'b0 ;
  assign y24543 = ~1'b0 ;
  assign y24544 = 1'b0 ;
  assign y24545 = n37243 ;
  assign y24546 = ~n29567 ;
  assign y24547 = n37244 ;
  assign y24548 = ~n37246 ;
  assign y24549 = ~1'b0 ;
  assign y24550 = ~n18105 ;
  assign y24551 = ~n37248 ;
  assign y24552 = ~n37249 ;
  assign y24553 = ~1'b0 ;
  assign y24554 = ~n37252 ;
  assign y24555 = ~1'b0 ;
  assign y24556 = n37255 ;
  assign y24557 = n37262 ;
  assign y24558 = ~n37264 ;
  assign y24559 = ~1'b0 ;
  assign y24560 = ~n24821 ;
  assign y24561 = ~n37265 ;
  assign y24562 = n37267 ;
  assign y24563 = ~n37269 ;
  assign y24564 = ~n37274 ;
  assign y24565 = ~1'b0 ;
  assign y24566 = ~1'b0 ;
  assign y24567 = ~1'b0 ;
  assign y24568 = n37279 ;
  assign y24569 = ~1'b0 ;
  assign y24570 = ~n37281 ;
  assign y24571 = ~n37284 ;
  assign y24572 = n37285 ;
  assign y24573 = ~n37286 ;
  assign y24574 = ~n37288 ;
  assign y24575 = ~1'b0 ;
  assign y24576 = n37291 ;
  assign y24577 = ~1'b0 ;
  assign y24578 = ~n37293 ;
  assign y24579 = ~n37294 ;
  assign y24580 = ~1'b0 ;
  assign y24581 = ~n37296 ;
  assign y24582 = ~n37300 ;
  assign y24583 = ~1'b0 ;
  assign y24584 = ~1'b0 ;
  assign y24585 = ~1'b0 ;
  assign y24586 = n37302 ;
  assign y24587 = ~1'b0 ;
  assign y24588 = ~1'b0 ;
  assign y24589 = ~n37303 ;
  assign y24590 = n37304 ;
  assign y24591 = 1'b0 ;
  assign y24592 = ~n37306 ;
  assign y24593 = n37307 ;
  assign y24594 = ~1'b0 ;
  assign y24595 = ~n37308 ;
  assign y24596 = n37310 ;
  assign y24597 = ~n37311 ;
  assign y24598 = ~1'b0 ;
  assign y24599 = ~n37313 ;
  assign y24600 = 1'b0 ;
  assign y24601 = ~n37322 ;
  assign y24602 = ~n37326 ;
  assign y24603 = ~1'b0 ;
  assign y24604 = n37328 ;
  assign y24605 = ~n37329 ;
  assign y24606 = n37330 ;
  assign y24607 = ~n37341 ;
  assign y24608 = n37342 ;
  assign y24609 = ~1'b0 ;
  assign y24610 = n37344 ;
  assign y24611 = ~n37347 ;
  assign y24612 = ~n27104 ;
  assign y24613 = ~n37349 ;
  assign y24614 = n37352 ;
  assign y24615 = n4301 ;
  assign y24616 = ~n37354 ;
  assign y24617 = ~n14238 ;
  assign y24618 = n37356 ;
  assign y24619 = ~1'b0 ;
  assign y24620 = ~n37358 ;
  assign y24621 = ~n37359 ;
  assign y24622 = ~n37360 ;
  assign y24623 = n37026 ;
  assign y24624 = n37361 ;
  assign y24625 = ~1'b0 ;
  assign y24626 = n8750 ;
  assign y24627 = ~n37362 ;
  assign y24628 = ~1'b0 ;
  assign y24629 = ~n37366 ;
  assign y24630 = ~n37367 ;
  assign y24631 = n37370 ;
  assign y24632 = n37371 ;
  assign y24633 = ~n37376 ;
  assign y24634 = ~n37378 ;
  assign y24635 = ~1'b0 ;
  assign y24636 = 1'b0 ;
  assign y24637 = n37380 ;
  assign y24638 = ~1'b0 ;
  assign y24639 = n37382 ;
  assign y24640 = ~n37384 ;
  assign y24641 = ~n37385 ;
  assign y24642 = ~n7522 ;
  assign y24643 = ~1'b0 ;
  assign y24644 = n37391 ;
  assign y24645 = ~n1521 ;
  assign y24646 = n37392 ;
  assign y24647 = ~n37393 ;
  assign y24648 = n15363 ;
  assign y24649 = n37395 ;
  assign y24650 = n37396 ;
  assign y24651 = ~n6850 ;
  assign y24652 = ~1'b0 ;
  assign y24653 = ~1'b0 ;
  assign y24654 = 1'b0 ;
  assign y24655 = n37402 ;
  assign y24656 = ~n37404 ;
  assign y24657 = ~n31139 ;
  assign y24658 = ~1'b0 ;
  assign y24659 = ~1'b0 ;
  assign y24660 = 1'b0 ;
  assign y24661 = ~n37409 ;
  assign y24662 = ~1'b0 ;
  assign y24663 = 1'b0 ;
  assign y24664 = n37414 ;
  assign y24665 = n37415 ;
  assign y24666 = ~n37416 ;
  assign y24667 = ~n37420 ;
  assign y24668 = ~n37429 ;
  assign y24669 = n3776 ;
  assign y24670 = ~1'b0 ;
  assign y24671 = n17209 ;
  assign y24672 = n11689 ;
  assign y24673 = ~n37432 ;
  assign y24674 = 1'b0 ;
  assign y24675 = ~1'b0 ;
  assign y24676 = ~1'b0 ;
  assign y24677 = n37437 ;
  assign y24678 = n37438 ;
  assign y24679 = ~1'b0 ;
  assign y24680 = ~1'b0 ;
  assign y24681 = n37439 ;
  assign y24682 = ~1'b0 ;
  assign y24683 = n37441 ;
  assign y24684 = ~n37442 ;
  assign y24685 = ~1'b0 ;
  assign y24686 = ~n16015 ;
  assign y24687 = ~1'b0 ;
  assign y24688 = ~n37443 ;
  assign y24689 = n37447 ;
  assign y24690 = ~n37448 ;
  assign y24691 = n37449 ;
  assign y24692 = ~n37450 ;
  assign y24693 = ~1'b0 ;
  assign y24694 = ~1'b0 ;
  assign y24695 = ~1'b0 ;
  assign y24696 = n37452 ;
  assign y24697 = n33801 ;
  assign y24698 = ~n37454 ;
  assign y24699 = ~n37457 ;
  assign y24700 = n37460 ;
  assign y24701 = ~1'b0 ;
  assign y24702 = ~1'b0 ;
  assign y24703 = n37462 ;
  assign y24704 = ~n37463 ;
  assign y24705 = ~1'b0 ;
  assign y24706 = ~1'b0 ;
  assign y24707 = n37464 ;
  assign y24708 = ~n37466 ;
  assign y24709 = 1'b0 ;
  assign y24710 = n37469 ;
  assign y24711 = ~1'b0 ;
  assign y24712 = ~1'b0 ;
  assign y24713 = ~n37471 ;
  assign y24714 = 1'b0 ;
  assign y24715 = ~1'b0 ;
  assign y24716 = ~1'b0 ;
  assign y24717 = ~n37474 ;
  assign y24718 = n14997 ;
  assign y24719 = n37475 ;
  assign y24720 = ~n37477 ;
  assign y24721 = ~n37479 ;
  assign y24722 = ~n5106 ;
  assign y24723 = ~n37481 ;
  assign y24724 = ~n37482 ;
  assign y24725 = ~1'b0 ;
  assign y24726 = ~n37484 ;
  assign y24727 = ~n37485 ;
  assign y24728 = n37486 ;
  assign y24729 = n11695 ;
  assign y24730 = ~1'b0 ;
  assign y24731 = n37489 ;
  assign y24732 = n37490 ;
  assign y24733 = ~n37491 ;
  assign y24734 = ~n37492 ;
  assign y24735 = ~n37493 ;
  assign y24736 = ~1'b0 ;
  assign y24737 = ~n37495 ;
  assign y24738 = ~n37496 ;
  assign y24739 = ~n37502 ;
  assign y24740 = n37504 ;
  assign y24741 = ~n37512 ;
  assign y24742 = n37513 ;
  assign y24743 = n16101 ;
  assign y24744 = ~1'b0 ;
  assign y24745 = ~1'b0 ;
  assign y24746 = 1'b0 ;
  assign y24747 = n37518 ;
  assign y24748 = ~n37520 ;
  assign y24749 = ~1'b0 ;
  assign y24750 = 1'b0 ;
  assign y24751 = ~1'b0 ;
  assign y24752 = ~n37522 ;
  assign y24753 = ~1'b0 ;
  assign y24754 = ~1'b0 ;
  assign y24755 = ~1'b0 ;
  assign y24756 = n37524 ;
  assign y24757 = n37525 ;
  assign y24758 = ~1'b0 ;
  assign y24759 = ~n37527 ;
  assign y24760 = ~n37530 ;
  assign y24761 = ~1'b0 ;
  assign y24762 = ~1'b0 ;
  assign y24763 = n37531 ;
  assign y24764 = n37532 ;
  assign y24765 = ~n20194 ;
  assign y24766 = n37534 ;
  assign y24767 = n37537 ;
  assign y24768 = n10965 ;
  assign y24769 = n37539 ;
  assign y24770 = n37541 ;
  assign y24771 = n37543 ;
  assign y24772 = ~n37545 ;
  assign y24773 = ~n37546 ;
  assign y24774 = n37547 ;
  assign y24775 = ~1'b0 ;
  assign y24776 = n26277 ;
  assign y24777 = ~1'b0 ;
  assign y24778 = n37548 ;
  assign y24779 = n37549 ;
  assign y24780 = ~n37557 ;
  assign y24781 = ~1'b0 ;
  assign y24782 = ~n5996 ;
  assign y24783 = n14112 ;
  assign y24784 = ~n37559 ;
  assign y24785 = n37561 ;
  assign y24786 = ~n36669 ;
  assign y24787 = ~n32521 ;
  assign y24788 = n37563 ;
  assign y24789 = n36330 ;
  assign y24790 = n37564 ;
  assign y24791 = n37565 ;
  assign y24792 = n37566 ;
  assign y24793 = ~n37567 ;
  assign y24794 = n37570 ;
  assign y24795 = 1'b0 ;
  assign y24796 = n29329 ;
  assign y24797 = n37571 ;
  assign y24798 = ~1'b0 ;
  assign y24799 = n37576 ;
  assign y24800 = ~n37577 ;
  assign y24801 = ~n37578 ;
  assign y24802 = n37579 ;
  assign y24803 = ~1'b0 ;
  assign y24804 = ~1'b0 ;
  assign y24805 = ~n37581 ;
  assign y24806 = ~1'b0 ;
  assign y24807 = ~1'b0 ;
  assign y24808 = n37582 ;
  assign y24809 = ~1'b0 ;
  assign y24810 = n37584 ;
  assign y24811 = ~n37585 ;
  assign y24812 = n37587 ;
  assign y24813 = ~1'b0 ;
  assign y24814 = ~n37588 ;
  assign y24815 = ~n37589 ;
  assign y24816 = ~n529 ;
  assign y24817 = ~1'b0 ;
  assign y24818 = ~n37591 ;
  assign y24819 = ~n1158 ;
  assign y24820 = ~n12797 ;
  assign y24821 = ~1'b0 ;
  assign y24822 = n30931 ;
  assign y24823 = n37592 ;
  assign y24824 = n37593 ;
  assign y24825 = ~n37595 ;
  assign y24826 = n11724 ;
  assign y24827 = ~1'b0 ;
  assign y24828 = n37597 ;
  assign y24829 = ~n37600 ;
  assign y24830 = ~n24898 ;
  assign y24831 = n37603 ;
  assign y24832 = ~n18994 ;
  assign y24833 = n37606 ;
  assign y24834 = n37608 ;
  assign y24835 = ~1'b0 ;
  assign y24836 = n37612 ;
  assign y24837 = ~1'b0 ;
  assign y24838 = n37613 ;
  assign y24839 = ~1'b0 ;
  assign y24840 = ~1'b0 ;
  assign y24841 = 1'b0 ;
  assign y24842 = ~n22408 ;
  assign y24843 = n37616 ;
  assign y24844 = n37617 ;
  assign y24845 = ~n37620 ;
  assign y24846 = n37622 ;
  assign y24847 = ~n37627 ;
  assign y24848 = n37628 ;
  assign y24849 = ~n37629 ;
  assign y24850 = n37633 ;
  assign y24851 = n37635 ;
  assign y24852 = ~n37637 ;
  assign y24853 = ~1'b0 ;
  assign y24854 = ~1'b0 ;
  assign y24855 = ~n37639 ;
  assign y24856 = ~1'b0 ;
  assign y24857 = ~n37640 ;
  assign y24858 = ~n37642 ;
  assign y24859 = ~1'b0 ;
  assign y24860 = ~n37644 ;
  assign y24861 = ~1'b0 ;
  assign y24862 = ~n37645 ;
  assign y24863 = ~1'b0 ;
  assign y24864 = n37647 ;
  assign y24865 = ~1'b0 ;
  assign y24866 = ~n3013 ;
  assign y24867 = n37648 ;
  assign y24868 = ~n37649 ;
  assign y24869 = ~1'b0 ;
  assign y24870 = ~n37651 ;
  assign y24871 = n37652 ;
  assign y24872 = n37654 ;
  assign y24873 = n37657 ;
  assign y24874 = ~n37662 ;
  assign y24875 = ~n37664 ;
  assign y24876 = n37666 ;
  assign y24877 = ~1'b0 ;
  assign y24878 = ~1'b0 ;
  assign y24879 = n37669 ;
  assign y24880 = n37673 ;
  assign y24881 = ~n37675 ;
  assign y24882 = ~n37676 ;
  assign y24883 = ~1'b0 ;
  assign y24884 = n37678 ;
  assign y24885 = ~n37682 ;
  assign y24886 = ~1'b0 ;
  assign y24887 = ~1'b0 ;
  assign y24888 = n37690 ;
  assign y24889 = ~1'b0 ;
  assign y24890 = ~1'b0 ;
  assign y24891 = 1'b0 ;
  assign y24892 = ~1'b0 ;
  assign y24893 = n2322 ;
  assign y24894 = ~1'b0 ;
  assign y24895 = ~1'b0 ;
  assign y24896 = ~n37693 ;
  assign y24897 = n17226 ;
  assign y24898 = ~1'b0 ;
  assign y24899 = n37697 ;
  assign y24900 = n37700 ;
  assign y24901 = n37704 ;
  assign y24902 = ~1'b0 ;
  assign y24903 = n37706 ;
  assign y24904 = n37709 ;
  assign y24905 = ~n37711 ;
  assign y24906 = n37713 ;
  assign y24907 = ~1'b0 ;
  assign y24908 = ~n37716 ;
  assign y24909 = ~n37718 ;
  assign y24910 = ~1'b0 ;
  assign y24911 = ~n37720 ;
  assign y24912 = ~1'b0 ;
  assign y24913 = ~n37723 ;
  assign y24914 = ~1'b0 ;
  assign y24915 = ~n37724 ;
  assign y24916 = n37728 ;
  assign y24917 = ~1'b0 ;
  assign y24918 = n37730 ;
  assign y24919 = ~1'b0 ;
  assign y24920 = n9652 ;
  assign y24921 = ~1'b0 ;
  assign y24922 = n37732 ;
endmodule
